
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h1f858708;
    ram_cell[       1] = 32'h0;  // 32'h2a9fb276;
    ram_cell[       2] = 32'h0;  // 32'h33634e48;
    ram_cell[       3] = 32'h0;  // 32'hdd19a913;
    ram_cell[       4] = 32'h0;  // 32'h0dcc0027;
    ram_cell[       5] = 32'h0;  // 32'h746ca6a6;
    ram_cell[       6] = 32'h0;  // 32'h85aec632;
    ram_cell[       7] = 32'h0;  // 32'h1a9b0ff1;
    ram_cell[       8] = 32'h0;  // 32'h28ab8708;
    ram_cell[       9] = 32'h0;  // 32'h54486e5a;
    ram_cell[      10] = 32'h0;  // 32'h6cef3c90;
    ram_cell[      11] = 32'h0;  // 32'hfd70577e;
    ram_cell[      12] = 32'h0;  // 32'ha43d3024;
    ram_cell[      13] = 32'h0;  // 32'he133ee6d;
    ram_cell[      14] = 32'h0;  // 32'h5e36ce1b;
    ram_cell[      15] = 32'h0;  // 32'h3d880172;
    ram_cell[      16] = 32'h0;  // 32'h7bd09799;
    ram_cell[      17] = 32'h0;  // 32'h8933ddbd;
    ram_cell[      18] = 32'h0;  // 32'h395ec8d6;
    ram_cell[      19] = 32'h0;  // 32'h652ffe5d;
    ram_cell[      20] = 32'h0;  // 32'h29dff6c4;
    ram_cell[      21] = 32'h0;  // 32'hd49da5be;
    ram_cell[      22] = 32'h0;  // 32'h64d56989;
    ram_cell[      23] = 32'h0;  // 32'hee72efbd;
    ram_cell[      24] = 32'h0;  // 32'h44ab3afa;
    ram_cell[      25] = 32'h0;  // 32'h800570a5;
    ram_cell[      26] = 32'h0;  // 32'hb70bf48a;
    ram_cell[      27] = 32'h0;  // 32'h5a2925e3;
    ram_cell[      28] = 32'h0;  // 32'h1119be85;
    ram_cell[      29] = 32'h0;  // 32'haadcaca7;
    ram_cell[      30] = 32'h0;  // 32'h9681af6f;
    ram_cell[      31] = 32'h0;  // 32'h17676c52;
    ram_cell[      32] = 32'h0;  // 32'hee07ab3a;
    ram_cell[      33] = 32'h0;  // 32'h483f6bfa;
    ram_cell[      34] = 32'h0;  // 32'h9734c419;
    ram_cell[      35] = 32'h0;  // 32'h3522708a;
    ram_cell[      36] = 32'h0;  // 32'h691c3d98;
    ram_cell[      37] = 32'h0;  // 32'hc57b3748;
    ram_cell[      38] = 32'h0;  // 32'h8ed7504f;
    ram_cell[      39] = 32'h0;  // 32'h4c7c0b2e;
    ram_cell[      40] = 32'h0;  // 32'h3b4b50b1;
    ram_cell[      41] = 32'h0;  // 32'h2d36ac42;
    ram_cell[      42] = 32'h0;  // 32'hef5a08b8;
    ram_cell[      43] = 32'h0;  // 32'ha6745686;
    ram_cell[      44] = 32'h0;  // 32'hcee49c0d;
    ram_cell[      45] = 32'h0;  // 32'h821ed5d4;
    ram_cell[      46] = 32'h0;  // 32'h6ebf9300;
    ram_cell[      47] = 32'h0;  // 32'h5f77db99;
    ram_cell[      48] = 32'h0;  // 32'h4c9c6305;
    ram_cell[      49] = 32'h0;  // 32'h22e63964;
    ram_cell[      50] = 32'h0;  // 32'hecfc3823;
    ram_cell[      51] = 32'h0;  // 32'hdbba52af;
    ram_cell[      52] = 32'h0;  // 32'h27426745;
    ram_cell[      53] = 32'h0;  // 32'hec91e82a;
    ram_cell[      54] = 32'h0;  // 32'h3c717b07;
    ram_cell[      55] = 32'h0;  // 32'hbcf5ac45;
    ram_cell[      56] = 32'h0;  // 32'h000cf119;
    ram_cell[      57] = 32'h0;  // 32'h289d9f37;
    ram_cell[      58] = 32'h0;  // 32'h41708524;
    ram_cell[      59] = 32'h0;  // 32'h658432a9;
    ram_cell[      60] = 32'h0;  // 32'hb6690e53;
    ram_cell[      61] = 32'h0;  // 32'h03c374c3;
    ram_cell[      62] = 32'h0;  // 32'h25a6eea3;
    ram_cell[      63] = 32'h0;  // 32'he88efeaf;
    ram_cell[      64] = 32'h0;  // 32'h817891b3;
    ram_cell[      65] = 32'h0;  // 32'h60db3a73;
    ram_cell[      66] = 32'h0;  // 32'he36fe980;
    ram_cell[      67] = 32'h0;  // 32'ha7421e55;
    ram_cell[      68] = 32'h0;  // 32'haac59018;
    ram_cell[      69] = 32'h0;  // 32'hab5cb5e6;
    ram_cell[      70] = 32'h0;  // 32'habfe34f2;
    ram_cell[      71] = 32'h0;  // 32'he207b6ed;
    ram_cell[      72] = 32'h0;  // 32'h60d36d25;
    ram_cell[      73] = 32'h0;  // 32'hbbc72548;
    ram_cell[      74] = 32'h0;  // 32'h9fb276b7;
    ram_cell[      75] = 32'h0;  // 32'hc3fa9806;
    ram_cell[      76] = 32'h0;  // 32'h238fa943;
    ram_cell[      77] = 32'h0;  // 32'hbc669815;
    ram_cell[      78] = 32'h0;  // 32'hc86124c5;
    ram_cell[      79] = 32'h0;  // 32'h785cf631;
    ram_cell[      80] = 32'h0;  // 32'h39947dc6;
    ram_cell[      81] = 32'h0;  // 32'hfab3d3c2;
    ram_cell[      82] = 32'h0;  // 32'h1de628b6;
    ram_cell[      83] = 32'h0;  // 32'h3e2ab314;
    ram_cell[      84] = 32'h0;  // 32'hc5dc2112;
    ram_cell[      85] = 32'h0;  // 32'h8794145b;
    ram_cell[      86] = 32'h0;  // 32'hfba5d4f3;
    ram_cell[      87] = 32'h0;  // 32'h20d0dc29;
    ram_cell[      88] = 32'h0;  // 32'h883f5bc6;
    ram_cell[      89] = 32'h0;  // 32'h49aa9e9a;
    ram_cell[      90] = 32'h0;  // 32'h616ca4e1;
    ram_cell[      91] = 32'h0;  // 32'hba093aa4;
    ram_cell[      92] = 32'h0;  // 32'he7974fbf;
    ram_cell[      93] = 32'h0;  // 32'h4251ef08;
    ram_cell[      94] = 32'h0;  // 32'hf2add520;
    ram_cell[      95] = 32'h0;  // 32'h49d89105;
    ram_cell[      96] = 32'h0;  // 32'h65c03f92;
    ram_cell[      97] = 32'h0;  // 32'haefb33be;
    ram_cell[      98] = 32'h0;  // 32'h3b7e8ee7;
    ram_cell[      99] = 32'h0;  // 32'h503b3415;
    ram_cell[     100] = 32'h0;  // 32'h469e596d;
    ram_cell[     101] = 32'h0;  // 32'h246872b6;
    ram_cell[     102] = 32'h0;  // 32'h5a25e720;
    ram_cell[     103] = 32'h0;  // 32'hf736e753;
    ram_cell[     104] = 32'h0;  // 32'h3619bf57;
    ram_cell[     105] = 32'h0;  // 32'hb9c45919;
    ram_cell[     106] = 32'h0;  // 32'h8b422463;
    ram_cell[     107] = 32'h0;  // 32'h657d44e3;
    ram_cell[     108] = 32'h0;  // 32'h49f5209b;
    ram_cell[     109] = 32'h0;  // 32'h96a66d48;
    ram_cell[     110] = 32'h0;  // 32'hcd6c5b0c;
    ram_cell[     111] = 32'h0;  // 32'h32f2217a;
    ram_cell[     112] = 32'h0;  // 32'he52c32bf;
    ram_cell[     113] = 32'h0;  // 32'h744f47fd;
    ram_cell[     114] = 32'h0;  // 32'hd78c63fb;
    ram_cell[     115] = 32'h0;  // 32'h8cc4ba26;
    ram_cell[     116] = 32'h0;  // 32'ha0cf7a66;
    ram_cell[     117] = 32'h0;  // 32'h3dcf14fa;
    ram_cell[     118] = 32'h0;  // 32'h5cddacd4;
    ram_cell[     119] = 32'h0;  // 32'ha325b232;
    ram_cell[     120] = 32'h0;  // 32'hee32f321;
    ram_cell[     121] = 32'h0;  // 32'h81fa2055;
    ram_cell[     122] = 32'h0;  // 32'h642598e7;
    ram_cell[     123] = 32'h0;  // 32'hbcb207a9;
    ram_cell[     124] = 32'h0;  // 32'h8e733675;
    ram_cell[     125] = 32'h0;  // 32'h855942f8;
    ram_cell[     126] = 32'h0;  // 32'h6b175d94;
    ram_cell[     127] = 32'h0;  // 32'h2c25ef9d;
    ram_cell[     128] = 32'h0;  // 32'hf40212b4;
    ram_cell[     129] = 32'h0;  // 32'h889b000c;
    ram_cell[     130] = 32'h0;  // 32'ha60f503e;
    ram_cell[     131] = 32'h0;  // 32'h4aca0454;
    ram_cell[     132] = 32'h0;  // 32'ha7a88412;
    ram_cell[     133] = 32'h0;  // 32'hf8ff75d2;
    ram_cell[     134] = 32'h0;  // 32'he1be2e42;
    ram_cell[     135] = 32'h0;  // 32'h1d4eb0cc;
    ram_cell[     136] = 32'h0;  // 32'hbc8574b2;
    ram_cell[     137] = 32'h0;  // 32'h7493decd;
    ram_cell[     138] = 32'h0;  // 32'heae33b7a;
    ram_cell[     139] = 32'h0;  // 32'h991f5b6c;
    ram_cell[     140] = 32'h0;  // 32'hae512b7b;
    ram_cell[     141] = 32'h0;  // 32'h5fe09f70;
    ram_cell[     142] = 32'h0;  // 32'h8580e4ab;
    ram_cell[     143] = 32'h0;  // 32'h4fda4ddc;
    ram_cell[     144] = 32'h0;  // 32'h99c4a00a;
    ram_cell[     145] = 32'h0;  // 32'h8e74eda8;
    ram_cell[     146] = 32'h0;  // 32'he33015d8;
    ram_cell[     147] = 32'h0;  // 32'hbfe4044a;
    ram_cell[     148] = 32'h0;  // 32'hf354152d;
    ram_cell[     149] = 32'h0;  // 32'h536db453;
    ram_cell[     150] = 32'h0;  // 32'h129d3ba7;
    ram_cell[     151] = 32'h0;  // 32'h0bbcd055;
    ram_cell[     152] = 32'h0;  // 32'h74bbd7ea;
    ram_cell[     153] = 32'h0;  // 32'ha660e662;
    ram_cell[     154] = 32'h0;  // 32'hd31a4eb3;
    ram_cell[     155] = 32'h0;  // 32'h1a2efd83;
    ram_cell[     156] = 32'h0;  // 32'h15e6e9f5;
    ram_cell[     157] = 32'h0;  // 32'h2c5af7d8;
    ram_cell[     158] = 32'h0;  // 32'h53629967;
    ram_cell[     159] = 32'h0;  // 32'h60b37612;
    ram_cell[     160] = 32'h0;  // 32'h27c24ac3;
    ram_cell[     161] = 32'h0;  // 32'h11f01390;
    ram_cell[     162] = 32'h0;  // 32'h043e11e6;
    ram_cell[     163] = 32'h0;  // 32'h2194f4fc;
    ram_cell[     164] = 32'h0;  // 32'h9561ff24;
    ram_cell[     165] = 32'h0;  // 32'h95d34540;
    ram_cell[     166] = 32'h0;  // 32'h6bc62636;
    ram_cell[     167] = 32'h0;  // 32'ha0c5b0f8;
    ram_cell[     168] = 32'h0;  // 32'hb6dbe572;
    ram_cell[     169] = 32'h0;  // 32'h9380af2e;
    ram_cell[     170] = 32'h0;  // 32'h54ca4275;
    ram_cell[     171] = 32'h0;  // 32'h19dbc8bc;
    ram_cell[     172] = 32'h0;  // 32'h76651e9d;
    ram_cell[     173] = 32'h0;  // 32'h72868f84;
    ram_cell[     174] = 32'h0;  // 32'h1ce47ff5;
    ram_cell[     175] = 32'h0;  // 32'h048b31ac;
    ram_cell[     176] = 32'h0;  // 32'h0d456e12;
    ram_cell[     177] = 32'h0;  // 32'h652c0ddc;
    ram_cell[     178] = 32'h0;  // 32'hc56c6b40;
    ram_cell[     179] = 32'h0;  // 32'hd2c00427;
    ram_cell[     180] = 32'h0;  // 32'hcf24808a;
    ram_cell[     181] = 32'h0;  // 32'h4bbf9e6a;
    ram_cell[     182] = 32'h0;  // 32'h2218a386;
    ram_cell[     183] = 32'h0;  // 32'hc7ee5bbf;
    ram_cell[     184] = 32'h0;  // 32'h93257797;
    ram_cell[     185] = 32'h0;  // 32'h99e6e38b;
    ram_cell[     186] = 32'h0;  // 32'h7de70bd4;
    ram_cell[     187] = 32'h0;  // 32'h2d20c9b7;
    ram_cell[     188] = 32'h0;  // 32'h96f18a3e;
    ram_cell[     189] = 32'h0;  // 32'h2cdf153b;
    ram_cell[     190] = 32'h0;  // 32'h0b8ecba6;
    ram_cell[     191] = 32'h0;  // 32'h91b61a26;
    ram_cell[     192] = 32'h0;  // 32'he64255ea;
    ram_cell[     193] = 32'h0;  // 32'hdcad5195;
    ram_cell[     194] = 32'h0;  // 32'h24a51684;
    ram_cell[     195] = 32'h0;  // 32'h98dabdee;
    ram_cell[     196] = 32'h0;  // 32'h48405ea5;
    ram_cell[     197] = 32'h0;  // 32'ha505a49c;
    ram_cell[     198] = 32'h0;  // 32'h2102e1f6;
    ram_cell[     199] = 32'h0;  // 32'h04669b51;
    ram_cell[     200] = 32'h0;  // 32'h8f21620d;
    ram_cell[     201] = 32'h0;  // 32'had3227af;
    ram_cell[     202] = 32'h0;  // 32'h21ae503a;
    ram_cell[     203] = 32'h0;  // 32'h04ea378a;
    ram_cell[     204] = 32'h0;  // 32'h126d1d6a;
    ram_cell[     205] = 32'h0;  // 32'h26268d70;
    ram_cell[     206] = 32'h0;  // 32'hefac8772;
    ram_cell[     207] = 32'h0;  // 32'h1d9d4f04;
    ram_cell[     208] = 32'h0;  // 32'hc89eb82b;
    ram_cell[     209] = 32'h0;  // 32'h1ddee48a;
    ram_cell[     210] = 32'h0;  // 32'h4672cb1c;
    ram_cell[     211] = 32'h0;  // 32'h68e34a4d;
    ram_cell[     212] = 32'h0;  // 32'h6a1025aa;
    ram_cell[     213] = 32'h0;  // 32'h724a4673;
    ram_cell[     214] = 32'h0;  // 32'h08503c17;
    ram_cell[     215] = 32'h0;  // 32'hdd3c2cee;
    ram_cell[     216] = 32'h0;  // 32'h68dd93e4;
    ram_cell[     217] = 32'h0;  // 32'ha7754671;
    ram_cell[     218] = 32'h0;  // 32'h0a1a4f4b;
    ram_cell[     219] = 32'h0;  // 32'he687c570;
    ram_cell[     220] = 32'h0;  // 32'h8d2b0a54;
    ram_cell[     221] = 32'h0;  // 32'h838a0a83;
    ram_cell[     222] = 32'h0;  // 32'ha802595f;
    ram_cell[     223] = 32'h0;  // 32'hb3971bf5;
    ram_cell[     224] = 32'h0;  // 32'h1421f6b7;
    ram_cell[     225] = 32'h0;  // 32'h0a4fc8a7;
    ram_cell[     226] = 32'h0;  // 32'h202d62e6;
    ram_cell[     227] = 32'h0;  // 32'h23e434b0;
    ram_cell[     228] = 32'h0;  // 32'h0227df78;
    ram_cell[     229] = 32'h0;  // 32'h226b48d0;
    ram_cell[     230] = 32'h0;  // 32'hcf95f190;
    ram_cell[     231] = 32'h0;  // 32'h81c5df81;
    ram_cell[     232] = 32'h0;  // 32'h0282797f;
    ram_cell[     233] = 32'h0;  // 32'hef3b0c82;
    ram_cell[     234] = 32'h0;  // 32'h34914769;
    ram_cell[     235] = 32'h0;  // 32'h855d479d;
    ram_cell[     236] = 32'h0;  // 32'h4f1fed7a;
    ram_cell[     237] = 32'h0;  // 32'h1145bee9;
    ram_cell[     238] = 32'h0;  // 32'h1e7be6c1;
    ram_cell[     239] = 32'h0;  // 32'ha8863473;
    ram_cell[     240] = 32'h0;  // 32'h10c2328b;
    ram_cell[     241] = 32'h0;  // 32'hd8de53fc;
    ram_cell[     242] = 32'h0;  // 32'h1395c22a;
    ram_cell[     243] = 32'h0;  // 32'h828fa930;
    ram_cell[     244] = 32'h0;  // 32'hb560ea1f;
    ram_cell[     245] = 32'h0;  // 32'h7612a7b6;
    ram_cell[     246] = 32'h0;  // 32'hf38e2376;
    ram_cell[     247] = 32'h0;  // 32'hd5f0c9a9;
    ram_cell[     248] = 32'h0;  // 32'hb90fa738;
    ram_cell[     249] = 32'h0;  // 32'hb94265c8;
    ram_cell[     250] = 32'h0;  // 32'h3e0d034d;
    ram_cell[     251] = 32'h0;  // 32'h3f30d7e4;
    ram_cell[     252] = 32'h0;  // 32'h4803a52d;
    ram_cell[     253] = 32'h0;  // 32'h420d457e;
    ram_cell[     254] = 32'h0;  // 32'hceaac279;
    ram_cell[     255] = 32'h0;  // 32'hd49bfc60;
    // src matrix A
    ram_cell[     256] = 32'h422845d1;
    ram_cell[     257] = 32'h8fa2c9dc;
    ram_cell[     258] = 32'h6ea92762;
    ram_cell[     259] = 32'h40dba90b;
    ram_cell[     260] = 32'hd55d49bf;
    ram_cell[     261] = 32'h8e6edbfb;
    ram_cell[     262] = 32'h4bb83d21;
    ram_cell[     263] = 32'h5d7878d1;
    ram_cell[     264] = 32'h50abf79c;
    ram_cell[     265] = 32'h765e8097;
    ram_cell[     266] = 32'hbb44b5d2;
    ram_cell[     267] = 32'h1b022b69;
    ram_cell[     268] = 32'h06eabff8;
    ram_cell[     269] = 32'he243b7d2;
    ram_cell[     270] = 32'hed3d58a1;
    ram_cell[     271] = 32'h5981938d;
    ram_cell[     272] = 32'h6cb877e7;
    ram_cell[     273] = 32'h349a12a7;
    ram_cell[     274] = 32'h0d91de6a;
    ram_cell[     275] = 32'ha3f00953;
    ram_cell[     276] = 32'hd6442566;
    ram_cell[     277] = 32'h4e08b69f;
    ram_cell[     278] = 32'h759a0749;
    ram_cell[     279] = 32'he13ed256;
    ram_cell[     280] = 32'h748d4f4f;
    ram_cell[     281] = 32'h13d1b066;
    ram_cell[     282] = 32'h88a167c1;
    ram_cell[     283] = 32'hf7a9110c;
    ram_cell[     284] = 32'h539d0642;
    ram_cell[     285] = 32'h88a3af76;
    ram_cell[     286] = 32'h8865e328;
    ram_cell[     287] = 32'h34d86515;
    ram_cell[     288] = 32'h52c5fefa;
    ram_cell[     289] = 32'h25d0b9f9;
    ram_cell[     290] = 32'h718deb3c;
    ram_cell[     291] = 32'h3ee6eaa4;
    ram_cell[     292] = 32'hbff68c3d;
    ram_cell[     293] = 32'h309778b5;
    ram_cell[     294] = 32'hb347ab2d;
    ram_cell[     295] = 32'h76d2fffb;
    ram_cell[     296] = 32'h41f34359;
    ram_cell[     297] = 32'h2339024c;
    ram_cell[     298] = 32'h08bc15ba;
    ram_cell[     299] = 32'h620d4ff8;
    ram_cell[     300] = 32'hd2709882;
    ram_cell[     301] = 32'h6cec4607;
    ram_cell[     302] = 32'h136bf513;
    ram_cell[     303] = 32'h5f5adcc6;
    ram_cell[     304] = 32'h04aaa837;
    ram_cell[     305] = 32'h182a2670;
    ram_cell[     306] = 32'hcbb08182;
    ram_cell[     307] = 32'hdd9854a7;
    ram_cell[     308] = 32'h5db8e687;
    ram_cell[     309] = 32'hc176154a;
    ram_cell[     310] = 32'h79090a07;
    ram_cell[     311] = 32'h26bab0ce;
    ram_cell[     312] = 32'h9e964ff1;
    ram_cell[     313] = 32'h9ac9d093;
    ram_cell[     314] = 32'h60c3b4d8;
    ram_cell[     315] = 32'ha60d11ea;
    ram_cell[     316] = 32'h2b50ae6c;
    ram_cell[     317] = 32'h1cd557f9;
    ram_cell[     318] = 32'h25bc10cd;
    ram_cell[     319] = 32'h15c7f7cb;
    ram_cell[     320] = 32'he072db68;
    ram_cell[     321] = 32'h5675f4f1;
    ram_cell[     322] = 32'hdb35d908;
    ram_cell[     323] = 32'h58fa73fe;
    ram_cell[     324] = 32'h68796669;
    ram_cell[     325] = 32'hab156c2c;
    ram_cell[     326] = 32'h2f42d38f;
    ram_cell[     327] = 32'h62c26f1c;
    ram_cell[     328] = 32'h8333d726;
    ram_cell[     329] = 32'hdc73ccdc;
    ram_cell[     330] = 32'h5a3e3082;
    ram_cell[     331] = 32'h7343e7d4;
    ram_cell[     332] = 32'hb64b7bfc;
    ram_cell[     333] = 32'hd4d78b53;
    ram_cell[     334] = 32'hbc220025;
    ram_cell[     335] = 32'h72a21de4;
    ram_cell[     336] = 32'h6f157b5f;
    ram_cell[     337] = 32'ha6f410f0;
    ram_cell[     338] = 32'h4270d9b6;
    ram_cell[     339] = 32'hed27946f;
    ram_cell[     340] = 32'hd2b96b39;
    ram_cell[     341] = 32'h675c9668;
    ram_cell[     342] = 32'hd64916f9;
    ram_cell[     343] = 32'hc72601b8;
    ram_cell[     344] = 32'h8ddf8d8e;
    ram_cell[     345] = 32'h94c7aaba;
    ram_cell[     346] = 32'h5b4705d4;
    ram_cell[     347] = 32'hc8928325;
    ram_cell[     348] = 32'hfdb8792a;
    ram_cell[     349] = 32'h44a78fcc;
    ram_cell[     350] = 32'hf3d3eb2c;
    ram_cell[     351] = 32'h1eef0416;
    ram_cell[     352] = 32'hc1d0d82c;
    ram_cell[     353] = 32'hd72fe1e0;
    ram_cell[     354] = 32'h5be07ac9;
    ram_cell[     355] = 32'h99e47f84;
    ram_cell[     356] = 32'he84abb92;
    ram_cell[     357] = 32'h6c14e4b8;
    ram_cell[     358] = 32'hcbdd2fa8;
    ram_cell[     359] = 32'h491a456a;
    ram_cell[     360] = 32'h2a10c4d6;
    ram_cell[     361] = 32'h0cfaafd6;
    ram_cell[     362] = 32'h38457a28;
    ram_cell[     363] = 32'h3ed0640c;
    ram_cell[     364] = 32'hcc624b4d;
    ram_cell[     365] = 32'h07edad78;
    ram_cell[     366] = 32'h57a9cb83;
    ram_cell[     367] = 32'hab33896a;
    ram_cell[     368] = 32'h69f798e1;
    ram_cell[     369] = 32'h530cd3c4;
    ram_cell[     370] = 32'hede998b7;
    ram_cell[     371] = 32'hec1686cc;
    ram_cell[     372] = 32'h1dfe0cb7;
    ram_cell[     373] = 32'hfe5f8ad7;
    ram_cell[     374] = 32'hfda60474;
    ram_cell[     375] = 32'h4a5988dc;
    ram_cell[     376] = 32'h9060a4b0;
    ram_cell[     377] = 32'ha3aa011d;
    ram_cell[     378] = 32'h5a47c467;
    ram_cell[     379] = 32'h408cd11f;
    ram_cell[     380] = 32'hcbed8d12;
    ram_cell[     381] = 32'h423ea334;
    ram_cell[     382] = 32'h57047a2a;
    ram_cell[     383] = 32'h956e3a61;
    ram_cell[     384] = 32'hdefbd5a2;
    ram_cell[     385] = 32'hed86b598;
    ram_cell[     386] = 32'hec66f9ef;
    ram_cell[     387] = 32'h8b41b24b;
    ram_cell[     388] = 32'h774f6d3c;
    ram_cell[     389] = 32'h098e5848;
    ram_cell[     390] = 32'h377d9323;
    ram_cell[     391] = 32'hab2b96f0;
    ram_cell[     392] = 32'h1a832174;
    ram_cell[     393] = 32'h84c9e579;
    ram_cell[     394] = 32'h18d36222;
    ram_cell[     395] = 32'hcd4d99bd;
    ram_cell[     396] = 32'h6f18ed0b;
    ram_cell[     397] = 32'h6f4430e4;
    ram_cell[     398] = 32'h2449b96b;
    ram_cell[     399] = 32'h76ae34ba;
    ram_cell[     400] = 32'h04a8954a;
    ram_cell[     401] = 32'hb285c179;
    ram_cell[     402] = 32'h0778a5d0;
    ram_cell[     403] = 32'h22ceab44;
    ram_cell[     404] = 32'h149fe07c;
    ram_cell[     405] = 32'ha0d306bb;
    ram_cell[     406] = 32'h37989e0c;
    ram_cell[     407] = 32'hacceaa8d;
    ram_cell[     408] = 32'hcd2e1d58;
    ram_cell[     409] = 32'h3ac93fd2;
    ram_cell[     410] = 32'hb6b808ba;
    ram_cell[     411] = 32'h962eb268;
    ram_cell[     412] = 32'h8893aed7;
    ram_cell[     413] = 32'h7eeea1f6;
    ram_cell[     414] = 32'h0428ea0f;
    ram_cell[     415] = 32'hd729ae58;
    ram_cell[     416] = 32'h295754e6;
    ram_cell[     417] = 32'h1d6f9797;
    ram_cell[     418] = 32'h797b9f93;
    ram_cell[     419] = 32'hf582d8c1;
    ram_cell[     420] = 32'h6ca84bc0;
    ram_cell[     421] = 32'hf7519727;
    ram_cell[     422] = 32'h363e8e0e;
    ram_cell[     423] = 32'h734fa244;
    ram_cell[     424] = 32'h1a87cf97;
    ram_cell[     425] = 32'h41ebb5a3;
    ram_cell[     426] = 32'h070bdee6;
    ram_cell[     427] = 32'h0607a5e7;
    ram_cell[     428] = 32'ha80bf5a4;
    ram_cell[     429] = 32'hb3645297;
    ram_cell[     430] = 32'hc048caad;
    ram_cell[     431] = 32'h9f24efac;
    ram_cell[     432] = 32'hc7043eec;
    ram_cell[     433] = 32'h7a8fe1ab;
    ram_cell[     434] = 32'h30a45c90;
    ram_cell[     435] = 32'h1a5af16f;
    ram_cell[     436] = 32'h3e64b4e8;
    ram_cell[     437] = 32'h2ce98b30;
    ram_cell[     438] = 32'h1407de7c;
    ram_cell[     439] = 32'hd5700560;
    ram_cell[     440] = 32'h97a1d1bb;
    ram_cell[     441] = 32'h286c4d9d;
    ram_cell[     442] = 32'h19ec98c7;
    ram_cell[     443] = 32'h9ea21566;
    ram_cell[     444] = 32'h3700f258;
    ram_cell[     445] = 32'h4a24523b;
    ram_cell[     446] = 32'h345d7575;
    ram_cell[     447] = 32'hf0c0abde;
    ram_cell[     448] = 32'h64074f1c;
    ram_cell[     449] = 32'h027c389f;
    ram_cell[     450] = 32'h58b890d6;
    ram_cell[     451] = 32'h8d267612;
    ram_cell[     452] = 32'hfc330161;
    ram_cell[     453] = 32'hc3d643aa;
    ram_cell[     454] = 32'h76885bec;
    ram_cell[     455] = 32'hf08971de;
    ram_cell[     456] = 32'h89b21539;
    ram_cell[     457] = 32'hb5e4f88f;
    ram_cell[     458] = 32'h2d3f4b64;
    ram_cell[     459] = 32'h1fc03742;
    ram_cell[     460] = 32'h3d4d2a9b;
    ram_cell[     461] = 32'h9e2cf51f;
    ram_cell[     462] = 32'habe12e3e;
    ram_cell[     463] = 32'hb71c51b9;
    ram_cell[     464] = 32'he37235db;
    ram_cell[     465] = 32'h1ed641d9;
    ram_cell[     466] = 32'h1cdf6863;
    ram_cell[     467] = 32'hb805fb3e;
    ram_cell[     468] = 32'ha55bb743;
    ram_cell[     469] = 32'h364a3248;
    ram_cell[     470] = 32'h37f85110;
    ram_cell[     471] = 32'h119df0ab;
    ram_cell[     472] = 32'haf1ffd73;
    ram_cell[     473] = 32'h218eaf61;
    ram_cell[     474] = 32'h6a96250c;
    ram_cell[     475] = 32'h2b5df1f6;
    ram_cell[     476] = 32'h90341f45;
    ram_cell[     477] = 32'h58c8b126;
    ram_cell[     478] = 32'h3c369a55;
    ram_cell[     479] = 32'ha28444ca;
    ram_cell[     480] = 32'h49b0c22c;
    ram_cell[     481] = 32'h5e1d1c0f;
    ram_cell[     482] = 32'h13aab7dc;
    ram_cell[     483] = 32'h3f2cd37f;
    ram_cell[     484] = 32'h0660f2a8;
    ram_cell[     485] = 32'hb687afeb;
    ram_cell[     486] = 32'h5d3f2919;
    ram_cell[     487] = 32'h974706e8;
    ram_cell[     488] = 32'h0a10e197;
    ram_cell[     489] = 32'hfec68dc0;
    ram_cell[     490] = 32'h11d99f9a;
    ram_cell[     491] = 32'h39a3dca4;
    ram_cell[     492] = 32'h2a1b11a3;
    ram_cell[     493] = 32'hce9b975f;
    ram_cell[     494] = 32'h93016994;
    ram_cell[     495] = 32'h21fef287;
    ram_cell[     496] = 32'hdebba339;
    ram_cell[     497] = 32'h8ca9ef62;
    ram_cell[     498] = 32'hf42e90fd;
    ram_cell[     499] = 32'h4f9ee48b;
    ram_cell[     500] = 32'h7cff2170;
    ram_cell[     501] = 32'h5ca1d52d;
    ram_cell[     502] = 32'hd18b4f20;
    ram_cell[     503] = 32'ha6c2cc28;
    ram_cell[     504] = 32'h43cd1e0e;
    ram_cell[     505] = 32'h6da61eb1;
    ram_cell[     506] = 32'he68e6728;
    ram_cell[     507] = 32'h544f8872;
    ram_cell[     508] = 32'h76c45e0f;
    ram_cell[     509] = 32'ha61c2852;
    ram_cell[     510] = 32'h51f33f56;
    ram_cell[     511] = 32'hbb2a2405;
    // src matrix B
    ram_cell[     512] = 32'he651e029;
    ram_cell[     513] = 32'hf00d6513;
    ram_cell[     514] = 32'hc7b35891;
    ram_cell[     515] = 32'h32108e56;
    ram_cell[     516] = 32'hc8f59979;
    ram_cell[     517] = 32'hbcd42b7c;
    ram_cell[     518] = 32'haecaf813;
    ram_cell[     519] = 32'hf1bd15b7;
    ram_cell[     520] = 32'h43f09a44;
    ram_cell[     521] = 32'h5474d3e9;
    ram_cell[     522] = 32'hbbdd943f;
    ram_cell[     523] = 32'h0a149677;
    ram_cell[     524] = 32'h997a28b1;
    ram_cell[     525] = 32'hcb002af5;
    ram_cell[     526] = 32'h465abc33;
    ram_cell[     527] = 32'h0483b3d3;
    ram_cell[     528] = 32'h3f64fa6e;
    ram_cell[     529] = 32'h25b6fbe1;
    ram_cell[     530] = 32'h58365862;
    ram_cell[     531] = 32'h2fa82142;
    ram_cell[     532] = 32'h753da530;
    ram_cell[     533] = 32'h01b28e6a;
    ram_cell[     534] = 32'h95b3b144;
    ram_cell[     535] = 32'h137dd37a;
    ram_cell[     536] = 32'he8f8a2b7;
    ram_cell[     537] = 32'hd32d4acf;
    ram_cell[     538] = 32'h89baa8e2;
    ram_cell[     539] = 32'h485a3bd6;
    ram_cell[     540] = 32'h87879fde;
    ram_cell[     541] = 32'hd9de7a12;
    ram_cell[     542] = 32'h7cf115ba;
    ram_cell[     543] = 32'he83cadb5;
    ram_cell[     544] = 32'hb981c864;
    ram_cell[     545] = 32'h3beec1e2;
    ram_cell[     546] = 32'h0c874d66;
    ram_cell[     547] = 32'h3e68e89f;
    ram_cell[     548] = 32'h8316c92f;
    ram_cell[     549] = 32'h5376108d;
    ram_cell[     550] = 32'hdf937c9f;
    ram_cell[     551] = 32'hd94274e3;
    ram_cell[     552] = 32'h4ef3f35c;
    ram_cell[     553] = 32'he437e55a;
    ram_cell[     554] = 32'hecb722c7;
    ram_cell[     555] = 32'h3ee342a0;
    ram_cell[     556] = 32'h0047aaf9;
    ram_cell[     557] = 32'he5436068;
    ram_cell[     558] = 32'h37891376;
    ram_cell[     559] = 32'h0351a3b9;
    ram_cell[     560] = 32'he8f10634;
    ram_cell[     561] = 32'hca2cce82;
    ram_cell[     562] = 32'hf2b63620;
    ram_cell[     563] = 32'h69c31118;
    ram_cell[     564] = 32'h65931353;
    ram_cell[     565] = 32'h21ee8bc1;
    ram_cell[     566] = 32'h822ece4b;
    ram_cell[     567] = 32'h0e6c087a;
    ram_cell[     568] = 32'h9869120e;
    ram_cell[     569] = 32'h435935ed;
    ram_cell[     570] = 32'h324c12ba;
    ram_cell[     571] = 32'h55ed7fd2;
    ram_cell[     572] = 32'h2dcc5a83;
    ram_cell[     573] = 32'hd9d0e1d8;
    ram_cell[     574] = 32'h947df66d;
    ram_cell[     575] = 32'h7e364b09;
    ram_cell[     576] = 32'h61452167;
    ram_cell[     577] = 32'hbe2c1be3;
    ram_cell[     578] = 32'h5bd8b2e2;
    ram_cell[     579] = 32'hb27d6768;
    ram_cell[     580] = 32'hf4cf4e3d;
    ram_cell[     581] = 32'h134d9a05;
    ram_cell[     582] = 32'h4b90ee47;
    ram_cell[     583] = 32'h9ad297af;
    ram_cell[     584] = 32'h08c70603;
    ram_cell[     585] = 32'h96c541df;
    ram_cell[     586] = 32'h5874cdb7;
    ram_cell[     587] = 32'h287c150d;
    ram_cell[     588] = 32'hfce8782a;
    ram_cell[     589] = 32'h2f4a366e;
    ram_cell[     590] = 32'hb0d16250;
    ram_cell[     591] = 32'hc0527a6b;
    ram_cell[     592] = 32'h504750a2;
    ram_cell[     593] = 32'h2df8f496;
    ram_cell[     594] = 32'hfb952689;
    ram_cell[     595] = 32'ha2bae61e;
    ram_cell[     596] = 32'hf050f194;
    ram_cell[     597] = 32'h79dd6922;
    ram_cell[     598] = 32'h6bf25695;
    ram_cell[     599] = 32'he35bd5a4;
    ram_cell[     600] = 32'hc6195df9;
    ram_cell[     601] = 32'h1b54000d;
    ram_cell[     602] = 32'hdd9ba121;
    ram_cell[     603] = 32'h781e7edc;
    ram_cell[     604] = 32'h20a74fec;
    ram_cell[     605] = 32'h4d424a58;
    ram_cell[     606] = 32'hd2d06255;
    ram_cell[     607] = 32'h5846ed55;
    ram_cell[     608] = 32'h46a3c47a;
    ram_cell[     609] = 32'h24ff32f1;
    ram_cell[     610] = 32'h233b1401;
    ram_cell[     611] = 32'h1935b0ef;
    ram_cell[     612] = 32'haaea066e;
    ram_cell[     613] = 32'h8385b198;
    ram_cell[     614] = 32'h72f28cf2;
    ram_cell[     615] = 32'hd1140c49;
    ram_cell[     616] = 32'ha5d448d8;
    ram_cell[     617] = 32'h4ef0565c;
    ram_cell[     618] = 32'hb5f58bc3;
    ram_cell[     619] = 32'hdc8c12db;
    ram_cell[     620] = 32'h79f5d353;
    ram_cell[     621] = 32'h0098a222;
    ram_cell[     622] = 32'hdc474453;
    ram_cell[     623] = 32'ha48190f5;
    ram_cell[     624] = 32'hb7f7834a;
    ram_cell[     625] = 32'he0dcf6d3;
    ram_cell[     626] = 32'he94e5e1c;
    ram_cell[     627] = 32'hb57a5ac8;
    ram_cell[     628] = 32'hd87ecf5f;
    ram_cell[     629] = 32'hea1bd9b4;
    ram_cell[     630] = 32'h63df0395;
    ram_cell[     631] = 32'hee52ddad;
    ram_cell[     632] = 32'h088cec3f;
    ram_cell[     633] = 32'h6db55951;
    ram_cell[     634] = 32'hb633477a;
    ram_cell[     635] = 32'h451ac508;
    ram_cell[     636] = 32'hafe6cb1d;
    ram_cell[     637] = 32'hc2ac5e6e;
    ram_cell[     638] = 32'h6e390588;
    ram_cell[     639] = 32'h5b2111e5;
    ram_cell[     640] = 32'hb06fa453;
    ram_cell[     641] = 32'ha0b9e178;
    ram_cell[     642] = 32'h8cbcf860;
    ram_cell[     643] = 32'hc24baf13;
    ram_cell[     644] = 32'h91a9204f;
    ram_cell[     645] = 32'hc36413de;
    ram_cell[     646] = 32'hfaf0e5d3;
    ram_cell[     647] = 32'hed54a8a8;
    ram_cell[     648] = 32'h478846ca;
    ram_cell[     649] = 32'hab874ae6;
    ram_cell[     650] = 32'h4824465c;
    ram_cell[     651] = 32'h099b4376;
    ram_cell[     652] = 32'hb4331663;
    ram_cell[     653] = 32'hc036afc5;
    ram_cell[     654] = 32'hf7722cb8;
    ram_cell[     655] = 32'h56257ddc;
    ram_cell[     656] = 32'hf26041a0;
    ram_cell[     657] = 32'h4706d676;
    ram_cell[     658] = 32'he424507a;
    ram_cell[     659] = 32'h332b7c51;
    ram_cell[     660] = 32'hdf3eeb85;
    ram_cell[     661] = 32'he9ae143e;
    ram_cell[     662] = 32'h21755897;
    ram_cell[     663] = 32'h4430637a;
    ram_cell[     664] = 32'he6335448;
    ram_cell[     665] = 32'hcf3db570;
    ram_cell[     666] = 32'h9050cb52;
    ram_cell[     667] = 32'h432077fd;
    ram_cell[     668] = 32'h1bb56544;
    ram_cell[     669] = 32'h853db15d;
    ram_cell[     670] = 32'h7209d88a;
    ram_cell[     671] = 32'hdf201b4b;
    ram_cell[     672] = 32'h609bced3;
    ram_cell[     673] = 32'h11a0cf09;
    ram_cell[     674] = 32'hb86d87a3;
    ram_cell[     675] = 32'ha9712aad;
    ram_cell[     676] = 32'h723600ee;
    ram_cell[     677] = 32'h8a42797a;
    ram_cell[     678] = 32'h399d4c0c;
    ram_cell[     679] = 32'h33a026cc;
    ram_cell[     680] = 32'hd666ac03;
    ram_cell[     681] = 32'h74e6abab;
    ram_cell[     682] = 32'hab24ad2d;
    ram_cell[     683] = 32'h33a7b6fe;
    ram_cell[     684] = 32'h750891c8;
    ram_cell[     685] = 32'hc265f094;
    ram_cell[     686] = 32'hd52fb485;
    ram_cell[     687] = 32'h62758125;
    ram_cell[     688] = 32'h30aa35b0;
    ram_cell[     689] = 32'h797cdb15;
    ram_cell[     690] = 32'h6fd99128;
    ram_cell[     691] = 32'hef35a619;
    ram_cell[     692] = 32'h75a26bad;
    ram_cell[     693] = 32'h439ad923;
    ram_cell[     694] = 32'he701ff34;
    ram_cell[     695] = 32'hf11ca922;
    ram_cell[     696] = 32'h23ecd6c9;
    ram_cell[     697] = 32'ha292f3dd;
    ram_cell[     698] = 32'h1d8355d0;
    ram_cell[     699] = 32'h547a3e01;
    ram_cell[     700] = 32'h7a843bc4;
    ram_cell[     701] = 32'h9b501977;
    ram_cell[     702] = 32'h2482e05b;
    ram_cell[     703] = 32'h8367f3c5;
    ram_cell[     704] = 32'hfa94fb0c;
    ram_cell[     705] = 32'hbb32dd4c;
    ram_cell[     706] = 32'h2d4d8eca;
    ram_cell[     707] = 32'h6934d384;
    ram_cell[     708] = 32'h734cae2a;
    ram_cell[     709] = 32'h0b27a835;
    ram_cell[     710] = 32'h6cf66652;
    ram_cell[     711] = 32'hd61a52ba;
    ram_cell[     712] = 32'hcfa64d80;
    ram_cell[     713] = 32'hfa8b6ffb;
    ram_cell[     714] = 32'h4e90efb0;
    ram_cell[     715] = 32'h8d226431;
    ram_cell[     716] = 32'hac2e416b;
    ram_cell[     717] = 32'hfbcc7ca1;
    ram_cell[     718] = 32'h4abcfe4c;
    ram_cell[     719] = 32'hda1e3a85;
    ram_cell[     720] = 32'he28de1ac;
    ram_cell[     721] = 32'hbce2d00e;
    ram_cell[     722] = 32'h6ade90d0;
    ram_cell[     723] = 32'hef6f6784;
    ram_cell[     724] = 32'h9da27e9b;
    ram_cell[     725] = 32'h8612e801;
    ram_cell[     726] = 32'h8f04adca;
    ram_cell[     727] = 32'hde660895;
    ram_cell[     728] = 32'hbd2cb5a8;
    ram_cell[     729] = 32'h19826632;
    ram_cell[     730] = 32'hd3137c81;
    ram_cell[     731] = 32'h39430184;
    ram_cell[     732] = 32'h5ce8ae63;
    ram_cell[     733] = 32'ha164c33e;
    ram_cell[     734] = 32'h253ac5f6;
    ram_cell[     735] = 32'h0b252286;
    ram_cell[     736] = 32'hecc585be;
    ram_cell[     737] = 32'h956a01e6;
    ram_cell[     738] = 32'h8ff69f95;
    ram_cell[     739] = 32'h312655f2;
    ram_cell[     740] = 32'h613373ea;
    ram_cell[     741] = 32'hdbd81748;
    ram_cell[     742] = 32'h7ea0f225;
    ram_cell[     743] = 32'h5ff253ca;
    ram_cell[     744] = 32'h461bfb9d;
    ram_cell[     745] = 32'hfb3294f4;
    ram_cell[     746] = 32'h5d62b8f2;
    ram_cell[     747] = 32'h04c11ffe;
    ram_cell[     748] = 32'h3f2814d3;
    ram_cell[     749] = 32'h814aa711;
    ram_cell[     750] = 32'hd684753c;
    ram_cell[     751] = 32'h286a1078;
    ram_cell[     752] = 32'hcca5acaa;
    ram_cell[     753] = 32'h22f2e433;
    ram_cell[     754] = 32'h5af88676;
    ram_cell[     755] = 32'ha1b8452c;
    ram_cell[     756] = 32'h61627fff;
    ram_cell[     757] = 32'hf2505751;
    ram_cell[     758] = 32'h4657843d;
    ram_cell[     759] = 32'h3583f2c9;
    ram_cell[     760] = 32'h7ea674d9;
    ram_cell[     761] = 32'hf78529c0;
    ram_cell[     762] = 32'h7c373c2e;
    ram_cell[     763] = 32'hc4391987;
    ram_cell[     764] = 32'hb1ca2f03;
    ram_cell[     765] = 32'h9b68e863;
    ram_cell[     766] = 32'hae0df40a;
    ram_cell[     767] = 32'hddebdc84;
end

endmodule

