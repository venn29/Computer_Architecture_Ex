
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hf8a29831;
    ram_cell[       1] = 32'h0;  // 32'hccc4f6b6;
    ram_cell[       2] = 32'h0;  // 32'h376d85ae;
    ram_cell[       3] = 32'h0;  // 32'h8b972b43;
    ram_cell[       4] = 32'h0;  // 32'h5596c4cf;
    ram_cell[       5] = 32'h0;  // 32'hdc803125;
    ram_cell[       6] = 32'h0;  // 32'h90e97d2b;
    ram_cell[       7] = 32'h0;  // 32'h510a3303;
    ram_cell[       8] = 32'h0;  // 32'h19a5a37a;
    ram_cell[       9] = 32'h0;  // 32'hfe20c023;
    ram_cell[      10] = 32'h0;  // 32'hf66e8d98;
    ram_cell[      11] = 32'h0;  // 32'h01ecff3c;
    ram_cell[      12] = 32'h0;  // 32'he95297e2;
    ram_cell[      13] = 32'h0;  // 32'ha51be022;
    ram_cell[      14] = 32'h0;  // 32'hfc22a6a9;
    ram_cell[      15] = 32'h0;  // 32'hf294b6f2;
    ram_cell[      16] = 32'h0;  // 32'h579015a7;
    ram_cell[      17] = 32'h0;  // 32'hcbb1dba8;
    ram_cell[      18] = 32'h0;  // 32'h3b6699de;
    ram_cell[      19] = 32'h0;  // 32'hcc656ea8;
    ram_cell[      20] = 32'h0;  // 32'h4a9f044b;
    ram_cell[      21] = 32'h0;  // 32'hbe44804c;
    ram_cell[      22] = 32'h0;  // 32'h6614c047;
    ram_cell[      23] = 32'h0;  // 32'h2278e45a;
    ram_cell[      24] = 32'h0;  // 32'h3d363e04;
    ram_cell[      25] = 32'h0;  // 32'h17930a06;
    ram_cell[      26] = 32'h0;  // 32'h8f42fdc5;
    ram_cell[      27] = 32'h0;  // 32'h48b110d8;
    ram_cell[      28] = 32'h0;  // 32'h3adfe6b9;
    ram_cell[      29] = 32'h0;  // 32'h795b7548;
    ram_cell[      30] = 32'h0;  // 32'hcb149081;
    ram_cell[      31] = 32'h0;  // 32'hce69dcef;
    ram_cell[      32] = 32'h0;  // 32'he6c00adc;
    ram_cell[      33] = 32'h0;  // 32'h3e9224f1;
    ram_cell[      34] = 32'h0;  // 32'h796c62c2;
    ram_cell[      35] = 32'h0;  // 32'h85f78f66;
    ram_cell[      36] = 32'h0;  // 32'h78b42140;
    ram_cell[      37] = 32'h0;  // 32'hcb5cacd5;
    ram_cell[      38] = 32'h0;  // 32'h57eb424a;
    ram_cell[      39] = 32'h0;  // 32'h4ebe1480;
    ram_cell[      40] = 32'h0;  // 32'hd16e4e59;
    ram_cell[      41] = 32'h0;  // 32'hd2f4f42d;
    ram_cell[      42] = 32'h0;  // 32'hbc2d87e3;
    ram_cell[      43] = 32'h0;  // 32'h23ccedcb;
    ram_cell[      44] = 32'h0;  // 32'hfb1e51cb;
    ram_cell[      45] = 32'h0;  // 32'hd7ffe749;
    ram_cell[      46] = 32'h0;  // 32'h730071ac;
    ram_cell[      47] = 32'h0;  // 32'hc68ff6ab;
    ram_cell[      48] = 32'h0;  // 32'ha7000d83;
    ram_cell[      49] = 32'h0;  // 32'h67e59f9a;
    ram_cell[      50] = 32'h0;  // 32'h3d51aaac;
    ram_cell[      51] = 32'h0;  // 32'ha0249cc1;
    ram_cell[      52] = 32'h0;  // 32'hf6a4f25f;
    ram_cell[      53] = 32'h0;  // 32'h289cca85;
    ram_cell[      54] = 32'h0;  // 32'he924d7ba;
    ram_cell[      55] = 32'h0;  // 32'hcd6cc9dc;
    ram_cell[      56] = 32'h0;  // 32'hcb270ef7;
    ram_cell[      57] = 32'h0;  // 32'h67c5902a;
    ram_cell[      58] = 32'h0;  // 32'h7bed43a0;
    ram_cell[      59] = 32'h0;  // 32'h067b4bfb;
    ram_cell[      60] = 32'h0;  // 32'hc9e9a0fb;
    ram_cell[      61] = 32'h0;  // 32'hc4fcd880;
    ram_cell[      62] = 32'h0;  // 32'hbfba6612;
    ram_cell[      63] = 32'h0;  // 32'h3a9114f8;
    ram_cell[      64] = 32'h0;  // 32'hed933bb7;
    ram_cell[      65] = 32'h0;  // 32'hb87ca46b;
    ram_cell[      66] = 32'h0;  // 32'h18dce0d8;
    ram_cell[      67] = 32'h0;  // 32'hdef87e89;
    ram_cell[      68] = 32'h0;  // 32'h5c6db246;
    ram_cell[      69] = 32'h0;  // 32'h68680cd9;
    ram_cell[      70] = 32'h0;  // 32'h492aed8f;
    ram_cell[      71] = 32'h0;  // 32'h2fd9c3f5;
    ram_cell[      72] = 32'h0;  // 32'h8490057a;
    ram_cell[      73] = 32'h0;  // 32'h0c61c7ad;
    ram_cell[      74] = 32'h0;  // 32'he8f3741f;
    ram_cell[      75] = 32'h0;  // 32'hb85e5856;
    ram_cell[      76] = 32'h0;  // 32'h754de21b;
    ram_cell[      77] = 32'h0;  // 32'h9d36628b;
    ram_cell[      78] = 32'h0;  // 32'h05443974;
    ram_cell[      79] = 32'h0;  // 32'hf754a45d;
    ram_cell[      80] = 32'h0;  // 32'h0dfce3a9;
    ram_cell[      81] = 32'h0;  // 32'hb950703d;
    ram_cell[      82] = 32'h0;  // 32'h18625662;
    ram_cell[      83] = 32'h0;  // 32'h986bd8de;
    ram_cell[      84] = 32'h0;  // 32'h7e25e4a6;
    ram_cell[      85] = 32'h0;  // 32'hd4710fac;
    ram_cell[      86] = 32'h0;  // 32'h436273b2;
    ram_cell[      87] = 32'h0;  // 32'h0d62be21;
    ram_cell[      88] = 32'h0;  // 32'h6cff3d49;
    ram_cell[      89] = 32'h0;  // 32'h82701177;
    ram_cell[      90] = 32'h0;  // 32'hb2bbfb06;
    ram_cell[      91] = 32'h0;  // 32'he796821e;
    ram_cell[      92] = 32'h0;  // 32'h87a62a62;
    ram_cell[      93] = 32'h0;  // 32'h7e566a75;
    ram_cell[      94] = 32'h0;  // 32'h569777b8;
    ram_cell[      95] = 32'h0;  // 32'h07b59cc9;
    ram_cell[      96] = 32'h0;  // 32'hb8306036;
    ram_cell[      97] = 32'h0;  // 32'h2a6c4e74;
    ram_cell[      98] = 32'h0;  // 32'h85a2ac2b;
    ram_cell[      99] = 32'h0;  // 32'h49f623e2;
    ram_cell[     100] = 32'h0;  // 32'he5d7fa40;
    ram_cell[     101] = 32'h0;  // 32'h86b86d90;
    ram_cell[     102] = 32'h0;  // 32'h817ca79b;
    ram_cell[     103] = 32'h0;  // 32'h92b2e995;
    ram_cell[     104] = 32'h0;  // 32'h3c4240c1;
    ram_cell[     105] = 32'h0;  // 32'hbc0b7d58;
    ram_cell[     106] = 32'h0;  // 32'h0f4ab100;
    ram_cell[     107] = 32'h0;  // 32'h82566847;
    ram_cell[     108] = 32'h0;  // 32'hb0928604;
    ram_cell[     109] = 32'h0;  // 32'h48f07370;
    ram_cell[     110] = 32'h0;  // 32'ha6877548;
    ram_cell[     111] = 32'h0;  // 32'hbfff6a8c;
    ram_cell[     112] = 32'h0;  // 32'h0efb9d67;
    ram_cell[     113] = 32'h0;  // 32'h32145375;
    ram_cell[     114] = 32'h0;  // 32'h55f486d5;
    ram_cell[     115] = 32'h0;  // 32'hef56fc54;
    ram_cell[     116] = 32'h0;  // 32'h89c0f0da;
    ram_cell[     117] = 32'h0;  // 32'h3286ae20;
    ram_cell[     118] = 32'h0;  // 32'hfa459fd0;
    ram_cell[     119] = 32'h0;  // 32'h196ebdb7;
    ram_cell[     120] = 32'h0;  // 32'he62258eb;
    ram_cell[     121] = 32'h0;  // 32'hb8783a2e;
    ram_cell[     122] = 32'h0;  // 32'h1eb309f8;
    ram_cell[     123] = 32'h0;  // 32'hdb62668f;
    ram_cell[     124] = 32'h0;  // 32'hf338d2e9;
    ram_cell[     125] = 32'h0;  // 32'hb6b9155d;
    ram_cell[     126] = 32'h0;  // 32'h0e6d3add;
    ram_cell[     127] = 32'h0;  // 32'hda8b0a01;
    ram_cell[     128] = 32'h0;  // 32'h0bd1756f;
    ram_cell[     129] = 32'h0;  // 32'hcc2406cf;
    ram_cell[     130] = 32'h0;  // 32'hc80a905d;
    ram_cell[     131] = 32'h0;  // 32'hf01e1233;
    ram_cell[     132] = 32'h0;  // 32'h62c5dfbd;
    ram_cell[     133] = 32'h0;  // 32'h86dee14d;
    ram_cell[     134] = 32'h0;  // 32'h4fca01a5;
    ram_cell[     135] = 32'h0;  // 32'h13ab1367;
    ram_cell[     136] = 32'h0;  // 32'h17dc9ab3;
    ram_cell[     137] = 32'h0;  // 32'he9ffec1e;
    ram_cell[     138] = 32'h0;  // 32'hf314e1e8;
    ram_cell[     139] = 32'h0;  // 32'hf77451f8;
    ram_cell[     140] = 32'h0;  // 32'h004d0b79;
    ram_cell[     141] = 32'h0;  // 32'h4b30c86e;
    ram_cell[     142] = 32'h0;  // 32'h07554be0;
    ram_cell[     143] = 32'h0;  // 32'hecb50ba6;
    ram_cell[     144] = 32'h0;  // 32'h20e83ac2;
    ram_cell[     145] = 32'h0;  // 32'h7e62aa69;
    ram_cell[     146] = 32'h0;  // 32'ha5d33801;
    ram_cell[     147] = 32'h0;  // 32'h89405761;
    ram_cell[     148] = 32'h0;  // 32'h6bc68606;
    ram_cell[     149] = 32'h0;  // 32'ha9da25f4;
    ram_cell[     150] = 32'h0;  // 32'hf25f5976;
    ram_cell[     151] = 32'h0;  // 32'h36c8ac47;
    ram_cell[     152] = 32'h0;  // 32'hfc4a7117;
    ram_cell[     153] = 32'h0;  // 32'h4f114d12;
    ram_cell[     154] = 32'h0;  // 32'hfe52fe16;
    ram_cell[     155] = 32'h0;  // 32'h734a39b2;
    ram_cell[     156] = 32'h0;  // 32'haf81c15f;
    ram_cell[     157] = 32'h0;  // 32'h08a92a89;
    ram_cell[     158] = 32'h0;  // 32'h4fc9044b;
    ram_cell[     159] = 32'h0;  // 32'h6bba5908;
    ram_cell[     160] = 32'h0;  // 32'he25beb1e;
    ram_cell[     161] = 32'h0;  // 32'h9c13b722;
    ram_cell[     162] = 32'h0;  // 32'h16b46a52;
    ram_cell[     163] = 32'h0;  // 32'hed65acb0;
    ram_cell[     164] = 32'h0;  // 32'h1962ae40;
    ram_cell[     165] = 32'h0;  // 32'h0c4f78e9;
    ram_cell[     166] = 32'h0;  // 32'h2d172b7e;
    ram_cell[     167] = 32'h0;  // 32'hbf5690c4;
    ram_cell[     168] = 32'h0;  // 32'h23179298;
    ram_cell[     169] = 32'h0;  // 32'he34fe80f;
    ram_cell[     170] = 32'h0;  // 32'h9fedef8b;
    ram_cell[     171] = 32'h0;  // 32'h1969508d;
    ram_cell[     172] = 32'h0;  // 32'h64e73035;
    ram_cell[     173] = 32'h0;  // 32'hf5b5e923;
    ram_cell[     174] = 32'h0;  // 32'h355e55b8;
    ram_cell[     175] = 32'h0;  // 32'h4d68e1e8;
    ram_cell[     176] = 32'h0;  // 32'hcbf56960;
    ram_cell[     177] = 32'h0;  // 32'h47252923;
    ram_cell[     178] = 32'h0;  // 32'hfac76fa2;
    ram_cell[     179] = 32'h0;  // 32'h2e6bd915;
    ram_cell[     180] = 32'h0;  // 32'h9cea0fa5;
    ram_cell[     181] = 32'h0;  // 32'he3a699e0;
    ram_cell[     182] = 32'h0;  // 32'hbeafa676;
    ram_cell[     183] = 32'h0;  // 32'hbdfb47e3;
    ram_cell[     184] = 32'h0;  // 32'hb161dde2;
    ram_cell[     185] = 32'h0;  // 32'h483bece9;
    ram_cell[     186] = 32'h0;  // 32'hd87c2ef3;
    ram_cell[     187] = 32'h0;  // 32'h277056e3;
    ram_cell[     188] = 32'h0;  // 32'hf1304b35;
    ram_cell[     189] = 32'h0;  // 32'h126725d5;
    ram_cell[     190] = 32'h0;  // 32'ha56b0c7e;
    ram_cell[     191] = 32'h0;  // 32'h32614251;
    ram_cell[     192] = 32'h0;  // 32'hb7b34ea4;
    ram_cell[     193] = 32'h0;  // 32'haa5d8642;
    ram_cell[     194] = 32'h0;  // 32'h6761c922;
    ram_cell[     195] = 32'h0;  // 32'h06920b25;
    ram_cell[     196] = 32'h0;  // 32'h3e4fd098;
    ram_cell[     197] = 32'h0;  // 32'h3f9846f2;
    ram_cell[     198] = 32'h0;  // 32'he4715051;
    ram_cell[     199] = 32'h0;  // 32'h92f0e0bd;
    ram_cell[     200] = 32'h0;  // 32'h5372521a;
    ram_cell[     201] = 32'h0;  // 32'h6905b83c;
    ram_cell[     202] = 32'h0;  // 32'h8f7f23e9;
    ram_cell[     203] = 32'h0;  // 32'h3f0cc48d;
    ram_cell[     204] = 32'h0;  // 32'h80db6a94;
    ram_cell[     205] = 32'h0;  // 32'h8e300367;
    ram_cell[     206] = 32'h0;  // 32'h89c09671;
    ram_cell[     207] = 32'h0;  // 32'h5ba95a16;
    ram_cell[     208] = 32'h0;  // 32'he7b5d74a;
    ram_cell[     209] = 32'h0;  // 32'hda3e4bdc;
    ram_cell[     210] = 32'h0;  // 32'h0c35d443;
    ram_cell[     211] = 32'h0;  // 32'h39009cb4;
    ram_cell[     212] = 32'h0;  // 32'hd314d622;
    ram_cell[     213] = 32'h0;  // 32'h9cede50f;
    ram_cell[     214] = 32'h0;  // 32'h3ecc3850;
    ram_cell[     215] = 32'h0;  // 32'h87965cad;
    ram_cell[     216] = 32'h0;  // 32'hdafbfb85;
    ram_cell[     217] = 32'h0;  // 32'heaae22b3;
    ram_cell[     218] = 32'h0;  // 32'h88f766cf;
    ram_cell[     219] = 32'h0;  // 32'hde8a5517;
    ram_cell[     220] = 32'h0;  // 32'h56eddc29;
    ram_cell[     221] = 32'h0;  // 32'hdb071e31;
    ram_cell[     222] = 32'h0;  // 32'ha28de746;
    ram_cell[     223] = 32'h0;  // 32'hcfb5c840;
    ram_cell[     224] = 32'h0;  // 32'hafdd712b;
    ram_cell[     225] = 32'h0;  // 32'h4c8aae3a;
    ram_cell[     226] = 32'h0;  // 32'h534fc31c;
    ram_cell[     227] = 32'h0;  // 32'hd8b3b0fe;
    ram_cell[     228] = 32'h0;  // 32'h58b05957;
    ram_cell[     229] = 32'h0;  // 32'haddb73ce;
    ram_cell[     230] = 32'h0;  // 32'he566efe1;
    ram_cell[     231] = 32'h0;  // 32'h7146dc33;
    ram_cell[     232] = 32'h0;  // 32'h47e6c1fb;
    ram_cell[     233] = 32'h0;  // 32'h18fff972;
    ram_cell[     234] = 32'h0;  // 32'h7fe4b4ec;
    ram_cell[     235] = 32'h0;  // 32'h10e94f2a;
    ram_cell[     236] = 32'h0;  // 32'h29b4c918;
    ram_cell[     237] = 32'h0;  // 32'h22998618;
    ram_cell[     238] = 32'h0;  // 32'h33f528f1;
    ram_cell[     239] = 32'h0;  // 32'h845a6680;
    ram_cell[     240] = 32'h0;  // 32'hf08f4413;
    ram_cell[     241] = 32'h0;  // 32'hf9512147;
    ram_cell[     242] = 32'h0;  // 32'h1bd81586;
    ram_cell[     243] = 32'h0;  // 32'h49884eef;
    ram_cell[     244] = 32'h0;  // 32'hf8ac1d11;
    ram_cell[     245] = 32'h0;  // 32'h0bcd7bed;
    ram_cell[     246] = 32'h0;  // 32'h9acbde4a;
    ram_cell[     247] = 32'h0;  // 32'h5ddfcb5f;
    ram_cell[     248] = 32'h0;  // 32'h3983f738;
    ram_cell[     249] = 32'h0;  // 32'hf7ea8edb;
    ram_cell[     250] = 32'h0;  // 32'h182ce0ab;
    ram_cell[     251] = 32'h0;  // 32'h13ee2d27;
    ram_cell[     252] = 32'h0;  // 32'hbb331da1;
    ram_cell[     253] = 32'h0;  // 32'h7f5da2c7;
    ram_cell[     254] = 32'h0;  // 32'h3c5da478;
    ram_cell[     255] = 32'h0;  // 32'hace7f473;
    ram_cell[     256] = 32'h0;  // 32'h1123772e;
    ram_cell[     257] = 32'h0;  // 32'h777d2b81;
    ram_cell[     258] = 32'h0;  // 32'h939aaa68;
    ram_cell[     259] = 32'h0;  // 32'h909c97f7;
    ram_cell[     260] = 32'h0;  // 32'h195bcdd9;
    ram_cell[     261] = 32'h0;  // 32'h4cf0aea0;
    ram_cell[     262] = 32'h0;  // 32'h88a96c05;
    ram_cell[     263] = 32'h0;  // 32'h90e0f935;
    ram_cell[     264] = 32'h0;  // 32'h59c31ea0;
    ram_cell[     265] = 32'h0;  // 32'hfe2bff14;
    ram_cell[     266] = 32'h0;  // 32'hb95e210e;
    ram_cell[     267] = 32'h0;  // 32'hbcaeb5d7;
    ram_cell[     268] = 32'h0;  // 32'hcf53b874;
    ram_cell[     269] = 32'h0;  // 32'hb96276dd;
    ram_cell[     270] = 32'h0;  // 32'h6f1e82a1;
    ram_cell[     271] = 32'h0;  // 32'h1356a14b;
    ram_cell[     272] = 32'h0;  // 32'h2ac3bf1a;
    ram_cell[     273] = 32'h0;  // 32'h41127b2c;
    ram_cell[     274] = 32'h0;  // 32'h13678c71;
    ram_cell[     275] = 32'h0;  // 32'h19409544;
    ram_cell[     276] = 32'h0;  // 32'h83dba674;
    ram_cell[     277] = 32'h0;  // 32'hadc1fa49;
    ram_cell[     278] = 32'h0;  // 32'h3bd8af3d;
    ram_cell[     279] = 32'h0;  // 32'h3ee99df8;
    ram_cell[     280] = 32'h0;  // 32'h65098b28;
    ram_cell[     281] = 32'h0;  // 32'hf43089f8;
    ram_cell[     282] = 32'h0;  // 32'hb01ac2df;
    ram_cell[     283] = 32'h0;  // 32'hddebcf2e;
    ram_cell[     284] = 32'h0;  // 32'h5d943796;
    ram_cell[     285] = 32'h0;  // 32'h4d04b22e;
    ram_cell[     286] = 32'h0;  // 32'h69ccd7d0;
    ram_cell[     287] = 32'h0;  // 32'hf140fa57;
    ram_cell[     288] = 32'h0;  // 32'h1532ffb7;
    ram_cell[     289] = 32'h0;  // 32'h7a3f38f9;
    ram_cell[     290] = 32'h0;  // 32'h9cb8b68f;
    ram_cell[     291] = 32'h0;  // 32'h4e413d81;
    ram_cell[     292] = 32'h0;  // 32'hacac36fe;
    ram_cell[     293] = 32'h0;  // 32'h3a016d85;
    ram_cell[     294] = 32'h0;  // 32'h1fbee14f;
    ram_cell[     295] = 32'h0;  // 32'h06b3f9a1;
    ram_cell[     296] = 32'h0;  // 32'hcd763185;
    ram_cell[     297] = 32'h0;  // 32'hed475699;
    ram_cell[     298] = 32'h0;  // 32'haf30acb0;
    ram_cell[     299] = 32'h0;  // 32'hf103e634;
    ram_cell[     300] = 32'h0;  // 32'h12bb514b;
    ram_cell[     301] = 32'h0;  // 32'h8b882652;
    ram_cell[     302] = 32'h0;  // 32'h2c27665c;
    ram_cell[     303] = 32'h0;  // 32'h1cee2551;
    ram_cell[     304] = 32'h0;  // 32'h9cae573e;
    ram_cell[     305] = 32'h0;  // 32'haef2bd8c;
    ram_cell[     306] = 32'h0;  // 32'h99414d69;
    ram_cell[     307] = 32'h0;  // 32'h9567a07b;
    ram_cell[     308] = 32'h0;  // 32'hed409dce;
    ram_cell[     309] = 32'h0;  // 32'hbe6d3acb;
    ram_cell[     310] = 32'h0;  // 32'h445df543;
    ram_cell[     311] = 32'h0;  // 32'hb455ce00;
    ram_cell[     312] = 32'h0;  // 32'h223f95f3;
    ram_cell[     313] = 32'h0;  // 32'ha3f109d3;
    ram_cell[     314] = 32'h0;  // 32'hce9e57a4;
    ram_cell[     315] = 32'h0;  // 32'h2250dfd1;
    ram_cell[     316] = 32'h0;  // 32'h4dfbe8c4;
    ram_cell[     317] = 32'h0;  // 32'h0fbfe357;
    ram_cell[     318] = 32'h0;  // 32'h22ae5697;
    ram_cell[     319] = 32'h0;  // 32'h6b8f3ea6;
    ram_cell[     320] = 32'h0;  // 32'h03ae3b3d;
    ram_cell[     321] = 32'h0;  // 32'h6697ae37;
    ram_cell[     322] = 32'h0;  // 32'h3aedb74e;
    ram_cell[     323] = 32'h0;  // 32'h93bbfc02;
    ram_cell[     324] = 32'h0;  // 32'h00c24090;
    ram_cell[     325] = 32'h0;  // 32'hcedfa1b0;
    ram_cell[     326] = 32'h0;  // 32'hfa09c55b;
    ram_cell[     327] = 32'h0;  // 32'h81e744a6;
    ram_cell[     328] = 32'h0;  // 32'h2711bc99;
    ram_cell[     329] = 32'h0;  // 32'hf660f7a1;
    ram_cell[     330] = 32'h0;  // 32'h15cd96ab;
    ram_cell[     331] = 32'h0;  // 32'h2f9ad876;
    ram_cell[     332] = 32'h0;  // 32'h2ccbcf1f;
    ram_cell[     333] = 32'h0;  // 32'hb60ddfa3;
    ram_cell[     334] = 32'h0;  // 32'h2ea0efcd;
    ram_cell[     335] = 32'h0;  // 32'h3ce9c6fd;
    ram_cell[     336] = 32'h0;  // 32'hbc7d2dc9;
    ram_cell[     337] = 32'h0;  // 32'h13d563fb;
    ram_cell[     338] = 32'h0;  // 32'h09300577;
    ram_cell[     339] = 32'h0;  // 32'h2160f169;
    ram_cell[     340] = 32'h0;  // 32'hce691a07;
    ram_cell[     341] = 32'h0;  // 32'h7d230768;
    ram_cell[     342] = 32'h0;  // 32'haf2b1187;
    ram_cell[     343] = 32'h0;  // 32'hb5c4e25a;
    ram_cell[     344] = 32'h0;  // 32'ha9431b0e;
    ram_cell[     345] = 32'h0;  // 32'h2408ad1e;
    ram_cell[     346] = 32'h0;  // 32'h4c5cd54f;
    ram_cell[     347] = 32'h0;  // 32'h0c3fc41e;
    ram_cell[     348] = 32'h0;  // 32'hdd6ec9bd;
    ram_cell[     349] = 32'h0;  // 32'h8f7f18cd;
    ram_cell[     350] = 32'h0;  // 32'hd31ea5d4;
    ram_cell[     351] = 32'h0;  // 32'hf61729cf;
    ram_cell[     352] = 32'h0;  // 32'hef41640c;
    ram_cell[     353] = 32'h0;  // 32'h66fd3fe0;
    ram_cell[     354] = 32'h0;  // 32'hda7d2d5b;
    ram_cell[     355] = 32'h0;  // 32'hc3da83dd;
    ram_cell[     356] = 32'h0;  // 32'h137e1e0b;
    ram_cell[     357] = 32'h0;  // 32'he06ffcf0;
    ram_cell[     358] = 32'h0;  // 32'hc58ab59a;
    ram_cell[     359] = 32'h0;  // 32'he7501833;
    ram_cell[     360] = 32'h0;  // 32'hc2effeb5;
    ram_cell[     361] = 32'h0;  // 32'hf753552f;
    ram_cell[     362] = 32'h0;  // 32'h4572f99d;
    ram_cell[     363] = 32'h0;  // 32'hca0e17c5;
    ram_cell[     364] = 32'h0;  // 32'h7505dd30;
    ram_cell[     365] = 32'h0;  // 32'h5dd39594;
    ram_cell[     366] = 32'h0;  // 32'h5f76c1d7;
    ram_cell[     367] = 32'h0;  // 32'hf85c84a0;
    ram_cell[     368] = 32'h0;  // 32'hc2b4c6ca;
    ram_cell[     369] = 32'h0;  // 32'hf5cd92dd;
    ram_cell[     370] = 32'h0;  // 32'ha20083fe;
    ram_cell[     371] = 32'h0;  // 32'h06497ef1;
    ram_cell[     372] = 32'h0;  // 32'h5705cd8d;
    ram_cell[     373] = 32'h0;  // 32'h5a60ea86;
    ram_cell[     374] = 32'h0;  // 32'h2232bd50;
    ram_cell[     375] = 32'h0;  // 32'h46d55d03;
    ram_cell[     376] = 32'h0;  // 32'h2061e84f;
    ram_cell[     377] = 32'h0;  // 32'hb493c7ae;
    ram_cell[     378] = 32'h0;  // 32'h81cd3760;
    ram_cell[     379] = 32'h0;  // 32'h542953b7;
    ram_cell[     380] = 32'h0;  // 32'h2c8ae397;
    ram_cell[     381] = 32'h0;  // 32'h08388a63;
    ram_cell[     382] = 32'h0;  // 32'hea56bdaf;
    ram_cell[     383] = 32'h0;  // 32'hf7113404;
    ram_cell[     384] = 32'h0;  // 32'h651a43ed;
    ram_cell[     385] = 32'h0;  // 32'hd115e497;
    ram_cell[     386] = 32'h0;  // 32'h1675b0d2;
    ram_cell[     387] = 32'h0;  // 32'h4a7c7ef7;
    ram_cell[     388] = 32'h0;  // 32'h5fd28538;
    ram_cell[     389] = 32'h0;  // 32'h1d0e9225;
    ram_cell[     390] = 32'h0;  // 32'hdde68188;
    ram_cell[     391] = 32'h0;  // 32'h63010b42;
    ram_cell[     392] = 32'h0;  // 32'h54efd51e;
    ram_cell[     393] = 32'h0;  // 32'hd56305a9;
    ram_cell[     394] = 32'h0;  // 32'h051caaf5;
    ram_cell[     395] = 32'h0;  // 32'hb1021b58;
    ram_cell[     396] = 32'h0;  // 32'h252f37b8;
    ram_cell[     397] = 32'h0;  // 32'he6a776fe;
    ram_cell[     398] = 32'h0;  // 32'h253be8d1;
    ram_cell[     399] = 32'h0;  // 32'h99879f2f;
    ram_cell[     400] = 32'h0;  // 32'h6f8e1303;
    ram_cell[     401] = 32'h0;  // 32'hbd987ad7;
    ram_cell[     402] = 32'h0;  // 32'h41e0e7c2;
    ram_cell[     403] = 32'h0;  // 32'h7d9e4dfe;
    ram_cell[     404] = 32'h0;  // 32'h94922845;
    ram_cell[     405] = 32'h0;  // 32'h59fade63;
    ram_cell[     406] = 32'h0;  // 32'h1dfbe461;
    ram_cell[     407] = 32'h0;  // 32'h3f7e2524;
    ram_cell[     408] = 32'h0;  // 32'hf164e49f;
    ram_cell[     409] = 32'h0;  // 32'h89227fd4;
    ram_cell[     410] = 32'h0;  // 32'hde1e6d63;
    ram_cell[     411] = 32'h0;  // 32'h14292298;
    ram_cell[     412] = 32'h0;  // 32'h1a889b30;
    ram_cell[     413] = 32'h0;  // 32'h748206a1;
    ram_cell[     414] = 32'h0;  // 32'hf669ce6b;
    ram_cell[     415] = 32'h0;  // 32'h9ecfb7a3;
    ram_cell[     416] = 32'h0;  // 32'hfeabf102;
    ram_cell[     417] = 32'h0;  // 32'h63556838;
    ram_cell[     418] = 32'h0;  // 32'h2a1bebc1;
    ram_cell[     419] = 32'h0;  // 32'h05f56788;
    ram_cell[     420] = 32'h0;  // 32'h8e23e571;
    ram_cell[     421] = 32'h0;  // 32'ha2fd9202;
    ram_cell[     422] = 32'h0;  // 32'h8f5df672;
    ram_cell[     423] = 32'h0;  // 32'h146dc976;
    ram_cell[     424] = 32'h0;  // 32'hd1e96b86;
    ram_cell[     425] = 32'h0;  // 32'h461473ba;
    ram_cell[     426] = 32'h0;  // 32'h634d45e4;
    ram_cell[     427] = 32'h0;  // 32'hf8fa1b2d;
    ram_cell[     428] = 32'h0;  // 32'h18c73763;
    ram_cell[     429] = 32'h0;  // 32'h51323efd;
    ram_cell[     430] = 32'h0;  // 32'hef67f32f;
    ram_cell[     431] = 32'h0;  // 32'he8305d3c;
    ram_cell[     432] = 32'h0;  // 32'h5d7d19b9;
    ram_cell[     433] = 32'h0;  // 32'hb06577c9;
    ram_cell[     434] = 32'h0;  // 32'he7432ad7;
    ram_cell[     435] = 32'h0;  // 32'h7cb61c2f;
    ram_cell[     436] = 32'h0;  // 32'hdf682a12;
    ram_cell[     437] = 32'h0;  // 32'h2d1218a0;
    ram_cell[     438] = 32'h0;  // 32'h44f07f19;
    ram_cell[     439] = 32'h0;  // 32'h8fce5d98;
    ram_cell[     440] = 32'h0;  // 32'he573dfee;
    ram_cell[     441] = 32'h0;  // 32'h5c281cf4;
    ram_cell[     442] = 32'h0;  // 32'h9bf91fb6;
    ram_cell[     443] = 32'h0;  // 32'hfa7ce087;
    ram_cell[     444] = 32'h0;  // 32'h6057d0d3;
    ram_cell[     445] = 32'h0;  // 32'h70bcdc9e;
    ram_cell[     446] = 32'h0;  // 32'hc2258558;
    ram_cell[     447] = 32'h0;  // 32'h1dc23528;
    ram_cell[     448] = 32'h0;  // 32'hf396b1d5;
    ram_cell[     449] = 32'h0;  // 32'h8cd27c2f;
    ram_cell[     450] = 32'h0;  // 32'hb523be5c;
    ram_cell[     451] = 32'h0;  // 32'h7a804af9;
    ram_cell[     452] = 32'h0;  // 32'hece144dd;
    ram_cell[     453] = 32'h0;  // 32'hed262bc5;
    ram_cell[     454] = 32'h0;  // 32'h6397bb3a;
    ram_cell[     455] = 32'h0;  // 32'h60ca834e;
    ram_cell[     456] = 32'h0;  // 32'h3fef3954;
    ram_cell[     457] = 32'h0;  // 32'h6fb39cb6;
    ram_cell[     458] = 32'h0;  // 32'hf0593040;
    ram_cell[     459] = 32'h0;  // 32'hf298dced;
    ram_cell[     460] = 32'h0;  // 32'ha24a2c32;
    ram_cell[     461] = 32'h0;  // 32'h79a2aa00;
    ram_cell[     462] = 32'h0;  // 32'h9a492304;
    ram_cell[     463] = 32'h0;  // 32'h4b15bed0;
    ram_cell[     464] = 32'h0;  // 32'h6fc7b6ef;
    ram_cell[     465] = 32'h0;  // 32'h7e55faa1;
    ram_cell[     466] = 32'h0;  // 32'hceb7cee2;
    ram_cell[     467] = 32'h0;  // 32'h05f8395c;
    ram_cell[     468] = 32'h0;  // 32'h83d10664;
    ram_cell[     469] = 32'h0;  // 32'h46f29e6d;
    ram_cell[     470] = 32'h0;  // 32'h5cc9de45;
    ram_cell[     471] = 32'h0;  // 32'h0a37c96c;
    ram_cell[     472] = 32'h0;  // 32'hb1fc825a;
    ram_cell[     473] = 32'h0;  // 32'h41b96ea9;
    ram_cell[     474] = 32'h0;  // 32'h349f4eb0;
    ram_cell[     475] = 32'h0;  // 32'hbc1f8c75;
    ram_cell[     476] = 32'h0;  // 32'hfa02266d;
    ram_cell[     477] = 32'h0;  // 32'h0f106a40;
    ram_cell[     478] = 32'h0;  // 32'h34fc3d1a;
    ram_cell[     479] = 32'h0;  // 32'h2713d55b;
    ram_cell[     480] = 32'h0;  // 32'h6856e694;
    ram_cell[     481] = 32'h0;  // 32'ha8f0b9f5;
    ram_cell[     482] = 32'h0;  // 32'h312b1797;
    ram_cell[     483] = 32'h0;  // 32'h465b8aac;
    ram_cell[     484] = 32'h0;  // 32'h0656692d;
    ram_cell[     485] = 32'h0;  // 32'hb4620c8c;
    ram_cell[     486] = 32'h0;  // 32'h8a66cfd1;
    ram_cell[     487] = 32'h0;  // 32'h84589065;
    ram_cell[     488] = 32'h0;  // 32'h1ae4ce1f;
    ram_cell[     489] = 32'h0;  // 32'h66eb5f4a;
    ram_cell[     490] = 32'h0;  // 32'h2e793291;
    ram_cell[     491] = 32'h0;  // 32'habc8f6bf;
    ram_cell[     492] = 32'h0;  // 32'h700b0860;
    ram_cell[     493] = 32'h0;  // 32'h27a13c94;
    ram_cell[     494] = 32'h0;  // 32'h978405d9;
    ram_cell[     495] = 32'h0;  // 32'h16cefc97;
    ram_cell[     496] = 32'h0;  // 32'h3253e85e;
    ram_cell[     497] = 32'h0;  // 32'hba5168f4;
    ram_cell[     498] = 32'h0;  // 32'h084493ae;
    ram_cell[     499] = 32'h0;  // 32'hd1303989;
    ram_cell[     500] = 32'h0;  // 32'h81ac17f3;
    ram_cell[     501] = 32'h0;  // 32'h4ea38ebd;
    ram_cell[     502] = 32'h0;  // 32'heafa77f6;
    ram_cell[     503] = 32'h0;  // 32'h28b0c733;
    ram_cell[     504] = 32'h0;  // 32'h3dc9dde3;
    ram_cell[     505] = 32'h0;  // 32'h20516c07;
    ram_cell[     506] = 32'h0;  // 32'hea70a703;
    ram_cell[     507] = 32'h0;  // 32'h4654bdf5;
    ram_cell[     508] = 32'h0;  // 32'had6bea27;
    ram_cell[     509] = 32'h0;  // 32'h48b8ede8;
    ram_cell[     510] = 32'h0;  // 32'h40562a71;
    ram_cell[     511] = 32'h0;  // 32'h36729ec1;
    ram_cell[     512] = 32'h0;  // 32'h5c1c01d9;
    ram_cell[     513] = 32'h0;  // 32'h74e6fa1d;
    ram_cell[     514] = 32'h0;  // 32'hf1ea5a5a;
    ram_cell[     515] = 32'h0;  // 32'h163a9690;
    ram_cell[     516] = 32'h0;  // 32'h451bd3e9;
    ram_cell[     517] = 32'h0;  // 32'h620070ba;
    ram_cell[     518] = 32'h0;  // 32'ha2e2a519;
    ram_cell[     519] = 32'h0;  // 32'hb482a982;
    ram_cell[     520] = 32'h0;  // 32'h2ece3478;
    ram_cell[     521] = 32'h0;  // 32'ha62f3f57;
    ram_cell[     522] = 32'h0;  // 32'hfa170f5b;
    ram_cell[     523] = 32'h0;  // 32'h4e0593e9;
    ram_cell[     524] = 32'h0;  // 32'hbcfdc2fb;
    ram_cell[     525] = 32'h0;  // 32'hb8c7b737;
    ram_cell[     526] = 32'h0;  // 32'h4a289160;
    ram_cell[     527] = 32'h0;  // 32'hf93ce36c;
    ram_cell[     528] = 32'h0;  // 32'h8340400c;
    ram_cell[     529] = 32'h0;  // 32'h269f437f;
    ram_cell[     530] = 32'h0;  // 32'hb1767b5f;
    ram_cell[     531] = 32'h0;  // 32'h4a158ef0;
    ram_cell[     532] = 32'h0;  // 32'hf4020995;
    ram_cell[     533] = 32'h0;  // 32'hf9befa20;
    ram_cell[     534] = 32'h0;  // 32'h9cadfa66;
    ram_cell[     535] = 32'h0;  // 32'h09dd6bd6;
    ram_cell[     536] = 32'h0;  // 32'h4c392fd8;
    ram_cell[     537] = 32'h0;  // 32'hf7e6d527;
    ram_cell[     538] = 32'h0;  // 32'h20bac34d;
    ram_cell[     539] = 32'h0;  // 32'h252cbec2;
    ram_cell[     540] = 32'h0;  // 32'he8bdefdb;
    ram_cell[     541] = 32'h0;  // 32'hb848ea3f;
    ram_cell[     542] = 32'h0;  // 32'ha7f583bc;
    ram_cell[     543] = 32'h0;  // 32'h3b51e9bb;
    ram_cell[     544] = 32'h0;  // 32'h2023d7d1;
    ram_cell[     545] = 32'h0;  // 32'h2eb6de2d;
    ram_cell[     546] = 32'h0;  // 32'hc298f0bf;
    ram_cell[     547] = 32'h0;  // 32'hae8e32a3;
    ram_cell[     548] = 32'h0;  // 32'h0e50f25c;
    ram_cell[     549] = 32'h0;  // 32'hcb7291ac;
    ram_cell[     550] = 32'h0;  // 32'he4f63fa4;
    ram_cell[     551] = 32'h0;  // 32'hcfba9ae0;
    ram_cell[     552] = 32'h0;  // 32'h1bb62fb9;
    ram_cell[     553] = 32'h0;  // 32'hc8e34eda;
    ram_cell[     554] = 32'h0;  // 32'h86a19042;
    ram_cell[     555] = 32'h0;  // 32'hf561b70e;
    ram_cell[     556] = 32'h0;  // 32'hb15ebc30;
    ram_cell[     557] = 32'h0;  // 32'hb41a6d2f;
    ram_cell[     558] = 32'h0;  // 32'h06c5e321;
    ram_cell[     559] = 32'h0;  // 32'h645b2a80;
    ram_cell[     560] = 32'h0;  // 32'h74fb4af7;
    ram_cell[     561] = 32'h0;  // 32'h22702c07;
    ram_cell[     562] = 32'h0;  // 32'h2feee2f7;
    ram_cell[     563] = 32'h0;  // 32'h6e76667f;
    ram_cell[     564] = 32'h0;  // 32'h4d534ff0;
    ram_cell[     565] = 32'h0;  // 32'h67f3b1e5;
    ram_cell[     566] = 32'h0;  // 32'h1916f63a;
    ram_cell[     567] = 32'h0;  // 32'h511b56d7;
    ram_cell[     568] = 32'h0;  // 32'hb81088ab;
    ram_cell[     569] = 32'h0;  // 32'h265164da;
    ram_cell[     570] = 32'h0;  // 32'hc8225004;
    ram_cell[     571] = 32'h0;  // 32'h704e9a51;
    ram_cell[     572] = 32'h0;  // 32'h883fae5d;
    ram_cell[     573] = 32'h0;  // 32'hddb4b71f;
    ram_cell[     574] = 32'h0;  // 32'h8b44be06;
    ram_cell[     575] = 32'h0;  // 32'haa24ede6;
    ram_cell[     576] = 32'h0;  // 32'h6adf0df9;
    ram_cell[     577] = 32'h0;  // 32'h30efb44e;
    ram_cell[     578] = 32'h0;  // 32'h22912ba8;
    ram_cell[     579] = 32'h0;  // 32'hbbb543ea;
    ram_cell[     580] = 32'h0;  // 32'h6af1cd9f;
    ram_cell[     581] = 32'h0;  // 32'h1ea2cd96;
    ram_cell[     582] = 32'h0;  // 32'he000508a;
    ram_cell[     583] = 32'h0;  // 32'haa6b5f97;
    ram_cell[     584] = 32'h0;  // 32'h18093cb5;
    ram_cell[     585] = 32'h0;  // 32'hab49ab1e;
    ram_cell[     586] = 32'h0;  // 32'h36aa6b94;
    ram_cell[     587] = 32'h0;  // 32'hdf7584f6;
    ram_cell[     588] = 32'h0;  // 32'h3889abd8;
    ram_cell[     589] = 32'h0;  // 32'hbbcfe1b2;
    ram_cell[     590] = 32'h0;  // 32'h518127bc;
    ram_cell[     591] = 32'h0;  // 32'h24962558;
    ram_cell[     592] = 32'h0;  // 32'h8ae6cdde;
    ram_cell[     593] = 32'h0;  // 32'h133ac2c2;
    ram_cell[     594] = 32'h0;  // 32'h6ee17fd6;
    ram_cell[     595] = 32'h0;  // 32'h900eb331;
    ram_cell[     596] = 32'h0;  // 32'h5c610620;
    ram_cell[     597] = 32'h0;  // 32'h1304b099;
    ram_cell[     598] = 32'h0;  // 32'hab65c768;
    ram_cell[     599] = 32'h0;  // 32'h2885ff4d;
    ram_cell[     600] = 32'h0;  // 32'hcc3efacc;
    ram_cell[     601] = 32'h0;  // 32'h7953ec15;
    ram_cell[     602] = 32'h0;  // 32'hf88273bd;
    ram_cell[     603] = 32'h0;  // 32'h54a256ce;
    ram_cell[     604] = 32'h0;  // 32'hf63af9a2;
    ram_cell[     605] = 32'h0;  // 32'h80546947;
    ram_cell[     606] = 32'h0;  // 32'h5dc9eaee;
    ram_cell[     607] = 32'h0;  // 32'h77378828;
    ram_cell[     608] = 32'h0;  // 32'h615d4ef9;
    ram_cell[     609] = 32'h0;  // 32'hb2b89559;
    ram_cell[     610] = 32'h0;  // 32'hb4e2a849;
    ram_cell[     611] = 32'h0;  // 32'h93b262ac;
    ram_cell[     612] = 32'h0;  // 32'h537610d6;
    ram_cell[     613] = 32'h0;  // 32'h9a7f1a9a;
    ram_cell[     614] = 32'h0;  // 32'ha3006a69;
    ram_cell[     615] = 32'h0;  // 32'he11f76c9;
    ram_cell[     616] = 32'h0;  // 32'hb287558a;
    ram_cell[     617] = 32'h0;  // 32'h896706b7;
    ram_cell[     618] = 32'h0;  // 32'he77dad12;
    ram_cell[     619] = 32'h0;  // 32'hf44bad7c;
    ram_cell[     620] = 32'h0;  // 32'h68da1298;
    ram_cell[     621] = 32'h0;  // 32'h4c431ce3;
    ram_cell[     622] = 32'h0;  // 32'h39ba19c4;
    ram_cell[     623] = 32'h0;  // 32'h01e9ce69;
    ram_cell[     624] = 32'h0;  // 32'h67d3e3a5;
    ram_cell[     625] = 32'h0;  // 32'hed33c8b0;
    ram_cell[     626] = 32'h0;  // 32'hc4899511;
    ram_cell[     627] = 32'h0;  // 32'h6d4982dc;
    ram_cell[     628] = 32'h0;  // 32'he6473465;
    ram_cell[     629] = 32'h0;  // 32'h0ab14696;
    ram_cell[     630] = 32'h0;  // 32'h6b47db84;
    ram_cell[     631] = 32'h0;  // 32'hdcf8dbb2;
    ram_cell[     632] = 32'h0;  // 32'h74a93d95;
    ram_cell[     633] = 32'h0;  // 32'h6d14eff5;
    ram_cell[     634] = 32'h0;  // 32'h43c07780;
    ram_cell[     635] = 32'h0;  // 32'h193cae63;
    ram_cell[     636] = 32'h0;  // 32'haf6cd0c8;
    ram_cell[     637] = 32'h0;  // 32'he1ccadbc;
    ram_cell[     638] = 32'h0;  // 32'h24718a39;
    ram_cell[     639] = 32'h0;  // 32'h79bd80fc;
    ram_cell[     640] = 32'h0;  // 32'h90ef650b;
    ram_cell[     641] = 32'h0;  // 32'h044855f7;
    ram_cell[     642] = 32'h0;  // 32'he9528c56;
    ram_cell[     643] = 32'h0;  // 32'hf25e98a6;
    ram_cell[     644] = 32'h0;  // 32'h24941b7a;
    ram_cell[     645] = 32'h0;  // 32'h1ea9350f;
    ram_cell[     646] = 32'h0;  // 32'hbab599cc;
    ram_cell[     647] = 32'h0;  // 32'hfd1620db;
    ram_cell[     648] = 32'h0;  // 32'h74beb6dc;
    ram_cell[     649] = 32'h0;  // 32'hca0bef5a;
    ram_cell[     650] = 32'h0;  // 32'hc1fd7b3f;
    ram_cell[     651] = 32'h0;  // 32'hea418db1;
    ram_cell[     652] = 32'h0;  // 32'hfe60e97f;
    ram_cell[     653] = 32'h0;  // 32'hc869f0b5;
    ram_cell[     654] = 32'h0;  // 32'h3bc940cf;
    ram_cell[     655] = 32'h0;  // 32'h199b0338;
    ram_cell[     656] = 32'h0;  // 32'hce54542d;
    ram_cell[     657] = 32'h0;  // 32'h830c8a55;
    ram_cell[     658] = 32'h0;  // 32'h13316c63;
    ram_cell[     659] = 32'h0;  // 32'hb007b027;
    ram_cell[     660] = 32'h0;  // 32'ha23182b8;
    ram_cell[     661] = 32'h0;  // 32'h95cfa8b7;
    ram_cell[     662] = 32'h0;  // 32'h814ab769;
    ram_cell[     663] = 32'h0;  // 32'h6c3383a2;
    ram_cell[     664] = 32'h0;  // 32'hbcda0f68;
    ram_cell[     665] = 32'h0;  // 32'hf183bfae;
    ram_cell[     666] = 32'h0;  // 32'hbc8a420c;
    ram_cell[     667] = 32'h0;  // 32'h7aa4894d;
    ram_cell[     668] = 32'h0;  // 32'he1f6d34f;
    ram_cell[     669] = 32'h0;  // 32'h442b31a3;
    ram_cell[     670] = 32'h0;  // 32'h1562a562;
    ram_cell[     671] = 32'h0;  // 32'h5d15922f;
    ram_cell[     672] = 32'h0;  // 32'h71641640;
    ram_cell[     673] = 32'h0;  // 32'hba6b3be3;
    ram_cell[     674] = 32'h0;  // 32'h6bc673d0;
    ram_cell[     675] = 32'h0;  // 32'h24195d68;
    ram_cell[     676] = 32'h0;  // 32'h754439a1;
    ram_cell[     677] = 32'h0;  // 32'h7b6d79c9;
    ram_cell[     678] = 32'h0;  // 32'h1712c2eb;
    ram_cell[     679] = 32'h0;  // 32'hf257eb2f;
    ram_cell[     680] = 32'h0;  // 32'h7ee26d08;
    ram_cell[     681] = 32'h0;  // 32'h8928b63a;
    ram_cell[     682] = 32'h0;  // 32'hdb9e292f;
    ram_cell[     683] = 32'h0;  // 32'ha6cc86ab;
    ram_cell[     684] = 32'h0;  // 32'h2fccab46;
    ram_cell[     685] = 32'h0;  // 32'h4bd8d27f;
    ram_cell[     686] = 32'h0;  // 32'h801b4fce;
    ram_cell[     687] = 32'h0;  // 32'h6c4631a8;
    ram_cell[     688] = 32'h0;  // 32'hc1e7246f;
    ram_cell[     689] = 32'h0;  // 32'hf567ba43;
    ram_cell[     690] = 32'h0;  // 32'hc165d928;
    ram_cell[     691] = 32'h0;  // 32'hf30365e1;
    ram_cell[     692] = 32'h0;  // 32'hd20392b2;
    ram_cell[     693] = 32'h0;  // 32'h0b4a0734;
    ram_cell[     694] = 32'h0;  // 32'h1fa84570;
    ram_cell[     695] = 32'h0;  // 32'hb29206fe;
    ram_cell[     696] = 32'h0;  // 32'he61aaa55;
    ram_cell[     697] = 32'h0;  // 32'h12e75359;
    ram_cell[     698] = 32'h0;  // 32'h3a4afea9;
    ram_cell[     699] = 32'h0;  // 32'h0725360e;
    ram_cell[     700] = 32'h0;  // 32'hee60183c;
    ram_cell[     701] = 32'h0;  // 32'h8092eea2;
    ram_cell[     702] = 32'h0;  // 32'h25d5c592;
    ram_cell[     703] = 32'h0;  // 32'h4d8f53ee;
    ram_cell[     704] = 32'h0;  // 32'h179eb602;
    ram_cell[     705] = 32'h0;  // 32'hbb1a2ac7;
    ram_cell[     706] = 32'h0;  // 32'h998a3b15;
    ram_cell[     707] = 32'h0;  // 32'h1bdf2ba0;
    ram_cell[     708] = 32'h0;  // 32'haab1892d;
    ram_cell[     709] = 32'h0;  // 32'h84a7f421;
    ram_cell[     710] = 32'h0;  // 32'h9bbd33d4;
    ram_cell[     711] = 32'h0;  // 32'h79123128;
    ram_cell[     712] = 32'h0;  // 32'h552a9f0c;
    ram_cell[     713] = 32'h0;  // 32'ha64b708f;
    ram_cell[     714] = 32'h0;  // 32'ha6d88298;
    ram_cell[     715] = 32'h0;  // 32'h8b41b2f3;
    ram_cell[     716] = 32'h0;  // 32'h859ecdfc;
    ram_cell[     717] = 32'h0;  // 32'hb92c7b60;
    ram_cell[     718] = 32'h0;  // 32'h6d92cd2a;
    ram_cell[     719] = 32'h0;  // 32'h6ae64430;
    ram_cell[     720] = 32'h0;  // 32'hf8e1b176;
    ram_cell[     721] = 32'h0;  // 32'h011c6b01;
    ram_cell[     722] = 32'h0;  // 32'h20e7e018;
    ram_cell[     723] = 32'h0;  // 32'hc032e754;
    ram_cell[     724] = 32'h0;  // 32'h1270a053;
    ram_cell[     725] = 32'h0;  // 32'h28e2e6cc;
    ram_cell[     726] = 32'h0;  // 32'hf22170d1;
    ram_cell[     727] = 32'h0;  // 32'h08488a5c;
    ram_cell[     728] = 32'h0;  // 32'hf461fdbc;
    ram_cell[     729] = 32'h0;  // 32'h95d44075;
    ram_cell[     730] = 32'h0;  // 32'h363b64c7;
    ram_cell[     731] = 32'h0;  // 32'hd75bbdd6;
    ram_cell[     732] = 32'h0;  // 32'h1f2ca247;
    ram_cell[     733] = 32'h0;  // 32'h5537bcab;
    ram_cell[     734] = 32'h0;  // 32'h19b43813;
    ram_cell[     735] = 32'h0;  // 32'h0144af8c;
    ram_cell[     736] = 32'h0;  // 32'hd6d0a98b;
    ram_cell[     737] = 32'h0;  // 32'h47227140;
    ram_cell[     738] = 32'h0;  // 32'h85cc247c;
    ram_cell[     739] = 32'h0;  // 32'hf70bb385;
    ram_cell[     740] = 32'h0;  // 32'h00983932;
    ram_cell[     741] = 32'h0;  // 32'h2b407c9e;
    ram_cell[     742] = 32'h0;  // 32'h44f27d7c;
    ram_cell[     743] = 32'h0;  // 32'h84a73e49;
    ram_cell[     744] = 32'h0;  // 32'h7c7b2421;
    ram_cell[     745] = 32'h0;  // 32'h9df049f1;
    ram_cell[     746] = 32'h0;  // 32'hff45dcea;
    ram_cell[     747] = 32'h0;  // 32'h7ad7bc6b;
    ram_cell[     748] = 32'h0;  // 32'h3e25c810;
    ram_cell[     749] = 32'h0;  // 32'hb314150f;
    ram_cell[     750] = 32'h0;  // 32'h09238aa4;
    ram_cell[     751] = 32'h0;  // 32'hc25b1d92;
    ram_cell[     752] = 32'h0;  // 32'h4d3655f9;
    ram_cell[     753] = 32'h0;  // 32'hc5da4bff;
    ram_cell[     754] = 32'h0;  // 32'h55a40961;
    ram_cell[     755] = 32'h0;  // 32'hbccdbe95;
    ram_cell[     756] = 32'h0;  // 32'h4be8d119;
    ram_cell[     757] = 32'h0;  // 32'h79ea5dfb;
    ram_cell[     758] = 32'h0;  // 32'h8743d405;
    ram_cell[     759] = 32'h0;  // 32'h385aa7e7;
    ram_cell[     760] = 32'h0;  // 32'ha8757d2f;
    ram_cell[     761] = 32'h0;  // 32'he20c7527;
    ram_cell[     762] = 32'h0;  // 32'h42cc96d8;
    ram_cell[     763] = 32'h0;  // 32'h04584364;
    ram_cell[     764] = 32'h0;  // 32'h494df7c7;
    ram_cell[     765] = 32'h0;  // 32'ha07e7e25;
    ram_cell[     766] = 32'h0;  // 32'hc6deb7e4;
    ram_cell[     767] = 32'h0;  // 32'h4076464c;
    ram_cell[     768] = 32'h0;  // 32'h964e3e86;
    ram_cell[     769] = 32'h0;  // 32'h5f751316;
    ram_cell[     770] = 32'h0;  // 32'h9686cc14;
    ram_cell[     771] = 32'h0;  // 32'hcab8e928;
    ram_cell[     772] = 32'h0;  // 32'hf89fb334;
    ram_cell[     773] = 32'h0;  // 32'hdd007eb5;
    ram_cell[     774] = 32'h0;  // 32'h1ac5070d;
    ram_cell[     775] = 32'h0;  // 32'h4cfd365a;
    ram_cell[     776] = 32'h0;  // 32'hc82c6d6c;
    ram_cell[     777] = 32'h0;  // 32'h95977139;
    ram_cell[     778] = 32'h0;  // 32'h66f287da;
    ram_cell[     779] = 32'h0;  // 32'h97e83608;
    ram_cell[     780] = 32'h0;  // 32'h530110d2;
    ram_cell[     781] = 32'h0;  // 32'h35f265b1;
    ram_cell[     782] = 32'h0;  // 32'h4f53d469;
    ram_cell[     783] = 32'h0;  // 32'h86b26b62;
    ram_cell[     784] = 32'h0;  // 32'h7032be9f;
    ram_cell[     785] = 32'h0;  // 32'hee71bc25;
    ram_cell[     786] = 32'h0;  // 32'hb6e0d006;
    ram_cell[     787] = 32'h0;  // 32'hf1889d6c;
    ram_cell[     788] = 32'h0;  // 32'h2f82c397;
    ram_cell[     789] = 32'h0;  // 32'h3cb51ea6;
    ram_cell[     790] = 32'h0;  // 32'h27db9e20;
    ram_cell[     791] = 32'h0;  // 32'hd2969e13;
    ram_cell[     792] = 32'h0;  // 32'h323ea740;
    ram_cell[     793] = 32'h0;  // 32'h7e4ba222;
    ram_cell[     794] = 32'h0;  // 32'hcba9e5f7;
    ram_cell[     795] = 32'h0;  // 32'he31ad8fb;
    ram_cell[     796] = 32'h0;  // 32'h838bb2ec;
    ram_cell[     797] = 32'h0;  // 32'hc643d7d6;
    ram_cell[     798] = 32'h0;  // 32'ha33db138;
    ram_cell[     799] = 32'h0;  // 32'ha219b49f;
    ram_cell[     800] = 32'h0;  // 32'h144d3a04;
    ram_cell[     801] = 32'h0;  // 32'he390bf1a;
    ram_cell[     802] = 32'h0;  // 32'h0ccefb56;
    ram_cell[     803] = 32'h0;  // 32'h88a926a2;
    ram_cell[     804] = 32'h0;  // 32'h233e27e0;
    ram_cell[     805] = 32'h0;  // 32'h95b0548d;
    ram_cell[     806] = 32'h0;  // 32'ha755ae93;
    ram_cell[     807] = 32'h0;  // 32'he5e4b5c0;
    ram_cell[     808] = 32'h0;  // 32'h41b0ce7d;
    ram_cell[     809] = 32'h0;  // 32'h6e1a2dbc;
    ram_cell[     810] = 32'h0;  // 32'h68ee99cf;
    ram_cell[     811] = 32'h0;  // 32'hdc7919cc;
    ram_cell[     812] = 32'h0;  // 32'h4f1de42a;
    ram_cell[     813] = 32'h0;  // 32'h8b1631b0;
    ram_cell[     814] = 32'h0;  // 32'ha8237758;
    ram_cell[     815] = 32'h0;  // 32'h133e8e07;
    ram_cell[     816] = 32'h0;  // 32'hf69911d5;
    ram_cell[     817] = 32'h0;  // 32'heb7f628b;
    ram_cell[     818] = 32'h0;  // 32'h596f8422;
    ram_cell[     819] = 32'h0;  // 32'h9eecf94a;
    ram_cell[     820] = 32'h0;  // 32'hcdc3cafb;
    ram_cell[     821] = 32'h0;  // 32'h7f202fcc;
    ram_cell[     822] = 32'h0;  // 32'h1d3a5623;
    ram_cell[     823] = 32'h0;  // 32'ha95da0b1;
    ram_cell[     824] = 32'h0;  // 32'h8e41d725;
    ram_cell[     825] = 32'h0;  // 32'h6684b1a4;
    ram_cell[     826] = 32'h0;  // 32'h6388c3f6;
    ram_cell[     827] = 32'h0;  // 32'h2e232763;
    ram_cell[     828] = 32'h0;  // 32'hef56a911;
    ram_cell[     829] = 32'h0;  // 32'h8a7bb589;
    ram_cell[     830] = 32'h0;  // 32'h41c82166;
    ram_cell[     831] = 32'h0;  // 32'ha3721f9b;
    ram_cell[     832] = 32'h0;  // 32'h079e4ba2;
    ram_cell[     833] = 32'h0;  // 32'h4385a20b;
    ram_cell[     834] = 32'h0;  // 32'hd2ea2215;
    ram_cell[     835] = 32'h0;  // 32'hb025a2d9;
    ram_cell[     836] = 32'h0;  // 32'hb8792317;
    ram_cell[     837] = 32'h0;  // 32'h0c2958fe;
    ram_cell[     838] = 32'h0;  // 32'h4b56991e;
    ram_cell[     839] = 32'h0;  // 32'h0a2cf201;
    ram_cell[     840] = 32'h0;  // 32'h027b535a;
    ram_cell[     841] = 32'h0;  // 32'h3c4783fa;
    ram_cell[     842] = 32'h0;  // 32'h4dde677a;
    ram_cell[     843] = 32'h0;  // 32'h2b0aa494;
    ram_cell[     844] = 32'h0;  // 32'hb2c42ff9;
    ram_cell[     845] = 32'h0;  // 32'h6b64955e;
    ram_cell[     846] = 32'h0;  // 32'he5cd9898;
    ram_cell[     847] = 32'h0;  // 32'hc39a6ee5;
    ram_cell[     848] = 32'h0;  // 32'h9772e7d5;
    ram_cell[     849] = 32'h0;  // 32'hd10a82cf;
    ram_cell[     850] = 32'h0;  // 32'h37696df1;
    ram_cell[     851] = 32'h0;  // 32'hfc78f9b8;
    ram_cell[     852] = 32'h0;  // 32'hc808419f;
    ram_cell[     853] = 32'h0;  // 32'hc759c891;
    ram_cell[     854] = 32'h0;  // 32'h4eca227a;
    ram_cell[     855] = 32'h0;  // 32'hd4bde57f;
    ram_cell[     856] = 32'h0;  // 32'hf38e6192;
    ram_cell[     857] = 32'h0;  // 32'hc905be6e;
    ram_cell[     858] = 32'h0;  // 32'hfbd5e269;
    ram_cell[     859] = 32'h0;  // 32'h41153c8e;
    ram_cell[     860] = 32'h0;  // 32'hfbd48883;
    ram_cell[     861] = 32'h0;  // 32'hc43a6352;
    ram_cell[     862] = 32'h0;  // 32'hd1ebb042;
    ram_cell[     863] = 32'h0;  // 32'h0eb303a2;
    ram_cell[     864] = 32'h0;  // 32'h327a79f5;
    ram_cell[     865] = 32'h0;  // 32'he2a1bf5d;
    ram_cell[     866] = 32'h0;  // 32'hfafe0469;
    ram_cell[     867] = 32'h0;  // 32'h3cac6a5c;
    ram_cell[     868] = 32'h0;  // 32'h6b8eb11e;
    ram_cell[     869] = 32'h0;  // 32'hbb53876c;
    ram_cell[     870] = 32'h0;  // 32'h70810247;
    ram_cell[     871] = 32'h0;  // 32'hb056b7b0;
    ram_cell[     872] = 32'h0;  // 32'h1ba3f2a0;
    ram_cell[     873] = 32'h0;  // 32'h5ea1bc7f;
    ram_cell[     874] = 32'h0;  // 32'hc3db8998;
    ram_cell[     875] = 32'h0;  // 32'h236fcf6a;
    ram_cell[     876] = 32'h0;  // 32'h210e13f7;
    ram_cell[     877] = 32'h0;  // 32'hb06154e4;
    ram_cell[     878] = 32'h0;  // 32'hd499604d;
    ram_cell[     879] = 32'h0;  // 32'hc458a71d;
    ram_cell[     880] = 32'h0;  // 32'hf1d4f29f;
    ram_cell[     881] = 32'h0;  // 32'h306df2e3;
    ram_cell[     882] = 32'h0;  // 32'hd3b7c1cd;
    ram_cell[     883] = 32'h0;  // 32'h13eb4abf;
    ram_cell[     884] = 32'h0;  // 32'h64a62e23;
    ram_cell[     885] = 32'h0;  // 32'h7c1257ac;
    ram_cell[     886] = 32'h0;  // 32'h0ee25731;
    ram_cell[     887] = 32'h0;  // 32'hb1141eec;
    ram_cell[     888] = 32'h0;  // 32'he2881ce0;
    ram_cell[     889] = 32'h0;  // 32'h9b8bd1a6;
    ram_cell[     890] = 32'h0;  // 32'h25f680b7;
    ram_cell[     891] = 32'h0;  // 32'had1b4a3c;
    ram_cell[     892] = 32'h0;  // 32'hfd6ae631;
    ram_cell[     893] = 32'h0;  // 32'h4c6c7a2f;
    ram_cell[     894] = 32'h0;  // 32'hafe15cc3;
    ram_cell[     895] = 32'h0;  // 32'h19cac404;
    ram_cell[     896] = 32'h0;  // 32'ha0e78307;
    ram_cell[     897] = 32'h0;  // 32'h776ca76f;
    ram_cell[     898] = 32'h0;  // 32'h9c8b2b98;
    ram_cell[     899] = 32'h0;  // 32'h88a6702d;
    ram_cell[     900] = 32'h0;  // 32'h8cb8033a;
    ram_cell[     901] = 32'h0;  // 32'h39a82df2;
    ram_cell[     902] = 32'h0;  // 32'h0420b824;
    ram_cell[     903] = 32'h0;  // 32'hb3fb2e2d;
    ram_cell[     904] = 32'h0;  // 32'hf435e8d1;
    ram_cell[     905] = 32'h0;  // 32'he3ff6eeb;
    ram_cell[     906] = 32'h0;  // 32'h4b814454;
    ram_cell[     907] = 32'h0;  // 32'h621fb3c6;
    ram_cell[     908] = 32'h0;  // 32'hc7f292ee;
    ram_cell[     909] = 32'h0;  // 32'he676a481;
    ram_cell[     910] = 32'h0;  // 32'h171ca91c;
    ram_cell[     911] = 32'h0;  // 32'h81a474bc;
    ram_cell[     912] = 32'h0;  // 32'hd028b833;
    ram_cell[     913] = 32'h0;  // 32'ha0c1d2ea;
    ram_cell[     914] = 32'h0;  // 32'h3ee630db;
    ram_cell[     915] = 32'h0;  // 32'h11cae788;
    ram_cell[     916] = 32'h0;  // 32'h5af729e7;
    ram_cell[     917] = 32'h0;  // 32'h6b52643c;
    ram_cell[     918] = 32'h0;  // 32'h893423b1;
    ram_cell[     919] = 32'h0;  // 32'h59e1609a;
    ram_cell[     920] = 32'h0;  // 32'hbd397e57;
    ram_cell[     921] = 32'h0;  // 32'h5501fd93;
    ram_cell[     922] = 32'h0;  // 32'h813a6636;
    ram_cell[     923] = 32'h0;  // 32'he9bd7ff6;
    ram_cell[     924] = 32'h0;  // 32'h5a907008;
    ram_cell[     925] = 32'h0;  // 32'h9483b7b0;
    ram_cell[     926] = 32'h0;  // 32'h249c818b;
    ram_cell[     927] = 32'h0;  // 32'hb103095a;
    ram_cell[     928] = 32'h0;  // 32'h03ce202b;
    ram_cell[     929] = 32'h0;  // 32'hab1c0b66;
    ram_cell[     930] = 32'h0;  // 32'h97ee484c;
    ram_cell[     931] = 32'h0;  // 32'h10aa2a47;
    ram_cell[     932] = 32'h0;  // 32'he9e8e48d;
    ram_cell[     933] = 32'h0;  // 32'h90cdcc58;
    ram_cell[     934] = 32'h0;  // 32'h4f108a3e;
    ram_cell[     935] = 32'h0;  // 32'he25cde68;
    ram_cell[     936] = 32'h0;  // 32'h8a89fb6d;
    ram_cell[     937] = 32'h0;  // 32'hef98c0e4;
    ram_cell[     938] = 32'h0;  // 32'h32a72b6c;
    ram_cell[     939] = 32'h0;  // 32'h02b0f72b;
    ram_cell[     940] = 32'h0;  // 32'h902cbb78;
    ram_cell[     941] = 32'h0;  // 32'hcb429ebc;
    ram_cell[     942] = 32'h0;  // 32'h0859c3e9;
    ram_cell[     943] = 32'h0;  // 32'h52c3dc03;
    ram_cell[     944] = 32'h0;  // 32'hb039d82a;
    ram_cell[     945] = 32'h0;  // 32'hfb8450de;
    ram_cell[     946] = 32'h0;  // 32'h529026af;
    ram_cell[     947] = 32'h0;  // 32'hc2c66695;
    ram_cell[     948] = 32'h0;  // 32'hee3800bf;
    ram_cell[     949] = 32'h0;  // 32'h9327b457;
    ram_cell[     950] = 32'h0;  // 32'hc17014b7;
    ram_cell[     951] = 32'h0;  // 32'h6d8d379c;
    ram_cell[     952] = 32'h0;  // 32'hebf3f15b;
    ram_cell[     953] = 32'h0;  // 32'hb404d9d1;
    ram_cell[     954] = 32'h0;  // 32'hcfbc8235;
    ram_cell[     955] = 32'h0;  // 32'h999e150a;
    ram_cell[     956] = 32'h0;  // 32'h21c6b528;
    ram_cell[     957] = 32'h0;  // 32'h3c56903e;
    ram_cell[     958] = 32'h0;  // 32'h9a25c8ee;
    ram_cell[     959] = 32'h0;  // 32'h2480dd46;
    ram_cell[     960] = 32'h0;  // 32'h445b4b91;
    ram_cell[     961] = 32'h0;  // 32'h05369b8f;
    ram_cell[     962] = 32'h0;  // 32'ha4f2008f;
    ram_cell[     963] = 32'h0;  // 32'hbd0f0308;
    ram_cell[     964] = 32'h0;  // 32'ha93c5457;
    ram_cell[     965] = 32'h0;  // 32'h11aa8d56;
    ram_cell[     966] = 32'h0;  // 32'h10f53e67;
    ram_cell[     967] = 32'h0;  // 32'hfcb3c5d3;
    ram_cell[     968] = 32'h0;  // 32'h79cdb55e;
    ram_cell[     969] = 32'h0;  // 32'hda84a75f;
    ram_cell[     970] = 32'h0;  // 32'hbaf9f985;
    ram_cell[     971] = 32'h0;  // 32'h93f68ef3;
    ram_cell[     972] = 32'h0;  // 32'hb94565f8;
    ram_cell[     973] = 32'h0;  // 32'h42952160;
    ram_cell[     974] = 32'h0;  // 32'h5ed194fb;
    ram_cell[     975] = 32'h0;  // 32'hf0557d2e;
    ram_cell[     976] = 32'h0;  // 32'ha29584e4;
    ram_cell[     977] = 32'h0;  // 32'hd7c58b3b;
    ram_cell[     978] = 32'h0;  // 32'h98dd3212;
    ram_cell[     979] = 32'h0;  // 32'hd76c970e;
    ram_cell[     980] = 32'h0;  // 32'h104a76bc;
    ram_cell[     981] = 32'h0;  // 32'h8edc3e50;
    ram_cell[     982] = 32'h0;  // 32'h1379cc7e;
    ram_cell[     983] = 32'h0;  // 32'h771cb130;
    ram_cell[     984] = 32'h0;  // 32'h2163be22;
    ram_cell[     985] = 32'h0;  // 32'ha3b15172;
    ram_cell[     986] = 32'h0;  // 32'hf16c3a76;
    ram_cell[     987] = 32'h0;  // 32'h2c3d9aee;
    ram_cell[     988] = 32'h0;  // 32'hfcac824a;
    ram_cell[     989] = 32'h0;  // 32'h9fa806c4;
    ram_cell[     990] = 32'h0;  // 32'hfec964f8;
    ram_cell[     991] = 32'h0;  // 32'h613d66fa;
    ram_cell[     992] = 32'h0;  // 32'h5f63f104;
    ram_cell[     993] = 32'h0;  // 32'h8ac34e6e;
    ram_cell[     994] = 32'h0;  // 32'h273df5db;
    ram_cell[     995] = 32'h0;  // 32'heb3132c1;
    ram_cell[     996] = 32'h0;  // 32'h00090e40;
    ram_cell[     997] = 32'h0;  // 32'hdf6c8ac7;
    ram_cell[     998] = 32'h0;  // 32'h4a22f45f;
    ram_cell[     999] = 32'h0;  // 32'hfe1259c7;
    ram_cell[    1000] = 32'h0;  // 32'h99cf519c;
    ram_cell[    1001] = 32'h0;  // 32'h818644a6;
    ram_cell[    1002] = 32'h0;  // 32'h0e949afa;
    ram_cell[    1003] = 32'h0;  // 32'hc2b417e2;
    ram_cell[    1004] = 32'h0;  // 32'h29688288;
    ram_cell[    1005] = 32'h0;  // 32'h4b2bb48b;
    ram_cell[    1006] = 32'h0;  // 32'h359b4044;
    ram_cell[    1007] = 32'h0;  // 32'hf114c969;
    ram_cell[    1008] = 32'h0;  // 32'h9687ad85;
    ram_cell[    1009] = 32'h0;  // 32'h3d95f2ad;
    ram_cell[    1010] = 32'h0;  // 32'had850664;
    ram_cell[    1011] = 32'h0;  // 32'h03e84b91;
    ram_cell[    1012] = 32'h0;  // 32'h9135c0ea;
    ram_cell[    1013] = 32'h0;  // 32'h725eb307;
    ram_cell[    1014] = 32'h0;  // 32'h53bc802a;
    ram_cell[    1015] = 32'h0;  // 32'h5e9f5b2e;
    ram_cell[    1016] = 32'h0;  // 32'h079c65c6;
    ram_cell[    1017] = 32'h0;  // 32'h27193899;
    ram_cell[    1018] = 32'h0;  // 32'h6f091c22;
    ram_cell[    1019] = 32'h0;  // 32'ha1a2424e;
    ram_cell[    1020] = 32'h0;  // 32'h50fda19e;
    ram_cell[    1021] = 32'h0;  // 32'h08ec60c3;
    ram_cell[    1022] = 32'h0;  // 32'h4140f12e;
    ram_cell[    1023] = 32'h0;  // 32'hfc804446;
    ram_cell[    1024] = 32'h0;  // 32'hda247e31;
    ram_cell[    1025] = 32'h0;  // 32'hd2d99da3;
    ram_cell[    1026] = 32'h0;  // 32'h62e322d1;
    ram_cell[    1027] = 32'h0;  // 32'hfbd86e73;
    ram_cell[    1028] = 32'h0;  // 32'he135bb4f;
    ram_cell[    1029] = 32'h0;  // 32'hf10451ac;
    ram_cell[    1030] = 32'h0;  // 32'h8d484fa4;
    ram_cell[    1031] = 32'h0;  // 32'h94ff857f;
    ram_cell[    1032] = 32'h0;  // 32'h1ba19934;
    ram_cell[    1033] = 32'h0;  // 32'h59bef329;
    ram_cell[    1034] = 32'h0;  // 32'h49e480d8;
    ram_cell[    1035] = 32'h0;  // 32'h81f7c810;
    ram_cell[    1036] = 32'h0;  // 32'h0a309b96;
    ram_cell[    1037] = 32'h0;  // 32'ha07592fe;
    ram_cell[    1038] = 32'h0;  // 32'h6dae306a;
    ram_cell[    1039] = 32'h0;  // 32'hb243cc3b;
    ram_cell[    1040] = 32'h0;  // 32'hca5fa0d3;
    ram_cell[    1041] = 32'h0;  // 32'h41b8be1c;
    ram_cell[    1042] = 32'h0;  // 32'h5249de64;
    ram_cell[    1043] = 32'h0;  // 32'h22045b3b;
    ram_cell[    1044] = 32'h0;  // 32'hbd3405dd;
    ram_cell[    1045] = 32'h0;  // 32'h7051e172;
    ram_cell[    1046] = 32'h0;  // 32'h32ff7e1f;
    ram_cell[    1047] = 32'h0;  // 32'h49bd57e2;
    ram_cell[    1048] = 32'h0;  // 32'hf3cae9f0;
    ram_cell[    1049] = 32'h0;  // 32'hb5510bb1;
    ram_cell[    1050] = 32'h0;  // 32'h0099a909;
    ram_cell[    1051] = 32'h0;  // 32'hd24ee3c8;
    ram_cell[    1052] = 32'h0;  // 32'hb70a196b;
    ram_cell[    1053] = 32'h0;  // 32'h90c15084;
    ram_cell[    1054] = 32'h0;  // 32'h89dccb2f;
    ram_cell[    1055] = 32'h0;  // 32'h720cb5db;
    ram_cell[    1056] = 32'h0;  // 32'hefb8d4d2;
    ram_cell[    1057] = 32'h0;  // 32'hb1864de0;
    ram_cell[    1058] = 32'h0;  // 32'h8cdb9100;
    ram_cell[    1059] = 32'h0;  // 32'h56c04f9f;
    ram_cell[    1060] = 32'h0;  // 32'h183b8c80;
    ram_cell[    1061] = 32'h0;  // 32'h3c9fa89b;
    ram_cell[    1062] = 32'h0;  // 32'hff4030cc;
    ram_cell[    1063] = 32'h0;  // 32'h900ac951;
    ram_cell[    1064] = 32'h0;  // 32'h8ce3ec7a;
    ram_cell[    1065] = 32'h0;  // 32'h77e0bb25;
    ram_cell[    1066] = 32'h0;  // 32'hbf63ccf7;
    ram_cell[    1067] = 32'h0;  // 32'hef58780e;
    ram_cell[    1068] = 32'h0;  // 32'hc09ccb5c;
    ram_cell[    1069] = 32'h0;  // 32'h4c63c2c6;
    ram_cell[    1070] = 32'h0;  // 32'h5bcdbb1f;
    ram_cell[    1071] = 32'h0;  // 32'hd70c6d81;
    ram_cell[    1072] = 32'h0;  // 32'h028188c3;
    ram_cell[    1073] = 32'h0;  // 32'h576a1e79;
    ram_cell[    1074] = 32'h0;  // 32'h2a5fd2ce;
    ram_cell[    1075] = 32'h0;  // 32'hbf29927e;
    ram_cell[    1076] = 32'h0;  // 32'h1b98a2da;
    ram_cell[    1077] = 32'h0;  // 32'hcd652d87;
    ram_cell[    1078] = 32'h0;  // 32'h616c22a6;
    ram_cell[    1079] = 32'h0;  // 32'h71b52477;
    ram_cell[    1080] = 32'h0;  // 32'h21fe825e;
    ram_cell[    1081] = 32'h0;  // 32'h6699bb95;
    ram_cell[    1082] = 32'h0;  // 32'h048a0964;
    ram_cell[    1083] = 32'h0;  // 32'h6befd088;
    ram_cell[    1084] = 32'h0;  // 32'h23410233;
    ram_cell[    1085] = 32'h0;  // 32'h23b5f39a;
    ram_cell[    1086] = 32'h0;  // 32'hedfa35ff;
    ram_cell[    1087] = 32'h0;  // 32'h8c824458;
    ram_cell[    1088] = 32'h0;  // 32'hc5bbdc68;
    ram_cell[    1089] = 32'h0;  // 32'ha938c7c7;
    ram_cell[    1090] = 32'h0;  // 32'h12130bb7;
    ram_cell[    1091] = 32'h0;  // 32'h77652fe8;
    ram_cell[    1092] = 32'h0;  // 32'h7553975d;
    ram_cell[    1093] = 32'h0;  // 32'h5919ad8c;
    ram_cell[    1094] = 32'h0;  // 32'hf5a48b43;
    ram_cell[    1095] = 32'h0;  // 32'hf7d21ed8;
    ram_cell[    1096] = 32'h0;  // 32'h0b929255;
    ram_cell[    1097] = 32'h0;  // 32'h1344981a;
    ram_cell[    1098] = 32'h0;  // 32'h0707e67d;
    ram_cell[    1099] = 32'h0;  // 32'hefe26039;
    ram_cell[    1100] = 32'h0;  // 32'h641e1233;
    ram_cell[    1101] = 32'h0;  // 32'h2ced16e5;
    ram_cell[    1102] = 32'h0;  // 32'h4816ad79;
    ram_cell[    1103] = 32'h0;  // 32'h80198926;
    ram_cell[    1104] = 32'h0;  // 32'h51544b06;
    ram_cell[    1105] = 32'h0;  // 32'h3626b893;
    ram_cell[    1106] = 32'h0;  // 32'ha3d7b2b7;
    ram_cell[    1107] = 32'h0;  // 32'h61137a53;
    ram_cell[    1108] = 32'h0;  // 32'h6664cabf;
    ram_cell[    1109] = 32'h0;  // 32'ha315c914;
    ram_cell[    1110] = 32'h0;  // 32'hada21f0b;
    ram_cell[    1111] = 32'h0;  // 32'h43a75602;
    ram_cell[    1112] = 32'h0;  // 32'h06652392;
    ram_cell[    1113] = 32'h0;  // 32'hc43a989e;
    ram_cell[    1114] = 32'h0;  // 32'hfe379232;
    ram_cell[    1115] = 32'h0;  // 32'hae47f41e;
    ram_cell[    1116] = 32'h0;  // 32'h0dd69110;
    ram_cell[    1117] = 32'h0;  // 32'hdf1f81ef;
    ram_cell[    1118] = 32'h0;  // 32'hf9c8a364;
    ram_cell[    1119] = 32'h0;  // 32'hfd569603;
    ram_cell[    1120] = 32'h0;  // 32'hcb08dea4;
    ram_cell[    1121] = 32'h0;  // 32'had9f3949;
    ram_cell[    1122] = 32'h0;  // 32'hbd79cdd2;
    ram_cell[    1123] = 32'h0;  // 32'h6f2344b1;
    ram_cell[    1124] = 32'h0;  // 32'h30f6c7be;
    ram_cell[    1125] = 32'h0;  // 32'h6eae4276;
    ram_cell[    1126] = 32'h0;  // 32'hf1406f69;
    ram_cell[    1127] = 32'h0;  // 32'h62536722;
    ram_cell[    1128] = 32'h0;  // 32'h62d4c541;
    ram_cell[    1129] = 32'h0;  // 32'hf9d493f6;
    ram_cell[    1130] = 32'h0;  // 32'ha9c4cae0;
    ram_cell[    1131] = 32'h0;  // 32'h72e68b82;
    ram_cell[    1132] = 32'h0;  // 32'h8dba106f;
    ram_cell[    1133] = 32'h0;  // 32'h8620bd29;
    ram_cell[    1134] = 32'h0;  // 32'hdcb21957;
    ram_cell[    1135] = 32'h0;  // 32'h7baa235c;
    ram_cell[    1136] = 32'h0;  // 32'hf3c2d157;
    ram_cell[    1137] = 32'h0;  // 32'hc1200dfe;
    ram_cell[    1138] = 32'h0;  // 32'hce9606f6;
    ram_cell[    1139] = 32'h0;  // 32'h1169a5b5;
    ram_cell[    1140] = 32'h0;  // 32'h5c87aa08;
    ram_cell[    1141] = 32'h0;  // 32'h31f5eed1;
    ram_cell[    1142] = 32'h0;  // 32'h72ddc00f;
    ram_cell[    1143] = 32'h0;  // 32'h1e232ed2;
    ram_cell[    1144] = 32'h0;  // 32'h59905c8c;
    ram_cell[    1145] = 32'h0;  // 32'h93eccb83;
    ram_cell[    1146] = 32'h0;  // 32'h950932c1;
    ram_cell[    1147] = 32'h0;  // 32'h4ac92a12;
    ram_cell[    1148] = 32'h0;  // 32'hba5d2c84;
    ram_cell[    1149] = 32'h0;  // 32'hf04c372b;
    ram_cell[    1150] = 32'h0;  // 32'h68c9ab76;
    ram_cell[    1151] = 32'h0;  // 32'h09823647;
    ram_cell[    1152] = 32'h0;  // 32'h0a457dff;
    ram_cell[    1153] = 32'h0;  // 32'hd0c1eed6;
    ram_cell[    1154] = 32'h0;  // 32'hb8a10a12;
    ram_cell[    1155] = 32'h0;  // 32'h01475cfd;
    ram_cell[    1156] = 32'h0;  // 32'h955ccf69;
    ram_cell[    1157] = 32'h0;  // 32'h29d7affb;
    ram_cell[    1158] = 32'h0;  // 32'hb48c5aa6;
    ram_cell[    1159] = 32'h0;  // 32'h940e246a;
    ram_cell[    1160] = 32'h0;  // 32'h204be4ac;
    ram_cell[    1161] = 32'h0;  // 32'h2bf42c6e;
    ram_cell[    1162] = 32'h0;  // 32'h9b7921a9;
    ram_cell[    1163] = 32'h0;  // 32'h5b2dd798;
    ram_cell[    1164] = 32'h0;  // 32'hf6a3c395;
    ram_cell[    1165] = 32'h0;  // 32'ha3c674ba;
    ram_cell[    1166] = 32'h0;  // 32'hb3c10c92;
    ram_cell[    1167] = 32'h0;  // 32'h39c36a85;
    ram_cell[    1168] = 32'h0;  // 32'hbb55e7d4;
    ram_cell[    1169] = 32'h0;  // 32'hd5d2a9e9;
    ram_cell[    1170] = 32'h0;  // 32'heb8a5fd9;
    ram_cell[    1171] = 32'h0;  // 32'h275dca75;
    ram_cell[    1172] = 32'h0;  // 32'h56b293b2;
    ram_cell[    1173] = 32'h0;  // 32'h03b889bc;
    ram_cell[    1174] = 32'h0;  // 32'h84d69e8e;
    ram_cell[    1175] = 32'h0;  // 32'hfef643b6;
    ram_cell[    1176] = 32'h0;  // 32'h34b96fe5;
    ram_cell[    1177] = 32'h0;  // 32'h8f872db1;
    ram_cell[    1178] = 32'h0;  // 32'h420fca7b;
    ram_cell[    1179] = 32'h0;  // 32'h639578f1;
    ram_cell[    1180] = 32'h0;  // 32'h9f146b39;
    ram_cell[    1181] = 32'h0;  // 32'hdd3bcb77;
    ram_cell[    1182] = 32'h0;  // 32'h26d6b47d;
    ram_cell[    1183] = 32'h0;  // 32'h10ed5672;
    ram_cell[    1184] = 32'h0;  // 32'hf419162b;
    ram_cell[    1185] = 32'h0;  // 32'h32bb0ce4;
    ram_cell[    1186] = 32'h0;  // 32'h81deab9c;
    ram_cell[    1187] = 32'h0;  // 32'hdd8cc51f;
    ram_cell[    1188] = 32'h0;  // 32'h8c8e3156;
    ram_cell[    1189] = 32'h0;  // 32'hb7d5638f;
    ram_cell[    1190] = 32'h0;  // 32'h46f721ff;
    ram_cell[    1191] = 32'h0;  // 32'h220a03f8;
    ram_cell[    1192] = 32'h0;  // 32'h8c9da1d1;
    ram_cell[    1193] = 32'h0;  // 32'h21a9763b;
    ram_cell[    1194] = 32'h0;  // 32'ha777f747;
    ram_cell[    1195] = 32'h0;  // 32'hcc860c40;
    ram_cell[    1196] = 32'h0;  // 32'he1f81766;
    ram_cell[    1197] = 32'h0;  // 32'h02f54a8a;
    ram_cell[    1198] = 32'h0;  // 32'hd1bab517;
    ram_cell[    1199] = 32'h0;  // 32'hc0e2b7a0;
    ram_cell[    1200] = 32'h0;  // 32'h722d8f75;
    ram_cell[    1201] = 32'h0;  // 32'hc6233ecb;
    ram_cell[    1202] = 32'h0;  // 32'hb0e6183c;
    ram_cell[    1203] = 32'h0;  // 32'hac5b9a11;
    ram_cell[    1204] = 32'h0;  // 32'hf974b027;
    ram_cell[    1205] = 32'h0;  // 32'h6763825a;
    ram_cell[    1206] = 32'h0;  // 32'h922f56f2;
    ram_cell[    1207] = 32'h0;  // 32'h8757d550;
    ram_cell[    1208] = 32'h0;  // 32'ha038bb79;
    ram_cell[    1209] = 32'h0;  // 32'hcd10d9ae;
    ram_cell[    1210] = 32'h0;  // 32'h5ee0555c;
    ram_cell[    1211] = 32'h0;  // 32'h086b5096;
    ram_cell[    1212] = 32'h0;  // 32'h0d59ce36;
    ram_cell[    1213] = 32'h0;  // 32'h564b7433;
    ram_cell[    1214] = 32'h0;  // 32'hff03a604;
    ram_cell[    1215] = 32'h0;  // 32'h99075ddc;
    ram_cell[    1216] = 32'h0;  // 32'h64c61a8a;
    ram_cell[    1217] = 32'h0;  // 32'h0386c04b;
    ram_cell[    1218] = 32'h0;  // 32'he6fcfbcf;
    ram_cell[    1219] = 32'h0;  // 32'h15bbb0a9;
    ram_cell[    1220] = 32'h0;  // 32'hc306aa65;
    ram_cell[    1221] = 32'h0;  // 32'h777ca51d;
    ram_cell[    1222] = 32'h0;  // 32'he068d91d;
    ram_cell[    1223] = 32'h0;  // 32'h5a776075;
    ram_cell[    1224] = 32'h0;  // 32'hcd9d4d30;
    ram_cell[    1225] = 32'h0;  // 32'hc5c58189;
    ram_cell[    1226] = 32'h0;  // 32'h6e7c0bcd;
    ram_cell[    1227] = 32'h0;  // 32'ha6169d02;
    ram_cell[    1228] = 32'h0;  // 32'hc75ccfaa;
    ram_cell[    1229] = 32'h0;  // 32'h4e673380;
    ram_cell[    1230] = 32'h0;  // 32'h5500eec1;
    ram_cell[    1231] = 32'h0;  // 32'hf7bf5fda;
    ram_cell[    1232] = 32'h0;  // 32'h357fd240;
    ram_cell[    1233] = 32'h0;  // 32'h54720aee;
    ram_cell[    1234] = 32'h0;  // 32'h93c38ed2;
    ram_cell[    1235] = 32'h0;  // 32'hdc955b27;
    ram_cell[    1236] = 32'h0;  // 32'h1d2063cf;
    ram_cell[    1237] = 32'h0;  // 32'h87bf7be7;
    ram_cell[    1238] = 32'h0;  // 32'hadda7091;
    ram_cell[    1239] = 32'h0;  // 32'h49e417de;
    ram_cell[    1240] = 32'h0;  // 32'h78b94061;
    ram_cell[    1241] = 32'h0;  // 32'h39cd0ccf;
    ram_cell[    1242] = 32'h0;  // 32'h9aa80641;
    ram_cell[    1243] = 32'h0;  // 32'h0ffc9cb4;
    ram_cell[    1244] = 32'h0;  // 32'h374a697d;
    ram_cell[    1245] = 32'h0;  // 32'hb071dd61;
    ram_cell[    1246] = 32'h0;  // 32'h6cf13fb1;
    ram_cell[    1247] = 32'h0;  // 32'ha6616dfd;
    ram_cell[    1248] = 32'h0;  // 32'hf39ad673;
    ram_cell[    1249] = 32'h0;  // 32'hf393b2aa;
    ram_cell[    1250] = 32'h0;  // 32'he34a225b;
    ram_cell[    1251] = 32'h0;  // 32'h1a2c8505;
    ram_cell[    1252] = 32'h0;  // 32'ha2393106;
    ram_cell[    1253] = 32'h0;  // 32'h3c9be45d;
    ram_cell[    1254] = 32'h0;  // 32'h98caa282;
    ram_cell[    1255] = 32'h0;  // 32'h89427f5a;
    ram_cell[    1256] = 32'h0;  // 32'h082a3b76;
    ram_cell[    1257] = 32'h0;  // 32'h8b95a1fc;
    ram_cell[    1258] = 32'h0;  // 32'h46da5484;
    ram_cell[    1259] = 32'h0;  // 32'habf54b99;
    ram_cell[    1260] = 32'h0;  // 32'h88e4c415;
    ram_cell[    1261] = 32'h0;  // 32'h1c13cced;
    ram_cell[    1262] = 32'h0;  // 32'h1a712983;
    ram_cell[    1263] = 32'h0;  // 32'he65f95c8;
    ram_cell[    1264] = 32'h0;  // 32'h882bdba0;
    ram_cell[    1265] = 32'h0;  // 32'h39e7aea5;
    ram_cell[    1266] = 32'h0;  // 32'hf9ff0d24;
    ram_cell[    1267] = 32'h0;  // 32'hae505188;
    ram_cell[    1268] = 32'h0;  // 32'hc93a8ec9;
    ram_cell[    1269] = 32'h0;  // 32'hbaaaf908;
    ram_cell[    1270] = 32'h0;  // 32'hab8868f4;
    ram_cell[    1271] = 32'h0;  // 32'he49a3346;
    ram_cell[    1272] = 32'h0;  // 32'h371c8e60;
    ram_cell[    1273] = 32'h0;  // 32'h3597a0ff;
    ram_cell[    1274] = 32'h0;  // 32'h7f25969a;
    ram_cell[    1275] = 32'h0;  // 32'h2ad287b4;
    ram_cell[    1276] = 32'h0;  // 32'hc1f0ea0a;
    ram_cell[    1277] = 32'h0;  // 32'h1ddd5a1f;
    ram_cell[    1278] = 32'h0;  // 32'hc7e0061c;
    ram_cell[    1279] = 32'h0;  // 32'h2c2919f6;
    ram_cell[    1280] = 32'h0;  // 32'h4ebfae00;
    ram_cell[    1281] = 32'h0;  // 32'hc67a572d;
    ram_cell[    1282] = 32'h0;  // 32'h8a884663;
    ram_cell[    1283] = 32'h0;  // 32'h29a2a445;
    ram_cell[    1284] = 32'h0;  // 32'h573b1a0c;
    ram_cell[    1285] = 32'h0;  // 32'h7a0038c4;
    ram_cell[    1286] = 32'h0;  // 32'h3f2d704b;
    ram_cell[    1287] = 32'h0;  // 32'hf0bf39b0;
    ram_cell[    1288] = 32'h0;  // 32'h59d39395;
    ram_cell[    1289] = 32'h0;  // 32'hca9c4b45;
    ram_cell[    1290] = 32'h0;  // 32'h3588177c;
    ram_cell[    1291] = 32'h0;  // 32'hb0052e3b;
    ram_cell[    1292] = 32'h0;  // 32'hae0ac1c9;
    ram_cell[    1293] = 32'h0;  // 32'h9e267b22;
    ram_cell[    1294] = 32'h0;  // 32'hce86b946;
    ram_cell[    1295] = 32'h0;  // 32'h753aaaee;
    ram_cell[    1296] = 32'h0;  // 32'h892101bb;
    ram_cell[    1297] = 32'h0;  // 32'hb137dfb2;
    ram_cell[    1298] = 32'h0;  // 32'h18ae1454;
    ram_cell[    1299] = 32'h0;  // 32'hfef492e4;
    ram_cell[    1300] = 32'h0;  // 32'h48225973;
    ram_cell[    1301] = 32'h0;  // 32'hbe6a4e3a;
    ram_cell[    1302] = 32'h0;  // 32'had8aa657;
    ram_cell[    1303] = 32'h0;  // 32'heece95a2;
    ram_cell[    1304] = 32'h0;  // 32'h73d5d3fb;
    ram_cell[    1305] = 32'h0;  // 32'h87a2f2e1;
    ram_cell[    1306] = 32'h0;  // 32'h25c2f435;
    ram_cell[    1307] = 32'h0;  // 32'h34bc795f;
    ram_cell[    1308] = 32'h0;  // 32'hfd276196;
    ram_cell[    1309] = 32'h0;  // 32'h07170067;
    ram_cell[    1310] = 32'h0;  // 32'h30913d8d;
    ram_cell[    1311] = 32'h0;  // 32'h4731e631;
    ram_cell[    1312] = 32'h0;  // 32'hc2928a6e;
    ram_cell[    1313] = 32'h0;  // 32'h52146786;
    ram_cell[    1314] = 32'h0;  // 32'hc384c1d3;
    ram_cell[    1315] = 32'h0;  // 32'ha6c292fb;
    ram_cell[    1316] = 32'h0;  // 32'h67eebcd9;
    ram_cell[    1317] = 32'h0;  // 32'h104d97ff;
    ram_cell[    1318] = 32'h0;  // 32'h7b669e95;
    ram_cell[    1319] = 32'h0;  // 32'hffa3f38f;
    ram_cell[    1320] = 32'h0;  // 32'h718ad383;
    ram_cell[    1321] = 32'h0;  // 32'h9eab0d5b;
    ram_cell[    1322] = 32'h0;  // 32'h5a6e478d;
    ram_cell[    1323] = 32'h0;  // 32'hbb121d02;
    ram_cell[    1324] = 32'h0;  // 32'he74fa7f1;
    ram_cell[    1325] = 32'h0;  // 32'h4f82ebc6;
    ram_cell[    1326] = 32'h0;  // 32'ha9a72a24;
    ram_cell[    1327] = 32'h0;  // 32'h3ee404df;
    ram_cell[    1328] = 32'h0;  // 32'hf48bc028;
    ram_cell[    1329] = 32'h0;  // 32'hf6e3d7ae;
    ram_cell[    1330] = 32'h0;  // 32'he81c7593;
    ram_cell[    1331] = 32'h0;  // 32'hfb0134c6;
    ram_cell[    1332] = 32'h0;  // 32'h9d7f96f9;
    ram_cell[    1333] = 32'h0;  // 32'h7fc8d611;
    ram_cell[    1334] = 32'h0;  // 32'h6f358b0c;
    ram_cell[    1335] = 32'h0;  // 32'ha3b1a629;
    ram_cell[    1336] = 32'h0;  // 32'h5a2dcf4d;
    ram_cell[    1337] = 32'h0;  // 32'h4380a9a3;
    ram_cell[    1338] = 32'h0;  // 32'h40a57047;
    ram_cell[    1339] = 32'h0;  // 32'he1357590;
    ram_cell[    1340] = 32'h0;  // 32'h94e89eab;
    ram_cell[    1341] = 32'h0;  // 32'h3da19ba9;
    ram_cell[    1342] = 32'h0;  // 32'hc27a4b8d;
    ram_cell[    1343] = 32'h0;  // 32'h5bcaaf01;
    ram_cell[    1344] = 32'h0;  // 32'h4c031068;
    ram_cell[    1345] = 32'h0;  // 32'he9ae4c62;
    ram_cell[    1346] = 32'h0;  // 32'h6f77b1b6;
    ram_cell[    1347] = 32'h0;  // 32'h9d051503;
    ram_cell[    1348] = 32'h0;  // 32'haf3965b3;
    ram_cell[    1349] = 32'h0;  // 32'h8aca67ab;
    ram_cell[    1350] = 32'h0;  // 32'h711ba6f5;
    ram_cell[    1351] = 32'h0;  // 32'hc4817bea;
    ram_cell[    1352] = 32'h0;  // 32'hcc17ef79;
    ram_cell[    1353] = 32'h0;  // 32'h54213eb4;
    ram_cell[    1354] = 32'h0;  // 32'h0c788c00;
    ram_cell[    1355] = 32'h0;  // 32'hca783e67;
    ram_cell[    1356] = 32'h0;  // 32'hdb6001cc;
    ram_cell[    1357] = 32'h0;  // 32'h1d291b08;
    ram_cell[    1358] = 32'h0;  // 32'hd94a747b;
    ram_cell[    1359] = 32'h0;  // 32'h9bbbfad4;
    ram_cell[    1360] = 32'h0;  // 32'h746affad;
    ram_cell[    1361] = 32'h0;  // 32'he9d46fbc;
    ram_cell[    1362] = 32'h0;  // 32'h1fbd9d12;
    ram_cell[    1363] = 32'h0;  // 32'h41868e48;
    ram_cell[    1364] = 32'h0;  // 32'h6ace89bc;
    ram_cell[    1365] = 32'h0;  // 32'hccc5d920;
    ram_cell[    1366] = 32'h0;  // 32'h04dd623c;
    ram_cell[    1367] = 32'h0;  // 32'h35d10610;
    ram_cell[    1368] = 32'h0;  // 32'h39ec48e6;
    ram_cell[    1369] = 32'h0;  // 32'h0bcd804b;
    ram_cell[    1370] = 32'h0;  // 32'hbafc6cb9;
    ram_cell[    1371] = 32'h0;  // 32'h588c1607;
    ram_cell[    1372] = 32'h0;  // 32'h8f90d02f;
    ram_cell[    1373] = 32'h0;  // 32'h3fdfaed6;
    ram_cell[    1374] = 32'h0;  // 32'h3dee3312;
    ram_cell[    1375] = 32'h0;  // 32'h5bc8e968;
    ram_cell[    1376] = 32'h0;  // 32'hd4887217;
    ram_cell[    1377] = 32'h0;  // 32'h8a9ba5ca;
    ram_cell[    1378] = 32'h0;  // 32'hc86e3336;
    ram_cell[    1379] = 32'h0;  // 32'he0a89724;
    ram_cell[    1380] = 32'h0;  // 32'hc6a16553;
    ram_cell[    1381] = 32'h0;  // 32'hf7e5cba5;
    ram_cell[    1382] = 32'h0;  // 32'hc849e544;
    ram_cell[    1383] = 32'h0;  // 32'hc8f43720;
    ram_cell[    1384] = 32'h0;  // 32'hc137b25c;
    ram_cell[    1385] = 32'h0;  // 32'hadeaff30;
    ram_cell[    1386] = 32'h0;  // 32'he48287f3;
    ram_cell[    1387] = 32'h0;  // 32'h3eea81cd;
    ram_cell[    1388] = 32'h0;  // 32'h937ec355;
    ram_cell[    1389] = 32'h0;  // 32'h314134ba;
    ram_cell[    1390] = 32'h0;  // 32'h543a058f;
    ram_cell[    1391] = 32'h0;  // 32'h837a45dc;
    ram_cell[    1392] = 32'h0;  // 32'hd09b4b35;
    ram_cell[    1393] = 32'h0;  // 32'hf5f7908a;
    ram_cell[    1394] = 32'h0;  // 32'h06d5c89c;
    ram_cell[    1395] = 32'h0;  // 32'hb6d22999;
    ram_cell[    1396] = 32'h0;  // 32'ha59cd64a;
    ram_cell[    1397] = 32'h0;  // 32'h9305628e;
    ram_cell[    1398] = 32'h0;  // 32'h60e1d1f0;
    ram_cell[    1399] = 32'h0;  // 32'h65e640a6;
    ram_cell[    1400] = 32'h0;  // 32'h279de8c5;
    ram_cell[    1401] = 32'h0;  // 32'hc7fcf2eb;
    ram_cell[    1402] = 32'h0;  // 32'h0243d2f1;
    ram_cell[    1403] = 32'h0;  // 32'h01983b08;
    ram_cell[    1404] = 32'h0;  // 32'h416ef3c5;
    ram_cell[    1405] = 32'h0;  // 32'h7807a494;
    ram_cell[    1406] = 32'h0;  // 32'hb53d76ca;
    ram_cell[    1407] = 32'h0;  // 32'hb141a678;
    ram_cell[    1408] = 32'h0;  // 32'hcf01e323;
    ram_cell[    1409] = 32'h0;  // 32'he3f8ea1b;
    ram_cell[    1410] = 32'h0;  // 32'h5da251ea;
    ram_cell[    1411] = 32'h0;  // 32'h785356eb;
    ram_cell[    1412] = 32'h0;  // 32'h719c6725;
    ram_cell[    1413] = 32'h0;  // 32'h8b0a64b6;
    ram_cell[    1414] = 32'h0;  // 32'hd08eb7b9;
    ram_cell[    1415] = 32'h0;  // 32'he621c9fc;
    ram_cell[    1416] = 32'h0;  // 32'h0c131bf5;
    ram_cell[    1417] = 32'h0;  // 32'h54d8cf8d;
    ram_cell[    1418] = 32'h0;  // 32'h2630ad07;
    ram_cell[    1419] = 32'h0;  // 32'hd4f67ab6;
    ram_cell[    1420] = 32'h0;  // 32'hb3b54dd6;
    ram_cell[    1421] = 32'h0;  // 32'h93490f2c;
    ram_cell[    1422] = 32'h0;  // 32'heb36739d;
    ram_cell[    1423] = 32'h0;  // 32'h19df57ae;
    ram_cell[    1424] = 32'h0;  // 32'h83db8f83;
    ram_cell[    1425] = 32'h0;  // 32'h9e7554bc;
    ram_cell[    1426] = 32'h0;  // 32'hf5eeadfd;
    ram_cell[    1427] = 32'h0;  // 32'hf5113cfe;
    ram_cell[    1428] = 32'h0;  // 32'h51718403;
    ram_cell[    1429] = 32'h0;  // 32'h7ef634da;
    ram_cell[    1430] = 32'h0;  // 32'h8c0b25dd;
    ram_cell[    1431] = 32'h0;  // 32'h6ecee6a6;
    ram_cell[    1432] = 32'h0;  // 32'hc58c2a1c;
    ram_cell[    1433] = 32'h0;  // 32'h5359d7d5;
    ram_cell[    1434] = 32'h0;  // 32'h4b734732;
    ram_cell[    1435] = 32'h0;  // 32'h1458e3d5;
    ram_cell[    1436] = 32'h0;  // 32'h89f468bb;
    ram_cell[    1437] = 32'h0;  // 32'h83ea8a4e;
    ram_cell[    1438] = 32'h0;  // 32'h26e4429f;
    ram_cell[    1439] = 32'h0;  // 32'h80b884b1;
    ram_cell[    1440] = 32'h0;  // 32'hbcd7c3e7;
    ram_cell[    1441] = 32'h0;  // 32'hafbc8688;
    ram_cell[    1442] = 32'h0;  // 32'hc31cd92e;
    ram_cell[    1443] = 32'h0;  // 32'h0364b820;
    ram_cell[    1444] = 32'h0;  // 32'ha1d496d7;
    ram_cell[    1445] = 32'h0;  // 32'hb319247c;
    ram_cell[    1446] = 32'h0;  // 32'h9249be0c;
    ram_cell[    1447] = 32'h0;  // 32'h6234afcf;
    ram_cell[    1448] = 32'h0;  // 32'h966c30a7;
    ram_cell[    1449] = 32'h0;  // 32'hf688c846;
    ram_cell[    1450] = 32'h0;  // 32'h74b6ea91;
    ram_cell[    1451] = 32'h0;  // 32'ha69078b5;
    ram_cell[    1452] = 32'h0;  // 32'h3dac26d2;
    ram_cell[    1453] = 32'h0;  // 32'h7748e1d2;
    ram_cell[    1454] = 32'h0;  // 32'h653d7286;
    ram_cell[    1455] = 32'h0;  // 32'h4d9a3871;
    ram_cell[    1456] = 32'h0;  // 32'h07c505dc;
    ram_cell[    1457] = 32'h0;  // 32'h38c3cef7;
    ram_cell[    1458] = 32'h0;  // 32'hcf7b23d5;
    ram_cell[    1459] = 32'h0;  // 32'h066bef1e;
    ram_cell[    1460] = 32'h0;  // 32'h1516cda9;
    ram_cell[    1461] = 32'h0;  // 32'h6edb0344;
    ram_cell[    1462] = 32'h0;  // 32'h6bf2bd2f;
    ram_cell[    1463] = 32'h0;  // 32'hf8dcf20f;
    ram_cell[    1464] = 32'h0;  // 32'ha7639666;
    ram_cell[    1465] = 32'h0;  // 32'h35752e3e;
    ram_cell[    1466] = 32'h0;  // 32'h3085333a;
    ram_cell[    1467] = 32'h0;  // 32'h4ecada78;
    ram_cell[    1468] = 32'h0;  // 32'h334e8779;
    ram_cell[    1469] = 32'h0;  // 32'hf8524d64;
    ram_cell[    1470] = 32'h0;  // 32'h7b5c497b;
    ram_cell[    1471] = 32'h0;  // 32'h65ece242;
    ram_cell[    1472] = 32'h0;  // 32'haa121730;
    ram_cell[    1473] = 32'h0;  // 32'hfc8a40d6;
    ram_cell[    1474] = 32'h0;  // 32'heba7157f;
    ram_cell[    1475] = 32'h0;  // 32'h48d551fb;
    ram_cell[    1476] = 32'h0;  // 32'hbdd77527;
    ram_cell[    1477] = 32'h0;  // 32'h67dea4b7;
    ram_cell[    1478] = 32'h0;  // 32'h1383f949;
    ram_cell[    1479] = 32'h0;  // 32'h6fed0468;
    ram_cell[    1480] = 32'h0;  // 32'he9d4761d;
    ram_cell[    1481] = 32'h0;  // 32'hd1f72552;
    ram_cell[    1482] = 32'h0;  // 32'h3228c33b;
    ram_cell[    1483] = 32'h0;  // 32'h8945b854;
    ram_cell[    1484] = 32'h0;  // 32'h980bc45c;
    ram_cell[    1485] = 32'h0;  // 32'h83d265ba;
    ram_cell[    1486] = 32'h0;  // 32'he37c1bb9;
    ram_cell[    1487] = 32'h0;  // 32'h37994757;
    ram_cell[    1488] = 32'h0;  // 32'he68c8006;
    ram_cell[    1489] = 32'h0;  // 32'he20e30c1;
    ram_cell[    1490] = 32'h0;  // 32'h2627ff00;
    ram_cell[    1491] = 32'h0;  // 32'h6a3f105e;
    ram_cell[    1492] = 32'h0;  // 32'hbcf9eee0;
    ram_cell[    1493] = 32'h0;  // 32'h619990a9;
    ram_cell[    1494] = 32'h0;  // 32'hbeea0dcd;
    ram_cell[    1495] = 32'h0;  // 32'h4f89b179;
    ram_cell[    1496] = 32'h0;  // 32'h81cfe0a5;
    ram_cell[    1497] = 32'h0;  // 32'h2aefa644;
    ram_cell[    1498] = 32'h0;  // 32'hd137647e;
    ram_cell[    1499] = 32'h0;  // 32'h9a7d07c8;
    ram_cell[    1500] = 32'h0;  // 32'h2bfb726a;
    ram_cell[    1501] = 32'h0;  // 32'h75f04d49;
    ram_cell[    1502] = 32'h0;  // 32'h7a3aff13;
    ram_cell[    1503] = 32'h0;  // 32'hdabdfe1d;
    ram_cell[    1504] = 32'h0;  // 32'h6d61e92d;
    ram_cell[    1505] = 32'h0;  // 32'hd13276d6;
    ram_cell[    1506] = 32'h0;  // 32'h2a2aa137;
    ram_cell[    1507] = 32'h0;  // 32'h55f5d48d;
    ram_cell[    1508] = 32'h0;  // 32'ha84a0d34;
    ram_cell[    1509] = 32'h0;  // 32'hc2889fee;
    ram_cell[    1510] = 32'h0;  // 32'hc098c708;
    ram_cell[    1511] = 32'h0;  // 32'h3aaabf70;
    ram_cell[    1512] = 32'h0;  // 32'h12170d5d;
    ram_cell[    1513] = 32'h0;  // 32'h8d627ac0;
    ram_cell[    1514] = 32'h0;  // 32'h5c15fd9c;
    ram_cell[    1515] = 32'h0;  // 32'hf61fec53;
    ram_cell[    1516] = 32'h0;  // 32'h964b6f75;
    ram_cell[    1517] = 32'h0;  // 32'h0791ea6e;
    ram_cell[    1518] = 32'h0;  // 32'h6cbec8a2;
    ram_cell[    1519] = 32'h0;  // 32'h8bdca4d0;
    ram_cell[    1520] = 32'h0;  // 32'he48efe07;
    ram_cell[    1521] = 32'h0;  // 32'hcce49713;
    ram_cell[    1522] = 32'h0;  // 32'h98e8fdbc;
    ram_cell[    1523] = 32'h0;  // 32'h30a2b276;
    ram_cell[    1524] = 32'h0;  // 32'h3f65c377;
    ram_cell[    1525] = 32'h0;  // 32'h403a2d73;
    ram_cell[    1526] = 32'h0;  // 32'hfbad23db;
    ram_cell[    1527] = 32'h0;  // 32'he967143b;
    ram_cell[    1528] = 32'h0;  // 32'h098c6a33;
    ram_cell[    1529] = 32'h0;  // 32'h9f58303f;
    ram_cell[    1530] = 32'h0;  // 32'h0b1dc1a0;
    ram_cell[    1531] = 32'h0;  // 32'hb57028d7;
    ram_cell[    1532] = 32'h0;  // 32'h380bb433;
    ram_cell[    1533] = 32'h0;  // 32'h0e518d21;
    ram_cell[    1534] = 32'h0;  // 32'h4569dd6c;
    ram_cell[    1535] = 32'h0;  // 32'h26f4c5a7;
    ram_cell[    1536] = 32'h0;  // 32'he9b6b070;
    ram_cell[    1537] = 32'h0;  // 32'hcd53ce27;
    ram_cell[    1538] = 32'h0;  // 32'h0c92b672;
    ram_cell[    1539] = 32'h0;  // 32'h30ba5f48;
    ram_cell[    1540] = 32'h0;  // 32'h3bbdd28d;
    ram_cell[    1541] = 32'h0;  // 32'h1a9f6d96;
    ram_cell[    1542] = 32'h0;  // 32'h6373bc87;
    ram_cell[    1543] = 32'h0;  // 32'h48aad4cb;
    ram_cell[    1544] = 32'h0;  // 32'h2a2c82f3;
    ram_cell[    1545] = 32'h0;  // 32'h6f8aea73;
    ram_cell[    1546] = 32'h0;  // 32'h213fcb6b;
    ram_cell[    1547] = 32'h0;  // 32'h0d3f3c25;
    ram_cell[    1548] = 32'h0;  // 32'h1b7e497a;
    ram_cell[    1549] = 32'h0;  // 32'hd96306e0;
    ram_cell[    1550] = 32'h0;  // 32'h40097cdb;
    ram_cell[    1551] = 32'h0;  // 32'h2c3a9824;
    ram_cell[    1552] = 32'h0;  // 32'ha45a0311;
    ram_cell[    1553] = 32'h0;  // 32'h57d1b1d1;
    ram_cell[    1554] = 32'h0;  // 32'haa2b762f;
    ram_cell[    1555] = 32'h0;  // 32'h8602ca7c;
    ram_cell[    1556] = 32'h0;  // 32'h3b795bdb;
    ram_cell[    1557] = 32'h0;  // 32'h4eb94fac;
    ram_cell[    1558] = 32'h0;  // 32'h7bb5d95d;
    ram_cell[    1559] = 32'h0;  // 32'h100fb067;
    ram_cell[    1560] = 32'h0;  // 32'h558fe166;
    ram_cell[    1561] = 32'h0;  // 32'hb567167f;
    ram_cell[    1562] = 32'h0;  // 32'h5cf5a199;
    ram_cell[    1563] = 32'h0;  // 32'h02c3ba16;
    ram_cell[    1564] = 32'h0;  // 32'hb60661ec;
    ram_cell[    1565] = 32'h0;  // 32'h13580b74;
    ram_cell[    1566] = 32'h0;  // 32'hb40bcc7b;
    ram_cell[    1567] = 32'h0;  // 32'he7e22c5d;
    ram_cell[    1568] = 32'h0;  // 32'hb0bdbc3e;
    ram_cell[    1569] = 32'h0;  // 32'h89637ab2;
    ram_cell[    1570] = 32'h0;  // 32'h82e91d7d;
    ram_cell[    1571] = 32'h0;  // 32'h3c9811b1;
    ram_cell[    1572] = 32'h0;  // 32'h9f4a5368;
    ram_cell[    1573] = 32'h0;  // 32'hee0154b8;
    ram_cell[    1574] = 32'h0;  // 32'h4640a97c;
    ram_cell[    1575] = 32'h0;  // 32'h193468f4;
    ram_cell[    1576] = 32'h0;  // 32'h4872ec37;
    ram_cell[    1577] = 32'h0;  // 32'h92a1f403;
    ram_cell[    1578] = 32'h0;  // 32'h0908f80c;
    ram_cell[    1579] = 32'h0;  // 32'h014943bf;
    ram_cell[    1580] = 32'h0;  // 32'hd3b0016d;
    ram_cell[    1581] = 32'h0;  // 32'hf47c05e9;
    ram_cell[    1582] = 32'h0;  // 32'hf91d06a2;
    ram_cell[    1583] = 32'h0;  // 32'h6e034171;
    ram_cell[    1584] = 32'h0;  // 32'h0dda8e3b;
    ram_cell[    1585] = 32'h0;  // 32'h752384f8;
    ram_cell[    1586] = 32'h0;  // 32'h6bb8b9b8;
    ram_cell[    1587] = 32'h0;  // 32'h233b06dc;
    ram_cell[    1588] = 32'h0;  // 32'hd9446e68;
    ram_cell[    1589] = 32'h0;  // 32'hc6dd324f;
    ram_cell[    1590] = 32'h0;  // 32'h3290f352;
    ram_cell[    1591] = 32'h0;  // 32'hd14a32bf;
    ram_cell[    1592] = 32'h0;  // 32'h121cd405;
    ram_cell[    1593] = 32'h0;  // 32'he5114021;
    ram_cell[    1594] = 32'h0;  // 32'h5a57c107;
    ram_cell[    1595] = 32'h0;  // 32'hcfefd049;
    ram_cell[    1596] = 32'h0;  // 32'h18832f6a;
    ram_cell[    1597] = 32'h0;  // 32'hab47020f;
    ram_cell[    1598] = 32'h0;  // 32'hddcbdc18;
    ram_cell[    1599] = 32'h0;  // 32'h0d8d3f9b;
    ram_cell[    1600] = 32'h0;  // 32'h021c54e4;
    ram_cell[    1601] = 32'h0;  // 32'hbeae62af;
    ram_cell[    1602] = 32'h0;  // 32'h63904b86;
    ram_cell[    1603] = 32'h0;  // 32'h09a76be3;
    ram_cell[    1604] = 32'h0;  // 32'h2d9535e5;
    ram_cell[    1605] = 32'h0;  // 32'hd3b721d6;
    ram_cell[    1606] = 32'h0;  // 32'h649ed2eb;
    ram_cell[    1607] = 32'h0;  // 32'h4dae4902;
    ram_cell[    1608] = 32'h0;  // 32'h1fd3ccfa;
    ram_cell[    1609] = 32'h0;  // 32'hb209adbd;
    ram_cell[    1610] = 32'h0;  // 32'h70fc8fd3;
    ram_cell[    1611] = 32'h0;  // 32'he2408a49;
    ram_cell[    1612] = 32'h0;  // 32'h9015bce7;
    ram_cell[    1613] = 32'h0;  // 32'ha7ac00b3;
    ram_cell[    1614] = 32'h0;  // 32'h124a3ecb;
    ram_cell[    1615] = 32'h0;  // 32'haa1f1239;
    ram_cell[    1616] = 32'h0;  // 32'h45679735;
    ram_cell[    1617] = 32'h0;  // 32'h2bb67d83;
    ram_cell[    1618] = 32'h0;  // 32'h0e1f1064;
    ram_cell[    1619] = 32'h0;  // 32'h764c1b1e;
    ram_cell[    1620] = 32'h0;  // 32'h045b9d17;
    ram_cell[    1621] = 32'h0;  // 32'h601b78e4;
    ram_cell[    1622] = 32'h0;  // 32'hf477a224;
    ram_cell[    1623] = 32'h0;  // 32'hf3b2caea;
    ram_cell[    1624] = 32'h0;  // 32'h397c8bb7;
    ram_cell[    1625] = 32'h0;  // 32'h72c346ee;
    ram_cell[    1626] = 32'h0;  // 32'h1249f91c;
    ram_cell[    1627] = 32'h0;  // 32'h2009ec7a;
    ram_cell[    1628] = 32'h0;  // 32'h07f7102a;
    ram_cell[    1629] = 32'h0;  // 32'hb325a266;
    ram_cell[    1630] = 32'h0;  // 32'h10e9f01e;
    ram_cell[    1631] = 32'h0;  // 32'h75b9348a;
    ram_cell[    1632] = 32'h0;  // 32'h0e0b032c;
    ram_cell[    1633] = 32'h0;  // 32'h978a6432;
    ram_cell[    1634] = 32'h0;  // 32'h9ed17f4e;
    ram_cell[    1635] = 32'h0;  // 32'hd7aa4568;
    ram_cell[    1636] = 32'h0;  // 32'h33162a14;
    ram_cell[    1637] = 32'h0;  // 32'h90ae0df3;
    ram_cell[    1638] = 32'h0;  // 32'h512273eb;
    ram_cell[    1639] = 32'h0;  // 32'h02b5a8ae;
    ram_cell[    1640] = 32'h0;  // 32'h303e8e1a;
    ram_cell[    1641] = 32'h0;  // 32'h200fb050;
    ram_cell[    1642] = 32'h0;  // 32'hd8f73fac;
    ram_cell[    1643] = 32'h0;  // 32'h0145a020;
    ram_cell[    1644] = 32'h0;  // 32'hf330b648;
    ram_cell[    1645] = 32'h0;  // 32'hede0f642;
    ram_cell[    1646] = 32'h0;  // 32'he06972db;
    ram_cell[    1647] = 32'h0;  // 32'h2b2c7361;
    ram_cell[    1648] = 32'h0;  // 32'h52fecf70;
    ram_cell[    1649] = 32'h0;  // 32'h36503c10;
    ram_cell[    1650] = 32'h0;  // 32'h8351d2f7;
    ram_cell[    1651] = 32'h0;  // 32'h13d1f173;
    ram_cell[    1652] = 32'h0;  // 32'hf788aa21;
    ram_cell[    1653] = 32'h0;  // 32'h7501732a;
    ram_cell[    1654] = 32'h0;  // 32'hc285ab08;
    ram_cell[    1655] = 32'h0;  // 32'hc6f427dd;
    ram_cell[    1656] = 32'h0;  // 32'h113a97ee;
    ram_cell[    1657] = 32'h0;  // 32'hb4376e7d;
    ram_cell[    1658] = 32'h0;  // 32'h92ebe47b;
    ram_cell[    1659] = 32'h0;  // 32'hea8f2f86;
    ram_cell[    1660] = 32'h0;  // 32'h6d11f8be;
    ram_cell[    1661] = 32'h0;  // 32'h00266e85;
    ram_cell[    1662] = 32'h0;  // 32'hc35541ed;
    ram_cell[    1663] = 32'h0;  // 32'h8c1da20d;
    ram_cell[    1664] = 32'h0;  // 32'h7a4812e7;
    ram_cell[    1665] = 32'h0;  // 32'hd380b9ff;
    ram_cell[    1666] = 32'h0;  // 32'h3546d0e8;
    ram_cell[    1667] = 32'h0;  // 32'hd37f03d3;
    ram_cell[    1668] = 32'h0;  // 32'hff101c93;
    ram_cell[    1669] = 32'h0;  // 32'hb8d94354;
    ram_cell[    1670] = 32'h0;  // 32'ha739c16b;
    ram_cell[    1671] = 32'h0;  // 32'hecea66d4;
    ram_cell[    1672] = 32'h0;  // 32'h5e7c8cf2;
    ram_cell[    1673] = 32'h0;  // 32'h10ef6163;
    ram_cell[    1674] = 32'h0;  // 32'h783c3d63;
    ram_cell[    1675] = 32'h0;  // 32'h4b17b847;
    ram_cell[    1676] = 32'h0;  // 32'h0550e72e;
    ram_cell[    1677] = 32'h0;  // 32'h819f27db;
    ram_cell[    1678] = 32'h0;  // 32'h31040c62;
    ram_cell[    1679] = 32'h0;  // 32'hca1777d1;
    ram_cell[    1680] = 32'h0;  // 32'hd0bf4f21;
    ram_cell[    1681] = 32'h0;  // 32'h76d210a5;
    ram_cell[    1682] = 32'h0;  // 32'h0ca776b5;
    ram_cell[    1683] = 32'h0;  // 32'h65899b60;
    ram_cell[    1684] = 32'h0;  // 32'h225f9a22;
    ram_cell[    1685] = 32'h0;  // 32'hb980530e;
    ram_cell[    1686] = 32'h0;  // 32'hff2c642a;
    ram_cell[    1687] = 32'h0;  // 32'h937c8344;
    ram_cell[    1688] = 32'h0;  // 32'hedaaba84;
    ram_cell[    1689] = 32'h0;  // 32'h613bd740;
    ram_cell[    1690] = 32'h0;  // 32'h4c6ff300;
    ram_cell[    1691] = 32'h0;  // 32'hd781dc30;
    ram_cell[    1692] = 32'h0;  // 32'hc383089f;
    ram_cell[    1693] = 32'h0;  // 32'hb1b6d540;
    ram_cell[    1694] = 32'h0;  // 32'h04d19983;
    ram_cell[    1695] = 32'h0;  // 32'h258efe5b;
    ram_cell[    1696] = 32'h0;  // 32'hf38069ee;
    ram_cell[    1697] = 32'h0;  // 32'h4204d81d;
    ram_cell[    1698] = 32'h0;  // 32'hcc0c6df1;
    ram_cell[    1699] = 32'h0;  // 32'ha1a5cb96;
    ram_cell[    1700] = 32'h0;  // 32'hf1552b6b;
    ram_cell[    1701] = 32'h0;  // 32'hf07fe542;
    ram_cell[    1702] = 32'h0;  // 32'haf1056bf;
    ram_cell[    1703] = 32'h0;  // 32'h88f322d3;
    ram_cell[    1704] = 32'h0;  // 32'hc8ca5556;
    ram_cell[    1705] = 32'h0;  // 32'hc52a79e4;
    ram_cell[    1706] = 32'h0;  // 32'h0e622438;
    ram_cell[    1707] = 32'h0;  // 32'hbb4ca33a;
    ram_cell[    1708] = 32'h0;  // 32'h50170f15;
    ram_cell[    1709] = 32'h0;  // 32'h16383375;
    ram_cell[    1710] = 32'h0;  // 32'h2a4ec55e;
    ram_cell[    1711] = 32'h0;  // 32'h27b3cf56;
    ram_cell[    1712] = 32'h0;  // 32'h3b527184;
    ram_cell[    1713] = 32'h0;  // 32'h67066d80;
    ram_cell[    1714] = 32'h0;  // 32'hb085a141;
    ram_cell[    1715] = 32'h0;  // 32'h73e196cb;
    ram_cell[    1716] = 32'h0;  // 32'ha566b6d0;
    ram_cell[    1717] = 32'h0;  // 32'he1fc7ee4;
    ram_cell[    1718] = 32'h0;  // 32'hb9b0c304;
    ram_cell[    1719] = 32'h0;  // 32'h7bae5b2d;
    ram_cell[    1720] = 32'h0;  // 32'h155bcd8d;
    ram_cell[    1721] = 32'h0;  // 32'hd9cf7b39;
    ram_cell[    1722] = 32'h0;  // 32'h3ebda0da;
    ram_cell[    1723] = 32'h0;  // 32'h2b3f3cc9;
    ram_cell[    1724] = 32'h0;  // 32'h7fb864c9;
    ram_cell[    1725] = 32'h0;  // 32'hc942d009;
    ram_cell[    1726] = 32'h0;  // 32'h9dc7f816;
    ram_cell[    1727] = 32'h0;  // 32'he0029dc8;
    ram_cell[    1728] = 32'h0;  // 32'h48c32ec0;
    ram_cell[    1729] = 32'h0;  // 32'hec9bcfc6;
    ram_cell[    1730] = 32'h0;  // 32'h185f6f68;
    ram_cell[    1731] = 32'h0;  // 32'he8dd1df7;
    ram_cell[    1732] = 32'h0;  // 32'h4b7ceb5e;
    ram_cell[    1733] = 32'h0;  // 32'h3b1f5127;
    ram_cell[    1734] = 32'h0;  // 32'h176eaa4f;
    ram_cell[    1735] = 32'h0;  // 32'hfa7157a4;
    ram_cell[    1736] = 32'h0;  // 32'h22eccd58;
    ram_cell[    1737] = 32'h0;  // 32'hfc7adea3;
    ram_cell[    1738] = 32'h0;  // 32'h6de9c70c;
    ram_cell[    1739] = 32'h0;  // 32'h4a99836b;
    ram_cell[    1740] = 32'h0;  // 32'h9328f76d;
    ram_cell[    1741] = 32'h0;  // 32'h718f5b19;
    ram_cell[    1742] = 32'h0;  // 32'h1846435c;
    ram_cell[    1743] = 32'h0;  // 32'h54e17c36;
    ram_cell[    1744] = 32'h0;  // 32'h236e2ecd;
    ram_cell[    1745] = 32'h0;  // 32'he61b7821;
    ram_cell[    1746] = 32'h0;  // 32'h57721bc9;
    ram_cell[    1747] = 32'h0;  // 32'h490ef471;
    ram_cell[    1748] = 32'h0;  // 32'hf979a296;
    ram_cell[    1749] = 32'h0;  // 32'hacdca1bc;
    ram_cell[    1750] = 32'h0;  // 32'hc678ee1b;
    ram_cell[    1751] = 32'h0;  // 32'h1efd40b8;
    ram_cell[    1752] = 32'h0;  // 32'h492fcf9a;
    ram_cell[    1753] = 32'h0;  // 32'h025fa7ca;
    ram_cell[    1754] = 32'h0;  // 32'h19f459be;
    ram_cell[    1755] = 32'h0;  // 32'h5885d949;
    ram_cell[    1756] = 32'h0;  // 32'h50c9a31d;
    ram_cell[    1757] = 32'h0;  // 32'haa306289;
    ram_cell[    1758] = 32'h0;  // 32'h2a6ab2f2;
    ram_cell[    1759] = 32'h0;  // 32'h0ed6464f;
    ram_cell[    1760] = 32'h0;  // 32'hbd5564b9;
    ram_cell[    1761] = 32'h0;  // 32'hc3d1922b;
    ram_cell[    1762] = 32'h0;  // 32'h92997f24;
    ram_cell[    1763] = 32'h0;  // 32'h5df56800;
    ram_cell[    1764] = 32'h0;  // 32'h1d528655;
    ram_cell[    1765] = 32'h0;  // 32'h8c101f4a;
    ram_cell[    1766] = 32'h0;  // 32'h3fe287b5;
    ram_cell[    1767] = 32'h0;  // 32'hf01af8e8;
    ram_cell[    1768] = 32'h0;  // 32'hbe238f13;
    ram_cell[    1769] = 32'h0;  // 32'h07110b61;
    ram_cell[    1770] = 32'h0;  // 32'hc8472a2f;
    ram_cell[    1771] = 32'h0;  // 32'h249fc1dd;
    ram_cell[    1772] = 32'h0;  // 32'h4ede798c;
    ram_cell[    1773] = 32'h0;  // 32'hb22498da;
    ram_cell[    1774] = 32'h0;  // 32'h7f8b4826;
    ram_cell[    1775] = 32'h0;  // 32'h4b1bd2f2;
    ram_cell[    1776] = 32'h0;  // 32'had65c307;
    ram_cell[    1777] = 32'h0;  // 32'h1d2b089f;
    ram_cell[    1778] = 32'h0;  // 32'h392a428f;
    ram_cell[    1779] = 32'h0;  // 32'hcd27ce60;
    ram_cell[    1780] = 32'h0;  // 32'h32e0d1e6;
    ram_cell[    1781] = 32'h0;  // 32'hcd8132ec;
    ram_cell[    1782] = 32'h0;  // 32'ha25636a7;
    ram_cell[    1783] = 32'h0;  // 32'h2bd933e8;
    ram_cell[    1784] = 32'h0;  // 32'h67ea8d02;
    ram_cell[    1785] = 32'h0;  // 32'h42e320e9;
    ram_cell[    1786] = 32'h0;  // 32'hf2c05b14;
    ram_cell[    1787] = 32'h0;  // 32'hb4e70143;
    ram_cell[    1788] = 32'h0;  // 32'h3bba385e;
    ram_cell[    1789] = 32'h0;  // 32'hf2264373;
    ram_cell[    1790] = 32'h0;  // 32'hab24cc97;
    ram_cell[    1791] = 32'h0;  // 32'h741d9fc0;
    ram_cell[    1792] = 32'h0;  // 32'h7f0909b8;
    ram_cell[    1793] = 32'h0;  // 32'ha211243f;
    ram_cell[    1794] = 32'h0;  // 32'h1468aea5;
    ram_cell[    1795] = 32'h0;  // 32'h884cae4a;
    ram_cell[    1796] = 32'h0;  // 32'he9b11cc3;
    ram_cell[    1797] = 32'h0;  // 32'ha8e9abfa;
    ram_cell[    1798] = 32'h0;  // 32'ha9420eb2;
    ram_cell[    1799] = 32'h0;  // 32'hba497f9a;
    ram_cell[    1800] = 32'h0;  // 32'h25c02c96;
    ram_cell[    1801] = 32'h0;  // 32'h8dd22c16;
    ram_cell[    1802] = 32'h0;  // 32'h089021ee;
    ram_cell[    1803] = 32'h0;  // 32'hc774a7f5;
    ram_cell[    1804] = 32'h0;  // 32'h745217f8;
    ram_cell[    1805] = 32'h0;  // 32'he64e85d0;
    ram_cell[    1806] = 32'h0;  // 32'h10b1541b;
    ram_cell[    1807] = 32'h0;  // 32'h5858c420;
    ram_cell[    1808] = 32'h0;  // 32'h6761abd6;
    ram_cell[    1809] = 32'h0;  // 32'h4922ff28;
    ram_cell[    1810] = 32'h0;  // 32'h35769226;
    ram_cell[    1811] = 32'h0;  // 32'ha2d37b63;
    ram_cell[    1812] = 32'h0;  // 32'h84b1d9cb;
    ram_cell[    1813] = 32'h0;  // 32'h1f4614ac;
    ram_cell[    1814] = 32'h0;  // 32'h137c13d6;
    ram_cell[    1815] = 32'h0;  // 32'h37a4774b;
    ram_cell[    1816] = 32'h0;  // 32'hd71b1dfa;
    ram_cell[    1817] = 32'h0;  // 32'hebed5bdd;
    ram_cell[    1818] = 32'h0;  // 32'h6546e941;
    ram_cell[    1819] = 32'h0;  // 32'hd203be47;
    ram_cell[    1820] = 32'h0;  // 32'h98ab8d3b;
    ram_cell[    1821] = 32'h0;  // 32'h71f7e658;
    ram_cell[    1822] = 32'h0;  // 32'hcd8c6790;
    ram_cell[    1823] = 32'h0;  // 32'h7e82b37f;
    ram_cell[    1824] = 32'h0;  // 32'h0e53cae9;
    ram_cell[    1825] = 32'h0;  // 32'hb3f5eac1;
    ram_cell[    1826] = 32'h0;  // 32'he3e9f919;
    ram_cell[    1827] = 32'h0;  // 32'h98c99010;
    ram_cell[    1828] = 32'h0;  // 32'ha5792402;
    ram_cell[    1829] = 32'h0;  // 32'hd0f796ee;
    ram_cell[    1830] = 32'h0;  // 32'h4f13fac7;
    ram_cell[    1831] = 32'h0;  // 32'h98577ada;
    ram_cell[    1832] = 32'h0;  // 32'hbe211bb1;
    ram_cell[    1833] = 32'h0;  // 32'hbaba267a;
    ram_cell[    1834] = 32'h0;  // 32'h5519f856;
    ram_cell[    1835] = 32'h0;  // 32'hbf2f4216;
    ram_cell[    1836] = 32'h0;  // 32'he66b3fe5;
    ram_cell[    1837] = 32'h0;  // 32'h664cf4f2;
    ram_cell[    1838] = 32'h0;  // 32'h3c512c8f;
    ram_cell[    1839] = 32'h0;  // 32'h3eeea20c;
    ram_cell[    1840] = 32'h0;  // 32'h58c522de;
    ram_cell[    1841] = 32'h0;  // 32'h0be40245;
    ram_cell[    1842] = 32'h0;  // 32'h06507d66;
    ram_cell[    1843] = 32'h0;  // 32'h4f65026c;
    ram_cell[    1844] = 32'h0;  // 32'h46ffb08f;
    ram_cell[    1845] = 32'h0;  // 32'hc849f6e2;
    ram_cell[    1846] = 32'h0;  // 32'h2de71c53;
    ram_cell[    1847] = 32'h0;  // 32'h31c724b1;
    ram_cell[    1848] = 32'h0;  // 32'hdd0f0978;
    ram_cell[    1849] = 32'h0;  // 32'heffbf2f0;
    ram_cell[    1850] = 32'h0;  // 32'h4b1183a2;
    ram_cell[    1851] = 32'h0;  // 32'hd9d31cd9;
    ram_cell[    1852] = 32'h0;  // 32'hcce44acb;
    ram_cell[    1853] = 32'h0;  // 32'hc874a365;
    ram_cell[    1854] = 32'h0;  // 32'h4a1831c0;
    ram_cell[    1855] = 32'h0;  // 32'hd6ac3602;
    ram_cell[    1856] = 32'h0;  // 32'hcbe62a57;
    ram_cell[    1857] = 32'h0;  // 32'h64424906;
    ram_cell[    1858] = 32'h0;  // 32'h6688c37d;
    ram_cell[    1859] = 32'h0;  // 32'he5d8f33d;
    ram_cell[    1860] = 32'h0;  // 32'h336d0cf3;
    ram_cell[    1861] = 32'h0;  // 32'h8c87467d;
    ram_cell[    1862] = 32'h0;  // 32'he946c5f9;
    ram_cell[    1863] = 32'h0;  // 32'h5832262b;
    ram_cell[    1864] = 32'h0;  // 32'hc5e9baeb;
    ram_cell[    1865] = 32'h0;  // 32'h8572e706;
    ram_cell[    1866] = 32'h0;  // 32'h11947939;
    ram_cell[    1867] = 32'h0;  // 32'h4895f943;
    ram_cell[    1868] = 32'h0;  // 32'h3e369717;
    ram_cell[    1869] = 32'h0;  // 32'hdaad85df;
    ram_cell[    1870] = 32'h0;  // 32'h98cfa5ce;
    ram_cell[    1871] = 32'h0;  // 32'ha6a39df4;
    ram_cell[    1872] = 32'h0;  // 32'h7b75a90b;
    ram_cell[    1873] = 32'h0;  // 32'hb88e6551;
    ram_cell[    1874] = 32'h0;  // 32'h6bfe72f1;
    ram_cell[    1875] = 32'h0;  // 32'hf3db1d0a;
    ram_cell[    1876] = 32'h0;  // 32'h599bf03a;
    ram_cell[    1877] = 32'h0;  // 32'h642c06c7;
    ram_cell[    1878] = 32'h0;  // 32'h6e6d98a0;
    ram_cell[    1879] = 32'h0;  // 32'h2a170f48;
    ram_cell[    1880] = 32'h0;  // 32'hce51546b;
    ram_cell[    1881] = 32'h0;  // 32'h5fbc0ebc;
    ram_cell[    1882] = 32'h0;  // 32'h09220069;
    ram_cell[    1883] = 32'h0;  // 32'h423a3362;
    ram_cell[    1884] = 32'h0;  // 32'h8c231cfb;
    ram_cell[    1885] = 32'h0;  // 32'h1e46b0cb;
    ram_cell[    1886] = 32'h0;  // 32'h1af6940b;
    ram_cell[    1887] = 32'h0;  // 32'h0806c74c;
    ram_cell[    1888] = 32'h0;  // 32'h439534c9;
    ram_cell[    1889] = 32'h0;  // 32'h1dac20e2;
    ram_cell[    1890] = 32'h0;  // 32'hdffb417e;
    ram_cell[    1891] = 32'h0;  // 32'h867bcad6;
    ram_cell[    1892] = 32'h0;  // 32'hc7c76716;
    ram_cell[    1893] = 32'h0;  // 32'h62e63c70;
    ram_cell[    1894] = 32'h0;  // 32'h95a75cfa;
    ram_cell[    1895] = 32'h0;  // 32'h13c2e46a;
    ram_cell[    1896] = 32'h0;  // 32'hcfd9f23e;
    ram_cell[    1897] = 32'h0;  // 32'he81589ac;
    ram_cell[    1898] = 32'h0;  // 32'h5d532aad;
    ram_cell[    1899] = 32'h0;  // 32'h00064e82;
    ram_cell[    1900] = 32'h0;  // 32'h53857f2b;
    ram_cell[    1901] = 32'h0;  // 32'he1542c66;
    ram_cell[    1902] = 32'h0;  // 32'h94738397;
    ram_cell[    1903] = 32'h0;  // 32'hb4fe595f;
    ram_cell[    1904] = 32'h0;  // 32'h7cdbe74f;
    ram_cell[    1905] = 32'h0;  // 32'hcbfc90d4;
    ram_cell[    1906] = 32'h0;  // 32'h5917af0b;
    ram_cell[    1907] = 32'h0;  // 32'hd30bb7bc;
    ram_cell[    1908] = 32'h0;  // 32'h137c008a;
    ram_cell[    1909] = 32'h0;  // 32'h363fa4e3;
    ram_cell[    1910] = 32'h0;  // 32'hd50598ea;
    ram_cell[    1911] = 32'h0;  // 32'h3f13a66b;
    ram_cell[    1912] = 32'h0;  // 32'h2721699a;
    ram_cell[    1913] = 32'h0;  // 32'h200348ef;
    ram_cell[    1914] = 32'h0;  // 32'h5f25c637;
    ram_cell[    1915] = 32'h0;  // 32'h95b50873;
    ram_cell[    1916] = 32'h0;  // 32'hdf04bd73;
    ram_cell[    1917] = 32'h0;  // 32'hfecaf201;
    ram_cell[    1918] = 32'h0;  // 32'haa6b3e4a;
    ram_cell[    1919] = 32'h0;  // 32'hfefd3770;
    ram_cell[    1920] = 32'h0;  // 32'h3e290aae;
    ram_cell[    1921] = 32'h0;  // 32'hd86c2b96;
    ram_cell[    1922] = 32'h0;  // 32'hfb1682b7;
    ram_cell[    1923] = 32'h0;  // 32'he6b72d06;
    ram_cell[    1924] = 32'h0;  // 32'hd6510938;
    ram_cell[    1925] = 32'h0;  // 32'h6cddb4bd;
    ram_cell[    1926] = 32'h0;  // 32'h329ba8e9;
    ram_cell[    1927] = 32'h0;  // 32'hcc5e171b;
    ram_cell[    1928] = 32'h0;  // 32'h73bcbde9;
    ram_cell[    1929] = 32'h0;  // 32'h5e8ebe72;
    ram_cell[    1930] = 32'h0;  // 32'h6e21c766;
    ram_cell[    1931] = 32'h0;  // 32'hbed98f14;
    ram_cell[    1932] = 32'h0;  // 32'h1b43da18;
    ram_cell[    1933] = 32'h0;  // 32'h913e5a9e;
    ram_cell[    1934] = 32'h0;  // 32'haebf3b17;
    ram_cell[    1935] = 32'h0;  // 32'h44e2132a;
    ram_cell[    1936] = 32'h0;  // 32'hb7ec4f63;
    ram_cell[    1937] = 32'h0;  // 32'h66e3e57a;
    ram_cell[    1938] = 32'h0;  // 32'ha65eef18;
    ram_cell[    1939] = 32'h0;  // 32'hd079d162;
    ram_cell[    1940] = 32'h0;  // 32'h0e87f0f6;
    ram_cell[    1941] = 32'h0;  // 32'h8332797b;
    ram_cell[    1942] = 32'h0;  // 32'h9b0195d8;
    ram_cell[    1943] = 32'h0;  // 32'h355a217b;
    ram_cell[    1944] = 32'h0;  // 32'hbf37203c;
    ram_cell[    1945] = 32'h0;  // 32'h29baf4c6;
    ram_cell[    1946] = 32'h0;  // 32'h47f5a838;
    ram_cell[    1947] = 32'h0;  // 32'h07bc23c3;
    ram_cell[    1948] = 32'h0;  // 32'hab01668e;
    ram_cell[    1949] = 32'h0;  // 32'h12776355;
    ram_cell[    1950] = 32'h0;  // 32'ha40d4c48;
    ram_cell[    1951] = 32'h0;  // 32'h91a74f9d;
    ram_cell[    1952] = 32'h0;  // 32'h0d23c055;
    ram_cell[    1953] = 32'h0;  // 32'haccf6a52;
    ram_cell[    1954] = 32'h0;  // 32'h8536b534;
    ram_cell[    1955] = 32'h0;  // 32'h52cfef58;
    ram_cell[    1956] = 32'h0;  // 32'h7fd558ab;
    ram_cell[    1957] = 32'h0;  // 32'h6376b04c;
    ram_cell[    1958] = 32'h0;  // 32'h2866ff0f;
    ram_cell[    1959] = 32'h0;  // 32'h12647867;
    ram_cell[    1960] = 32'h0;  // 32'h02425e58;
    ram_cell[    1961] = 32'h0;  // 32'hcaa5e97e;
    ram_cell[    1962] = 32'h0;  // 32'he3b2c95f;
    ram_cell[    1963] = 32'h0;  // 32'h2ccbc03f;
    ram_cell[    1964] = 32'h0;  // 32'he607988c;
    ram_cell[    1965] = 32'h0;  // 32'h13e3dc01;
    ram_cell[    1966] = 32'h0;  // 32'ha85d2546;
    ram_cell[    1967] = 32'h0;  // 32'hbe62e88a;
    ram_cell[    1968] = 32'h0;  // 32'h19ad265d;
    ram_cell[    1969] = 32'h0;  // 32'h74baaede;
    ram_cell[    1970] = 32'h0;  // 32'hedcf8061;
    ram_cell[    1971] = 32'h0;  // 32'h535e1f18;
    ram_cell[    1972] = 32'h0;  // 32'h1688deb8;
    ram_cell[    1973] = 32'h0;  // 32'h83477bf6;
    ram_cell[    1974] = 32'h0;  // 32'h0d72700c;
    ram_cell[    1975] = 32'h0;  // 32'h7d3f323e;
    ram_cell[    1976] = 32'h0;  // 32'h4638fd7f;
    ram_cell[    1977] = 32'h0;  // 32'hf7376ae3;
    ram_cell[    1978] = 32'h0;  // 32'h1b76b9e8;
    ram_cell[    1979] = 32'h0;  // 32'h38a65fee;
    ram_cell[    1980] = 32'h0;  // 32'h2eb0cd7a;
    ram_cell[    1981] = 32'h0;  // 32'h11d196dc;
    ram_cell[    1982] = 32'h0;  // 32'h24ce8ce9;
    ram_cell[    1983] = 32'h0;  // 32'hfff01af7;
    ram_cell[    1984] = 32'h0;  // 32'he6f7abc4;
    ram_cell[    1985] = 32'h0;  // 32'h7e867cf1;
    ram_cell[    1986] = 32'h0;  // 32'hd2091cd7;
    ram_cell[    1987] = 32'h0;  // 32'ha663cc61;
    ram_cell[    1988] = 32'h0;  // 32'hcddaaf6b;
    ram_cell[    1989] = 32'h0;  // 32'hdf206dab;
    ram_cell[    1990] = 32'h0;  // 32'h3c4f8420;
    ram_cell[    1991] = 32'h0;  // 32'h814d5085;
    ram_cell[    1992] = 32'h0;  // 32'h6d9e1c49;
    ram_cell[    1993] = 32'h0;  // 32'h6911eec5;
    ram_cell[    1994] = 32'h0;  // 32'h0f6c8c18;
    ram_cell[    1995] = 32'h0;  // 32'h3cb4076d;
    ram_cell[    1996] = 32'h0;  // 32'h53c55fe9;
    ram_cell[    1997] = 32'h0;  // 32'hb6a363e9;
    ram_cell[    1998] = 32'h0;  // 32'hfd3382c4;
    ram_cell[    1999] = 32'h0;  // 32'hc25fb5a5;
    ram_cell[    2000] = 32'h0;  // 32'h97dab281;
    ram_cell[    2001] = 32'h0;  // 32'h2a9e46b3;
    ram_cell[    2002] = 32'h0;  // 32'hf39f1ff4;
    ram_cell[    2003] = 32'h0;  // 32'hb7ddbca8;
    ram_cell[    2004] = 32'h0;  // 32'h0bc647ec;
    ram_cell[    2005] = 32'h0;  // 32'h8126e089;
    ram_cell[    2006] = 32'h0;  // 32'h369ce354;
    ram_cell[    2007] = 32'h0;  // 32'h794717d4;
    ram_cell[    2008] = 32'h0;  // 32'h7862338b;
    ram_cell[    2009] = 32'h0;  // 32'hedb2f942;
    ram_cell[    2010] = 32'h0;  // 32'h298e4cec;
    ram_cell[    2011] = 32'h0;  // 32'ha44eda57;
    ram_cell[    2012] = 32'h0;  // 32'h20c34ed2;
    ram_cell[    2013] = 32'h0;  // 32'hf9894f8f;
    ram_cell[    2014] = 32'h0;  // 32'he7895c09;
    ram_cell[    2015] = 32'h0;  // 32'habe80650;
    ram_cell[    2016] = 32'h0;  // 32'h3326dcaa;
    ram_cell[    2017] = 32'h0;  // 32'h2beb906c;
    ram_cell[    2018] = 32'h0;  // 32'hd153023b;
    ram_cell[    2019] = 32'h0;  // 32'hc324716f;
    ram_cell[    2020] = 32'h0;  // 32'h17b14f44;
    ram_cell[    2021] = 32'h0;  // 32'hfe60ce1f;
    ram_cell[    2022] = 32'h0;  // 32'hbba11821;
    ram_cell[    2023] = 32'h0;  // 32'h481ecd4a;
    ram_cell[    2024] = 32'h0;  // 32'h4846187f;
    ram_cell[    2025] = 32'h0;  // 32'h4a426419;
    ram_cell[    2026] = 32'h0;  // 32'h94dbaa02;
    ram_cell[    2027] = 32'h0;  // 32'hf9d86ac4;
    ram_cell[    2028] = 32'h0;  // 32'h95ff61c6;
    ram_cell[    2029] = 32'h0;  // 32'h6d2b66a2;
    ram_cell[    2030] = 32'h0;  // 32'hd3903d66;
    ram_cell[    2031] = 32'h0;  // 32'hbe34e61e;
    ram_cell[    2032] = 32'h0;  // 32'hebbdcafc;
    ram_cell[    2033] = 32'h0;  // 32'hd708f8fe;
    ram_cell[    2034] = 32'h0;  // 32'hc71f4455;
    ram_cell[    2035] = 32'h0;  // 32'h066ccd61;
    ram_cell[    2036] = 32'h0;  // 32'hfb0d910c;
    ram_cell[    2037] = 32'h0;  // 32'h87fec5c9;
    ram_cell[    2038] = 32'h0;  // 32'h38ac549c;
    ram_cell[    2039] = 32'h0;  // 32'hb83a687d;
    ram_cell[    2040] = 32'h0;  // 32'hc358b8fe;
    ram_cell[    2041] = 32'h0;  // 32'h87ab2e2b;
    ram_cell[    2042] = 32'h0;  // 32'hc55cf8fe;
    ram_cell[    2043] = 32'h0;  // 32'ha40d8a13;
    ram_cell[    2044] = 32'h0;  // 32'h1bdc71c1;
    ram_cell[    2045] = 32'h0;  // 32'h8bbb4738;
    ram_cell[    2046] = 32'h0;  // 32'h8153655c;
    ram_cell[    2047] = 32'h0;  // 32'hce5f2f9b;
    ram_cell[    2048] = 32'h0;  // 32'hcec20111;
    ram_cell[    2049] = 32'h0;  // 32'h04266818;
    ram_cell[    2050] = 32'h0;  // 32'hdb5f698b;
    ram_cell[    2051] = 32'h0;  // 32'hbb4d4ee8;
    ram_cell[    2052] = 32'h0;  // 32'h2a9b801c;
    ram_cell[    2053] = 32'h0;  // 32'hfa4cc8ae;
    ram_cell[    2054] = 32'h0;  // 32'h2f02668f;
    ram_cell[    2055] = 32'h0;  // 32'ha53f290e;
    ram_cell[    2056] = 32'h0;  // 32'hb1c1dd95;
    ram_cell[    2057] = 32'h0;  // 32'hd1f4976b;
    ram_cell[    2058] = 32'h0;  // 32'h4906f68c;
    ram_cell[    2059] = 32'h0;  // 32'he9f76556;
    ram_cell[    2060] = 32'h0;  // 32'h6e302f02;
    ram_cell[    2061] = 32'h0;  // 32'hab36e998;
    ram_cell[    2062] = 32'h0;  // 32'h2e3b9322;
    ram_cell[    2063] = 32'h0;  // 32'h801e1513;
    ram_cell[    2064] = 32'h0;  // 32'ha9d18e10;
    ram_cell[    2065] = 32'h0;  // 32'hbd6c34e3;
    ram_cell[    2066] = 32'h0;  // 32'h5d3e252d;
    ram_cell[    2067] = 32'h0;  // 32'h555a5d53;
    ram_cell[    2068] = 32'h0;  // 32'ha8707801;
    ram_cell[    2069] = 32'h0;  // 32'h14f704c2;
    ram_cell[    2070] = 32'h0;  // 32'hc4cf50ad;
    ram_cell[    2071] = 32'h0;  // 32'hcc2ad2f7;
    ram_cell[    2072] = 32'h0;  // 32'hdd857ffb;
    ram_cell[    2073] = 32'h0;  // 32'h83d186e7;
    ram_cell[    2074] = 32'h0;  // 32'h3834422d;
    ram_cell[    2075] = 32'h0;  // 32'h3f275501;
    ram_cell[    2076] = 32'h0;  // 32'haa1623d6;
    ram_cell[    2077] = 32'h0;  // 32'h658665dc;
    ram_cell[    2078] = 32'h0;  // 32'hebebf848;
    ram_cell[    2079] = 32'h0;  // 32'h4b803f04;
    ram_cell[    2080] = 32'h0;  // 32'h1eb2f7d2;
    ram_cell[    2081] = 32'h0;  // 32'h3c10fab6;
    ram_cell[    2082] = 32'h0;  // 32'h99ffc986;
    ram_cell[    2083] = 32'h0;  // 32'hf9e64a01;
    ram_cell[    2084] = 32'h0;  // 32'hc8162054;
    ram_cell[    2085] = 32'h0;  // 32'h3d1e0961;
    ram_cell[    2086] = 32'h0;  // 32'ha0b1816c;
    ram_cell[    2087] = 32'h0;  // 32'h474545d0;
    ram_cell[    2088] = 32'h0;  // 32'hf5feae52;
    ram_cell[    2089] = 32'h0;  // 32'h51bd67c0;
    ram_cell[    2090] = 32'h0;  // 32'he8273063;
    ram_cell[    2091] = 32'h0;  // 32'h0c86c6e5;
    ram_cell[    2092] = 32'h0;  // 32'hd592fac6;
    ram_cell[    2093] = 32'h0;  // 32'h6b818fad;
    ram_cell[    2094] = 32'h0;  // 32'h38af2a5b;
    ram_cell[    2095] = 32'h0;  // 32'hbf05934c;
    ram_cell[    2096] = 32'h0;  // 32'ha821d2fe;
    ram_cell[    2097] = 32'h0;  // 32'h35e5f0ff;
    ram_cell[    2098] = 32'h0;  // 32'h51124c0c;
    ram_cell[    2099] = 32'h0;  // 32'h54e1f1e3;
    ram_cell[    2100] = 32'h0;  // 32'h99cce913;
    ram_cell[    2101] = 32'h0;  // 32'h275c58d8;
    ram_cell[    2102] = 32'h0;  // 32'h0d046142;
    ram_cell[    2103] = 32'h0;  // 32'hc45d5cb3;
    ram_cell[    2104] = 32'h0;  // 32'hd887a412;
    ram_cell[    2105] = 32'h0;  // 32'h8dfe5493;
    ram_cell[    2106] = 32'h0;  // 32'hac0a43b0;
    ram_cell[    2107] = 32'h0;  // 32'hbd65833d;
    ram_cell[    2108] = 32'h0;  // 32'hb7ad89b6;
    ram_cell[    2109] = 32'h0;  // 32'hca75b704;
    ram_cell[    2110] = 32'h0;  // 32'h8d31e95a;
    ram_cell[    2111] = 32'h0;  // 32'hbbdcc4dc;
    ram_cell[    2112] = 32'h0;  // 32'h3b543cf1;
    ram_cell[    2113] = 32'h0;  // 32'h4d29cda5;
    ram_cell[    2114] = 32'h0;  // 32'h99bfbee2;
    ram_cell[    2115] = 32'h0;  // 32'h1790d722;
    ram_cell[    2116] = 32'h0;  // 32'h8d9fa281;
    ram_cell[    2117] = 32'h0;  // 32'hb4b8c67a;
    ram_cell[    2118] = 32'h0;  // 32'h6b1d708e;
    ram_cell[    2119] = 32'h0;  // 32'h1c4ad7a3;
    ram_cell[    2120] = 32'h0;  // 32'h2138a6b2;
    ram_cell[    2121] = 32'h0;  // 32'hdc8687f1;
    ram_cell[    2122] = 32'h0;  // 32'h3e7cc7a0;
    ram_cell[    2123] = 32'h0;  // 32'hf10ff173;
    ram_cell[    2124] = 32'h0;  // 32'h70356980;
    ram_cell[    2125] = 32'h0;  // 32'he4ae9030;
    ram_cell[    2126] = 32'h0;  // 32'h03521858;
    ram_cell[    2127] = 32'h0;  // 32'h8e9296b5;
    ram_cell[    2128] = 32'h0;  // 32'hfb65b727;
    ram_cell[    2129] = 32'h0;  // 32'h3f3a6214;
    ram_cell[    2130] = 32'h0;  // 32'h690101da;
    ram_cell[    2131] = 32'h0;  // 32'h3c04d86e;
    ram_cell[    2132] = 32'h0;  // 32'h7a66d869;
    ram_cell[    2133] = 32'h0;  // 32'h229d7a5d;
    ram_cell[    2134] = 32'h0;  // 32'h0df4ad36;
    ram_cell[    2135] = 32'h0;  // 32'heb5845f7;
    ram_cell[    2136] = 32'h0;  // 32'hfeadd3c4;
    ram_cell[    2137] = 32'h0;  // 32'hdbbc9783;
    ram_cell[    2138] = 32'h0;  // 32'h262c7922;
    ram_cell[    2139] = 32'h0;  // 32'hd19bd722;
    ram_cell[    2140] = 32'h0;  // 32'h8b30f67f;
    ram_cell[    2141] = 32'h0;  // 32'hdb9fbe01;
    ram_cell[    2142] = 32'h0;  // 32'hc9ac5bc8;
    ram_cell[    2143] = 32'h0;  // 32'hfe353587;
    ram_cell[    2144] = 32'h0;  // 32'h01b2c58c;
    ram_cell[    2145] = 32'h0;  // 32'h54516ef9;
    ram_cell[    2146] = 32'h0;  // 32'haf88e2dd;
    ram_cell[    2147] = 32'h0;  // 32'h91716fc6;
    ram_cell[    2148] = 32'h0;  // 32'h573a478c;
    ram_cell[    2149] = 32'h0;  // 32'h63ba4a5f;
    ram_cell[    2150] = 32'h0;  // 32'h2ab1cdb7;
    ram_cell[    2151] = 32'h0;  // 32'h5b81486f;
    ram_cell[    2152] = 32'h0;  // 32'h0cbe74d6;
    ram_cell[    2153] = 32'h0;  // 32'h84c5a001;
    ram_cell[    2154] = 32'h0;  // 32'hb3381b8f;
    ram_cell[    2155] = 32'h0;  // 32'h9500a2e6;
    ram_cell[    2156] = 32'h0;  // 32'hea864b45;
    ram_cell[    2157] = 32'h0;  // 32'hff0941c0;
    ram_cell[    2158] = 32'h0;  // 32'h73913639;
    ram_cell[    2159] = 32'h0;  // 32'h166c4391;
    ram_cell[    2160] = 32'h0;  // 32'hf43f7bee;
    ram_cell[    2161] = 32'h0;  // 32'he820c8b8;
    ram_cell[    2162] = 32'h0;  // 32'hee411c88;
    ram_cell[    2163] = 32'h0;  // 32'h8e859f88;
    ram_cell[    2164] = 32'h0;  // 32'h9a7b4dbd;
    ram_cell[    2165] = 32'h0;  // 32'h36499cb8;
    ram_cell[    2166] = 32'h0;  // 32'ha193e8fe;
    ram_cell[    2167] = 32'h0;  // 32'he762fb8b;
    ram_cell[    2168] = 32'h0;  // 32'h07776df1;
    ram_cell[    2169] = 32'h0;  // 32'h09385f94;
    ram_cell[    2170] = 32'h0;  // 32'hdab80b24;
    ram_cell[    2171] = 32'h0;  // 32'ha827d699;
    ram_cell[    2172] = 32'h0;  // 32'h1e7836af;
    ram_cell[    2173] = 32'h0;  // 32'h792f7869;
    ram_cell[    2174] = 32'h0;  // 32'h4dc72a6e;
    ram_cell[    2175] = 32'h0;  // 32'h025491b6;
    ram_cell[    2176] = 32'h0;  // 32'he1ec1b7f;
    ram_cell[    2177] = 32'h0;  // 32'h467b63f6;
    ram_cell[    2178] = 32'h0;  // 32'hd2be0419;
    ram_cell[    2179] = 32'h0;  // 32'hcc4b241c;
    ram_cell[    2180] = 32'h0;  // 32'hd647b6f1;
    ram_cell[    2181] = 32'h0;  // 32'h3c6188e0;
    ram_cell[    2182] = 32'h0;  // 32'h5db14f0a;
    ram_cell[    2183] = 32'h0;  // 32'h737f2989;
    ram_cell[    2184] = 32'h0;  // 32'h7a0191b9;
    ram_cell[    2185] = 32'h0;  // 32'h2aeedf62;
    ram_cell[    2186] = 32'h0;  // 32'h6fa2a74f;
    ram_cell[    2187] = 32'h0;  // 32'h04e4ec92;
    ram_cell[    2188] = 32'h0;  // 32'h56d14df6;
    ram_cell[    2189] = 32'h0;  // 32'h0320f647;
    ram_cell[    2190] = 32'h0;  // 32'h1bd5e99f;
    ram_cell[    2191] = 32'h0;  // 32'h0d067f39;
    ram_cell[    2192] = 32'h0;  // 32'h5a9f1f52;
    ram_cell[    2193] = 32'h0;  // 32'haebc0032;
    ram_cell[    2194] = 32'h0;  // 32'h1d95f310;
    ram_cell[    2195] = 32'h0;  // 32'h9e851144;
    ram_cell[    2196] = 32'h0;  // 32'he057bdf0;
    ram_cell[    2197] = 32'h0;  // 32'hf41c5e35;
    ram_cell[    2198] = 32'h0;  // 32'ha2fb2bf8;
    ram_cell[    2199] = 32'h0;  // 32'h5364bee8;
    ram_cell[    2200] = 32'h0;  // 32'h1c7e2f21;
    ram_cell[    2201] = 32'h0;  // 32'ha7568c27;
    ram_cell[    2202] = 32'h0;  // 32'h624369ce;
    ram_cell[    2203] = 32'h0;  // 32'hb9a451eb;
    ram_cell[    2204] = 32'h0;  // 32'h0d3e4b37;
    ram_cell[    2205] = 32'h0;  // 32'h13ea486a;
    ram_cell[    2206] = 32'h0;  // 32'h48ebaca1;
    ram_cell[    2207] = 32'h0;  // 32'ha87269e3;
    ram_cell[    2208] = 32'h0;  // 32'h04143ae9;
    ram_cell[    2209] = 32'h0;  // 32'heaae30ae;
    ram_cell[    2210] = 32'h0;  // 32'hdfe74508;
    ram_cell[    2211] = 32'h0;  // 32'haea97383;
    ram_cell[    2212] = 32'h0;  // 32'h97b710c9;
    ram_cell[    2213] = 32'h0;  // 32'h01f53d28;
    ram_cell[    2214] = 32'h0;  // 32'h6911eab1;
    ram_cell[    2215] = 32'h0;  // 32'h7fea1a76;
    ram_cell[    2216] = 32'h0;  // 32'h1f44b824;
    ram_cell[    2217] = 32'h0;  // 32'hccc03093;
    ram_cell[    2218] = 32'h0;  // 32'hf9f593b0;
    ram_cell[    2219] = 32'h0;  // 32'h39e4fc4b;
    ram_cell[    2220] = 32'h0;  // 32'h85293fd5;
    ram_cell[    2221] = 32'h0;  // 32'h57195540;
    ram_cell[    2222] = 32'h0;  // 32'h8316ede8;
    ram_cell[    2223] = 32'h0;  // 32'h24cd482f;
    ram_cell[    2224] = 32'h0;  // 32'h563ce767;
    ram_cell[    2225] = 32'h0;  // 32'h6096f1f5;
    ram_cell[    2226] = 32'h0;  // 32'hed340134;
    ram_cell[    2227] = 32'h0;  // 32'h5632ef34;
    ram_cell[    2228] = 32'h0;  // 32'h4477cbf0;
    ram_cell[    2229] = 32'h0;  // 32'hc79e10e9;
    ram_cell[    2230] = 32'h0;  // 32'h7f81ade6;
    ram_cell[    2231] = 32'h0;  // 32'h836cba04;
    ram_cell[    2232] = 32'h0;  // 32'h3831b6a0;
    ram_cell[    2233] = 32'h0;  // 32'hbc99fdd9;
    ram_cell[    2234] = 32'h0;  // 32'hb3a7c693;
    ram_cell[    2235] = 32'h0;  // 32'h10eb7885;
    ram_cell[    2236] = 32'h0;  // 32'h04f22926;
    ram_cell[    2237] = 32'h0;  // 32'h7c09af0f;
    ram_cell[    2238] = 32'h0;  // 32'hc4645e60;
    ram_cell[    2239] = 32'h0;  // 32'h5c472bf4;
    ram_cell[    2240] = 32'h0;  // 32'h947c60bb;
    ram_cell[    2241] = 32'h0;  // 32'he3233e7b;
    ram_cell[    2242] = 32'h0;  // 32'h82fdb534;
    ram_cell[    2243] = 32'h0;  // 32'hda368f89;
    ram_cell[    2244] = 32'h0;  // 32'hbe688134;
    ram_cell[    2245] = 32'h0;  // 32'h84c69881;
    ram_cell[    2246] = 32'h0;  // 32'hcdfb70ac;
    ram_cell[    2247] = 32'h0;  // 32'hb0496f1b;
    ram_cell[    2248] = 32'h0;  // 32'h989cfd59;
    ram_cell[    2249] = 32'h0;  // 32'hc8d45b14;
    ram_cell[    2250] = 32'h0;  // 32'h7bd535b3;
    ram_cell[    2251] = 32'h0;  // 32'ha4b0b497;
    ram_cell[    2252] = 32'h0;  // 32'hbbe5aa20;
    ram_cell[    2253] = 32'h0;  // 32'h86490621;
    ram_cell[    2254] = 32'h0;  // 32'ha793c970;
    ram_cell[    2255] = 32'h0;  // 32'h58f267c9;
    ram_cell[    2256] = 32'h0;  // 32'hc75bcda8;
    ram_cell[    2257] = 32'h0;  // 32'h108ced12;
    ram_cell[    2258] = 32'h0;  // 32'h12d4ba96;
    ram_cell[    2259] = 32'h0;  // 32'h543989ee;
    ram_cell[    2260] = 32'h0;  // 32'h2ea12fac;
    ram_cell[    2261] = 32'h0;  // 32'h75305626;
    ram_cell[    2262] = 32'h0;  // 32'h0c0cfbe9;
    ram_cell[    2263] = 32'h0;  // 32'he622c299;
    ram_cell[    2264] = 32'h0;  // 32'hf847f61a;
    ram_cell[    2265] = 32'h0;  // 32'hcb8fd2bd;
    ram_cell[    2266] = 32'h0;  // 32'h2bc8e197;
    ram_cell[    2267] = 32'h0;  // 32'hd1e0e756;
    ram_cell[    2268] = 32'h0;  // 32'h93dbdf9f;
    ram_cell[    2269] = 32'h0;  // 32'h1de818b6;
    ram_cell[    2270] = 32'h0;  // 32'hd1e22ae4;
    ram_cell[    2271] = 32'h0;  // 32'h783f0e6c;
    ram_cell[    2272] = 32'h0;  // 32'h5453a3d4;
    ram_cell[    2273] = 32'h0;  // 32'h8b16a20d;
    ram_cell[    2274] = 32'h0;  // 32'hc26c66bb;
    ram_cell[    2275] = 32'h0;  // 32'h9b94b841;
    ram_cell[    2276] = 32'h0;  // 32'h4e1a3725;
    ram_cell[    2277] = 32'h0;  // 32'hca2c0fef;
    ram_cell[    2278] = 32'h0;  // 32'hc8f30581;
    ram_cell[    2279] = 32'h0;  // 32'h67a7e83d;
    ram_cell[    2280] = 32'h0;  // 32'h335797d1;
    ram_cell[    2281] = 32'h0;  // 32'hde0e6059;
    ram_cell[    2282] = 32'h0;  // 32'hd6a42884;
    ram_cell[    2283] = 32'h0;  // 32'h6aed7331;
    ram_cell[    2284] = 32'h0;  // 32'ha5e6c60c;
    ram_cell[    2285] = 32'h0;  // 32'hf2254875;
    ram_cell[    2286] = 32'h0;  // 32'hd6a5f155;
    ram_cell[    2287] = 32'h0;  // 32'h799df49f;
    ram_cell[    2288] = 32'h0;  // 32'h7a2cccc3;
    ram_cell[    2289] = 32'h0;  // 32'hdf205582;
    ram_cell[    2290] = 32'h0;  // 32'h4c1b4f88;
    ram_cell[    2291] = 32'h0;  // 32'h16981a9d;
    ram_cell[    2292] = 32'h0;  // 32'hdd6adc1a;
    ram_cell[    2293] = 32'h0;  // 32'h70f33c90;
    ram_cell[    2294] = 32'h0;  // 32'hf5277867;
    ram_cell[    2295] = 32'h0;  // 32'h871f49a2;
    ram_cell[    2296] = 32'h0;  // 32'h6d510f81;
    ram_cell[    2297] = 32'h0;  // 32'h35c965dc;
    ram_cell[    2298] = 32'h0;  // 32'hb61ec7ff;
    ram_cell[    2299] = 32'h0;  // 32'he0a3e501;
    ram_cell[    2300] = 32'h0;  // 32'h053ccbfd;
    ram_cell[    2301] = 32'h0;  // 32'h8d28ba22;
    ram_cell[    2302] = 32'h0;  // 32'h196d5afe;
    ram_cell[    2303] = 32'h0;  // 32'h4b39eb84;
    ram_cell[    2304] = 32'h0;  // 32'h0859c475;
    ram_cell[    2305] = 32'h0;  // 32'h5b56097d;
    ram_cell[    2306] = 32'h0;  // 32'h75b03c18;
    ram_cell[    2307] = 32'h0;  // 32'hb5972ab2;
    ram_cell[    2308] = 32'h0;  // 32'h6aa647c7;
    ram_cell[    2309] = 32'h0;  // 32'ha67d2958;
    ram_cell[    2310] = 32'h0;  // 32'h7d88b30b;
    ram_cell[    2311] = 32'h0;  // 32'h0b53bbcf;
    ram_cell[    2312] = 32'h0;  // 32'h91848398;
    ram_cell[    2313] = 32'h0;  // 32'h305b7d4a;
    ram_cell[    2314] = 32'h0;  // 32'h1a3e9455;
    ram_cell[    2315] = 32'h0;  // 32'h006638dd;
    ram_cell[    2316] = 32'h0;  // 32'h712f6998;
    ram_cell[    2317] = 32'h0;  // 32'hd9522eb5;
    ram_cell[    2318] = 32'h0;  // 32'h67b999f3;
    ram_cell[    2319] = 32'h0;  // 32'h9b38fc01;
    ram_cell[    2320] = 32'h0;  // 32'h4bcda710;
    ram_cell[    2321] = 32'h0;  // 32'h7c773357;
    ram_cell[    2322] = 32'h0;  // 32'h61866ea3;
    ram_cell[    2323] = 32'h0;  // 32'h03f58b27;
    ram_cell[    2324] = 32'h0;  // 32'h87dc261e;
    ram_cell[    2325] = 32'h0;  // 32'ha6d3db9f;
    ram_cell[    2326] = 32'h0;  // 32'h8d52058c;
    ram_cell[    2327] = 32'h0;  // 32'h99682fdb;
    ram_cell[    2328] = 32'h0;  // 32'h5583e5ab;
    ram_cell[    2329] = 32'h0;  // 32'h000747c3;
    ram_cell[    2330] = 32'h0;  // 32'ha09092ed;
    ram_cell[    2331] = 32'h0;  // 32'hea19c4da;
    ram_cell[    2332] = 32'h0;  // 32'h65eefbe6;
    ram_cell[    2333] = 32'h0;  // 32'h6b96cd48;
    ram_cell[    2334] = 32'h0;  // 32'hfac236d2;
    ram_cell[    2335] = 32'h0;  // 32'h9472a876;
    ram_cell[    2336] = 32'h0;  // 32'hf6a42a23;
    ram_cell[    2337] = 32'h0;  // 32'h883f193b;
    ram_cell[    2338] = 32'h0;  // 32'hac8d2929;
    ram_cell[    2339] = 32'h0;  // 32'h05a2323e;
    ram_cell[    2340] = 32'h0;  // 32'h2b86aeb2;
    ram_cell[    2341] = 32'h0;  // 32'hfcc7176a;
    ram_cell[    2342] = 32'h0;  // 32'h7cd74746;
    ram_cell[    2343] = 32'h0;  // 32'h5451b0b7;
    ram_cell[    2344] = 32'h0;  // 32'h8579d3a9;
    ram_cell[    2345] = 32'h0;  // 32'ha7c4b9d2;
    ram_cell[    2346] = 32'h0;  // 32'hb889cfed;
    ram_cell[    2347] = 32'h0;  // 32'h6112a4cc;
    ram_cell[    2348] = 32'h0;  // 32'hae2e9aca;
    ram_cell[    2349] = 32'h0;  // 32'h980b9fb1;
    ram_cell[    2350] = 32'h0;  // 32'h6bc828a9;
    ram_cell[    2351] = 32'h0;  // 32'h7796c921;
    ram_cell[    2352] = 32'h0;  // 32'heedfb219;
    ram_cell[    2353] = 32'h0;  // 32'h0f42cb7c;
    ram_cell[    2354] = 32'h0;  // 32'h06f1b6ad;
    ram_cell[    2355] = 32'h0;  // 32'h75906ae8;
    ram_cell[    2356] = 32'h0;  // 32'h5fbb9b75;
    ram_cell[    2357] = 32'h0;  // 32'h74fd7205;
    ram_cell[    2358] = 32'h0;  // 32'hb80d4386;
    ram_cell[    2359] = 32'h0;  // 32'hb352ea84;
    ram_cell[    2360] = 32'h0;  // 32'h6760b2e7;
    ram_cell[    2361] = 32'h0;  // 32'h6aeffd4b;
    ram_cell[    2362] = 32'h0;  // 32'hc344f740;
    ram_cell[    2363] = 32'h0;  // 32'h06c6a85f;
    ram_cell[    2364] = 32'h0;  // 32'hf6896040;
    ram_cell[    2365] = 32'h0;  // 32'he2852664;
    ram_cell[    2366] = 32'h0;  // 32'h4a8f4a4e;
    ram_cell[    2367] = 32'h0;  // 32'hd3d31303;
    ram_cell[    2368] = 32'h0;  // 32'h7088b12a;
    ram_cell[    2369] = 32'h0;  // 32'hc6f323ce;
    ram_cell[    2370] = 32'h0;  // 32'h420087cb;
    ram_cell[    2371] = 32'h0;  // 32'h034783e4;
    ram_cell[    2372] = 32'h0;  // 32'h9d6d3ee2;
    ram_cell[    2373] = 32'h0;  // 32'h3992a719;
    ram_cell[    2374] = 32'h0;  // 32'h6f81ef50;
    ram_cell[    2375] = 32'h0;  // 32'h37fdff5f;
    ram_cell[    2376] = 32'h0;  // 32'h6f3d18c4;
    ram_cell[    2377] = 32'h0;  // 32'hfae35cea;
    ram_cell[    2378] = 32'h0;  // 32'h34b72d6d;
    ram_cell[    2379] = 32'h0;  // 32'h41291b1f;
    ram_cell[    2380] = 32'h0;  // 32'h9d202060;
    ram_cell[    2381] = 32'h0;  // 32'h17331d95;
    ram_cell[    2382] = 32'h0;  // 32'hfcf98fdb;
    ram_cell[    2383] = 32'h0;  // 32'h8bddd04b;
    ram_cell[    2384] = 32'h0;  // 32'h6a850bed;
    ram_cell[    2385] = 32'h0;  // 32'h72ab72b5;
    ram_cell[    2386] = 32'h0;  // 32'h04c014c8;
    ram_cell[    2387] = 32'h0;  // 32'h3df8b6b3;
    ram_cell[    2388] = 32'h0;  // 32'h83fd4487;
    ram_cell[    2389] = 32'h0;  // 32'hb6242d07;
    ram_cell[    2390] = 32'h0;  // 32'h9f61c440;
    ram_cell[    2391] = 32'h0;  // 32'hf9b738ab;
    ram_cell[    2392] = 32'h0;  // 32'h5e057367;
    ram_cell[    2393] = 32'h0;  // 32'haa881d3e;
    ram_cell[    2394] = 32'h0;  // 32'h47b3b980;
    ram_cell[    2395] = 32'h0;  // 32'h64889ced;
    ram_cell[    2396] = 32'h0;  // 32'he5c32837;
    ram_cell[    2397] = 32'h0;  // 32'hbdc03020;
    ram_cell[    2398] = 32'h0;  // 32'h2c02a55a;
    ram_cell[    2399] = 32'h0;  // 32'h545392de;
    ram_cell[    2400] = 32'h0;  // 32'h3b34a2c1;
    ram_cell[    2401] = 32'h0;  // 32'h9061f720;
    ram_cell[    2402] = 32'h0;  // 32'h23863818;
    ram_cell[    2403] = 32'h0;  // 32'h9fb8fb12;
    ram_cell[    2404] = 32'h0;  // 32'hdce24e12;
    ram_cell[    2405] = 32'h0;  // 32'h3d0fa2f8;
    ram_cell[    2406] = 32'h0;  // 32'h4add043d;
    ram_cell[    2407] = 32'h0;  // 32'h5d6ae62b;
    ram_cell[    2408] = 32'h0;  // 32'hbabb18f1;
    ram_cell[    2409] = 32'h0;  // 32'heaa8402d;
    ram_cell[    2410] = 32'h0;  // 32'hb53e6c40;
    ram_cell[    2411] = 32'h0;  // 32'he6d652d3;
    ram_cell[    2412] = 32'h0;  // 32'hbbbeda46;
    ram_cell[    2413] = 32'h0;  // 32'hf35f9057;
    ram_cell[    2414] = 32'h0;  // 32'h34a1c2af;
    ram_cell[    2415] = 32'h0;  // 32'hae455ed3;
    ram_cell[    2416] = 32'h0;  // 32'h070b642c;
    ram_cell[    2417] = 32'h0;  // 32'h33cd7799;
    ram_cell[    2418] = 32'h0;  // 32'he711bc8d;
    ram_cell[    2419] = 32'h0;  // 32'h8a520365;
    ram_cell[    2420] = 32'h0;  // 32'h2fabba2e;
    ram_cell[    2421] = 32'h0;  // 32'h473eaaa4;
    ram_cell[    2422] = 32'h0;  // 32'hed191de8;
    ram_cell[    2423] = 32'h0;  // 32'h8b411caf;
    ram_cell[    2424] = 32'h0;  // 32'hf01abe1a;
    ram_cell[    2425] = 32'h0;  // 32'h47796431;
    ram_cell[    2426] = 32'h0;  // 32'hfb72b864;
    ram_cell[    2427] = 32'h0;  // 32'h5deae654;
    ram_cell[    2428] = 32'h0;  // 32'h8ec27aaf;
    ram_cell[    2429] = 32'h0;  // 32'h73918a6f;
    ram_cell[    2430] = 32'h0;  // 32'h66affd27;
    ram_cell[    2431] = 32'h0;  // 32'h33dcf9e6;
    ram_cell[    2432] = 32'h0;  // 32'ha8a0f6a0;
    ram_cell[    2433] = 32'h0;  // 32'hbfd74eda;
    ram_cell[    2434] = 32'h0;  // 32'hae367c18;
    ram_cell[    2435] = 32'h0;  // 32'h1c9d40a9;
    ram_cell[    2436] = 32'h0;  // 32'h9fcd62b0;
    ram_cell[    2437] = 32'h0;  // 32'ha1c11aae;
    ram_cell[    2438] = 32'h0;  // 32'h4b72d98e;
    ram_cell[    2439] = 32'h0;  // 32'ha66c38ad;
    ram_cell[    2440] = 32'h0;  // 32'h98580d69;
    ram_cell[    2441] = 32'h0;  // 32'h40a40746;
    ram_cell[    2442] = 32'h0;  // 32'h6b862d6c;
    ram_cell[    2443] = 32'h0;  // 32'h16050830;
    ram_cell[    2444] = 32'h0;  // 32'h3065598a;
    ram_cell[    2445] = 32'h0;  // 32'ha9aafac0;
    ram_cell[    2446] = 32'h0;  // 32'h1cf42a2f;
    ram_cell[    2447] = 32'h0;  // 32'h39455985;
    ram_cell[    2448] = 32'h0;  // 32'h7ed9af94;
    ram_cell[    2449] = 32'h0;  // 32'haf309753;
    ram_cell[    2450] = 32'h0;  // 32'h2bacd72f;
    ram_cell[    2451] = 32'h0;  // 32'h8fb33992;
    ram_cell[    2452] = 32'h0;  // 32'h1f81c2af;
    ram_cell[    2453] = 32'h0;  // 32'ha7d8701c;
    ram_cell[    2454] = 32'h0;  // 32'he175e1de;
    ram_cell[    2455] = 32'h0;  // 32'h5cec1628;
    ram_cell[    2456] = 32'h0;  // 32'h6ef10867;
    ram_cell[    2457] = 32'h0;  // 32'hcd8bfb25;
    ram_cell[    2458] = 32'h0;  // 32'h37263357;
    ram_cell[    2459] = 32'h0;  // 32'hf02ffff5;
    ram_cell[    2460] = 32'h0;  // 32'hdb2be4cb;
    ram_cell[    2461] = 32'h0;  // 32'hc5f3d4a9;
    ram_cell[    2462] = 32'h0;  // 32'hafcac30a;
    ram_cell[    2463] = 32'h0;  // 32'hb6752270;
    ram_cell[    2464] = 32'h0;  // 32'h0ac8b51b;
    ram_cell[    2465] = 32'h0;  // 32'h562d05c7;
    ram_cell[    2466] = 32'h0;  // 32'h377cacb4;
    ram_cell[    2467] = 32'h0;  // 32'h2b74a42c;
    ram_cell[    2468] = 32'h0;  // 32'hd983a262;
    ram_cell[    2469] = 32'h0;  // 32'hc1517a51;
    ram_cell[    2470] = 32'h0;  // 32'h11272a56;
    ram_cell[    2471] = 32'h0;  // 32'h9d253c2c;
    ram_cell[    2472] = 32'h0;  // 32'hbe5f76be;
    ram_cell[    2473] = 32'h0;  // 32'h826bd097;
    ram_cell[    2474] = 32'h0;  // 32'hbd939e67;
    ram_cell[    2475] = 32'h0;  // 32'ha3709847;
    ram_cell[    2476] = 32'h0;  // 32'h9e72b1f2;
    ram_cell[    2477] = 32'h0;  // 32'hab41e208;
    ram_cell[    2478] = 32'h0;  // 32'hb9338f76;
    ram_cell[    2479] = 32'h0;  // 32'h1eab1c31;
    ram_cell[    2480] = 32'h0;  // 32'hae17dd5c;
    ram_cell[    2481] = 32'h0;  // 32'hbc82dff3;
    ram_cell[    2482] = 32'h0;  // 32'h3a1e9190;
    ram_cell[    2483] = 32'h0;  // 32'h61c93afa;
    ram_cell[    2484] = 32'h0;  // 32'h92b650b2;
    ram_cell[    2485] = 32'h0;  // 32'h67d8fba7;
    ram_cell[    2486] = 32'h0;  // 32'h3b6e4b89;
    ram_cell[    2487] = 32'h0;  // 32'h1f1b5554;
    ram_cell[    2488] = 32'h0;  // 32'hacb0b950;
    ram_cell[    2489] = 32'h0;  // 32'hd5c42c79;
    ram_cell[    2490] = 32'h0;  // 32'h419974ff;
    ram_cell[    2491] = 32'h0;  // 32'h8c2137a4;
    ram_cell[    2492] = 32'h0;  // 32'h394043de;
    ram_cell[    2493] = 32'h0;  // 32'h4b36ff45;
    ram_cell[    2494] = 32'h0;  // 32'h5487530e;
    ram_cell[    2495] = 32'h0;  // 32'h60f4f192;
    ram_cell[    2496] = 32'h0;  // 32'h4da44158;
    ram_cell[    2497] = 32'h0;  // 32'haf6f8e55;
    ram_cell[    2498] = 32'h0;  // 32'he14e42aa;
    ram_cell[    2499] = 32'h0;  // 32'ha5e8dc7e;
    ram_cell[    2500] = 32'h0;  // 32'h6a895631;
    ram_cell[    2501] = 32'h0;  // 32'h2691dbfb;
    ram_cell[    2502] = 32'h0;  // 32'hcc77e900;
    ram_cell[    2503] = 32'h0;  // 32'h99fb5999;
    ram_cell[    2504] = 32'h0;  // 32'hffca848e;
    ram_cell[    2505] = 32'h0;  // 32'h49971a09;
    ram_cell[    2506] = 32'h0;  // 32'h26349b7f;
    ram_cell[    2507] = 32'h0;  // 32'hc9ae18ed;
    ram_cell[    2508] = 32'h0;  // 32'h502914f8;
    ram_cell[    2509] = 32'h0;  // 32'h829bf238;
    ram_cell[    2510] = 32'h0;  // 32'h1fd03cf4;
    ram_cell[    2511] = 32'h0;  // 32'hc363c10a;
    ram_cell[    2512] = 32'h0;  // 32'hfa6377d9;
    ram_cell[    2513] = 32'h0;  // 32'h030b8a62;
    ram_cell[    2514] = 32'h0;  // 32'hfda2b014;
    ram_cell[    2515] = 32'h0;  // 32'hd5b2a8ff;
    ram_cell[    2516] = 32'h0;  // 32'hbc17e26e;
    ram_cell[    2517] = 32'h0;  // 32'h0546da01;
    ram_cell[    2518] = 32'h0;  // 32'he780bb43;
    ram_cell[    2519] = 32'h0;  // 32'h1c32feab;
    ram_cell[    2520] = 32'h0;  // 32'he43ff654;
    ram_cell[    2521] = 32'h0;  // 32'h95936235;
    ram_cell[    2522] = 32'h0;  // 32'hf33a8ef5;
    ram_cell[    2523] = 32'h0;  // 32'h653443b1;
    ram_cell[    2524] = 32'h0;  // 32'h84f9a416;
    ram_cell[    2525] = 32'h0;  // 32'hd5d62fdf;
    ram_cell[    2526] = 32'h0;  // 32'h385ad0a7;
    ram_cell[    2527] = 32'h0;  // 32'h6b2f2c7c;
    ram_cell[    2528] = 32'h0;  // 32'h25df28c1;
    ram_cell[    2529] = 32'h0;  // 32'hf5f00868;
    ram_cell[    2530] = 32'h0;  // 32'hf670ca5a;
    ram_cell[    2531] = 32'h0;  // 32'h0da8aa9a;
    ram_cell[    2532] = 32'h0;  // 32'h894ee93a;
    ram_cell[    2533] = 32'h0;  // 32'h3ec379ad;
    ram_cell[    2534] = 32'h0;  // 32'h51012551;
    ram_cell[    2535] = 32'h0;  // 32'h4033d1ce;
    ram_cell[    2536] = 32'h0;  // 32'h57292ef0;
    ram_cell[    2537] = 32'h0;  // 32'hb993c854;
    ram_cell[    2538] = 32'h0;  // 32'h920bb2c2;
    ram_cell[    2539] = 32'h0;  // 32'h60c273f5;
    ram_cell[    2540] = 32'h0;  // 32'h73ccb187;
    ram_cell[    2541] = 32'h0;  // 32'hf82d10f8;
    ram_cell[    2542] = 32'h0;  // 32'h0d41e9f4;
    ram_cell[    2543] = 32'h0;  // 32'hd8f3492a;
    ram_cell[    2544] = 32'h0;  // 32'h7a1db361;
    ram_cell[    2545] = 32'h0;  // 32'h14872658;
    ram_cell[    2546] = 32'h0;  // 32'h70d09b27;
    ram_cell[    2547] = 32'h0;  // 32'h0c147b5a;
    ram_cell[    2548] = 32'h0;  // 32'h2fc2ba0e;
    ram_cell[    2549] = 32'h0;  // 32'hdf78fb61;
    ram_cell[    2550] = 32'h0;  // 32'h5ffde277;
    ram_cell[    2551] = 32'h0;  // 32'h98fc3d4e;
    ram_cell[    2552] = 32'h0;  // 32'hc26e979a;
    ram_cell[    2553] = 32'h0;  // 32'hcc70b318;
    ram_cell[    2554] = 32'h0;  // 32'h6eab5946;
    ram_cell[    2555] = 32'h0;  // 32'heb204f58;
    ram_cell[    2556] = 32'h0;  // 32'h7a3f76e4;
    ram_cell[    2557] = 32'h0;  // 32'hca95add2;
    ram_cell[    2558] = 32'h0;  // 32'hea7b1ef0;
    ram_cell[    2559] = 32'h0;  // 32'h26c68c5c;
    ram_cell[    2560] = 32'h0;  // 32'h72d6960d;
    ram_cell[    2561] = 32'h0;  // 32'h7a53741e;
    ram_cell[    2562] = 32'h0;  // 32'hf441ce58;
    ram_cell[    2563] = 32'h0;  // 32'h4ad8e2d4;
    ram_cell[    2564] = 32'h0;  // 32'h4ceacf28;
    ram_cell[    2565] = 32'h0;  // 32'h5f2215fd;
    ram_cell[    2566] = 32'h0;  // 32'h3a71a96e;
    ram_cell[    2567] = 32'h0;  // 32'hbe784b8c;
    ram_cell[    2568] = 32'h0;  // 32'hb7a8e804;
    ram_cell[    2569] = 32'h0;  // 32'h6dd529ca;
    ram_cell[    2570] = 32'h0;  // 32'hd4de6228;
    ram_cell[    2571] = 32'h0;  // 32'hdbf32a99;
    ram_cell[    2572] = 32'h0;  // 32'h60c0327a;
    ram_cell[    2573] = 32'h0;  // 32'hdc8abe4c;
    ram_cell[    2574] = 32'h0;  // 32'h5250bff1;
    ram_cell[    2575] = 32'h0;  // 32'heb696377;
    ram_cell[    2576] = 32'h0;  // 32'he7c82273;
    ram_cell[    2577] = 32'h0;  // 32'hb9321d4b;
    ram_cell[    2578] = 32'h0;  // 32'h966a2e86;
    ram_cell[    2579] = 32'h0;  // 32'h7e28674b;
    ram_cell[    2580] = 32'h0;  // 32'he1263e6e;
    ram_cell[    2581] = 32'h0;  // 32'hcaab45ea;
    ram_cell[    2582] = 32'h0;  // 32'h2f1af3ca;
    ram_cell[    2583] = 32'h0;  // 32'h64e39eea;
    ram_cell[    2584] = 32'h0;  // 32'h75abb930;
    ram_cell[    2585] = 32'h0;  // 32'hf926b040;
    ram_cell[    2586] = 32'h0;  // 32'h065fcef0;
    ram_cell[    2587] = 32'h0;  // 32'h6e4dd685;
    ram_cell[    2588] = 32'h0;  // 32'h394a7f56;
    ram_cell[    2589] = 32'h0;  // 32'he6407678;
    ram_cell[    2590] = 32'h0;  // 32'h64d7a959;
    ram_cell[    2591] = 32'h0;  // 32'h1fb3d33d;
    ram_cell[    2592] = 32'h0;  // 32'h3efc8ed9;
    ram_cell[    2593] = 32'h0;  // 32'he7c87432;
    ram_cell[    2594] = 32'h0;  // 32'hd52a2afe;
    ram_cell[    2595] = 32'h0;  // 32'h8b0542ba;
    ram_cell[    2596] = 32'h0;  // 32'h6c4c3177;
    ram_cell[    2597] = 32'h0;  // 32'hde923f4f;
    ram_cell[    2598] = 32'h0;  // 32'heca45d04;
    ram_cell[    2599] = 32'h0;  // 32'h73e3f459;
    ram_cell[    2600] = 32'h0;  // 32'he381b457;
    ram_cell[    2601] = 32'h0;  // 32'h35c26587;
    ram_cell[    2602] = 32'h0;  // 32'h5ccac9cd;
    ram_cell[    2603] = 32'h0;  // 32'he96451aa;
    ram_cell[    2604] = 32'h0;  // 32'h0dabb5dd;
    ram_cell[    2605] = 32'h0;  // 32'h46005441;
    ram_cell[    2606] = 32'h0;  // 32'h890e77a4;
    ram_cell[    2607] = 32'h0;  // 32'hff2700dc;
    ram_cell[    2608] = 32'h0;  // 32'hd5ab3f71;
    ram_cell[    2609] = 32'h0;  // 32'ha3630003;
    ram_cell[    2610] = 32'h0;  // 32'h6440d255;
    ram_cell[    2611] = 32'h0;  // 32'h7680a544;
    ram_cell[    2612] = 32'h0;  // 32'hf39a9d45;
    ram_cell[    2613] = 32'h0;  // 32'he5a0b0bf;
    ram_cell[    2614] = 32'h0;  // 32'h232367e1;
    ram_cell[    2615] = 32'h0;  // 32'ha036fa9a;
    ram_cell[    2616] = 32'h0;  // 32'h94e74523;
    ram_cell[    2617] = 32'h0;  // 32'h97936f1d;
    ram_cell[    2618] = 32'h0;  // 32'hd077f1d6;
    ram_cell[    2619] = 32'h0;  // 32'h67f0af3b;
    ram_cell[    2620] = 32'h0;  // 32'h78b177b3;
    ram_cell[    2621] = 32'h0;  // 32'h8b57ca52;
    ram_cell[    2622] = 32'h0;  // 32'h20908297;
    ram_cell[    2623] = 32'h0;  // 32'h60a35b62;
    ram_cell[    2624] = 32'h0;  // 32'ha8267c84;
    ram_cell[    2625] = 32'h0;  // 32'h9a2bdd96;
    ram_cell[    2626] = 32'h0;  // 32'hc5924cbc;
    ram_cell[    2627] = 32'h0;  // 32'h9e2fed65;
    ram_cell[    2628] = 32'h0;  // 32'h86c4d9f4;
    ram_cell[    2629] = 32'h0;  // 32'h18d09d97;
    ram_cell[    2630] = 32'h0;  // 32'h89f36953;
    ram_cell[    2631] = 32'h0;  // 32'hd1e7c6b8;
    ram_cell[    2632] = 32'h0;  // 32'h6979b474;
    ram_cell[    2633] = 32'h0;  // 32'he181da12;
    ram_cell[    2634] = 32'h0;  // 32'hc1ee7316;
    ram_cell[    2635] = 32'h0;  // 32'h69bea922;
    ram_cell[    2636] = 32'h0;  // 32'h1244c8cb;
    ram_cell[    2637] = 32'h0;  // 32'h588b4bbb;
    ram_cell[    2638] = 32'h0;  // 32'hcb085334;
    ram_cell[    2639] = 32'h0;  // 32'h93ab7abf;
    ram_cell[    2640] = 32'h0;  // 32'hafe6f86a;
    ram_cell[    2641] = 32'h0;  // 32'h8af69402;
    ram_cell[    2642] = 32'h0;  // 32'he7df01dc;
    ram_cell[    2643] = 32'h0;  // 32'h6f1a2264;
    ram_cell[    2644] = 32'h0;  // 32'h7624998f;
    ram_cell[    2645] = 32'h0;  // 32'hc14b38d2;
    ram_cell[    2646] = 32'h0;  // 32'h762bc55d;
    ram_cell[    2647] = 32'h0;  // 32'hf98ac395;
    ram_cell[    2648] = 32'h0;  // 32'h269153d6;
    ram_cell[    2649] = 32'h0;  // 32'h90158e0c;
    ram_cell[    2650] = 32'h0;  // 32'h65197f3a;
    ram_cell[    2651] = 32'h0;  // 32'h395e68cd;
    ram_cell[    2652] = 32'h0;  // 32'h40c9bb39;
    ram_cell[    2653] = 32'h0;  // 32'hb9ca71e8;
    ram_cell[    2654] = 32'h0;  // 32'h1d890ca1;
    ram_cell[    2655] = 32'h0;  // 32'h6d544305;
    ram_cell[    2656] = 32'h0;  // 32'h060a9af6;
    ram_cell[    2657] = 32'h0;  // 32'h1baaf1de;
    ram_cell[    2658] = 32'h0;  // 32'h83597862;
    ram_cell[    2659] = 32'h0;  // 32'hc2a3021a;
    ram_cell[    2660] = 32'h0;  // 32'ha2f4fd90;
    ram_cell[    2661] = 32'h0;  // 32'hf646454e;
    ram_cell[    2662] = 32'h0;  // 32'h12c04820;
    ram_cell[    2663] = 32'h0;  // 32'h263f4f45;
    ram_cell[    2664] = 32'h0;  // 32'h74b29d09;
    ram_cell[    2665] = 32'h0;  // 32'h0dafa4f7;
    ram_cell[    2666] = 32'h0;  // 32'h2d8dde0f;
    ram_cell[    2667] = 32'h0;  // 32'h0172860e;
    ram_cell[    2668] = 32'h0;  // 32'hbc7adb0e;
    ram_cell[    2669] = 32'h0;  // 32'hb1ffda07;
    ram_cell[    2670] = 32'h0;  // 32'h474764ce;
    ram_cell[    2671] = 32'h0;  // 32'heb058a2b;
    ram_cell[    2672] = 32'h0;  // 32'he5fc9aaa;
    ram_cell[    2673] = 32'h0;  // 32'h6a10104a;
    ram_cell[    2674] = 32'h0;  // 32'h07cfa6a4;
    ram_cell[    2675] = 32'h0;  // 32'h50b23fb2;
    ram_cell[    2676] = 32'h0;  // 32'h9963081c;
    ram_cell[    2677] = 32'h0;  // 32'hda61623a;
    ram_cell[    2678] = 32'h0;  // 32'h90a5b358;
    ram_cell[    2679] = 32'h0;  // 32'hbec87bd0;
    ram_cell[    2680] = 32'h0;  // 32'h7fb2b912;
    ram_cell[    2681] = 32'h0;  // 32'h056c4213;
    ram_cell[    2682] = 32'h0;  // 32'h1f5164a8;
    ram_cell[    2683] = 32'h0;  // 32'h8607bc17;
    ram_cell[    2684] = 32'h0;  // 32'h7cb4b1a1;
    ram_cell[    2685] = 32'h0;  // 32'h16ca645b;
    ram_cell[    2686] = 32'h0;  // 32'h4ecc72c9;
    ram_cell[    2687] = 32'h0;  // 32'he2270bf6;
    ram_cell[    2688] = 32'h0;  // 32'h8f2c444d;
    ram_cell[    2689] = 32'h0;  // 32'h76e09868;
    ram_cell[    2690] = 32'h0;  // 32'hdc48e0f1;
    ram_cell[    2691] = 32'h0;  // 32'hae8d5c54;
    ram_cell[    2692] = 32'h0;  // 32'h28a4b207;
    ram_cell[    2693] = 32'h0;  // 32'h2c862549;
    ram_cell[    2694] = 32'h0;  // 32'h897998fd;
    ram_cell[    2695] = 32'h0;  // 32'h131c5f95;
    ram_cell[    2696] = 32'h0;  // 32'h54c92636;
    ram_cell[    2697] = 32'h0;  // 32'h05827ffb;
    ram_cell[    2698] = 32'h0;  // 32'h462888b8;
    ram_cell[    2699] = 32'h0;  // 32'h89d2bcd0;
    ram_cell[    2700] = 32'h0;  // 32'h0bb78df4;
    ram_cell[    2701] = 32'h0;  // 32'h8c298b81;
    ram_cell[    2702] = 32'h0;  // 32'h1e551c6b;
    ram_cell[    2703] = 32'h0;  // 32'h836d0028;
    ram_cell[    2704] = 32'h0;  // 32'he895955f;
    ram_cell[    2705] = 32'h0;  // 32'h8d57871e;
    ram_cell[    2706] = 32'h0;  // 32'he60927b4;
    ram_cell[    2707] = 32'h0;  // 32'hb9a090f1;
    ram_cell[    2708] = 32'h0;  // 32'h97625911;
    ram_cell[    2709] = 32'h0;  // 32'h17561287;
    ram_cell[    2710] = 32'h0;  // 32'h6e495271;
    ram_cell[    2711] = 32'h0;  // 32'hd9d27e60;
    ram_cell[    2712] = 32'h0;  // 32'h5d72b10d;
    ram_cell[    2713] = 32'h0;  // 32'h18c4faaf;
    ram_cell[    2714] = 32'h0;  // 32'h73be807d;
    ram_cell[    2715] = 32'h0;  // 32'hf02d401d;
    ram_cell[    2716] = 32'h0;  // 32'h2deb5846;
    ram_cell[    2717] = 32'h0;  // 32'h623e5789;
    ram_cell[    2718] = 32'h0;  // 32'hf73b4e74;
    ram_cell[    2719] = 32'h0;  // 32'h08e6ec22;
    ram_cell[    2720] = 32'h0;  // 32'hd374483f;
    ram_cell[    2721] = 32'h0;  // 32'hc35b0150;
    ram_cell[    2722] = 32'h0;  // 32'h45f1f617;
    ram_cell[    2723] = 32'h0;  // 32'h91d1bbdb;
    ram_cell[    2724] = 32'h0;  // 32'hdf11639d;
    ram_cell[    2725] = 32'h0;  // 32'hbe821501;
    ram_cell[    2726] = 32'h0;  // 32'hdc7861b9;
    ram_cell[    2727] = 32'h0;  // 32'h17f1078f;
    ram_cell[    2728] = 32'h0;  // 32'h443c6f07;
    ram_cell[    2729] = 32'h0;  // 32'h64626aa6;
    ram_cell[    2730] = 32'h0;  // 32'h6693f496;
    ram_cell[    2731] = 32'h0;  // 32'h3e99e3a3;
    ram_cell[    2732] = 32'h0;  // 32'h474de8dc;
    ram_cell[    2733] = 32'h0;  // 32'h322dd18a;
    ram_cell[    2734] = 32'h0;  // 32'hef527ba5;
    ram_cell[    2735] = 32'h0;  // 32'haac92f49;
    ram_cell[    2736] = 32'h0;  // 32'hdd52c416;
    ram_cell[    2737] = 32'h0;  // 32'h6cf31634;
    ram_cell[    2738] = 32'h0;  // 32'hf407db58;
    ram_cell[    2739] = 32'h0;  // 32'h424dbb5c;
    ram_cell[    2740] = 32'h0;  // 32'h31ba30c0;
    ram_cell[    2741] = 32'h0;  // 32'h19a10f1d;
    ram_cell[    2742] = 32'h0;  // 32'hb73a842a;
    ram_cell[    2743] = 32'h0;  // 32'h8b5907b3;
    ram_cell[    2744] = 32'h0;  // 32'he5fc71d5;
    ram_cell[    2745] = 32'h0;  // 32'hb6c32fe6;
    ram_cell[    2746] = 32'h0;  // 32'h5009a91c;
    ram_cell[    2747] = 32'h0;  // 32'hc8be5977;
    ram_cell[    2748] = 32'h0;  // 32'h4876e923;
    ram_cell[    2749] = 32'h0;  // 32'hcae5dfb5;
    ram_cell[    2750] = 32'h0;  // 32'h0bdbe9ec;
    ram_cell[    2751] = 32'h0;  // 32'ha7a710b1;
    ram_cell[    2752] = 32'h0;  // 32'hc95ba60f;
    ram_cell[    2753] = 32'h0;  // 32'h02a444b8;
    ram_cell[    2754] = 32'h0;  // 32'h496da1be;
    ram_cell[    2755] = 32'h0;  // 32'h0024f10e;
    ram_cell[    2756] = 32'h0;  // 32'h6ac7c0e9;
    ram_cell[    2757] = 32'h0;  // 32'hd36b584e;
    ram_cell[    2758] = 32'h0;  // 32'hf25ec678;
    ram_cell[    2759] = 32'h0;  // 32'hf55acde6;
    ram_cell[    2760] = 32'h0;  // 32'hefd7ba8b;
    ram_cell[    2761] = 32'h0;  // 32'h2334dd8c;
    ram_cell[    2762] = 32'h0;  // 32'h43f633a3;
    ram_cell[    2763] = 32'h0;  // 32'h3d608f03;
    ram_cell[    2764] = 32'h0;  // 32'h778378f9;
    ram_cell[    2765] = 32'h0;  // 32'h218b183b;
    ram_cell[    2766] = 32'h0;  // 32'h6bac0b45;
    ram_cell[    2767] = 32'h0;  // 32'h770710a6;
    ram_cell[    2768] = 32'h0;  // 32'h7b2e1f8a;
    ram_cell[    2769] = 32'h0;  // 32'hbd96338d;
    ram_cell[    2770] = 32'h0;  // 32'h7c816259;
    ram_cell[    2771] = 32'h0;  // 32'hb0609a4c;
    ram_cell[    2772] = 32'h0;  // 32'h3d21ee76;
    ram_cell[    2773] = 32'h0;  // 32'heaa4390c;
    ram_cell[    2774] = 32'h0;  // 32'h5df9eead;
    ram_cell[    2775] = 32'h0;  // 32'h5d8ed9cc;
    ram_cell[    2776] = 32'h0;  // 32'h5acea1ad;
    ram_cell[    2777] = 32'h0;  // 32'h7e3c5d02;
    ram_cell[    2778] = 32'h0;  // 32'h4b5ea513;
    ram_cell[    2779] = 32'h0;  // 32'he7391009;
    ram_cell[    2780] = 32'h0;  // 32'h5cfca342;
    ram_cell[    2781] = 32'h0;  // 32'hfb191fde;
    ram_cell[    2782] = 32'h0;  // 32'h30452a16;
    ram_cell[    2783] = 32'h0;  // 32'hb8376881;
    ram_cell[    2784] = 32'h0;  // 32'h9280fa31;
    ram_cell[    2785] = 32'h0;  // 32'h9b8c8931;
    ram_cell[    2786] = 32'h0;  // 32'h8a84f837;
    ram_cell[    2787] = 32'h0;  // 32'h4c96de69;
    ram_cell[    2788] = 32'h0;  // 32'h7372647e;
    ram_cell[    2789] = 32'h0;  // 32'he6830b8f;
    ram_cell[    2790] = 32'h0;  // 32'h7c1e17cd;
    ram_cell[    2791] = 32'h0;  // 32'h0155d85e;
    ram_cell[    2792] = 32'h0;  // 32'h6a264143;
    ram_cell[    2793] = 32'h0;  // 32'h54e255bd;
    ram_cell[    2794] = 32'h0;  // 32'h0e26d230;
    ram_cell[    2795] = 32'h0;  // 32'hfec53f23;
    ram_cell[    2796] = 32'h0;  // 32'h16408c69;
    ram_cell[    2797] = 32'h0;  // 32'ha394a801;
    ram_cell[    2798] = 32'h0;  // 32'hd13f42db;
    ram_cell[    2799] = 32'h0;  // 32'hd75ba819;
    ram_cell[    2800] = 32'h0;  // 32'hb7ed3b24;
    ram_cell[    2801] = 32'h0;  // 32'h6263add3;
    ram_cell[    2802] = 32'h0;  // 32'h37fef16d;
    ram_cell[    2803] = 32'h0;  // 32'h5c52afc2;
    ram_cell[    2804] = 32'h0;  // 32'ha76a9617;
    ram_cell[    2805] = 32'h0;  // 32'hc4692872;
    ram_cell[    2806] = 32'h0;  // 32'h29b6d68e;
    ram_cell[    2807] = 32'h0;  // 32'ha34e9be6;
    ram_cell[    2808] = 32'h0;  // 32'hd6c5acf3;
    ram_cell[    2809] = 32'h0;  // 32'h72f6eed5;
    ram_cell[    2810] = 32'h0;  // 32'h90d2e381;
    ram_cell[    2811] = 32'h0;  // 32'h02b41563;
    ram_cell[    2812] = 32'h0;  // 32'h1c5b7050;
    ram_cell[    2813] = 32'h0;  // 32'hacd89ff0;
    ram_cell[    2814] = 32'h0;  // 32'hb5ec14f4;
    ram_cell[    2815] = 32'h0;  // 32'hc72de4bf;
    ram_cell[    2816] = 32'h0;  // 32'hb6e6feb7;
    ram_cell[    2817] = 32'h0;  // 32'h16fac2cb;
    ram_cell[    2818] = 32'h0;  // 32'ha35782f7;
    ram_cell[    2819] = 32'h0;  // 32'h29855aa9;
    ram_cell[    2820] = 32'h0;  // 32'hd9ca9559;
    ram_cell[    2821] = 32'h0;  // 32'ha7a3364e;
    ram_cell[    2822] = 32'h0;  // 32'h5d1af8c0;
    ram_cell[    2823] = 32'h0;  // 32'h78bf0598;
    ram_cell[    2824] = 32'h0;  // 32'h38995053;
    ram_cell[    2825] = 32'h0;  // 32'ha5b86fd2;
    ram_cell[    2826] = 32'h0;  // 32'h5c32b5c3;
    ram_cell[    2827] = 32'h0;  // 32'haa0e22e9;
    ram_cell[    2828] = 32'h0;  // 32'hc905d0a8;
    ram_cell[    2829] = 32'h0;  // 32'h3d2bb07a;
    ram_cell[    2830] = 32'h0;  // 32'h433e56cb;
    ram_cell[    2831] = 32'h0;  // 32'h84ce6a56;
    ram_cell[    2832] = 32'h0;  // 32'h121eb13f;
    ram_cell[    2833] = 32'h0;  // 32'h0bcbbed4;
    ram_cell[    2834] = 32'h0;  // 32'h41d31fb0;
    ram_cell[    2835] = 32'h0;  // 32'hf3895b8a;
    ram_cell[    2836] = 32'h0;  // 32'h55449b96;
    ram_cell[    2837] = 32'h0;  // 32'h3c175dc7;
    ram_cell[    2838] = 32'h0;  // 32'hfc7522d5;
    ram_cell[    2839] = 32'h0;  // 32'h6d34026a;
    ram_cell[    2840] = 32'h0;  // 32'h2e1af5d2;
    ram_cell[    2841] = 32'h0;  // 32'hf03a99a1;
    ram_cell[    2842] = 32'h0;  // 32'hdf397a44;
    ram_cell[    2843] = 32'h0;  // 32'h36b78d02;
    ram_cell[    2844] = 32'h0;  // 32'hcbac66f6;
    ram_cell[    2845] = 32'h0;  // 32'h20d1b3e5;
    ram_cell[    2846] = 32'h0;  // 32'h134bfef6;
    ram_cell[    2847] = 32'h0;  // 32'h7a043072;
    ram_cell[    2848] = 32'h0;  // 32'h6b0e08d1;
    ram_cell[    2849] = 32'h0;  // 32'hc68e46db;
    ram_cell[    2850] = 32'h0;  // 32'h67e3b00f;
    ram_cell[    2851] = 32'h0;  // 32'h5234cc32;
    ram_cell[    2852] = 32'h0;  // 32'h22928c05;
    ram_cell[    2853] = 32'h0;  // 32'h174615fa;
    ram_cell[    2854] = 32'h0;  // 32'hea951711;
    ram_cell[    2855] = 32'h0;  // 32'h68709947;
    ram_cell[    2856] = 32'h0;  // 32'h9ceff50e;
    ram_cell[    2857] = 32'h0;  // 32'hb777cd05;
    ram_cell[    2858] = 32'h0;  // 32'hafddd8f3;
    ram_cell[    2859] = 32'h0;  // 32'h1302baa2;
    ram_cell[    2860] = 32'h0;  // 32'hfcdd0215;
    ram_cell[    2861] = 32'h0;  // 32'h45c81a88;
    ram_cell[    2862] = 32'h0;  // 32'h583db18e;
    ram_cell[    2863] = 32'h0;  // 32'hba798273;
    ram_cell[    2864] = 32'h0;  // 32'haf2b2597;
    ram_cell[    2865] = 32'h0;  // 32'hbee30fa7;
    ram_cell[    2866] = 32'h0;  // 32'h174256d9;
    ram_cell[    2867] = 32'h0;  // 32'h9bfb6dc6;
    ram_cell[    2868] = 32'h0;  // 32'hdb144564;
    ram_cell[    2869] = 32'h0;  // 32'h8af7c5a3;
    ram_cell[    2870] = 32'h0;  // 32'h1dafb539;
    ram_cell[    2871] = 32'h0;  // 32'h406b27a0;
    ram_cell[    2872] = 32'h0;  // 32'h7f6e1ee9;
    ram_cell[    2873] = 32'h0;  // 32'hca836ea9;
    ram_cell[    2874] = 32'h0;  // 32'h8240c2c6;
    ram_cell[    2875] = 32'h0;  // 32'hc6a4613c;
    ram_cell[    2876] = 32'h0;  // 32'hb9fc1808;
    ram_cell[    2877] = 32'h0;  // 32'hc11ec521;
    ram_cell[    2878] = 32'h0;  // 32'h4265645a;
    ram_cell[    2879] = 32'h0;  // 32'hcdbf24fe;
    ram_cell[    2880] = 32'h0;  // 32'h2c36a03d;
    ram_cell[    2881] = 32'h0;  // 32'h0236a2fc;
    ram_cell[    2882] = 32'h0;  // 32'h7f7fdff5;
    ram_cell[    2883] = 32'h0;  // 32'hbf02b292;
    ram_cell[    2884] = 32'h0;  // 32'hbf8f99c0;
    ram_cell[    2885] = 32'h0;  // 32'hf27e9e02;
    ram_cell[    2886] = 32'h0;  // 32'h0cc8efca;
    ram_cell[    2887] = 32'h0;  // 32'ha8e9f971;
    ram_cell[    2888] = 32'h0;  // 32'h0c422293;
    ram_cell[    2889] = 32'h0;  // 32'h3b52e193;
    ram_cell[    2890] = 32'h0;  // 32'h1b8944d7;
    ram_cell[    2891] = 32'h0;  // 32'hc2566723;
    ram_cell[    2892] = 32'h0;  // 32'h93266288;
    ram_cell[    2893] = 32'h0;  // 32'h99ff2240;
    ram_cell[    2894] = 32'h0;  // 32'h5a3b22dc;
    ram_cell[    2895] = 32'h0;  // 32'h62bc72ca;
    ram_cell[    2896] = 32'h0;  // 32'h549e7e9d;
    ram_cell[    2897] = 32'h0;  // 32'h61636d05;
    ram_cell[    2898] = 32'h0;  // 32'hb93f93f4;
    ram_cell[    2899] = 32'h0;  // 32'hac647c9d;
    ram_cell[    2900] = 32'h0;  // 32'hea869156;
    ram_cell[    2901] = 32'h0;  // 32'h6faba347;
    ram_cell[    2902] = 32'h0;  // 32'h18e0d056;
    ram_cell[    2903] = 32'h0;  // 32'hce6afce2;
    ram_cell[    2904] = 32'h0;  // 32'hd6e8f874;
    ram_cell[    2905] = 32'h0;  // 32'ha8751912;
    ram_cell[    2906] = 32'h0;  // 32'hd92ea72d;
    ram_cell[    2907] = 32'h0;  // 32'he105157f;
    ram_cell[    2908] = 32'h0;  // 32'h29666583;
    ram_cell[    2909] = 32'h0;  // 32'hfce22193;
    ram_cell[    2910] = 32'h0;  // 32'h83c3bef7;
    ram_cell[    2911] = 32'h0;  // 32'h9a20e468;
    ram_cell[    2912] = 32'h0;  // 32'h51f0788e;
    ram_cell[    2913] = 32'h0;  // 32'heefb256a;
    ram_cell[    2914] = 32'h0;  // 32'h6dbfb505;
    ram_cell[    2915] = 32'h0;  // 32'had2f50ff;
    ram_cell[    2916] = 32'h0;  // 32'hb1a119b5;
    ram_cell[    2917] = 32'h0;  // 32'ha5c828c1;
    ram_cell[    2918] = 32'h0;  // 32'h15868f45;
    ram_cell[    2919] = 32'h0;  // 32'h2baf8783;
    ram_cell[    2920] = 32'h0;  // 32'h38f217cb;
    ram_cell[    2921] = 32'h0;  // 32'h6c5fbbc8;
    ram_cell[    2922] = 32'h0;  // 32'h0364042f;
    ram_cell[    2923] = 32'h0;  // 32'h52a9c573;
    ram_cell[    2924] = 32'h0;  // 32'he5142bdd;
    ram_cell[    2925] = 32'h0;  // 32'h09a4d58b;
    ram_cell[    2926] = 32'h0;  // 32'h40ad4232;
    ram_cell[    2927] = 32'h0;  // 32'hf063bf3f;
    ram_cell[    2928] = 32'h0;  // 32'h407bd4ec;
    ram_cell[    2929] = 32'h0;  // 32'h23868214;
    ram_cell[    2930] = 32'h0;  // 32'h605b5d35;
    ram_cell[    2931] = 32'h0;  // 32'h8feb0f8f;
    ram_cell[    2932] = 32'h0;  // 32'h3d87e10b;
    ram_cell[    2933] = 32'h0;  // 32'h78cdb273;
    ram_cell[    2934] = 32'h0;  // 32'h1da73a28;
    ram_cell[    2935] = 32'h0;  // 32'hb83be7b5;
    ram_cell[    2936] = 32'h0;  // 32'h20c30026;
    ram_cell[    2937] = 32'h0;  // 32'h7bd61168;
    ram_cell[    2938] = 32'h0;  // 32'hbea55ee6;
    ram_cell[    2939] = 32'h0;  // 32'h3f2f1eda;
    ram_cell[    2940] = 32'h0;  // 32'hc2598ee8;
    ram_cell[    2941] = 32'h0;  // 32'h4fd69c43;
    ram_cell[    2942] = 32'h0;  // 32'h0fdc5320;
    ram_cell[    2943] = 32'h0;  // 32'h3d6baa17;
    ram_cell[    2944] = 32'h0;  // 32'h1478fa7d;
    ram_cell[    2945] = 32'h0;  // 32'h1f494af5;
    ram_cell[    2946] = 32'h0;  // 32'h1a487231;
    ram_cell[    2947] = 32'h0;  // 32'h3e0e40ad;
    ram_cell[    2948] = 32'h0;  // 32'h1eb521da;
    ram_cell[    2949] = 32'h0;  // 32'h6b2ed229;
    ram_cell[    2950] = 32'h0;  // 32'h0d55b3ed;
    ram_cell[    2951] = 32'h0;  // 32'he133fc24;
    ram_cell[    2952] = 32'h0;  // 32'he69ac5da;
    ram_cell[    2953] = 32'h0;  // 32'ha7a5589a;
    ram_cell[    2954] = 32'h0;  // 32'h0b77efb6;
    ram_cell[    2955] = 32'h0;  // 32'hbde0ac7f;
    ram_cell[    2956] = 32'h0;  // 32'h484193b7;
    ram_cell[    2957] = 32'h0;  // 32'h02618ab4;
    ram_cell[    2958] = 32'h0;  // 32'h2742ba60;
    ram_cell[    2959] = 32'h0;  // 32'h0d947070;
    ram_cell[    2960] = 32'h0;  // 32'had809feb;
    ram_cell[    2961] = 32'h0;  // 32'hb0b5427d;
    ram_cell[    2962] = 32'h0;  // 32'hd83516cc;
    ram_cell[    2963] = 32'h0;  // 32'hd24c2b3a;
    ram_cell[    2964] = 32'h0;  // 32'h90a1f585;
    ram_cell[    2965] = 32'h0;  // 32'h07d33daf;
    ram_cell[    2966] = 32'h0;  // 32'h28a87673;
    ram_cell[    2967] = 32'h0;  // 32'h15d85229;
    ram_cell[    2968] = 32'h0;  // 32'h37e7267e;
    ram_cell[    2969] = 32'h0;  // 32'hd5044752;
    ram_cell[    2970] = 32'h0;  // 32'he8164afb;
    ram_cell[    2971] = 32'h0;  // 32'h9eb8fc30;
    ram_cell[    2972] = 32'h0;  // 32'hdb87c14a;
    ram_cell[    2973] = 32'h0;  // 32'h871c471a;
    ram_cell[    2974] = 32'h0;  // 32'h1d96c371;
    ram_cell[    2975] = 32'h0;  // 32'h35dfe9b9;
    ram_cell[    2976] = 32'h0;  // 32'h78d7f582;
    ram_cell[    2977] = 32'h0;  // 32'h4c9386ee;
    ram_cell[    2978] = 32'h0;  // 32'h6efb609d;
    ram_cell[    2979] = 32'h0;  // 32'h28cc554a;
    ram_cell[    2980] = 32'h0;  // 32'h7d42569c;
    ram_cell[    2981] = 32'h0;  // 32'h9e22fa4a;
    ram_cell[    2982] = 32'h0;  // 32'h763ec523;
    ram_cell[    2983] = 32'h0;  // 32'hd069b8e9;
    ram_cell[    2984] = 32'h0;  // 32'h9b256a13;
    ram_cell[    2985] = 32'h0;  // 32'h758fb4ff;
    ram_cell[    2986] = 32'h0;  // 32'h515779d3;
    ram_cell[    2987] = 32'h0;  // 32'h8760f0f2;
    ram_cell[    2988] = 32'h0;  // 32'hb9228a04;
    ram_cell[    2989] = 32'h0;  // 32'h6cb58a8f;
    ram_cell[    2990] = 32'h0;  // 32'he01e6f7d;
    ram_cell[    2991] = 32'h0;  // 32'h851cc4da;
    ram_cell[    2992] = 32'h0;  // 32'h10b45aa7;
    ram_cell[    2993] = 32'h0;  // 32'h300f8eda;
    ram_cell[    2994] = 32'h0;  // 32'hc59028e3;
    ram_cell[    2995] = 32'h0;  // 32'h9ba58f66;
    ram_cell[    2996] = 32'h0;  // 32'h31041265;
    ram_cell[    2997] = 32'h0;  // 32'ha9262af4;
    ram_cell[    2998] = 32'h0;  // 32'h9ad007ac;
    ram_cell[    2999] = 32'h0;  // 32'h9783011f;
    ram_cell[    3000] = 32'h0;  // 32'h6c009b2a;
    ram_cell[    3001] = 32'h0;  // 32'h5dda7f4c;
    ram_cell[    3002] = 32'h0;  // 32'h73c77735;
    ram_cell[    3003] = 32'h0;  // 32'hc1277ccb;
    ram_cell[    3004] = 32'h0;  // 32'h3b145c53;
    ram_cell[    3005] = 32'h0;  // 32'h7a3194ca;
    ram_cell[    3006] = 32'h0;  // 32'hda5d3c1d;
    ram_cell[    3007] = 32'h0;  // 32'h8fd51b58;
    ram_cell[    3008] = 32'h0;  // 32'h488660a1;
    ram_cell[    3009] = 32'h0;  // 32'h714901f6;
    ram_cell[    3010] = 32'h0;  // 32'h411b4c8a;
    ram_cell[    3011] = 32'h0;  // 32'h23196345;
    ram_cell[    3012] = 32'h0;  // 32'h1cdb1384;
    ram_cell[    3013] = 32'h0;  // 32'hdafa44e1;
    ram_cell[    3014] = 32'h0;  // 32'h691393ea;
    ram_cell[    3015] = 32'h0;  // 32'h090aa029;
    ram_cell[    3016] = 32'h0;  // 32'h5be76f4c;
    ram_cell[    3017] = 32'h0;  // 32'h4a3dded0;
    ram_cell[    3018] = 32'h0;  // 32'he6c3876b;
    ram_cell[    3019] = 32'h0;  // 32'h0737a4db;
    ram_cell[    3020] = 32'h0;  // 32'h8c660119;
    ram_cell[    3021] = 32'h0;  // 32'hb1286ccc;
    ram_cell[    3022] = 32'h0;  // 32'h18e12f79;
    ram_cell[    3023] = 32'h0;  // 32'h9aebe130;
    ram_cell[    3024] = 32'h0;  // 32'hc66bd3ce;
    ram_cell[    3025] = 32'h0;  // 32'h81c8c9d6;
    ram_cell[    3026] = 32'h0;  // 32'h3b5dcd20;
    ram_cell[    3027] = 32'h0;  // 32'h2d3772d3;
    ram_cell[    3028] = 32'h0;  // 32'h9a878a6e;
    ram_cell[    3029] = 32'h0;  // 32'h1bb36a57;
    ram_cell[    3030] = 32'h0;  // 32'hdd09da2e;
    ram_cell[    3031] = 32'h0;  // 32'hcc757df2;
    ram_cell[    3032] = 32'h0;  // 32'hc90434b5;
    ram_cell[    3033] = 32'h0;  // 32'hcba85c5b;
    ram_cell[    3034] = 32'h0;  // 32'h7665c3cb;
    ram_cell[    3035] = 32'h0;  // 32'hf2ed6137;
    ram_cell[    3036] = 32'h0;  // 32'h4c611db2;
    ram_cell[    3037] = 32'h0;  // 32'hc187ac07;
    ram_cell[    3038] = 32'h0;  // 32'h5ed5dbd6;
    ram_cell[    3039] = 32'h0;  // 32'h3349021c;
    ram_cell[    3040] = 32'h0;  // 32'h6a51e8d7;
    ram_cell[    3041] = 32'h0;  // 32'hd3cedaee;
    ram_cell[    3042] = 32'h0;  // 32'ha0881272;
    ram_cell[    3043] = 32'h0;  // 32'h15e389fc;
    ram_cell[    3044] = 32'h0;  // 32'hb359e11f;
    ram_cell[    3045] = 32'h0;  // 32'h5c890712;
    ram_cell[    3046] = 32'h0;  // 32'he2467849;
    ram_cell[    3047] = 32'h0;  // 32'h8c3456f8;
    ram_cell[    3048] = 32'h0;  // 32'hfb527c50;
    ram_cell[    3049] = 32'h0;  // 32'hac21b4ef;
    ram_cell[    3050] = 32'h0;  // 32'h27071deb;
    ram_cell[    3051] = 32'h0;  // 32'h912c3f1a;
    ram_cell[    3052] = 32'h0;  // 32'h261db59a;
    ram_cell[    3053] = 32'h0;  // 32'h5ad65973;
    ram_cell[    3054] = 32'h0;  // 32'h2d6cc44e;
    ram_cell[    3055] = 32'h0;  // 32'ha735aab3;
    ram_cell[    3056] = 32'h0;  // 32'h6de366fc;
    ram_cell[    3057] = 32'h0;  // 32'h9a45b822;
    ram_cell[    3058] = 32'h0;  // 32'ha4e217e2;
    ram_cell[    3059] = 32'h0;  // 32'ha3770811;
    ram_cell[    3060] = 32'h0;  // 32'ha109aa9d;
    ram_cell[    3061] = 32'h0;  // 32'hdc582ad9;
    ram_cell[    3062] = 32'h0;  // 32'hadd1bdb3;
    ram_cell[    3063] = 32'h0;  // 32'h39f3ac16;
    ram_cell[    3064] = 32'h0;  // 32'h8a189aeb;
    ram_cell[    3065] = 32'h0;  // 32'hde235ec1;
    ram_cell[    3066] = 32'h0;  // 32'h578e219f;
    ram_cell[    3067] = 32'h0;  // 32'hf784e813;
    ram_cell[    3068] = 32'h0;  // 32'h98c32e2f;
    ram_cell[    3069] = 32'h0;  // 32'h69d9b82b;
    ram_cell[    3070] = 32'h0;  // 32'h2f9d7b1e;
    ram_cell[    3071] = 32'h0;  // 32'h9e54eda7;
    ram_cell[    3072] = 32'h0;  // 32'h594dd87a;
    ram_cell[    3073] = 32'h0;  // 32'hd0ad6ac4;
    ram_cell[    3074] = 32'h0;  // 32'h8d593127;
    ram_cell[    3075] = 32'h0;  // 32'h43adc0df;
    ram_cell[    3076] = 32'h0;  // 32'hb9fe67d5;
    ram_cell[    3077] = 32'h0;  // 32'h8a9eb0a9;
    ram_cell[    3078] = 32'h0;  // 32'h44fff159;
    ram_cell[    3079] = 32'h0;  // 32'h1a98f4e8;
    ram_cell[    3080] = 32'h0;  // 32'h2bf522f6;
    ram_cell[    3081] = 32'h0;  // 32'hf41b2197;
    ram_cell[    3082] = 32'h0;  // 32'h8bb75cb1;
    ram_cell[    3083] = 32'h0;  // 32'hdb3cf15a;
    ram_cell[    3084] = 32'h0;  // 32'h37c9e264;
    ram_cell[    3085] = 32'h0;  // 32'hc4e37333;
    ram_cell[    3086] = 32'h0;  // 32'hc7f23c24;
    ram_cell[    3087] = 32'h0;  // 32'hc8ffea3c;
    ram_cell[    3088] = 32'h0;  // 32'ha2f0758b;
    ram_cell[    3089] = 32'h0;  // 32'h0e8e98e6;
    ram_cell[    3090] = 32'h0;  // 32'h58132ebc;
    ram_cell[    3091] = 32'h0;  // 32'h35ffc47d;
    ram_cell[    3092] = 32'h0;  // 32'hbe8adeec;
    ram_cell[    3093] = 32'h0;  // 32'h022ee573;
    ram_cell[    3094] = 32'h0;  // 32'h4893df55;
    ram_cell[    3095] = 32'h0;  // 32'h44670f9f;
    ram_cell[    3096] = 32'h0;  // 32'hcbe181ed;
    ram_cell[    3097] = 32'h0;  // 32'h74c02fd7;
    ram_cell[    3098] = 32'h0;  // 32'ha8a8adda;
    ram_cell[    3099] = 32'h0;  // 32'h3bbfdf67;
    ram_cell[    3100] = 32'h0;  // 32'h532b28d9;
    ram_cell[    3101] = 32'h0;  // 32'h206a64e2;
    ram_cell[    3102] = 32'h0;  // 32'h9d954b72;
    ram_cell[    3103] = 32'h0;  // 32'hccdd3402;
    ram_cell[    3104] = 32'h0;  // 32'h02950755;
    ram_cell[    3105] = 32'h0;  // 32'h60386d6e;
    ram_cell[    3106] = 32'h0;  // 32'h7ce2b62b;
    ram_cell[    3107] = 32'h0;  // 32'hcb80b989;
    ram_cell[    3108] = 32'h0;  // 32'h13edef93;
    ram_cell[    3109] = 32'h0;  // 32'hcd6c78c2;
    ram_cell[    3110] = 32'h0;  // 32'h380c336b;
    ram_cell[    3111] = 32'h0;  // 32'h827a5759;
    ram_cell[    3112] = 32'h0;  // 32'h43d9be58;
    ram_cell[    3113] = 32'h0;  // 32'h1ae81b58;
    ram_cell[    3114] = 32'h0;  // 32'he5a90f27;
    ram_cell[    3115] = 32'h0;  // 32'hdd4707e6;
    ram_cell[    3116] = 32'h0;  // 32'hfd6d0e37;
    ram_cell[    3117] = 32'h0;  // 32'hf8fefaf6;
    ram_cell[    3118] = 32'h0;  // 32'hc1ab87da;
    ram_cell[    3119] = 32'h0;  // 32'hb088297b;
    ram_cell[    3120] = 32'h0;  // 32'h5bf0a188;
    ram_cell[    3121] = 32'h0;  // 32'h72d6f085;
    ram_cell[    3122] = 32'h0;  // 32'h5237b7e9;
    ram_cell[    3123] = 32'h0;  // 32'h7c4f7bd2;
    ram_cell[    3124] = 32'h0;  // 32'h1311decd;
    ram_cell[    3125] = 32'h0;  // 32'ha161684a;
    ram_cell[    3126] = 32'h0;  // 32'hd6b58b46;
    ram_cell[    3127] = 32'h0;  // 32'hd0e94b2b;
    ram_cell[    3128] = 32'h0;  // 32'h53226c95;
    ram_cell[    3129] = 32'h0;  // 32'h1bca2199;
    ram_cell[    3130] = 32'h0;  // 32'hcd46e533;
    ram_cell[    3131] = 32'h0;  // 32'h6e40ee5e;
    ram_cell[    3132] = 32'h0;  // 32'h2ba3ba00;
    ram_cell[    3133] = 32'h0;  // 32'h13e28268;
    ram_cell[    3134] = 32'h0;  // 32'hc098563d;
    ram_cell[    3135] = 32'h0;  // 32'hbf67d509;
    ram_cell[    3136] = 32'h0;  // 32'h8532cc9d;
    ram_cell[    3137] = 32'h0;  // 32'h4942b291;
    ram_cell[    3138] = 32'h0;  // 32'hb3028ffc;
    ram_cell[    3139] = 32'h0;  // 32'ha01f6783;
    ram_cell[    3140] = 32'h0;  // 32'hef246a8d;
    ram_cell[    3141] = 32'h0;  // 32'h1fe2dcaf;
    ram_cell[    3142] = 32'h0;  // 32'h4e1eba76;
    ram_cell[    3143] = 32'h0;  // 32'hef9844ee;
    ram_cell[    3144] = 32'h0;  // 32'h1356d969;
    ram_cell[    3145] = 32'h0;  // 32'h85a722fa;
    ram_cell[    3146] = 32'h0;  // 32'he996ff3e;
    ram_cell[    3147] = 32'h0;  // 32'h13b4c18d;
    ram_cell[    3148] = 32'h0;  // 32'h5db2762c;
    ram_cell[    3149] = 32'h0;  // 32'h85f4ae87;
    ram_cell[    3150] = 32'h0;  // 32'h81e747bd;
    ram_cell[    3151] = 32'h0;  // 32'h6a339a61;
    ram_cell[    3152] = 32'h0;  // 32'h1a463cca;
    ram_cell[    3153] = 32'h0;  // 32'hdf325d35;
    ram_cell[    3154] = 32'h0;  // 32'h61d2bb5c;
    ram_cell[    3155] = 32'h0;  // 32'h29d1ef67;
    ram_cell[    3156] = 32'h0;  // 32'h7eb2313e;
    ram_cell[    3157] = 32'h0;  // 32'hfe37b0bc;
    ram_cell[    3158] = 32'h0;  // 32'hcd1d9129;
    ram_cell[    3159] = 32'h0;  // 32'h256982f9;
    ram_cell[    3160] = 32'h0;  // 32'h0e43382a;
    ram_cell[    3161] = 32'h0;  // 32'h4b9b6f6f;
    ram_cell[    3162] = 32'h0;  // 32'h0a5b1891;
    ram_cell[    3163] = 32'h0;  // 32'h58cf4d47;
    ram_cell[    3164] = 32'h0;  // 32'he5d1f172;
    ram_cell[    3165] = 32'h0;  // 32'h9b5a581f;
    ram_cell[    3166] = 32'h0;  // 32'h34a552b9;
    ram_cell[    3167] = 32'h0;  // 32'hf00e1727;
    ram_cell[    3168] = 32'h0;  // 32'hb315f75f;
    ram_cell[    3169] = 32'h0;  // 32'hd832068f;
    ram_cell[    3170] = 32'h0;  // 32'hca1b17d3;
    ram_cell[    3171] = 32'h0;  // 32'ha4159dfe;
    ram_cell[    3172] = 32'h0;  // 32'h90fea072;
    ram_cell[    3173] = 32'h0;  // 32'h51a9d5f5;
    ram_cell[    3174] = 32'h0;  // 32'h6898cc24;
    ram_cell[    3175] = 32'h0;  // 32'h4b57a61e;
    ram_cell[    3176] = 32'h0;  // 32'h213dba08;
    ram_cell[    3177] = 32'h0;  // 32'hb70f027b;
    ram_cell[    3178] = 32'h0;  // 32'h8981eb6e;
    ram_cell[    3179] = 32'h0;  // 32'h3dfba68e;
    ram_cell[    3180] = 32'h0;  // 32'h3908f6d3;
    ram_cell[    3181] = 32'h0;  // 32'h4b7e7d30;
    ram_cell[    3182] = 32'h0;  // 32'h403df3ba;
    ram_cell[    3183] = 32'h0;  // 32'h26bdfb04;
    ram_cell[    3184] = 32'h0;  // 32'h5f495c7a;
    ram_cell[    3185] = 32'h0;  // 32'hafa1d36f;
    ram_cell[    3186] = 32'h0;  // 32'h36e6b3da;
    ram_cell[    3187] = 32'h0;  // 32'h5c081060;
    ram_cell[    3188] = 32'h0;  // 32'h773473ec;
    ram_cell[    3189] = 32'h0;  // 32'h578a801e;
    ram_cell[    3190] = 32'h0;  // 32'h7813620e;
    ram_cell[    3191] = 32'h0;  // 32'h9cbc8e8d;
    ram_cell[    3192] = 32'h0;  // 32'h2f246d7c;
    ram_cell[    3193] = 32'h0;  // 32'h34f2d438;
    ram_cell[    3194] = 32'h0;  // 32'hffa45ee4;
    ram_cell[    3195] = 32'h0;  // 32'hbe22f80a;
    ram_cell[    3196] = 32'h0;  // 32'h1f2d5044;
    ram_cell[    3197] = 32'h0;  // 32'h534aa3e6;
    ram_cell[    3198] = 32'h0;  // 32'hea1691bf;
    ram_cell[    3199] = 32'h0;  // 32'h20e52053;
    ram_cell[    3200] = 32'h0;  // 32'h714f66d9;
    ram_cell[    3201] = 32'h0;  // 32'hb4c3715b;
    ram_cell[    3202] = 32'h0;  // 32'h98ce3185;
    ram_cell[    3203] = 32'h0;  // 32'h88e74352;
    ram_cell[    3204] = 32'h0;  // 32'hc3eb248b;
    ram_cell[    3205] = 32'h0;  // 32'hd2325e1a;
    ram_cell[    3206] = 32'h0;  // 32'hbbebd434;
    ram_cell[    3207] = 32'h0;  // 32'h8c7f4fbb;
    ram_cell[    3208] = 32'h0;  // 32'h6a56d603;
    ram_cell[    3209] = 32'h0;  // 32'hc56f8697;
    ram_cell[    3210] = 32'h0;  // 32'hbdd80539;
    ram_cell[    3211] = 32'h0;  // 32'hc837a50a;
    ram_cell[    3212] = 32'h0;  // 32'hff73311f;
    ram_cell[    3213] = 32'h0;  // 32'hab060618;
    ram_cell[    3214] = 32'h0;  // 32'he4344592;
    ram_cell[    3215] = 32'h0;  // 32'hc8782bab;
    ram_cell[    3216] = 32'h0;  // 32'h22ee93c6;
    ram_cell[    3217] = 32'h0;  // 32'h35ce9f7c;
    ram_cell[    3218] = 32'h0;  // 32'h005d3d4b;
    ram_cell[    3219] = 32'h0;  // 32'hd205f2bd;
    ram_cell[    3220] = 32'h0;  // 32'hbfbc7522;
    ram_cell[    3221] = 32'h0;  // 32'ha1d1ea4d;
    ram_cell[    3222] = 32'h0;  // 32'h3ed03ac9;
    ram_cell[    3223] = 32'h0;  // 32'hc0844b53;
    ram_cell[    3224] = 32'h0;  // 32'hb2b144e7;
    ram_cell[    3225] = 32'h0;  // 32'hffd214d1;
    ram_cell[    3226] = 32'h0;  // 32'ha39c8c95;
    ram_cell[    3227] = 32'h0;  // 32'h96cd3d1d;
    ram_cell[    3228] = 32'h0;  // 32'h1c163d4b;
    ram_cell[    3229] = 32'h0;  // 32'hd241228a;
    ram_cell[    3230] = 32'h0;  // 32'ha11e8809;
    ram_cell[    3231] = 32'h0;  // 32'h8e01b789;
    ram_cell[    3232] = 32'h0;  // 32'he7ee4c34;
    ram_cell[    3233] = 32'h0;  // 32'h596e1863;
    ram_cell[    3234] = 32'h0;  // 32'h002aaa98;
    ram_cell[    3235] = 32'h0;  // 32'h3425ee09;
    ram_cell[    3236] = 32'h0;  // 32'h9d0e414a;
    ram_cell[    3237] = 32'h0;  // 32'heed5e791;
    ram_cell[    3238] = 32'h0;  // 32'hd0030255;
    ram_cell[    3239] = 32'h0;  // 32'ha4c42bf1;
    ram_cell[    3240] = 32'h0;  // 32'h68b0fc19;
    ram_cell[    3241] = 32'h0;  // 32'hdab662b0;
    ram_cell[    3242] = 32'h0;  // 32'h3eab7b7d;
    ram_cell[    3243] = 32'h0;  // 32'h22ab1050;
    ram_cell[    3244] = 32'h0;  // 32'h9ec27808;
    ram_cell[    3245] = 32'h0;  // 32'h40312a9f;
    ram_cell[    3246] = 32'h0;  // 32'h275303cd;
    ram_cell[    3247] = 32'h0;  // 32'ha28423b2;
    ram_cell[    3248] = 32'h0;  // 32'h12641f48;
    ram_cell[    3249] = 32'h0;  // 32'hdbca7620;
    ram_cell[    3250] = 32'h0;  // 32'h92ec302c;
    ram_cell[    3251] = 32'h0;  // 32'hf555c2eb;
    ram_cell[    3252] = 32'h0;  // 32'hf9ad090c;
    ram_cell[    3253] = 32'h0;  // 32'h40220b4d;
    ram_cell[    3254] = 32'h0;  // 32'ha6e2fa76;
    ram_cell[    3255] = 32'h0;  // 32'h0654629e;
    ram_cell[    3256] = 32'h0;  // 32'hd80650a9;
    ram_cell[    3257] = 32'h0;  // 32'h01061d96;
    ram_cell[    3258] = 32'h0;  // 32'h8ca8a9c9;
    ram_cell[    3259] = 32'h0;  // 32'h8b3d58a2;
    ram_cell[    3260] = 32'h0;  // 32'he789ac97;
    ram_cell[    3261] = 32'h0;  // 32'heb8bf2d6;
    ram_cell[    3262] = 32'h0;  // 32'h7200480e;
    ram_cell[    3263] = 32'h0;  // 32'h8ac72788;
    ram_cell[    3264] = 32'h0;  // 32'he4d90b43;
    ram_cell[    3265] = 32'h0;  // 32'h476e7fd3;
    ram_cell[    3266] = 32'h0;  // 32'ha24d4649;
    ram_cell[    3267] = 32'h0;  // 32'hace2dca1;
    ram_cell[    3268] = 32'h0;  // 32'h301e8a17;
    ram_cell[    3269] = 32'h0;  // 32'h2c1d15f2;
    ram_cell[    3270] = 32'h0;  // 32'h63ad8f64;
    ram_cell[    3271] = 32'h0;  // 32'heb16331c;
    ram_cell[    3272] = 32'h0;  // 32'h215d5326;
    ram_cell[    3273] = 32'h0;  // 32'h52f2398a;
    ram_cell[    3274] = 32'h0;  // 32'h40c5e491;
    ram_cell[    3275] = 32'h0;  // 32'h6ff88fa9;
    ram_cell[    3276] = 32'h0;  // 32'hc6afe2ac;
    ram_cell[    3277] = 32'h0;  // 32'h05d31946;
    ram_cell[    3278] = 32'h0;  // 32'ha461129e;
    ram_cell[    3279] = 32'h0;  // 32'h6ee83269;
    ram_cell[    3280] = 32'h0;  // 32'hb21691ee;
    ram_cell[    3281] = 32'h0;  // 32'ha6aa036d;
    ram_cell[    3282] = 32'h0;  // 32'habf70f5e;
    ram_cell[    3283] = 32'h0;  // 32'hafa3d5c5;
    ram_cell[    3284] = 32'h0;  // 32'h37849eaa;
    ram_cell[    3285] = 32'h0;  // 32'h2ff3ea68;
    ram_cell[    3286] = 32'h0;  // 32'hb5fb65b5;
    ram_cell[    3287] = 32'h0;  // 32'hecbcc0ad;
    ram_cell[    3288] = 32'h0;  // 32'hf5c3fcb3;
    ram_cell[    3289] = 32'h0;  // 32'h4deccf37;
    ram_cell[    3290] = 32'h0;  // 32'h86006af3;
    ram_cell[    3291] = 32'h0;  // 32'hf660c40d;
    ram_cell[    3292] = 32'h0;  // 32'hb327f8a4;
    ram_cell[    3293] = 32'h0;  // 32'h320564df;
    ram_cell[    3294] = 32'h0;  // 32'hea9f7509;
    ram_cell[    3295] = 32'h0;  // 32'h23b74386;
    ram_cell[    3296] = 32'h0;  // 32'hfcdbc090;
    ram_cell[    3297] = 32'h0;  // 32'h0f22aac8;
    ram_cell[    3298] = 32'h0;  // 32'h92b4f9cf;
    ram_cell[    3299] = 32'h0;  // 32'h97a50821;
    ram_cell[    3300] = 32'h0;  // 32'hc9762add;
    ram_cell[    3301] = 32'h0;  // 32'hd8686bc0;
    ram_cell[    3302] = 32'h0;  // 32'hf327f9d2;
    ram_cell[    3303] = 32'h0;  // 32'he6c00f16;
    ram_cell[    3304] = 32'h0;  // 32'heeaa5b2c;
    ram_cell[    3305] = 32'h0;  // 32'hd81fc9a6;
    ram_cell[    3306] = 32'h0;  // 32'h9cf49cc4;
    ram_cell[    3307] = 32'h0;  // 32'h0f0bc6c9;
    ram_cell[    3308] = 32'h0;  // 32'h7106ee49;
    ram_cell[    3309] = 32'h0;  // 32'h99f38a93;
    ram_cell[    3310] = 32'h0;  // 32'h66a17b3c;
    ram_cell[    3311] = 32'h0;  // 32'h265495ef;
    ram_cell[    3312] = 32'h0;  // 32'h53849e04;
    ram_cell[    3313] = 32'h0;  // 32'ha5b7c95d;
    ram_cell[    3314] = 32'h0;  // 32'h2f34c970;
    ram_cell[    3315] = 32'h0;  // 32'hdb8fc456;
    ram_cell[    3316] = 32'h0;  // 32'h4837f13e;
    ram_cell[    3317] = 32'h0;  // 32'he5dc4346;
    ram_cell[    3318] = 32'h0;  // 32'h46eee521;
    ram_cell[    3319] = 32'h0;  // 32'h1ece1019;
    ram_cell[    3320] = 32'h0;  // 32'hc37efe1e;
    ram_cell[    3321] = 32'h0;  // 32'hbd9580ad;
    ram_cell[    3322] = 32'h0;  // 32'hf5463109;
    ram_cell[    3323] = 32'h0;  // 32'h5b77b002;
    ram_cell[    3324] = 32'h0;  // 32'ha7d2a5ca;
    ram_cell[    3325] = 32'h0;  // 32'h5088d288;
    ram_cell[    3326] = 32'h0;  // 32'h1b6d0b07;
    ram_cell[    3327] = 32'h0;  // 32'h231a21ac;
    ram_cell[    3328] = 32'h0;  // 32'h1d2a58eb;
    ram_cell[    3329] = 32'h0;  // 32'h98e458e3;
    ram_cell[    3330] = 32'h0;  // 32'h0f6db84e;
    ram_cell[    3331] = 32'h0;  // 32'h9dbfac6b;
    ram_cell[    3332] = 32'h0;  // 32'hdc6f17a9;
    ram_cell[    3333] = 32'h0;  // 32'h280c9161;
    ram_cell[    3334] = 32'h0;  // 32'h2e2f827c;
    ram_cell[    3335] = 32'h0;  // 32'h3e619fae;
    ram_cell[    3336] = 32'h0;  // 32'h0b05ebaa;
    ram_cell[    3337] = 32'h0;  // 32'h1f6fbf48;
    ram_cell[    3338] = 32'h0;  // 32'h1dcc3b49;
    ram_cell[    3339] = 32'h0;  // 32'h7998b3f0;
    ram_cell[    3340] = 32'h0;  // 32'h8d5ed578;
    ram_cell[    3341] = 32'h0;  // 32'h0dbefd9c;
    ram_cell[    3342] = 32'h0;  // 32'ha1e3694b;
    ram_cell[    3343] = 32'h0;  // 32'hbfb690d0;
    ram_cell[    3344] = 32'h0;  // 32'h53280c2b;
    ram_cell[    3345] = 32'h0;  // 32'he8895f9e;
    ram_cell[    3346] = 32'h0;  // 32'h2e64a65c;
    ram_cell[    3347] = 32'h0;  // 32'hf02c2b6c;
    ram_cell[    3348] = 32'h0;  // 32'h9946e2c6;
    ram_cell[    3349] = 32'h0;  // 32'h26d4c1ba;
    ram_cell[    3350] = 32'h0;  // 32'h86feba86;
    ram_cell[    3351] = 32'h0;  // 32'h0736966f;
    ram_cell[    3352] = 32'h0;  // 32'h6b7cd588;
    ram_cell[    3353] = 32'h0;  // 32'hb6174d30;
    ram_cell[    3354] = 32'h0;  // 32'h4244b089;
    ram_cell[    3355] = 32'h0;  // 32'h2c2cb5e9;
    ram_cell[    3356] = 32'h0;  // 32'h6de04b8c;
    ram_cell[    3357] = 32'h0;  // 32'h6c9af1a0;
    ram_cell[    3358] = 32'h0;  // 32'h213c7753;
    ram_cell[    3359] = 32'h0;  // 32'h16c1cfca;
    ram_cell[    3360] = 32'h0;  // 32'h768e41bc;
    ram_cell[    3361] = 32'h0;  // 32'h04777603;
    ram_cell[    3362] = 32'h0;  // 32'h8a499190;
    ram_cell[    3363] = 32'h0;  // 32'h534907ce;
    ram_cell[    3364] = 32'h0;  // 32'h9e9aefb0;
    ram_cell[    3365] = 32'h0;  // 32'h04ec8581;
    ram_cell[    3366] = 32'h0;  // 32'h73eded2b;
    ram_cell[    3367] = 32'h0;  // 32'h590f2c71;
    ram_cell[    3368] = 32'h0;  // 32'ha6544803;
    ram_cell[    3369] = 32'h0;  // 32'h90b0e24b;
    ram_cell[    3370] = 32'h0;  // 32'h47fc157b;
    ram_cell[    3371] = 32'h0;  // 32'haad2ceb9;
    ram_cell[    3372] = 32'h0;  // 32'ha28d31a0;
    ram_cell[    3373] = 32'h0;  // 32'h0fd77d78;
    ram_cell[    3374] = 32'h0;  // 32'hdb56bdb6;
    ram_cell[    3375] = 32'h0;  // 32'h67d047b7;
    ram_cell[    3376] = 32'h0;  // 32'hd8c5285d;
    ram_cell[    3377] = 32'h0;  // 32'had08550b;
    ram_cell[    3378] = 32'h0;  // 32'hf423e8a9;
    ram_cell[    3379] = 32'h0;  // 32'h8bf93141;
    ram_cell[    3380] = 32'h0;  // 32'h41c027b2;
    ram_cell[    3381] = 32'h0;  // 32'hfa23d337;
    ram_cell[    3382] = 32'h0;  // 32'hf72daffb;
    ram_cell[    3383] = 32'h0;  // 32'h59845d5f;
    ram_cell[    3384] = 32'h0;  // 32'hab66b36a;
    ram_cell[    3385] = 32'h0;  // 32'ha847f09c;
    ram_cell[    3386] = 32'h0;  // 32'h93c8bf4e;
    ram_cell[    3387] = 32'h0;  // 32'h61fcd76f;
    ram_cell[    3388] = 32'h0;  // 32'h55d44f9e;
    ram_cell[    3389] = 32'h0;  // 32'h8d9adbbc;
    ram_cell[    3390] = 32'h0;  // 32'hb9e1cdf3;
    ram_cell[    3391] = 32'h0;  // 32'h7c69a724;
    ram_cell[    3392] = 32'h0;  // 32'hb79c102a;
    ram_cell[    3393] = 32'h0;  // 32'h38a5d238;
    ram_cell[    3394] = 32'h0;  // 32'h35d2269c;
    ram_cell[    3395] = 32'h0;  // 32'hf96905af;
    ram_cell[    3396] = 32'h0;  // 32'h69e4c181;
    ram_cell[    3397] = 32'h0;  // 32'h081e2774;
    ram_cell[    3398] = 32'h0;  // 32'hd0feac1a;
    ram_cell[    3399] = 32'h0;  // 32'hb0f94c48;
    ram_cell[    3400] = 32'h0;  // 32'hf9a7a3ca;
    ram_cell[    3401] = 32'h0;  // 32'hf3878192;
    ram_cell[    3402] = 32'h0;  // 32'h70367598;
    ram_cell[    3403] = 32'h0;  // 32'hca6e67e6;
    ram_cell[    3404] = 32'h0;  // 32'h124ec489;
    ram_cell[    3405] = 32'h0;  // 32'hb2e45359;
    ram_cell[    3406] = 32'h0;  // 32'h9dca91e1;
    ram_cell[    3407] = 32'h0;  // 32'h36ee4795;
    ram_cell[    3408] = 32'h0;  // 32'h7d150302;
    ram_cell[    3409] = 32'h0;  // 32'h2a407393;
    ram_cell[    3410] = 32'h0;  // 32'h91a4ff43;
    ram_cell[    3411] = 32'h0;  // 32'h4ab7c0bc;
    ram_cell[    3412] = 32'h0;  // 32'h74469268;
    ram_cell[    3413] = 32'h0;  // 32'he96cdc7f;
    ram_cell[    3414] = 32'h0;  // 32'ha7d00969;
    ram_cell[    3415] = 32'h0;  // 32'hbceddc04;
    ram_cell[    3416] = 32'h0;  // 32'h3952a22b;
    ram_cell[    3417] = 32'h0;  // 32'h672142b9;
    ram_cell[    3418] = 32'h0;  // 32'ha547366f;
    ram_cell[    3419] = 32'h0;  // 32'hbbb5f452;
    ram_cell[    3420] = 32'h0;  // 32'h590d3df8;
    ram_cell[    3421] = 32'h0;  // 32'ha3dc1c35;
    ram_cell[    3422] = 32'h0;  // 32'hedf6bee4;
    ram_cell[    3423] = 32'h0;  // 32'h1ae32462;
    ram_cell[    3424] = 32'h0;  // 32'ha5c80ea6;
    ram_cell[    3425] = 32'h0;  // 32'h34daba94;
    ram_cell[    3426] = 32'h0;  // 32'hcde6f6fe;
    ram_cell[    3427] = 32'h0;  // 32'h150b3d34;
    ram_cell[    3428] = 32'h0;  // 32'he566e927;
    ram_cell[    3429] = 32'h0;  // 32'h8dfe5229;
    ram_cell[    3430] = 32'h0;  // 32'haf8f0d81;
    ram_cell[    3431] = 32'h0;  // 32'hd48deae3;
    ram_cell[    3432] = 32'h0;  // 32'h7f2f09bb;
    ram_cell[    3433] = 32'h0;  // 32'hbcbc4173;
    ram_cell[    3434] = 32'h0;  // 32'h05f2158b;
    ram_cell[    3435] = 32'h0;  // 32'h9e5e913c;
    ram_cell[    3436] = 32'h0;  // 32'h07c3543b;
    ram_cell[    3437] = 32'h0;  // 32'hb0099538;
    ram_cell[    3438] = 32'h0;  // 32'h977c3853;
    ram_cell[    3439] = 32'h0;  // 32'h9c09c69f;
    ram_cell[    3440] = 32'h0;  // 32'h2df96af6;
    ram_cell[    3441] = 32'h0;  // 32'he120524f;
    ram_cell[    3442] = 32'h0;  // 32'haa311b17;
    ram_cell[    3443] = 32'h0;  // 32'h33857c74;
    ram_cell[    3444] = 32'h0;  // 32'hfeaaa00e;
    ram_cell[    3445] = 32'h0;  // 32'h38301181;
    ram_cell[    3446] = 32'h0;  // 32'h30d90a3e;
    ram_cell[    3447] = 32'h0;  // 32'hf2834384;
    ram_cell[    3448] = 32'h0;  // 32'h6bf5195f;
    ram_cell[    3449] = 32'h0;  // 32'hc3577d22;
    ram_cell[    3450] = 32'h0;  // 32'h1fdab248;
    ram_cell[    3451] = 32'h0;  // 32'hf8c3e009;
    ram_cell[    3452] = 32'h0;  // 32'ha8117b2f;
    ram_cell[    3453] = 32'h0;  // 32'h29131a2a;
    ram_cell[    3454] = 32'h0;  // 32'h6cc4b8eb;
    ram_cell[    3455] = 32'h0;  // 32'h6f3d6b9e;
    ram_cell[    3456] = 32'h0;  // 32'h2ba59cb6;
    ram_cell[    3457] = 32'h0;  // 32'h46205790;
    ram_cell[    3458] = 32'h0;  // 32'h060d8c05;
    ram_cell[    3459] = 32'h0;  // 32'h1b670915;
    ram_cell[    3460] = 32'h0;  // 32'h31671f0b;
    ram_cell[    3461] = 32'h0;  // 32'he7329595;
    ram_cell[    3462] = 32'h0;  // 32'h5f8311fb;
    ram_cell[    3463] = 32'h0;  // 32'hbe4eeaab;
    ram_cell[    3464] = 32'h0;  // 32'h871cd85b;
    ram_cell[    3465] = 32'h0;  // 32'h53c40134;
    ram_cell[    3466] = 32'h0;  // 32'hb1dee1c5;
    ram_cell[    3467] = 32'h0;  // 32'hf3519101;
    ram_cell[    3468] = 32'h0;  // 32'h07380f6f;
    ram_cell[    3469] = 32'h0;  // 32'hcc7d65f9;
    ram_cell[    3470] = 32'h0;  // 32'hf976c935;
    ram_cell[    3471] = 32'h0;  // 32'hfffe28ea;
    ram_cell[    3472] = 32'h0;  // 32'h53293f14;
    ram_cell[    3473] = 32'h0;  // 32'hb53c6a1d;
    ram_cell[    3474] = 32'h0;  // 32'h09dbec6e;
    ram_cell[    3475] = 32'h0;  // 32'h7551f959;
    ram_cell[    3476] = 32'h0;  // 32'h2e832e0f;
    ram_cell[    3477] = 32'h0;  // 32'he6a7f784;
    ram_cell[    3478] = 32'h0;  // 32'h7fb7b427;
    ram_cell[    3479] = 32'h0;  // 32'he8ceca53;
    ram_cell[    3480] = 32'h0;  // 32'h119d7f2a;
    ram_cell[    3481] = 32'h0;  // 32'hee7eda1a;
    ram_cell[    3482] = 32'h0;  // 32'hb885bb93;
    ram_cell[    3483] = 32'h0;  // 32'hbd1c7b6c;
    ram_cell[    3484] = 32'h0;  // 32'hc19e257e;
    ram_cell[    3485] = 32'h0;  // 32'h538f4bb7;
    ram_cell[    3486] = 32'h0;  // 32'h27a90718;
    ram_cell[    3487] = 32'h0;  // 32'hbdc11e56;
    ram_cell[    3488] = 32'h0;  // 32'h88f6698f;
    ram_cell[    3489] = 32'h0;  // 32'h6fe4839f;
    ram_cell[    3490] = 32'h0;  // 32'h11df4b65;
    ram_cell[    3491] = 32'h0;  // 32'h719f5927;
    ram_cell[    3492] = 32'h0;  // 32'hfb0642d9;
    ram_cell[    3493] = 32'h0;  // 32'hafe40d16;
    ram_cell[    3494] = 32'h0;  // 32'h7de3a297;
    ram_cell[    3495] = 32'h0;  // 32'hbcabdbd1;
    ram_cell[    3496] = 32'h0;  // 32'h84ae34e6;
    ram_cell[    3497] = 32'h0;  // 32'h047c0e16;
    ram_cell[    3498] = 32'h0;  // 32'hb1f99110;
    ram_cell[    3499] = 32'h0;  // 32'h5a770855;
    ram_cell[    3500] = 32'h0;  // 32'h8d0c923e;
    ram_cell[    3501] = 32'h0;  // 32'h05584397;
    ram_cell[    3502] = 32'h0;  // 32'h5e5b2a37;
    ram_cell[    3503] = 32'h0;  // 32'h0bf6dc21;
    ram_cell[    3504] = 32'h0;  // 32'h0efc76da;
    ram_cell[    3505] = 32'h0;  // 32'h0c49673c;
    ram_cell[    3506] = 32'h0;  // 32'he559925d;
    ram_cell[    3507] = 32'h0;  // 32'h5687e2dc;
    ram_cell[    3508] = 32'h0;  // 32'h74f89270;
    ram_cell[    3509] = 32'h0;  // 32'hdb16f00a;
    ram_cell[    3510] = 32'h0;  // 32'hc1cec2db;
    ram_cell[    3511] = 32'h0;  // 32'h2fcf68c0;
    ram_cell[    3512] = 32'h0;  // 32'h61f318b0;
    ram_cell[    3513] = 32'h0;  // 32'he65d4e3d;
    ram_cell[    3514] = 32'h0;  // 32'h0813aa97;
    ram_cell[    3515] = 32'h0;  // 32'h5fc967b7;
    ram_cell[    3516] = 32'h0;  // 32'h21c71c9a;
    ram_cell[    3517] = 32'h0;  // 32'h6b162ee8;
    ram_cell[    3518] = 32'h0;  // 32'h89a90a91;
    ram_cell[    3519] = 32'h0;  // 32'hbf2d8504;
    ram_cell[    3520] = 32'h0;  // 32'hcdd730dd;
    ram_cell[    3521] = 32'h0;  // 32'h96ffaa4f;
    ram_cell[    3522] = 32'h0;  // 32'h6f99b720;
    ram_cell[    3523] = 32'h0;  // 32'hf5631a72;
    ram_cell[    3524] = 32'h0;  // 32'hf8098b53;
    ram_cell[    3525] = 32'h0;  // 32'hdd3b97f6;
    ram_cell[    3526] = 32'h0;  // 32'h0696963c;
    ram_cell[    3527] = 32'h0;  // 32'h3822791b;
    ram_cell[    3528] = 32'h0;  // 32'h06964800;
    ram_cell[    3529] = 32'h0;  // 32'h140c4e67;
    ram_cell[    3530] = 32'h0;  // 32'h0ad65ca1;
    ram_cell[    3531] = 32'h0;  // 32'h64865f57;
    ram_cell[    3532] = 32'h0;  // 32'ha3aa3616;
    ram_cell[    3533] = 32'h0;  // 32'h0f7febb1;
    ram_cell[    3534] = 32'h0;  // 32'h7497c537;
    ram_cell[    3535] = 32'h0;  // 32'h1d53bedc;
    ram_cell[    3536] = 32'h0;  // 32'h13d90835;
    ram_cell[    3537] = 32'h0;  // 32'h3253a143;
    ram_cell[    3538] = 32'h0;  // 32'h0a33a53d;
    ram_cell[    3539] = 32'h0;  // 32'hde2c50e0;
    ram_cell[    3540] = 32'h0;  // 32'h4bd7c807;
    ram_cell[    3541] = 32'h0;  // 32'h0dfffae5;
    ram_cell[    3542] = 32'h0;  // 32'h9ec163e0;
    ram_cell[    3543] = 32'h0;  // 32'hed9483dc;
    ram_cell[    3544] = 32'h0;  // 32'h98f7da31;
    ram_cell[    3545] = 32'h0;  // 32'hf3a7f3cb;
    ram_cell[    3546] = 32'h0;  // 32'h1d9b4c68;
    ram_cell[    3547] = 32'h0;  // 32'h39098059;
    ram_cell[    3548] = 32'h0;  // 32'h015a6e08;
    ram_cell[    3549] = 32'h0;  // 32'hb3d14ea0;
    ram_cell[    3550] = 32'h0;  // 32'hf7152da9;
    ram_cell[    3551] = 32'h0;  // 32'hd5953945;
    ram_cell[    3552] = 32'h0;  // 32'hcdc9fbff;
    ram_cell[    3553] = 32'h0;  // 32'h4f968f6f;
    ram_cell[    3554] = 32'h0;  // 32'h151ba658;
    ram_cell[    3555] = 32'h0;  // 32'h71cdd034;
    ram_cell[    3556] = 32'h0;  // 32'h11f329eb;
    ram_cell[    3557] = 32'h0;  // 32'h6b03eb7a;
    ram_cell[    3558] = 32'h0;  // 32'hb372ea3b;
    ram_cell[    3559] = 32'h0;  // 32'h984b61df;
    ram_cell[    3560] = 32'h0;  // 32'h6a3abf66;
    ram_cell[    3561] = 32'h0;  // 32'he07620f8;
    ram_cell[    3562] = 32'h0;  // 32'h003304ca;
    ram_cell[    3563] = 32'h0;  // 32'h17a00dad;
    ram_cell[    3564] = 32'h0;  // 32'h6a584f63;
    ram_cell[    3565] = 32'h0;  // 32'hb0467cf5;
    ram_cell[    3566] = 32'h0;  // 32'h61307c50;
    ram_cell[    3567] = 32'h0;  // 32'h1de88720;
    ram_cell[    3568] = 32'h0;  // 32'hfa71c19a;
    ram_cell[    3569] = 32'h0;  // 32'h6f4ea38f;
    ram_cell[    3570] = 32'h0;  // 32'h3b82f747;
    ram_cell[    3571] = 32'h0;  // 32'he3918b06;
    ram_cell[    3572] = 32'h0;  // 32'h5db14b29;
    ram_cell[    3573] = 32'h0;  // 32'h466056a7;
    ram_cell[    3574] = 32'h0;  // 32'hff77f45e;
    ram_cell[    3575] = 32'h0;  // 32'hfbb9427b;
    ram_cell[    3576] = 32'h0;  // 32'h5e0b9faf;
    ram_cell[    3577] = 32'h0;  // 32'hfbbf9a5f;
    ram_cell[    3578] = 32'h0;  // 32'hefb3740b;
    ram_cell[    3579] = 32'h0;  // 32'h31f1ef04;
    ram_cell[    3580] = 32'h0;  // 32'h0d1f9326;
    ram_cell[    3581] = 32'h0;  // 32'hb66a2713;
    ram_cell[    3582] = 32'h0;  // 32'h43430b34;
    ram_cell[    3583] = 32'h0;  // 32'hc6f6b783;
    ram_cell[    3584] = 32'h0;  // 32'h48628a3a;
    ram_cell[    3585] = 32'h0;  // 32'h3973a9b4;
    ram_cell[    3586] = 32'h0;  // 32'heb4e31de;
    ram_cell[    3587] = 32'h0;  // 32'hfb789ad6;
    ram_cell[    3588] = 32'h0;  // 32'h0a7a24ee;
    ram_cell[    3589] = 32'h0;  // 32'hfd6fde24;
    ram_cell[    3590] = 32'h0;  // 32'he9e94e72;
    ram_cell[    3591] = 32'h0;  // 32'h73cac9d8;
    ram_cell[    3592] = 32'h0;  // 32'h2cfe096c;
    ram_cell[    3593] = 32'h0;  // 32'h8b230164;
    ram_cell[    3594] = 32'h0;  // 32'h25e235ce;
    ram_cell[    3595] = 32'h0;  // 32'h5fdb39cc;
    ram_cell[    3596] = 32'h0;  // 32'hd3c2192a;
    ram_cell[    3597] = 32'h0;  // 32'h8ae04fb1;
    ram_cell[    3598] = 32'h0;  // 32'h0593dcb7;
    ram_cell[    3599] = 32'h0;  // 32'h8d254583;
    ram_cell[    3600] = 32'h0;  // 32'h3356a26d;
    ram_cell[    3601] = 32'h0;  // 32'h8235cf6a;
    ram_cell[    3602] = 32'h0;  // 32'h49ca3880;
    ram_cell[    3603] = 32'h0;  // 32'hed63942c;
    ram_cell[    3604] = 32'h0;  // 32'hd73ed98d;
    ram_cell[    3605] = 32'h0;  // 32'h177dfd52;
    ram_cell[    3606] = 32'h0;  // 32'h965646f2;
    ram_cell[    3607] = 32'h0;  // 32'h6ff5a7b1;
    ram_cell[    3608] = 32'h0;  // 32'h51a2b1da;
    ram_cell[    3609] = 32'h0;  // 32'hb2620ffe;
    ram_cell[    3610] = 32'h0;  // 32'h39bc7268;
    ram_cell[    3611] = 32'h0;  // 32'h2c972bf4;
    ram_cell[    3612] = 32'h0;  // 32'h010f67bd;
    ram_cell[    3613] = 32'h0;  // 32'hc01df8f4;
    ram_cell[    3614] = 32'h0;  // 32'h49da1225;
    ram_cell[    3615] = 32'h0;  // 32'h1581211b;
    ram_cell[    3616] = 32'h0;  // 32'h5a7f49b8;
    ram_cell[    3617] = 32'h0;  // 32'h2f8af763;
    ram_cell[    3618] = 32'h0;  // 32'hed58d927;
    ram_cell[    3619] = 32'h0;  // 32'h1fc45bfe;
    ram_cell[    3620] = 32'h0;  // 32'h98688054;
    ram_cell[    3621] = 32'h0;  // 32'hc07c0592;
    ram_cell[    3622] = 32'h0;  // 32'hc76f28ca;
    ram_cell[    3623] = 32'h0;  // 32'hbf67c58f;
    ram_cell[    3624] = 32'h0;  // 32'h5d283fd1;
    ram_cell[    3625] = 32'h0;  // 32'ha8c9a2cd;
    ram_cell[    3626] = 32'h0;  // 32'hec688954;
    ram_cell[    3627] = 32'h0;  // 32'he5353262;
    ram_cell[    3628] = 32'h0;  // 32'he5ca5b26;
    ram_cell[    3629] = 32'h0;  // 32'hd7b360f7;
    ram_cell[    3630] = 32'h0;  // 32'h54d67c42;
    ram_cell[    3631] = 32'h0;  // 32'h29c7fcb2;
    ram_cell[    3632] = 32'h0;  // 32'hd29c3bc0;
    ram_cell[    3633] = 32'h0;  // 32'h1079813b;
    ram_cell[    3634] = 32'h0;  // 32'h0889cf7c;
    ram_cell[    3635] = 32'h0;  // 32'h0b8c0acf;
    ram_cell[    3636] = 32'h0;  // 32'h1d57d38c;
    ram_cell[    3637] = 32'h0;  // 32'he477f334;
    ram_cell[    3638] = 32'h0;  // 32'h5a64569b;
    ram_cell[    3639] = 32'h0;  // 32'h2b1433d9;
    ram_cell[    3640] = 32'h0;  // 32'h545860c8;
    ram_cell[    3641] = 32'h0;  // 32'hc63c370e;
    ram_cell[    3642] = 32'h0;  // 32'h34214adc;
    ram_cell[    3643] = 32'h0;  // 32'h835c2e08;
    ram_cell[    3644] = 32'h0;  // 32'h92ee88be;
    ram_cell[    3645] = 32'h0;  // 32'h808f8d8a;
    ram_cell[    3646] = 32'h0;  // 32'h608012d7;
    ram_cell[    3647] = 32'h0;  // 32'hf6467a41;
    ram_cell[    3648] = 32'h0;  // 32'h55f0f419;
    ram_cell[    3649] = 32'h0;  // 32'he9737d50;
    ram_cell[    3650] = 32'h0;  // 32'h53b3a428;
    ram_cell[    3651] = 32'h0;  // 32'had8862b5;
    ram_cell[    3652] = 32'h0;  // 32'h1d75a425;
    ram_cell[    3653] = 32'h0;  // 32'hf4298f0d;
    ram_cell[    3654] = 32'h0;  // 32'hd86f104d;
    ram_cell[    3655] = 32'h0;  // 32'h8abfa715;
    ram_cell[    3656] = 32'h0;  // 32'h5ab17ea4;
    ram_cell[    3657] = 32'h0;  // 32'hae8b6587;
    ram_cell[    3658] = 32'h0;  // 32'h26e1cb5f;
    ram_cell[    3659] = 32'h0;  // 32'heee9954d;
    ram_cell[    3660] = 32'h0;  // 32'h5b054bd3;
    ram_cell[    3661] = 32'h0;  // 32'he06410e6;
    ram_cell[    3662] = 32'h0;  // 32'h31c82701;
    ram_cell[    3663] = 32'h0;  // 32'h66524ca3;
    ram_cell[    3664] = 32'h0;  // 32'he3fb2d90;
    ram_cell[    3665] = 32'h0;  // 32'hf94657d6;
    ram_cell[    3666] = 32'h0;  // 32'h63360dc0;
    ram_cell[    3667] = 32'h0;  // 32'h5858daee;
    ram_cell[    3668] = 32'h0;  // 32'h38759701;
    ram_cell[    3669] = 32'h0;  // 32'h821048cd;
    ram_cell[    3670] = 32'h0;  // 32'h9b3aa315;
    ram_cell[    3671] = 32'h0;  // 32'h93979841;
    ram_cell[    3672] = 32'h0;  // 32'h580d24c1;
    ram_cell[    3673] = 32'h0;  // 32'h9c9417b8;
    ram_cell[    3674] = 32'h0;  // 32'hba408c75;
    ram_cell[    3675] = 32'h0;  // 32'hfb1bfac5;
    ram_cell[    3676] = 32'h0;  // 32'h1b98645f;
    ram_cell[    3677] = 32'h0;  // 32'h52120af9;
    ram_cell[    3678] = 32'h0;  // 32'hedcf2722;
    ram_cell[    3679] = 32'h0;  // 32'h91e31924;
    ram_cell[    3680] = 32'h0;  // 32'hc4420548;
    ram_cell[    3681] = 32'h0;  // 32'h4a8984d6;
    ram_cell[    3682] = 32'h0;  // 32'hcd96ff00;
    ram_cell[    3683] = 32'h0;  // 32'hc831f43d;
    ram_cell[    3684] = 32'h0;  // 32'h0fc9e14c;
    ram_cell[    3685] = 32'h0;  // 32'hd51e6acf;
    ram_cell[    3686] = 32'h0;  // 32'h129e4567;
    ram_cell[    3687] = 32'h0;  // 32'ha09ff778;
    ram_cell[    3688] = 32'h0;  // 32'h9e34ba06;
    ram_cell[    3689] = 32'h0;  // 32'h91fd26c7;
    ram_cell[    3690] = 32'h0;  // 32'ha22e434a;
    ram_cell[    3691] = 32'h0;  // 32'h9ba86d56;
    ram_cell[    3692] = 32'h0;  // 32'hb3317015;
    ram_cell[    3693] = 32'h0;  // 32'h09e6c6a0;
    ram_cell[    3694] = 32'h0;  // 32'hdcab0841;
    ram_cell[    3695] = 32'h0;  // 32'hffd9f486;
    ram_cell[    3696] = 32'h0;  // 32'h832f8832;
    ram_cell[    3697] = 32'h0;  // 32'hafec6642;
    ram_cell[    3698] = 32'h0;  // 32'ha923f32d;
    ram_cell[    3699] = 32'h0;  // 32'h50930a01;
    ram_cell[    3700] = 32'h0;  // 32'ha3718aaf;
    ram_cell[    3701] = 32'h0;  // 32'hee03030d;
    ram_cell[    3702] = 32'h0;  // 32'hcf351008;
    ram_cell[    3703] = 32'h0;  // 32'hec491993;
    ram_cell[    3704] = 32'h0;  // 32'hdcdb23ee;
    ram_cell[    3705] = 32'h0;  // 32'h07cd1be6;
    ram_cell[    3706] = 32'h0;  // 32'ha305449d;
    ram_cell[    3707] = 32'h0;  // 32'hef8b239b;
    ram_cell[    3708] = 32'h0;  // 32'hb46b177b;
    ram_cell[    3709] = 32'h0;  // 32'hfa9a083e;
    ram_cell[    3710] = 32'h0;  // 32'h1a3984a9;
    ram_cell[    3711] = 32'h0;  // 32'h0043c491;
    ram_cell[    3712] = 32'h0;  // 32'hc8c6384d;
    ram_cell[    3713] = 32'h0;  // 32'hc11f20e6;
    ram_cell[    3714] = 32'h0;  // 32'h1bc4d554;
    ram_cell[    3715] = 32'h0;  // 32'he8a04c72;
    ram_cell[    3716] = 32'h0;  // 32'h80319a90;
    ram_cell[    3717] = 32'h0;  // 32'hd43d7543;
    ram_cell[    3718] = 32'h0;  // 32'h08e5f029;
    ram_cell[    3719] = 32'h0;  // 32'hdad4102c;
    ram_cell[    3720] = 32'h0;  // 32'h6a6987d1;
    ram_cell[    3721] = 32'h0;  // 32'h9d18c0e4;
    ram_cell[    3722] = 32'h0;  // 32'h45ddc20f;
    ram_cell[    3723] = 32'h0;  // 32'h0a6843ce;
    ram_cell[    3724] = 32'h0;  // 32'h3a8899a3;
    ram_cell[    3725] = 32'h0;  // 32'h4230ca1d;
    ram_cell[    3726] = 32'h0;  // 32'hadc65c20;
    ram_cell[    3727] = 32'h0;  // 32'he110c683;
    ram_cell[    3728] = 32'h0;  // 32'h5790199f;
    ram_cell[    3729] = 32'h0;  // 32'hd2fffe36;
    ram_cell[    3730] = 32'h0;  // 32'h8e3512a9;
    ram_cell[    3731] = 32'h0;  // 32'hd0d67fba;
    ram_cell[    3732] = 32'h0;  // 32'hbba86d70;
    ram_cell[    3733] = 32'h0;  // 32'h09d2032e;
    ram_cell[    3734] = 32'h0;  // 32'he8e0414b;
    ram_cell[    3735] = 32'h0;  // 32'h4e6851cb;
    ram_cell[    3736] = 32'h0;  // 32'h2b1cb67e;
    ram_cell[    3737] = 32'h0;  // 32'h79eae17f;
    ram_cell[    3738] = 32'h0;  // 32'h1351faf0;
    ram_cell[    3739] = 32'h0;  // 32'h4963ac53;
    ram_cell[    3740] = 32'h0;  // 32'hfeb3e4b4;
    ram_cell[    3741] = 32'h0;  // 32'hcde415e3;
    ram_cell[    3742] = 32'h0;  // 32'h54cfc3e8;
    ram_cell[    3743] = 32'h0;  // 32'hcec9d641;
    ram_cell[    3744] = 32'h0;  // 32'h6f65764b;
    ram_cell[    3745] = 32'h0;  // 32'hde9cbd47;
    ram_cell[    3746] = 32'h0;  // 32'h73f9ddd3;
    ram_cell[    3747] = 32'h0;  // 32'hf4f2b175;
    ram_cell[    3748] = 32'h0;  // 32'h0096ce68;
    ram_cell[    3749] = 32'h0;  // 32'haf8867aa;
    ram_cell[    3750] = 32'h0;  // 32'hd3b90d7f;
    ram_cell[    3751] = 32'h0;  // 32'hd2b5a5a1;
    ram_cell[    3752] = 32'h0;  // 32'hc0d43477;
    ram_cell[    3753] = 32'h0;  // 32'h0ffe0cde;
    ram_cell[    3754] = 32'h0;  // 32'h4744cfa2;
    ram_cell[    3755] = 32'h0;  // 32'ha7d53109;
    ram_cell[    3756] = 32'h0;  // 32'h0489fda6;
    ram_cell[    3757] = 32'h0;  // 32'h5a516269;
    ram_cell[    3758] = 32'h0;  // 32'h89f3b251;
    ram_cell[    3759] = 32'h0;  // 32'hc42ed866;
    ram_cell[    3760] = 32'h0;  // 32'h56872382;
    ram_cell[    3761] = 32'h0;  // 32'h20178abf;
    ram_cell[    3762] = 32'h0;  // 32'hed3787aa;
    ram_cell[    3763] = 32'h0;  // 32'he68585e8;
    ram_cell[    3764] = 32'h0;  // 32'h4ca2240f;
    ram_cell[    3765] = 32'h0;  // 32'h480066de;
    ram_cell[    3766] = 32'h0;  // 32'h348ca6e6;
    ram_cell[    3767] = 32'h0;  // 32'hd88ef17c;
    ram_cell[    3768] = 32'h0;  // 32'h5a0516c2;
    ram_cell[    3769] = 32'h0;  // 32'h7db08d0f;
    ram_cell[    3770] = 32'h0;  // 32'h45f26390;
    ram_cell[    3771] = 32'h0;  // 32'h6b4d9a4e;
    ram_cell[    3772] = 32'h0;  // 32'h927faf3f;
    ram_cell[    3773] = 32'h0;  // 32'hc9786ecf;
    ram_cell[    3774] = 32'h0;  // 32'h4d42bcdd;
    ram_cell[    3775] = 32'h0;  // 32'h725e0721;
    ram_cell[    3776] = 32'h0;  // 32'hda0e8972;
    ram_cell[    3777] = 32'h0;  // 32'h44e88949;
    ram_cell[    3778] = 32'h0;  // 32'h47ede77c;
    ram_cell[    3779] = 32'h0;  // 32'h637c1cff;
    ram_cell[    3780] = 32'h0;  // 32'h7efc4bde;
    ram_cell[    3781] = 32'h0;  // 32'hb767e368;
    ram_cell[    3782] = 32'h0;  // 32'hfdcc422a;
    ram_cell[    3783] = 32'h0;  // 32'hb2d5e240;
    ram_cell[    3784] = 32'h0;  // 32'h9582d740;
    ram_cell[    3785] = 32'h0;  // 32'h305f79bc;
    ram_cell[    3786] = 32'h0;  // 32'hf3aadbd5;
    ram_cell[    3787] = 32'h0;  // 32'hcd61e059;
    ram_cell[    3788] = 32'h0;  // 32'haa77fd19;
    ram_cell[    3789] = 32'h0;  // 32'h8f3ab7f5;
    ram_cell[    3790] = 32'h0;  // 32'hd71f6385;
    ram_cell[    3791] = 32'h0;  // 32'h8b922003;
    ram_cell[    3792] = 32'h0;  // 32'hf8d26862;
    ram_cell[    3793] = 32'h0;  // 32'h5ed98568;
    ram_cell[    3794] = 32'h0;  // 32'h50379cf0;
    ram_cell[    3795] = 32'h0;  // 32'he06c13ac;
    ram_cell[    3796] = 32'h0;  // 32'h5f3e4b9e;
    ram_cell[    3797] = 32'h0;  // 32'h88563870;
    ram_cell[    3798] = 32'h0;  // 32'hef345b27;
    ram_cell[    3799] = 32'h0;  // 32'h4d34a4f9;
    ram_cell[    3800] = 32'h0;  // 32'h016273bc;
    ram_cell[    3801] = 32'h0;  // 32'h00eccabc;
    ram_cell[    3802] = 32'h0;  // 32'h4ae5eb99;
    ram_cell[    3803] = 32'h0;  // 32'hddc2b17f;
    ram_cell[    3804] = 32'h0;  // 32'h601f8aad;
    ram_cell[    3805] = 32'h0;  // 32'h71980671;
    ram_cell[    3806] = 32'h0;  // 32'h6475dafa;
    ram_cell[    3807] = 32'h0;  // 32'hec0d5ad5;
    ram_cell[    3808] = 32'h0;  // 32'h6a1ca6a6;
    ram_cell[    3809] = 32'h0;  // 32'hb8ed92ee;
    ram_cell[    3810] = 32'h0;  // 32'h07f5a7ef;
    ram_cell[    3811] = 32'h0;  // 32'h64ca4939;
    ram_cell[    3812] = 32'h0;  // 32'he472449f;
    ram_cell[    3813] = 32'h0;  // 32'h56e851dd;
    ram_cell[    3814] = 32'h0;  // 32'h2f71374d;
    ram_cell[    3815] = 32'h0;  // 32'h468c6def;
    ram_cell[    3816] = 32'h0;  // 32'he1e48c63;
    ram_cell[    3817] = 32'h0;  // 32'h7509792e;
    ram_cell[    3818] = 32'h0;  // 32'hc1ab5137;
    ram_cell[    3819] = 32'h0;  // 32'h5b9c6e20;
    ram_cell[    3820] = 32'h0;  // 32'hfcf9271d;
    ram_cell[    3821] = 32'h0;  // 32'h896ee29a;
    ram_cell[    3822] = 32'h0;  // 32'hbed78a49;
    ram_cell[    3823] = 32'h0;  // 32'hc46abb29;
    ram_cell[    3824] = 32'h0;  // 32'h9379311c;
    ram_cell[    3825] = 32'h0;  // 32'h44e1c20d;
    ram_cell[    3826] = 32'h0;  // 32'h948ff740;
    ram_cell[    3827] = 32'h0;  // 32'hdcb5248d;
    ram_cell[    3828] = 32'h0;  // 32'h2760fa65;
    ram_cell[    3829] = 32'h0;  // 32'hb63a3775;
    ram_cell[    3830] = 32'h0;  // 32'h4e6a36c2;
    ram_cell[    3831] = 32'h0;  // 32'h348b852c;
    ram_cell[    3832] = 32'h0;  // 32'hb079cc8a;
    ram_cell[    3833] = 32'h0;  // 32'heeaa852f;
    ram_cell[    3834] = 32'h0;  // 32'heefe2a9c;
    ram_cell[    3835] = 32'h0;  // 32'h89d6c691;
    ram_cell[    3836] = 32'h0;  // 32'hdfb60e0e;
    ram_cell[    3837] = 32'h0;  // 32'hb2102b38;
    ram_cell[    3838] = 32'h0;  // 32'hcdbc9441;
    ram_cell[    3839] = 32'h0;  // 32'h9db54038;
    ram_cell[    3840] = 32'h0;  // 32'h56de5cd2;
    ram_cell[    3841] = 32'h0;  // 32'h7d412f46;
    ram_cell[    3842] = 32'h0;  // 32'h95cef025;
    ram_cell[    3843] = 32'h0;  // 32'h5dc521e0;
    ram_cell[    3844] = 32'h0;  // 32'hd06c3097;
    ram_cell[    3845] = 32'h0;  // 32'h58a61bce;
    ram_cell[    3846] = 32'h0;  // 32'he73aeea8;
    ram_cell[    3847] = 32'h0;  // 32'h5f26c65a;
    ram_cell[    3848] = 32'h0;  // 32'h9a97ee0a;
    ram_cell[    3849] = 32'h0;  // 32'hc0fa4f44;
    ram_cell[    3850] = 32'h0;  // 32'h3caf8759;
    ram_cell[    3851] = 32'h0;  // 32'h6b0f292c;
    ram_cell[    3852] = 32'h0;  // 32'h0c9eb8b4;
    ram_cell[    3853] = 32'h0;  // 32'h841cd704;
    ram_cell[    3854] = 32'h0;  // 32'h5a91f2f0;
    ram_cell[    3855] = 32'h0;  // 32'hcfded02f;
    ram_cell[    3856] = 32'h0;  // 32'he3f6f145;
    ram_cell[    3857] = 32'h0;  // 32'hdb427056;
    ram_cell[    3858] = 32'h0;  // 32'h83732a0f;
    ram_cell[    3859] = 32'h0;  // 32'h0f8da133;
    ram_cell[    3860] = 32'h0;  // 32'h4f64d817;
    ram_cell[    3861] = 32'h0;  // 32'hcba4671a;
    ram_cell[    3862] = 32'h0;  // 32'h52b0617b;
    ram_cell[    3863] = 32'h0;  // 32'h301d8b63;
    ram_cell[    3864] = 32'h0;  // 32'h384aa1bb;
    ram_cell[    3865] = 32'h0;  // 32'h42e84042;
    ram_cell[    3866] = 32'h0;  // 32'ha0f51e4c;
    ram_cell[    3867] = 32'h0;  // 32'h02ae13f3;
    ram_cell[    3868] = 32'h0;  // 32'had311cc2;
    ram_cell[    3869] = 32'h0;  // 32'h01ea110b;
    ram_cell[    3870] = 32'h0;  // 32'ha12686c8;
    ram_cell[    3871] = 32'h0;  // 32'h836fb494;
    ram_cell[    3872] = 32'h0;  // 32'he4b0bbf2;
    ram_cell[    3873] = 32'h0;  // 32'hd4a6d4c8;
    ram_cell[    3874] = 32'h0;  // 32'h0299c2b0;
    ram_cell[    3875] = 32'h0;  // 32'h19c4045e;
    ram_cell[    3876] = 32'h0;  // 32'h861625b4;
    ram_cell[    3877] = 32'h0;  // 32'h8055f636;
    ram_cell[    3878] = 32'h0;  // 32'hcf869a99;
    ram_cell[    3879] = 32'h0;  // 32'h25e708eb;
    ram_cell[    3880] = 32'h0;  // 32'hf4d9f53a;
    ram_cell[    3881] = 32'h0;  // 32'h440ca1d7;
    ram_cell[    3882] = 32'h0;  // 32'hab0c8452;
    ram_cell[    3883] = 32'h0;  // 32'h4d9c04dc;
    ram_cell[    3884] = 32'h0;  // 32'h9473ce72;
    ram_cell[    3885] = 32'h0;  // 32'h6b8a47bd;
    ram_cell[    3886] = 32'h0;  // 32'h265ba322;
    ram_cell[    3887] = 32'h0;  // 32'h95730c3b;
    ram_cell[    3888] = 32'h0;  // 32'hf3d7418b;
    ram_cell[    3889] = 32'h0;  // 32'hf4ba5080;
    ram_cell[    3890] = 32'h0;  // 32'headf2efb;
    ram_cell[    3891] = 32'h0;  // 32'h2b81196d;
    ram_cell[    3892] = 32'h0;  // 32'hf7af433f;
    ram_cell[    3893] = 32'h0;  // 32'h46a75bf2;
    ram_cell[    3894] = 32'h0;  // 32'h134b3e62;
    ram_cell[    3895] = 32'h0;  // 32'hb64ed7df;
    ram_cell[    3896] = 32'h0;  // 32'h5a51addc;
    ram_cell[    3897] = 32'h0;  // 32'hb98714e4;
    ram_cell[    3898] = 32'h0;  // 32'h58d59a22;
    ram_cell[    3899] = 32'h0;  // 32'h886be2cf;
    ram_cell[    3900] = 32'h0;  // 32'h2aedb87e;
    ram_cell[    3901] = 32'h0;  // 32'he68dd8da;
    ram_cell[    3902] = 32'h0;  // 32'h772360b7;
    ram_cell[    3903] = 32'h0;  // 32'h43ceed71;
    ram_cell[    3904] = 32'h0;  // 32'hbecaeec1;
    ram_cell[    3905] = 32'h0;  // 32'hf8c3d993;
    ram_cell[    3906] = 32'h0;  // 32'h8ded8a9d;
    ram_cell[    3907] = 32'h0;  // 32'he75493c6;
    ram_cell[    3908] = 32'h0;  // 32'hb3df8d50;
    ram_cell[    3909] = 32'h0;  // 32'h8684ca4a;
    ram_cell[    3910] = 32'h0;  // 32'he1fb7232;
    ram_cell[    3911] = 32'h0;  // 32'he9c098a3;
    ram_cell[    3912] = 32'h0;  // 32'h0440f35b;
    ram_cell[    3913] = 32'h0;  // 32'h04c2c767;
    ram_cell[    3914] = 32'h0;  // 32'h2b888b2c;
    ram_cell[    3915] = 32'h0;  // 32'h3d36477e;
    ram_cell[    3916] = 32'h0;  // 32'h2645640a;
    ram_cell[    3917] = 32'h0;  // 32'hefbd0102;
    ram_cell[    3918] = 32'h0;  // 32'hb46b3a0f;
    ram_cell[    3919] = 32'h0;  // 32'hd0af4cb6;
    ram_cell[    3920] = 32'h0;  // 32'h621c60ee;
    ram_cell[    3921] = 32'h0;  // 32'hcd07c8c3;
    ram_cell[    3922] = 32'h0;  // 32'h5c671fed;
    ram_cell[    3923] = 32'h0;  // 32'h3b4c1ab5;
    ram_cell[    3924] = 32'h0;  // 32'h8ba6eda7;
    ram_cell[    3925] = 32'h0;  // 32'h750a35b2;
    ram_cell[    3926] = 32'h0;  // 32'h9d8d9319;
    ram_cell[    3927] = 32'h0;  // 32'h99e8c6bf;
    ram_cell[    3928] = 32'h0;  // 32'h9cd29782;
    ram_cell[    3929] = 32'h0;  // 32'h4b25c789;
    ram_cell[    3930] = 32'h0;  // 32'h151ee444;
    ram_cell[    3931] = 32'h0;  // 32'he6d2bf6f;
    ram_cell[    3932] = 32'h0;  // 32'h38c38266;
    ram_cell[    3933] = 32'h0;  // 32'h99b45471;
    ram_cell[    3934] = 32'h0;  // 32'h348ffc67;
    ram_cell[    3935] = 32'h0;  // 32'h1fc1045e;
    ram_cell[    3936] = 32'h0;  // 32'hf7236b95;
    ram_cell[    3937] = 32'h0;  // 32'h9c460c12;
    ram_cell[    3938] = 32'h0;  // 32'h1f817892;
    ram_cell[    3939] = 32'h0;  // 32'h9b197102;
    ram_cell[    3940] = 32'h0;  // 32'hbccfe193;
    ram_cell[    3941] = 32'h0;  // 32'h5b0c94a4;
    ram_cell[    3942] = 32'h0;  // 32'hf7f6df8d;
    ram_cell[    3943] = 32'h0;  // 32'habd84146;
    ram_cell[    3944] = 32'h0;  // 32'hb7a823de;
    ram_cell[    3945] = 32'h0;  // 32'ha542350b;
    ram_cell[    3946] = 32'h0;  // 32'hdb72f7ef;
    ram_cell[    3947] = 32'h0;  // 32'hc22ee796;
    ram_cell[    3948] = 32'h0;  // 32'hda12c016;
    ram_cell[    3949] = 32'h0;  // 32'h9b1473e7;
    ram_cell[    3950] = 32'h0;  // 32'hc2a17541;
    ram_cell[    3951] = 32'h0;  // 32'hb08d45e2;
    ram_cell[    3952] = 32'h0;  // 32'hfcf4534c;
    ram_cell[    3953] = 32'h0;  // 32'h8e81ef1d;
    ram_cell[    3954] = 32'h0;  // 32'hb49c2222;
    ram_cell[    3955] = 32'h0;  // 32'hea03f948;
    ram_cell[    3956] = 32'h0;  // 32'h0ec52529;
    ram_cell[    3957] = 32'h0;  // 32'h73c2437b;
    ram_cell[    3958] = 32'h0;  // 32'hfb5be422;
    ram_cell[    3959] = 32'h0;  // 32'h8e686fc6;
    ram_cell[    3960] = 32'h0;  // 32'hae46bc13;
    ram_cell[    3961] = 32'h0;  // 32'h708ebacd;
    ram_cell[    3962] = 32'h0;  // 32'h7aafad1f;
    ram_cell[    3963] = 32'h0;  // 32'he646e69c;
    ram_cell[    3964] = 32'h0;  // 32'h563ae90b;
    ram_cell[    3965] = 32'h0;  // 32'hc4d11a2e;
    ram_cell[    3966] = 32'h0;  // 32'h1399f95e;
    ram_cell[    3967] = 32'h0;  // 32'he9787e61;
    ram_cell[    3968] = 32'h0;  // 32'h832dabac;
    ram_cell[    3969] = 32'h0;  // 32'h0e258911;
    ram_cell[    3970] = 32'h0;  // 32'h2fff1e3d;
    ram_cell[    3971] = 32'h0;  // 32'h581de7fa;
    ram_cell[    3972] = 32'h0;  // 32'h691830d6;
    ram_cell[    3973] = 32'h0;  // 32'h0a6dae0a;
    ram_cell[    3974] = 32'h0;  // 32'h501927e4;
    ram_cell[    3975] = 32'h0;  // 32'h6541b3ee;
    ram_cell[    3976] = 32'h0;  // 32'h1b358155;
    ram_cell[    3977] = 32'h0;  // 32'hce2aa258;
    ram_cell[    3978] = 32'h0;  // 32'h228e3bc4;
    ram_cell[    3979] = 32'h0;  // 32'hef208b23;
    ram_cell[    3980] = 32'h0;  // 32'hd8eb0390;
    ram_cell[    3981] = 32'h0;  // 32'h518ee6bb;
    ram_cell[    3982] = 32'h0;  // 32'h9cce0e07;
    ram_cell[    3983] = 32'h0;  // 32'h75f5e620;
    ram_cell[    3984] = 32'h0;  // 32'h9e5090f2;
    ram_cell[    3985] = 32'h0;  // 32'ha7356cc6;
    ram_cell[    3986] = 32'h0;  // 32'h36d7919d;
    ram_cell[    3987] = 32'h0;  // 32'h04fbe54a;
    ram_cell[    3988] = 32'h0;  // 32'h9a2c6f6f;
    ram_cell[    3989] = 32'h0;  // 32'ha72c6bd9;
    ram_cell[    3990] = 32'h0;  // 32'h8a56fdf1;
    ram_cell[    3991] = 32'h0;  // 32'h0ab55dff;
    ram_cell[    3992] = 32'h0;  // 32'hbae419ed;
    ram_cell[    3993] = 32'h0;  // 32'hf25b5590;
    ram_cell[    3994] = 32'h0;  // 32'h74011d5d;
    ram_cell[    3995] = 32'h0;  // 32'h3413c885;
    ram_cell[    3996] = 32'h0;  // 32'h3b41637f;
    ram_cell[    3997] = 32'h0;  // 32'hce0b9b9e;
    ram_cell[    3998] = 32'h0;  // 32'he69e0ae6;
    ram_cell[    3999] = 32'h0;  // 32'h481030b1;
    ram_cell[    4000] = 32'h0;  // 32'h1d45571f;
    ram_cell[    4001] = 32'h0;  // 32'h07024d98;
    ram_cell[    4002] = 32'h0;  // 32'h62824304;
    ram_cell[    4003] = 32'h0;  // 32'h5bcdeeb4;
    ram_cell[    4004] = 32'h0;  // 32'hd6e4954a;
    ram_cell[    4005] = 32'h0;  // 32'had37d763;
    ram_cell[    4006] = 32'h0;  // 32'h9f7cdb3d;
    ram_cell[    4007] = 32'h0;  // 32'h1b8d2c8f;
    ram_cell[    4008] = 32'h0;  // 32'h3e881d93;
    ram_cell[    4009] = 32'h0;  // 32'h193ae8b4;
    ram_cell[    4010] = 32'h0;  // 32'h3837726d;
    ram_cell[    4011] = 32'h0;  // 32'hc3343fae;
    ram_cell[    4012] = 32'h0;  // 32'h6a86585b;
    ram_cell[    4013] = 32'h0;  // 32'h5a839f56;
    ram_cell[    4014] = 32'h0;  // 32'h1645c837;
    ram_cell[    4015] = 32'h0;  // 32'hf652bdc9;
    ram_cell[    4016] = 32'h0;  // 32'h591aa724;
    ram_cell[    4017] = 32'h0;  // 32'h5ce5e28f;
    ram_cell[    4018] = 32'h0;  // 32'he74ac934;
    ram_cell[    4019] = 32'h0;  // 32'h3c852ac4;
    ram_cell[    4020] = 32'h0;  // 32'haaaeadbc;
    ram_cell[    4021] = 32'h0;  // 32'hfb63fada;
    ram_cell[    4022] = 32'h0;  // 32'h7e024cf7;
    ram_cell[    4023] = 32'h0;  // 32'he1cef598;
    ram_cell[    4024] = 32'h0;  // 32'h31f2a5d2;
    ram_cell[    4025] = 32'h0;  // 32'h7293b981;
    ram_cell[    4026] = 32'h0;  // 32'hfd43dab2;
    ram_cell[    4027] = 32'h0;  // 32'he7e914b8;
    ram_cell[    4028] = 32'h0;  // 32'hf2699f75;
    ram_cell[    4029] = 32'h0;  // 32'hbb6fd016;
    ram_cell[    4030] = 32'h0;  // 32'he54dd763;
    ram_cell[    4031] = 32'h0;  // 32'h387e05fc;
    ram_cell[    4032] = 32'h0;  // 32'h19e78e63;
    ram_cell[    4033] = 32'h0;  // 32'h99e56e91;
    ram_cell[    4034] = 32'h0;  // 32'h208611e2;
    ram_cell[    4035] = 32'h0;  // 32'h3284d536;
    ram_cell[    4036] = 32'h0;  // 32'h359d8b15;
    ram_cell[    4037] = 32'h0;  // 32'he1a8b933;
    ram_cell[    4038] = 32'h0;  // 32'h03f0aca3;
    ram_cell[    4039] = 32'h0;  // 32'hc7c65904;
    ram_cell[    4040] = 32'h0;  // 32'h0ea8725e;
    ram_cell[    4041] = 32'h0;  // 32'h066319ae;
    ram_cell[    4042] = 32'h0;  // 32'h85620689;
    ram_cell[    4043] = 32'h0;  // 32'h2ee4a70e;
    ram_cell[    4044] = 32'h0;  // 32'h04accbf7;
    ram_cell[    4045] = 32'h0;  // 32'h6706e472;
    ram_cell[    4046] = 32'h0;  // 32'h30c52e0f;
    ram_cell[    4047] = 32'h0;  // 32'h722ef7ff;
    ram_cell[    4048] = 32'h0;  // 32'h29ce1d54;
    ram_cell[    4049] = 32'h0;  // 32'h2c3169f4;
    ram_cell[    4050] = 32'h0;  // 32'h82b28a17;
    ram_cell[    4051] = 32'h0;  // 32'he9fa6117;
    ram_cell[    4052] = 32'h0;  // 32'h67f63ebd;
    ram_cell[    4053] = 32'h0;  // 32'h514ef208;
    ram_cell[    4054] = 32'h0;  // 32'h4d510d83;
    ram_cell[    4055] = 32'h0;  // 32'hc41bb303;
    ram_cell[    4056] = 32'h0;  // 32'h0457e77e;
    ram_cell[    4057] = 32'h0;  // 32'h04fc8e7e;
    ram_cell[    4058] = 32'h0;  // 32'h68df1c0e;
    ram_cell[    4059] = 32'h0;  // 32'ha14617bc;
    ram_cell[    4060] = 32'h0;  // 32'h531eac3b;
    ram_cell[    4061] = 32'h0;  // 32'hf1e7ef0d;
    ram_cell[    4062] = 32'h0;  // 32'h04b7a6ca;
    ram_cell[    4063] = 32'h0;  // 32'h40e35fe1;
    ram_cell[    4064] = 32'h0;  // 32'ha936e5af;
    ram_cell[    4065] = 32'h0;  // 32'h8aa981c7;
    ram_cell[    4066] = 32'h0;  // 32'hb58ea5ea;
    ram_cell[    4067] = 32'h0;  // 32'h54fc9bcb;
    ram_cell[    4068] = 32'h0;  // 32'hc219f9a6;
    ram_cell[    4069] = 32'h0;  // 32'h2fa261f5;
    ram_cell[    4070] = 32'h0;  // 32'he0abeb81;
    ram_cell[    4071] = 32'h0;  // 32'hebfc90f5;
    ram_cell[    4072] = 32'h0;  // 32'h661d658f;
    ram_cell[    4073] = 32'h0;  // 32'h0b1801a8;
    ram_cell[    4074] = 32'h0;  // 32'h366390cb;
    ram_cell[    4075] = 32'h0;  // 32'hfa2d6026;
    ram_cell[    4076] = 32'h0;  // 32'h8dd53d3a;
    ram_cell[    4077] = 32'h0;  // 32'h1b1182fe;
    ram_cell[    4078] = 32'h0;  // 32'h114617fc;
    ram_cell[    4079] = 32'h0;  // 32'h5896812b;
    ram_cell[    4080] = 32'h0;  // 32'h41bc917d;
    ram_cell[    4081] = 32'h0;  // 32'h888615c0;
    ram_cell[    4082] = 32'h0;  // 32'hf1232246;
    ram_cell[    4083] = 32'h0;  // 32'h793e694f;
    ram_cell[    4084] = 32'h0;  // 32'h291760f6;
    ram_cell[    4085] = 32'h0;  // 32'h946f5f92;
    ram_cell[    4086] = 32'h0;  // 32'hab3a7b53;
    ram_cell[    4087] = 32'h0;  // 32'h097a7a79;
    ram_cell[    4088] = 32'h0;  // 32'h1b5565ec;
    ram_cell[    4089] = 32'h0;  // 32'hc8cca379;
    ram_cell[    4090] = 32'h0;  // 32'h2f87ed8a;
    ram_cell[    4091] = 32'h0;  // 32'hd0104160;
    ram_cell[    4092] = 32'h0;  // 32'h38a4c9cf;
    ram_cell[    4093] = 32'h0;  // 32'h60a17d5a;
    ram_cell[    4094] = 32'h0;  // 32'h7bc9b359;
    ram_cell[    4095] = 32'h0;  // 32'h8c380a75;
    // src matrix A
    ram_cell[    4096] = 32'ha7a1ef5a;
    ram_cell[    4097] = 32'h5beb79d9;
    ram_cell[    4098] = 32'he2ee8c0b;
    ram_cell[    4099] = 32'hc7560283;
    ram_cell[    4100] = 32'h7b3cde48;
    ram_cell[    4101] = 32'h189470ec;
    ram_cell[    4102] = 32'h372b0673;
    ram_cell[    4103] = 32'hc30c2748;
    ram_cell[    4104] = 32'h0cec4c9a;
    ram_cell[    4105] = 32'h8da5c4a5;
    ram_cell[    4106] = 32'h5ecca58d;
    ram_cell[    4107] = 32'h77c687da;
    ram_cell[    4108] = 32'h6682de9b;
    ram_cell[    4109] = 32'h296e5546;
    ram_cell[    4110] = 32'h783dd747;
    ram_cell[    4111] = 32'h4b7f5afa;
    ram_cell[    4112] = 32'h28c2276b;
    ram_cell[    4113] = 32'hdd5642d8;
    ram_cell[    4114] = 32'h5df44330;
    ram_cell[    4115] = 32'h4005780b;
    ram_cell[    4116] = 32'hb200334d;
    ram_cell[    4117] = 32'h11db681d;
    ram_cell[    4118] = 32'hc3514de1;
    ram_cell[    4119] = 32'he315ecc9;
    ram_cell[    4120] = 32'hd67c4e89;
    ram_cell[    4121] = 32'h6fef9009;
    ram_cell[    4122] = 32'h99be27ed;
    ram_cell[    4123] = 32'he50ab0f1;
    ram_cell[    4124] = 32'hc768b8d1;
    ram_cell[    4125] = 32'h1a839b07;
    ram_cell[    4126] = 32'h8454f26e;
    ram_cell[    4127] = 32'hdd6873b0;
    ram_cell[    4128] = 32'hea4053ac;
    ram_cell[    4129] = 32'h4b290a1c;
    ram_cell[    4130] = 32'h015072be;
    ram_cell[    4131] = 32'h613e785c;
    ram_cell[    4132] = 32'h1c908e0d;
    ram_cell[    4133] = 32'h76c25281;
    ram_cell[    4134] = 32'h3c3103cc;
    ram_cell[    4135] = 32'hd9802206;
    ram_cell[    4136] = 32'h86a93a5b;
    ram_cell[    4137] = 32'hd9d40071;
    ram_cell[    4138] = 32'h8184e8b1;
    ram_cell[    4139] = 32'hf9d8ef40;
    ram_cell[    4140] = 32'h44ca5f42;
    ram_cell[    4141] = 32'ha560b50c;
    ram_cell[    4142] = 32'hd10f0cc9;
    ram_cell[    4143] = 32'hbc8e63ff;
    ram_cell[    4144] = 32'hab14c380;
    ram_cell[    4145] = 32'h7b587c00;
    ram_cell[    4146] = 32'h4cf04106;
    ram_cell[    4147] = 32'h6b26dea5;
    ram_cell[    4148] = 32'h9f2b70e0;
    ram_cell[    4149] = 32'h84303ecc;
    ram_cell[    4150] = 32'h62ebf33a;
    ram_cell[    4151] = 32'h50f41a1d;
    ram_cell[    4152] = 32'haf7d32ae;
    ram_cell[    4153] = 32'h9337c39d;
    ram_cell[    4154] = 32'h30baaef5;
    ram_cell[    4155] = 32'h3a12a78d;
    ram_cell[    4156] = 32'h971fb05c;
    ram_cell[    4157] = 32'h578b3514;
    ram_cell[    4158] = 32'h80e0ccd9;
    ram_cell[    4159] = 32'h644a1f74;
    ram_cell[    4160] = 32'h4064f78a;
    ram_cell[    4161] = 32'h30d4bcc1;
    ram_cell[    4162] = 32'hf6f5232a;
    ram_cell[    4163] = 32'h54a2ff3a;
    ram_cell[    4164] = 32'hcac62e64;
    ram_cell[    4165] = 32'he2d3b2e2;
    ram_cell[    4166] = 32'hf50b4885;
    ram_cell[    4167] = 32'h2bbe0c41;
    ram_cell[    4168] = 32'h5aeb55cf;
    ram_cell[    4169] = 32'h4fc91892;
    ram_cell[    4170] = 32'hb0980f8d;
    ram_cell[    4171] = 32'h51774e16;
    ram_cell[    4172] = 32'h57e85499;
    ram_cell[    4173] = 32'h3183724a;
    ram_cell[    4174] = 32'h98fb22dc;
    ram_cell[    4175] = 32'hbd5f0449;
    ram_cell[    4176] = 32'h190a7d72;
    ram_cell[    4177] = 32'hde743de1;
    ram_cell[    4178] = 32'hbc07c393;
    ram_cell[    4179] = 32'h37eef69d;
    ram_cell[    4180] = 32'hff20a2c3;
    ram_cell[    4181] = 32'he24edc77;
    ram_cell[    4182] = 32'h21f400c0;
    ram_cell[    4183] = 32'hecd37526;
    ram_cell[    4184] = 32'haf1ca186;
    ram_cell[    4185] = 32'h5280e8c1;
    ram_cell[    4186] = 32'heb4676e5;
    ram_cell[    4187] = 32'h0c4ba573;
    ram_cell[    4188] = 32'hafdb2819;
    ram_cell[    4189] = 32'hd4e35abe;
    ram_cell[    4190] = 32'h9338c401;
    ram_cell[    4191] = 32'hbc3bb8df;
    ram_cell[    4192] = 32'hd8e4081b;
    ram_cell[    4193] = 32'h386a151a;
    ram_cell[    4194] = 32'h5b391505;
    ram_cell[    4195] = 32'h71a6a69a;
    ram_cell[    4196] = 32'hde892db6;
    ram_cell[    4197] = 32'hf3b3ec25;
    ram_cell[    4198] = 32'h52579d9e;
    ram_cell[    4199] = 32'h4c0524ad;
    ram_cell[    4200] = 32'h2bfda6b4;
    ram_cell[    4201] = 32'h888bddf9;
    ram_cell[    4202] = 32'hc8be2e27;
    ram_cell[    4203] = 32'h16ff2d8d;
    ram_cell[    4204] = 32'h3347c2fd;
    ram_cell[    4205] = 32'h633c706f;
    ram_cell[    4206] = 32'hecd98ff0;
    ram_cell[    4207] = 32'h36211ebc;
    ram_cell[    4208] = 32'hafdb7031;
    ram_cell[    4209] = 32'h6015e064;
    ram_cell[    4210] = 32'haad72034;
    ram_cell[    4211] = 32'h3a3f95cf;
    ram_cell[    4212] = 32'h9ea7245a;
    ram_cell[    4213] = 32'hdbdb8bf8;
    ram_cell[    4214] = 32'h3e202588;
    ram_cell[    4215] = 32'h481bc131;
    ram_cell[    4216] = 32'h22203371;
    ram_cell[    4217] = 32'heb3d0f3d;
    ram_cell[    4218] = 32'hde83ec55;
    ram_cell[    4219] = 32'h6238cc9f;
    ram_cell[    4220] = 32'h2c7d2911;
    ram_cell[    4221] = 32'he7bfa4bc;
    ram_cell[    4222] = 32'hebccb9fc;
    ram_cell[    4223] = 32'hb8c74f11;
    ram_cell[    4224] = 32'h8562cc25;
    ram_cell[    4225] = 32'h5f0b1460;
    ram_cell[    4226] = 32'h60f1c9b8;
    ram_cell[    4227] = 32'h2ce26f18;
    ram_cell[    4228] = 32'h1959a099;
    ram_cell[    4229] = 32'hc2f9ca6a;
    ram_cell[    4230] = 32'h5dd4402c;
    ram_cell[    4231] = 32'h3362bc33;
    ram_cell[    4232] = 32'hdbb48525;
    ram_cell[    4233] = 32'he5ee1c0c;
    ram_cell[    4234] = 32'h0c4c0035;
    ram_cell[    4235] = 32'hc9de8cd7;
    ram_cell[    4236] = 32'h342abfaa;
    ram_cell[    4237] = 32'hd094015b;
    ram_cell[    4238] = 32'hc1c04927;
    ram_cell[    4239] = 32'h94254005;
    ram_cell[    4240] = 32'hf99c1667;
    ram_cell[    4241] = 32'hee8a8f25;
    ram_cell[    4242] = 32'hbbb17dc4;
    ram_cell[    4243] = 32'h8e7d8df9;
    ram_cell[    4244] = 32'h7b3df979;
    ram_cell[    4245] = 32'hd4f3e543;
    ram_cell[    4246] = 32'h0114e02b;
    ram_cell[    4247] = 32'hf824b014;
    ram_cell[    4248] = 32'h0c2af2d2;
    ram_cell[    4249] = 32'hde960eea;
    ram_cell[    4250] = 32'he709087a;
    ram_cell[    4251] = 32'h007a9a03;
    ram_cell[    4252] = 32'h49eeaebb;
    ram_cell[    4253] = 32'h3f68160c;
    ram_cell[    4254] = 32'h05b8af39;
    ram_cell[    4255] = 32'h471bb25b;
    ram_cell[    4256] = 32'hcfc2cb8d;
    ram_cell[    4257] = 32'h67631fd6;
    ram_cell[    4258] = 32'h4ec10638;
    ram_cell[    4259] = 32'heed8731b;
    ram_cell[    4260] = 32'h8476793f;
    ram_cell[    4261] = 32'h2cd255ec;
    ram_cell[    4262] = 32'h93b68f62;
    ram_cell[    4263] = 32'hd93aa31c;
    ram_cell[    4264] = 32'h2d5a450e;
    ram_cell[    4265] = 32'h74e0bdc5;
    ram_cell[    4266] = 32'hf9724852;
    ram_cell[    4267] = 32'hb4fdbf4e;
    ram_cell[    4268] = 32'hb0cf3d3a;
    ram_cell[    4269] = 32'h984362cd;
    ram_cell[    4270] = 32'h9f942f5b;
    ram_cell[    4271] = 32'hd4e09ad5;
    ram_cell[    4272] = 32'hf2ec81ec;
    ram_cell[    4273] = 32'h767e13e7;
    ram_cell[    4274] = 32'hbaae158d;
    ram_cell[    4275] = 32'h63457b9b;
    ram_cell[    4276] = 32'h80aaca5d;
    ram_cell[    4277] = 32'hda5356b2;
    ram_cell[    4278] = 32'h674d314c;
    ram_cell[    4279] = 32'hf2489a6f;
    ram_cell[    4280] = 32'h2834e8c5;
    ram_cell[    4281] = 32'h33c90676;
    ram_cell[    4282] = 32'hf64b93fb;
    ram_cell[    4283] = 32'h63a5004a;
    ram_cell[    4284] = 32'h949ecb77;
    ram_cell[    4285] = 32'h53b27039;
    ram_cell[    4286] = 32'hc3e5573a;
    ram_cell[    4287] = 32'hb5ce8b21;
    ram_cell[    4288] = 32'h70141f64;
    ram_cell[    4289] = 32'h68a0ec93;
    ram_cell[    4290] = 32'h44302c49;
    ram_cell[    4291] = 32'h09521165;
    ram_cell[    4292] = 32'h5f8d5fb4;
    ram_cell[    4293] = 32'hd07d6bef;
    ram_cell[    4294] = 32'h5b268f7a;
    ram_cell[    4295] = 32'h2454a3f4;
    ram_cell[    4296] = 32'h6a6ef13d;
    ram_cell[    4297] = 32'hfb7966e5;
    ram_cell[    4298] = 32'h707c4b14;
    ram_cell[    4299] = 32'hb1e6ef40;
    ram_cell[    4300] = 32'h59e3ca49;
    ram_cell[    4301] = 32'h6749f3a0;
    ram_cell[    4302] = 32'heef49b3b;
    ram_cell[    4303] = 32'h323676d5;
    ram_cell[    4304] = 32'h206d2e79;
    ram_cell[    4305] = 32'h3ea62b63;
    ram_cell[    4306] = 32'h6152ff04;
    ram_cell[    4307] = 32'hb17e455f;
    ram_cell[    4308] = 32'hd07ae0da;
    ram_cell[    4309] = 32'h288534af;
    ram_cell[    4310] = 32'he7bd6275;
    ram_cell[    4311] = 32'h499f1814;
    ram_cell[    4312] = 32'hd27761cc;
    ram_cell[    4313] = 32'h14e870e1;
    ram_cell[    4314] = 32'h16283dd0;
    ram_cell[    4315] = 32'hccca4a6e;
    ram_cell[    4316] = 32'h7fb32629;
    ram_cell[    4317] = 32'hbac94107;
    ram_cell[    4318] = 32'hf1c30d2e;
    ram_cell[    4319] = 32'h65c6b9a5;
    ram_cell[    4320] = 32'h4ce5ff78;
    ram_cell[    4321] = 32'he712bba3;
    ram_cell[    4322] = 32'hc0c595aa;
    ram_cell[    4323] = 32'h8a8764c1;
    ram_cell[    4324] = 32'h083b12a3;
    ram_cell[    4325] = 32'he9a91293;
    ram_cell[    4326] = 32'h04eff6c7;
    ram_cell[    4327] = 32'h141e87a9;
    ram_cell[    4328] = 32'hf4b571ad;
    ram_cell[    4329] = 32'hdfe6ef56;
    ram_cell[    4330] = 32'he5fc757d;
    ram_cell[    4331] = 32'h9034d584;
    ram_cell[    4332] = 32'h26e1784e;
    ram_cell[    4333] = 32'h1de1663c;
    ram_cell[    4334] = 32'h6306920f;
    ram_cell[    4335] = 32'h17efd76f;
    ram_cell[    4336] = 32'h89c2da8b;
    ram_cell[    4337] = 32'hcda4e803;
    ram_cell[    4338] = 32'ha60e32b1;
    ram_cell[    4339] = 32'ha2686652;
    ram_cell[    4340] = 32'heba249bc;
    ram_cell[    4341] = 32'h3f52d358;
    ram_cell[    4342] = 32'hb5adeb2c;
    ram_cell[    4343] = 32'ha090ae84;
    ram_cell[    4344] = 32'h40360f30;
    ram_cell[    4345] = 32'hc553f21d;
    ram_cell[    4346] = 32'h9e01c576;
    ram_cell[    4347] = 32'hfb2a81a3;
    ram_cell[    4348] = 32'h0f9e0a3a;
    ram_cell[    4349] = 32'h023e4efc;
    ram_cell[    4350] = 32'hf1587e43;
    ram_cell[    4351] = 32'h449f42aa;
    ram_cell[    4352] = 32'h8b095b53;
    ram_cell[    4353] = 32'hcd1ed169;
    ram_cell[    4354] = 32'hdf47944c;
    ram_cell[    4355] = 32'hfca1d4d6;
    ram_cell[    4356] = 32'hffa64d75;
    ram_cell[    4357] = 32'h313ae481;
    ram_cell[    4358] = 32'h06c3202b;
    ram_cell[    4359] = 32'h42db5412;
    ram_cell[    4360] = 32'hd2aea796;
    ram_cell[    4361] = 32'h19df40e5;
    ram_cell[    4362] = 32'h4a1d3a66;
    ram_cell[    4363] = 32'hc12b038f;
    ram_cell[    4364] = 32'h2d4a3c53;
    ram_cell[    4365] = 32'h36c51fb9;
    ram_cell[    4366] = 32'h59e0a122;
    ram_cell[    4367] = 32'h4e7129e9;
    ram_cell[    4368] = 32'h15fcde2f;
    ram_cell[    4369] = 32'hc47ec6a3;
    ram_cell[    4370] = 32'h8a604ca9;
    ram_cell[    4371] = 32'ha10beafe;
    ram_cell[    4372] = 32'h17f65dd0;
    ram_cell[    4373] = 32'h4f0f7e68;
    ram_cell[    4374] = 32'h6f1deaa5;
    ram_cell[    4375] = 32'h5cc8de07;
    ram_cell[    4376] = 32'ha2a05ceb;
    ram_cell[    4377] = 32'h55b342f7;
    ram_cell[    4378] = 32'h796a44aa;
    ram_cell[    4379] = 32'h9b562f7a;
    ram_cell[    4380] = 32'hf5b73b38;
    ram_cell[    4381] = 32'h9f81655c;
    ram_cell[    4382] = 32'h41db9e49;
    ram_cell[    4383] = 32'h446f143d;
    ram_cell[    4384] = 32'h019ecdad;
    ram_cell[    4385] = 32'h5bda1342;
    ram_cell[    4386] = 32'h3ebb491f;
    ram_cell[    4387] = 32'h946addba;
    ram_cell[    4388] = 32'h98f028cf;
    ram_cell[    4389] = 32'h5412f37d;
    ram_cell[    4390] = 32'h03807507;
    ram_cell[    4391] = 32'h82dcf9a1;
    ram_cell[    4392] = 32'h543ca029;
    ram_cell[    4393] = 32'h4a9dd424;
    ram_cell[    4394] = 32'hf4fe7778;
    ram_cell[    4395] = 32'hbdceb64c;
    ram_cell[    4396] = 32'hf454b12f;
    ram_cell[    4397] = 32'hc4786cab;
    ram_cell[    4398] = 32'h3fa5aaee;
    ram_cell[    4399] = 32'h1fac4951;
    ram_cell[    4400] = 32'h44302f27;
    ram_cell[    4401] = 32'hb8a2154c;
    ram_cell[    4402] = 32'hb91708f0;
    ram_cell[    4403] = 32'hec72efde;
    ram_cell[    4404] = 32'h3cd9ae59;
    ram_cell[    4405] = 32'h44b6f48e;
    ram_cell[    4406] = 32'hb2ef7857;
    ram_cell[    4407] = 32'h3c365b32;
    ram_cell[    4408] = 32'h387bef87;
    ram_cell[    4409] = 32'h404fe091;
    ram_cell[    4410] = 32'h82f66881;
    ram_cell[    4411] = 32'he3165e7d;
    ram_cell[    4412] = 32'hd8f96afa;
    ram_cell[    4413] = 32'h20c4af3f;
    ram_cell[    4414] = 32'ha5ac6dbe;
    ram_cell[    4415] = 32'hdf824614;
    ram_cell[    4416] = 32'hf0189b0c;
    ram_cell[    4417] = 32'h97a0d56e;
    ram_cell[    4418] = 32'h4bf2acf7;
    ram_cell[    4419] = 32'h2904b43d;
    ram_cell[    4420] = 32'h9bfa4139;
    ram_cell[    4421] = 32'ha94af8a2;
    ram_cell[    4422] = 32'hf1d81f28;
    ram_cell[    4423] = 32'h4a837914;
    ram_cell[    4424] = 32'hfac1ecd5;
    ram_cell[    4425] = 32'h4a96297d;
    ram_cell[    4426] = 32'hf1d4fefb;
    ram_cell[    4427] = 32'h7a150d95;
    ram_cell[    4428] = 32'hf530b788;
    ram_cell[    4429] = 32'h5a1dde8b;
    ram_cell[    4430] = 32'hf8c40a5c;
    ram_cell[    4431] = 32'he2d7bb4d;
    ram_cell[    4432] = 32'h6d1c2925;
    ram_cell[    4433] = 32'h41309ea2;
    ram_cell[    4434] = 32'h387f43fe;
    ram_cell[    4435] = 32'h0ca607ec;
    ram_cell[    4436] = 32'h023d3350;
    ram_cell[    4437] = 32'h5ff2d266;
    ram_cell[    4438] = 32'h33e4158e;
    ram_cell[    4439] = 32'hb2e56341;
    ram_cell[    4440] = 32'hb25a1d58;
    ram_cell[    4441] = 32'hfa298ba4;
    ram_cell[    4442] = 32'h8307e99c;
    ram_cell[    4443] = 32'h7d138344;
    ram_cell[    4444] = 32'h0ea79908;
    ram_cell[    4445] = 32'hd28c1ae8;
    ram_cell[    4446] = 32'h59958e04;
    ram_cell[    4447] = 32'h19d0f1ad;
    ram_cell[    4448] = 32'h29097870;
    ram_cell[    4449] = 32'hdfd7b993;
    ram_cell[    4450] = 32'h8fd50304;
    ram_cell[    4451] = 32'h15b39bf3;
    ram_cell[    4452] = 32'h2cdb5cfe;
    ram_cell[    4453] = 32'h3cd9a0d2;
    ram_cell[    4454] = 32'h12f07e50;
    ram_cell[    4455] = 32'h60476e89;
    ram_cell[    4456] = 32'h5c32e599;
    ram_cell[    4457] = 32'h1c1d7305;
    ram_cell[    4458] = 32'hc068a479;
    ram_cell[    4459] = 32'hda1f97cf;
    ram_cell[    4460] = 32'hd1d606b2;
    ram_cell[    4461] = 32'h88abcf8b;
    ram_cell[    4462] = 32'h8c24a434;
    ram_cell[    4463] = 32'h05ffbafd;
    ram_cell[    4464] = 32'he9df612b;
    ram_cell[    4465] = 32'h1fa96c34;
    ram_cell[    4466] = 32'he07b1725;
    ram_cell[    4467] = 32'hb69cc487;
    ram_cell[    4468] = 32'h9338cee9;
    ram_cell[    4469] = 32'hbdd48d7d;
    ram_cell[    4470] = 32'he0ccfc3d;
    ram_cell[    4471] = 32'hefd758c6;
    ram_cell[    4472] = 32'h54f8ff0b;
    ram_cell[    4473] = 32'hc903df5d;
    ram_cell[    4474] = 32'h4d9bfa9e;
    ram_cell[    4475] = 32'h999462ea;
    ram_cell[    4476] = 32'h1eacef07;
    ram_cell[    4477] = 32'hf1af2f35;
    ram_cell[    4478] = 32'h367ccf00;
    ram_cell[    4479] = 32'h2e3ed72a;
    ram_cell[    4480] = 32'hd22fe504;
    ram_cell[    4481] = 32'ha568e8f2;
    ram_cell[    4482] = 32'h678fee98;
    ram_cell[    4483] = 32'hf2f180cb;
    ram_cell[    4484] = 32'hcfdeeff2;
    ram_cell[    4485] = 32'h9cf7c77d;
    ram_cell[    4486] = 32'h2d261ede;
    ram_cell[    4487] = 32'h87a1a852;
    ram_cell[    4488] = 32'h37e1518f;
    ram_cell[    4489] = 32'he445f520;
    ram_cell[    4490] = 32'h55b1e594;
    ram_cell[    4491] = 32'h3daf56d7;
    ram_cell[    4492] = 32'hd7d7ee97;
    ram_cell[    4493] = 32'h29a61451;
    ram_cell[    4494] = 32'h6f5ab722;
    ram_cell[    4495] = 32'hcd758a7e;
    ram_cell[    4496] = 32'hceecdc92;
    ram_cell[    4497] = 32'haf433b54;
    ram_cell[    4498] = 32'heb3aab19;
    ram_cell[    4499] = 32'h9eeaf84b;
    ram_cell[    4500] = 32'hee4098af;
    ram_cell[    4501] = 32'hfead47cf;
    ram_cell[    4502] = 32'ha2bcff4e;
    ram_cell[    4503] = 32'he87e2ba6;
    ram_cell[    4504] = 32'h48756be0;
    ram_cell[    4505] = 32'h0a28df16;
    ram_cell[    4506] = 32'hfec87be1;
    ram_cell[    4507] = 32'hd1125839;
    ram_cell[    4508] = 32'h0a31e122;
    ram_cell[    4509] = 32'h7ffc2570;
    ram_cell[    4510] = 32'h28c716f2;
    ram_cell[    4511] = 32'h5bf145d3;
    ram_cell[    4512] = 32'h5173bc1c;
    ram_cell[    4513] = 32'h087052eb;
    ram_cell[    4514] = 32'h51cab3ce;
    ram_cell[    4515] = 32'ha4402eaf;
    ram_cell[    4516] = 32'h4f0f32d3;
    ram_cell[    4517] = 32'hf9db9d39;
    ram_cell[    4518] = 32'h642ad752;
    ram_cell[    4519] = 32'hecaeb3be;
    ram_cell[    4520] = 32'hecaaa56f;
    ram_cell[    4521] = 32'h8a2fde03;
    ram_cell[    4522] = 32'h47767365;
    ram_cell[    4523] = 32'h6aa8e2d0;
    ram_cell[    4524] = 32'hc7672823;
    ram_cell[    4525] = 32'h5058cc39;
    ram_cell[    4526] = 32'h9f36017a;
    ram_cell[    4527] = 32'h0c2b5a03;
    ram_cell[    4528] = 32'h5934602b;
    ram_cell[    4529] = 32'hb230631b;
    ram_cell[    4530] = 32'h99b41c77;
    ram_cell[    4531] = 32'h703f3cd4;
    ram_cell[    4532] = 32'h349250b2;
    ram_cell[    4533] = 32'h83a4c3ca;
    ram_cell[    4534] = 32'h8bbb9c29;
    ram_cell[    4535] = 32'hb71a5dbd;
    ram_cell[    4536] = 32'hf7b1c639;
    ram_cell[    4537] = 32'hf22e65ed;
    ram_cell[    4538] = 32'hc9de0470;
    ram_cell[    4539] = 32'ha91b2300;
    ram_cell[    4540] = 32'h5c8427e1;
    ram_cell[    4541] = 32'hbd1d68a0;
    ram_cell[    4542] = 32'hfd60bd2c;
    ram_cell[    4543] = 32'h4708ce0b;
    ram_cell[    4544] = 32'haadd7828;
    ram_cell[    4545] = 32'ha81c8bce;
    ram_cell[    4546] = 32'hd49dc329;
    ram_cell[    4547] = 32'h97a44aee;
    ram_cell[    4548] = 32'h0df5f455;
    ram_cell[    4549] = 32'h61c8fd0d;
    ram_cell[    4550] = 32'ha48a5c60;
    ram_cell[    4551] = 32'h2ad3601f;
    ram_cell[    4552] = 32'h8c14d288;
    ram_cell[    4553] = 32'h45747c13;
    ram_cell[    4554] = 32'ha96d0cf5;
    ram_cell[    4555] = 32'h1469fb7c;
    ram_cell[    4556] = 32'hc55e60af;
    ram_cell[    4557] = 32'h8f1d903f;
    ram_cell[    4558] = 32'hf36513c4;
    ram_cell[    4559] = 32'hde68a8c6;
    ram_cell[    4560] = 32'h0757239c;
    ram_cell[    4561] = 32'hf237f059;
    ram_cell[    4562] = 32'hbd38ff0e;
    ram_cell[    4563] = 32'hc63f0cca;
    ram_cell[    4564] = 32'h54473e40;
    ram_cell[    4565] = 32'h1698cfa4;
    ram_cell[    4566] = 32'h6c497693;
    ram_cell[    4567] = 32'h2b98fde4;
    ram_cell[    4568] = 32'he4430b68;
    ram_cell[    4569] = 32'h91916767;
    ram_cell[    4570] = 32'h4ab6ad8f;
    ram_cell[    4571] = 32'h149d53bb;
    ram_cell[    4572] = 32'h11c7be49;
    ram_cell[    4573] = 32'h06a749ab;
    ram_cell[    4574] = 32'hbd6c15e0;
    ram_cell[    4575] = 32'hb43981f8;
    ram_cell[    4576] = 32'h278a578e;
    ram_cell[    4577] = 32'h046fadb2;
    ram_cell[    4578] = 32'h76030350;
    ram_cell[    4579] = 32'hee57f8e7;
    ram_cell[    4580] = 32'h5e7f79f8;
    ram_cell[    4581] = 32'h916d1426;
    ram_cell[    4582] = 32'hb75505ce;
    ram_cell[    4583] = 32'h1ac4aed8;
    ram_cell[    4584] = 32'hba56803e;
    ram_cell[    4585] = 32'hcf6bf28e;
    ram_cell[    4586] = 32'hefb11fe9;
    ram_cell[    4587] = 32'h33b6a84f;
    ram_cell[    4588] = 32'h4c6b2716;
    ram_cell[    4589] = 32'h722f3434;
    ram_cell[    4590] = 32'h6c1f2a5b;
    ram_cell[    4591] = 32'h84314f2c;
    ram_cell[    4592] = 32'h0972ebf8;
    ram_cell[    4593] = 32'hc6186669;
    ram_cell[    4594] = 32'hf5834dcd;
    ram_cell[    4595] = 32'h5d470dff;
    ram_cell[    4596] = 32'h002d4a0d;
    ram_cell[    4597] = 32'hcdcdf35f;
    ram_cell[    4598] = 32'h0bfe37ed;
    ram_cell[    4599] = 32'hf7d12c58;
    ram_cell[    4600] = 32'haee2172a;
    ram_cell[    4601] = 32'h98ef0c00;
    ram_cell[    4602] = 32'h9fe6c30b;
    ram_cell[    4603] = 32'h25c771ee;
    ram_cell[    4604] = 32'h516064bb;
    ram_cell[    4605] = 32'hab41568e;
    ram_cell[    4606] = 32'h09ffa993;
    ram_cell[    4607] = 32'hbf4b4313;
    ram_cell[    4608] = 32'hcf0f45b4;
    ram_cell[    4609] = 32'hd1b18f95;
    ram_cell[    4610] = 32'h8f874e02;
    ram_cell[    4611] = 32'h6f20039c;
    ram_cell[    4612] = 32'ha182e71e;
    ram_cell[    4613] = 32'h5c02cefb;
    ram_cell[    4614] = 32'hd630a070;
    ram_cell[    4615] = 32'he59b460d;
    ram_cell[    4616] = 32'h7ea79413;
    ram_cell[    4617] = 32'h43c4b76b;
    ram_cell[    4618] = 32'h6d06a2d8;
    ram_cell[    4619] = 32'h82a9d32e;
    ram_cell[    4620] = 32'hb9230d6e;
    ram_cell[    4621] = 32'hecf9312c;
    ram_cell[    4622] = 32'h0d7d6174;
    ram_cell[    4623] = 32'h62c9029e;
    ram_cell[    4624] = 32'hcf4f7aac;
    ram_cell[    4625] = 32'h815b772a;
    ram_cell[    4626] = 32'h3cddd093;
    ram_cell[    4627] = 32'h3a6ff2b6;
    ram_cell[    4628] = 32'h34d09c73;
    ram_cell[    4629] = 32'h65b572ea;
    ram_cell[    4630] = 32'ha7a38c71;
    ram_cell[    4631] = 32'h998548d9;
    ram_cell[    4632] = 32'h0ba1bbfc;
    ram_cell[    4633] = 32'hc1506d01;
    ram_cell[    4634] = 32'h0acaf279;
    ram_cell[    4635] = 32'hbd27f8a9;
    ram_cell[    4636] = 32'he1ffd763;
    ram_cell[    4637] = 32'h72c633df;
    ram_cell[    4638] = 32'h0fa53f0b;
    ram_cell[    4639] = 32'h3b386047;
    ram_cell[    4640] = 32'hb456f058;
    ram_cell[    4641] = 32'hf3cee5e5;
    ram_cell[    4642] = 32'h410cb5f9;
    ram_cell[    4643] = 32'h9f541dcf;
    ram_cell[    4644] = 32'h0bbc9672;
    ram_cell[    4645] = 32'h81d2e43c;
    ram_cell[    4646] = 32'h93a0628f;
    ram_cell[    4647] = 32'haec3a59e;
    ram_cell[    4648] = 32'h6990cf0e;
    ram_cell[    4649] = 32'h29647aea;
    ram_cell[    4650] = 32'h6d4fe09f;
    ram_cell[    4651] = 32'hd0b82dc6;
    ram_cell[    4652] = 32'h2950e839;
    ram_cell[    4653] = 32'h6a162ee8;
    ram_cell[    4654] = 32'heea882fa;
    ram_cell[    4655] = 32'h9a9f6360;
    ram_cell[    4656] = 32'h00c4fe1e;
    ram_cell[    4657] = 32'hf86f1fcd;
    ram_cell[    4658] = 32'h9ad787ff;
    ram_cell[    4659] = 32'hd15ba2c7;
    ram_cell[    4660] = 32'h9077f5bb;
    ram_cell[    4661] = 32'h276971e7;
    ram_cell[    4662] = 32'h5019638e;
    ram_cell[    4663] = 32'h891d35bd;
    ram_cell[    4664] = 32'h17552504;
    ram_cell[    4665] = 32'h924740e4;
    ram_cell[    4666] = 32'h2dcd0d76;
    ram_cell[    4667] = 32'h86f21de4;
    ram_cell[    4668] = 32'h81d6dd8a;
    ram_cell[    4669] = 32'h6e4aba4f;
    ram_cell[    4670] = 32'h96b838c6;
    ram_cell[    4671] = 32'h6b275eaa;
    ram_cell[    4672] = 32'hbd631008;
    ram_cell[    4673] = 32'hef103383;
    ram_cell[    4674] = 32'h6c75f71c;
    ram_cell[    4675] = 32'h489f7361;
    ram_cell[    4676] = 32'h000bc2a6;
    ram_cell[    4677] = 32'h2cc1ceb2;
    ram_cell[    4678] = 32'h23a2eee2;
    ram_cell[    4679] = 32'hb327ca62;
    ram_cell[    4680] = 32'h463afce9;
    ram_cell[    4681] = 32'hf1890fa1;
    ram_cell[    4682] = 32'hd2fca4bf;
    ram_cell[    4683] = 32'h6ab9fab5;
    ram_cell[    4684] = 32'h8d44d080;
    ram_cell[    4685] = 32'h7ddf9d86;
    ram_cell[    4686] = 32'h24b43dae;
    ram_cell[    4687] = 32'h173b987c;
    ram_cell[    4688] = 32'h67fe2d38;
    ram_cell[    4689] = 32'hbf310b37;
    ram_cell[    4690] = 32'h96866100;
    ram_cell[    4691] = 32'hd5a5cd97;
    ram_cell[    4692] = 32'he4a2a8d1;
    ram_cell[    4693] = 32'h3ce6872d;
    ram_cell[    4694] = 32'h0b23f8e9;
    ram_cell[    4695] = 32'h42f5e893;
    ram_cell[    4696] = 32'haa86579d;
    ram_cell[    4697] = 32'hf309e6d0;
    ram_cell[    4698] = 32'hfde04eb9;
    ram_cell[    4699] = 32'h2b4393a5;
    ram_cell[    4700] = 32'h13cdaa24;
    ram_cell[    4701] = 32'h1079db29;
    ram_cell[    4702] = 32'h22d80311;
    ram_cell[    4703] = 32'h58176135;
    ram_cell[    4704] = 32'h797b73b3;
    ram_cell[    4705] = 32'h691adbff;
    ram_cell[    4706] = 32'hc6dd9b57;
    ram_cell[    4707] = 32'h2fa986ad;
    ram_cell[    4708] = 32'hdb248926;
    ram_cell[    4709] = 32'h1b3b594b;
    ram_cell[    4710] = 32'h1401bb75;
    ram_cell[    4711] = 32'hf09051ff;
    ram_cell[    4712] = 32'he91cbcad;
    ram_cell[    4713] = 32'h62d6805e;
    ram_cell[    4714] = 32'hadac7450;
    ram_cell[    4715] = 32'h9b15b741;
    ram_cell[    4716] = 32'h451a9126;
    ram_cell[    4717] = 32'hd0e446d8;
    ram_cell[    4718] = 32'h8c67298d;
    ram_cell[    4719] = 32'hd91ab679;
    ram_cell[    4720] = 32'h25c9689c;
    ram_cell[    4721] = 32'h7e992906;
    ram_cell[    4722] = 32'h5a098fdd;
    ram_cell[    4723] = 32'h92d2ce68;
    ram_cell[    4724] = 32'h06f8f8b5;
    ram_cell[    4725] = 32'h80e18419;
    ram_cell[    4726] = 32'h58ecc64f;
    ram_cell[    4727] = 32'h769e7561;
    ram_cell[    4728] = 32'hc978745d;
    ram_cell[    4729] = 32'heba2503c;
    ram_cell[    4730] = 32'h2ff11c55;
    ram_cell[    4731] = 32'h2959eb3f;
    ram_cell[    4732] = 32'hdd08853e;
    ram_cell[    4733] = 32'h475c15e6;
    ram_cell[    4734] = 32'hced413a6;
    ram_cell[    4735] = 32'h8f0f8e56;
    ram_cell[    4736] = 32'h19a97341;
    ram_cell[    4737] = 32'h10dbb7ca;
    ram_cell[    4738] = 32'hd12ad4f5;
    ram_cell[    4739] = 32'hbe0feb72;
    ram_cell[    4740] = 32'h8218dd6a;
    ram_cell[    4741] = 32'hdf68ec51;
    ram_cell[    4742] = 32'h0b85b2e1;
    ram_cell[    4743] = 32'h851584a2;
    ram_cell[    4744] = 32'h3887f59f;
    ram_cell[    4745] = 32'h054389f3;
    ram_cell[    4746] = 32'h10018331;
    ram_cell[    4747] = 32'h70ff395e;
    ram_cell[    4748] = 32'h423bc6cf;
    ram_cell[    4749] = 32'he5b24d9d;
    ram_cell[    4750] = 32'h8db47d68;
    ram_cell[    4751] = 32'hb806a86f;
    ram_cell[    4752] = 32'h41c48b8f;
    ram_cell[    4753] = 32'ha337b6db;
    ram_cell[    4754] = 32'h05dcc055;
    ram_cell[    4755] = 32'h01e59ab8;
    ram_cell[    4756] = 32'h24c2ad69;
    ram_cell[    4757] = 32'hd83a0ffd;
    ram_cell[    4758] = 32'h748d7b99;
    ram_cell[    4759] = 32'hde4988ec;
    ram_cell[    4760] = 32'h58af2f0c;
    ram_cell[    4761] = 32'h16a1ba33;
    ram_cell[    4762] = 32'h7b5ec376;
    ram_cell[    4763] = 32'h4d98a7e9;
    ram_cell[    4764] = 32'h10839276;
    ram_cell[    4765] = 32'hc150f302;
    ram_cell[    4766] = 32'h759e8d0b;
    ram_cell[    4767] = 32'hcb2c887c;
    ram_cell[    4768] = 32'h80acb91d;
    ram_cell[    4769] = 32'h9ddc73d7;
    ram_cell[    4770] = 32'ha8ed4cbc;
    ram_cell[    4771] = 32'h8be0a237;
    ram_cell[    4772] = 32'h74d40ac2;
    ram_cell[    4773] = 32'h02bfd71a;
    ram_cell[    4774] = 32'h93f25651;
    ram_cell[    4775] = 32'hbcc7b6c2;
    ram_cell[    4776] = 32'h45b3242b;
    ram_cell[    4777] = 32'h8fcefd75;
    ram_cell[    4778] = 32'h625b62ac;
    ram_cell[    4779] = 32'hd8a9a7be;
    ram_cell[    4780] = 32'h40757058;
    ram_cell[    4781] = 32'h0084ac39;
    ram_cell[    4782] = 32'h08906c84;
    ram_cell[    4783] = 32'h3bcc9715;
    ram_cell[    4784] = 32'h26a30a2a;
    ram_cell[    4785] = 32'hc4914c38;
    ram_cell[    4786] = 32'hd7e2f8be;
    ram_cell[    4787] = 32'h4d3581f3;
    ram_cell[    4788] = 32'hd35e00e2;
    ram_cell[    4789] = 32'h89411fb1;
    ram_cell[    4790] = 32'h4d1fabe0;
    ram_cell[    4791] = 32'hdc8d5142;
    ram_cell[    4792] = 32'hfe566111;
    ram_cell[    4793] = 32'hf211fbd9;
    ram_cell[    4794] = 32'h4e747e6e;
    ram_cell[    4795] = 32'h8446ee9b;
    ram_cell[    4796] = 32'h8f53443f;
    ram_cell[    4797] = 32'h6ed1188d;
    ram_cell[    4798] = 32'h1d57854c;
    ram_cell[    4799] = 32'hc2e7a6bb;
    ram_cell[    4800] = 32'h0678b68a;
    ram_cell[    4801] = 32'hb1002906;
    ram_cell[    4802] = 32'hd4f6407f;
    ram_cell[    4803] = 32'h14545b6b;
    ram_cell[    4804] = 32'h5774df77;
    ram_cell[    4805] = 32'hc35f5f1a;
    ram_cell[    4806] = 32'ha689ca38;
    ram_cell[    4807] = 32'he35454fd;
    ram_cell[    4808] = 32'h929ff7a2;
    ram_cell[    4809] = 32'h8c3399bf;
    ram_cell[    4810] = 32'hea41fff0;
    ram_cell[    4811] = 32'he917599b;
    ram_cell[    4812] = 32'h7c49f7f4;
    ram_cell[    4813] = 32'h6e9145a7;
    ram_cell[    4814] = 32'h79739f4b;
    ram_cell[    4815] = 32'hff98cabe;
    ram_cell[    4816] = 32'h3e25bd1a;
    ram_cell[    4817] = 32'hc8320fa7;
    ram_cell[    4818] = 32'h1acc9317;
    ram_cell[    4819] = 32'h80900bde;
    ram_cell[    4820] = 32'h5a5b8d12;
    ram_cell[    4821] = 32'h42f84ce1;
    ram_cell[    4822] = 32'h581e5e7b;
    ram_cell[    4823] = 32'h23cc051d;
    ram_cell[    4824] = 32'h817293cc;
    ram_cell[    4825] = 32'hf7fe50ff;
    ram_cell[    4826] = 32'hc29e0a6e;
    ram_cell[    4827] = 32'h8bd42f4f;
    ram_cell[    4828] = 32'h96c72cdc;
    ram_cell[    4829] = 32'h4f36e44f;
    ram_cell[    4830] = 32'h941e2ad4;
    ram_cell[    4831] = 32'h8fab3a0f;
    ram_cell[    4832] = 32'h31c428e8;
    ram_cell[    4833] = 32'hb0c650aa;
    ram_cell[    4834] = 32'h4fe0f073;
    ram_cell[    4835] = 32'heea3571e;
    ram_cell[    4836] = 32'h43e74553;
    ram_cell[    4837] = 32'h2b014d49;
    ram_cell[    4838] = 32'hea5e467a;
    ram_cell[    4839] = 32'hbdd37ae9;
    ram_cell[    4840] = 32'h439b4b7e;
    ram_cell[    4841] = 32'h856cfa24;
    ram_cell[    4842] = 32'h84a581cd;
    ram_cell[    4843] = 32'hed030317;
    ram_cell[    4844] = 32'hf96a6602;
    ram_cell[    4845] = 32'h6dea2892;
    ram_cell[    4846] = 32'hfb866651;
    ram_cell[    4847] = 32'h4674c7d4;
    ram_cell[    4848] = 32'ha216eade;
    ram_cell[    4849] = 32'hf36a36c8;
    ram_cell[    4850] = 32'hd5d53ed0;
    ram_cell[    4851] = 32'hd1dcfbd2;
    ram_cell[    4852] = 32'h3fe1047f;
    ram_cell[    4853] = 32'h9ac640cd;
    ram_cell[    4854] = 32'h38c0e3a9;
    ram_cell[    4855] = 32'h7acc20d5;
    ram_cell[    4856] = 32'h922a91cf;
    ram_cell[    4857] = 32'hb65fb1b6;
    ram_cell[    4858] = 32'h89e46dfa;
    ram_cell[    4859] = 32'h0ccc18e2;
    ram_cell[    4860] = 32'he2ad8eb6;
    ram_cell[    4861] = 32'h61533831;
    ram_cell[    4862] = 32'h6d5803de;
    ram_cell[    4863] = 32'h638c3919;
    ram_cell[    4864] = 32'h788f295a;
    ram_cell[    4865] = 32'h5028c41b;
    ram_cell[    4866] = 32'hddf64622;
    ram_cell[    4867] = 32'hc3d373b0;
    ram_cell[    4868] = 32'h140211e9;
    ram_cell[    4869] = 32'h778bf93b;
    ram_cell[    4870] = 32'h1ecb2ed1;
    ram_cell[    4871] = 32'h838811ae;
    ram_cell[    4872] = 32'h501061c3;
    ram_cell[    4873] = 32'hf9a05fa0;
    ram_cell[    4874] = 32'haa59c686;
    ram_cell[    4875] = 32'hbfdfca0b;
    ram_cell[    4876] = 32'h7ad9a0a8;
    ram_cell[    4877] = 32'hcda5b896;
    ram_cell[    4878] = 32'h3caabc80;
    ram_cell[    4879] = 32'h937faa57;
    ram_cell[    4880] = 32'h5f7778ed;
    ram_cell[    4881] = 32'h96eac543;
    ram_cell[    4882] = 32'h1e7f3684;
    ram_cell[    4883] = 32'h838f9d40;
    ram_cell[    4884] = 32'hf2bba52a;
    ram_cell[    4885] = 32'h7588c87f;
    ram_cell[    4886] = 32'hb39c4e94;
    ram_cell[    4887] = 32'h7c0c79f8;
    ram_cell[    4888] = 32'hdd7c9205;
    ram_cell[    4889] = 32'h86c7d453;
    ram_cell[    4890] = 32'h0f4fa2ab;
    ram_cell[    4891] = 32'h40b6fc78;
    ram_cell[    4892] = 32'he0e7bc0b;
    ram_cell[    4893] = 32'he40e5a98;
    ram_cell[    4894] = 32'h84bcfed7;
    ram_cell[    4895] = 32'hf023390f;
    ram_cell[    4896] = 32'h6c3a6a71;
    ram_cell[    4897] = 32'hde3243ae;
    ram_cell[    4898] = 32'hae7211fe;
    ram_cell[    4899] = 32'hf786fe87;
    ram_cell[    4900] = 32'h9531fd16;
    ram_cell[    4901] = 32'ha2a2cb5c;
    ram_cell[    4902] = 32'hbba3f0a3;
    ram_cell[    4903] = 32'h0f255c21;
    ram_cell[    4904] = 32'h8e0e0723;
    ram_cell[    4905] = 32'h05ada4ea;
    ram_cell[    4906] = 32'hdecb7c83;
    ram_cell[    4907] = 32'h96190cfb;
    ram_cell[    4908] = 32'h6867b6cc;
    ram_cell[    4909] = 32'h67bcddf6;
    ram_cell[    4910] = 32'h419cb468;
    ram_cell[    4911] = 32'h521ce81e;
    ram_cell[    4912] = 32'h02bb2e47;
    ram_cell[    4913] = 32'hfbac7e60;
    ram_cell[    4914] = 32'hcb921a47;
    ram_cell[    4915] = 32'hc4c316bf;
    ram_cell[    4916] = 32'he9362eb7;
    ram_cell[    4917] = 32'haa5dd6cc;
    ram_cell[    4918] = 32'h878e5a87;
    ram_cell[    4919] = 32'h5d27b664;
    ram_cell[    4920] = 32'habe75c31;
    ram_cell[    4921] = 32'h23a14215;
    ram_cell[    4922] = 32'hb6fa7935;
    ram_cell[    4923] = 32'h3a13f6e3;
    ram_cell[    4924] = 32'ha80a2326;
    ram_cell[    4925] = 32'h1f15f7ec;
    ram_cell[    4926] = 32'hccf7af4a;
    ram_cell[    4927] = 32'h130c466d;
    ram_cell[    4928] = 32'hcfc44887;
    ram_cell[    4929] = 32'h9f5cf1a9;
    ram_cell[    4930] = 32'h5dc18fe4;
    ram_cell[    4931] = 32'hfcdaf356;
    ram_cell[    4932] = 32'hc4c1e918;
    ram_cell[    4933] = 32'h9c30a3a3;
    ram_cell[    4934] = 32'hfd7b9f8d;
    ram_cell[    4935] = 32'h9d7d4ea6;
    ram_cell[    4936] = 32'h4ec874aa;
    ram_cell[    4937] = 32'h776b00d8;
    ram_cell[    4938] = 32'h09e53a8b;
    ram_cell[    4939] = 32'hbd2e4531;
    ram_cell[    4940] = 32'hd6e77de0;
    ram_cell[    4941] = 32'h1848a1c9;
    ram_cell[    4942] = 32'h1351abda;
    ram_cell[    4943] = 32'hf0164ab5;
    ram_cell[    4944] = 32'h3c7ce7f8;
    ram_cell[    4945] = 32'hb945a742;
    ram_cell[    4946] = 32'ha42d4305;
    ram_cell[    4947] = 32'he84eb251;
    ram_cell[    4948] = 32'h4aa34ba0;
    ram_cell[    4949] = 32'hb2f5131e;
    ram_cell[    4950] = 32'h2852bc48;
    ram_cell[    4951] = 32'h5daeab1d;
    ram_cell[    4952] = 32'hd592ba1f;
    ram_cell[    4953] = 32'h4f0760f2;
    ram_cell[    4954] = 32'h42c67c7b;
    ram_cell[    4955] = 32'hcc19304d;
    ram_cell[    4956] = 32'h2e29fdd7;
    ram_cell[    4957] = 32'h30f5164a;
    ram_cell[    4958] = 32'hc2c12dd5;
    ram_cell[    4959] = 32'he1dbd793;
    ram_cell[    4960] = 32'h42a9411b;
    ram_cell[    4961] = 32'hc770fae0;
    ram_cell[    4962] = 32'h8193311e;
    ram_cell[    4963] = 32'h1f32b799;
    ram_cell[    4964] = 32'hd445fa01;
    ram_cell[    4965] = 32'h2ccf4486;
    ram_cell[    4966] = 32'h7a80c0c2;
    ram_cell[    4967] = 32'haad456c2;
    ram_cell[    4968] = 32'hc3e6f7c5;
    ram_cell[    4969] = 32'h515b148d;
    ram_cell[    4970] = 32'hfe6c6d71;
    ram_cell[    4971] = 32'hb8e335ef;
    ram_cell[    4972] = 32'hec4f3861;
    ram_cell[    4973] = 32'hceea3313;
    ram_cell[    4974] = 32'h75536816;
    ram_cell[    4975] = 32'h515e4733;
    ram_cell[    4976] = 32'h55ff4dbc;
    ram_cell[    4977] = 32'h7b87612a;
    ram_cell[    4978] = 32'h913284cf;
    ram_cell[    4979] = 32'h7589f4b3;
    ram_cell[    4980] = 32'hb177a948;
    ram_cell[    4981] = 32'h0aa4ac9e;
    ram_cell[    4982] = 32'h14da236a;
    ram_cell[    4983] = 32'h0f04c66f;
    ram_cell[    4984] = 32'hd29777cf;
    ram_cell[    4985] = 32'h044ab02b;
    ram_cell[    4986] = 32'h0969ee88;
    ram_cell[    4987] = 32'hc62fbcac;
    ram_cell[    4988] = 32'hce5ad717;
    ram_cell[    4989] = 32'h4571f9bd;
    ram_cell[    4990] = 32'h3bfa3650;
    ram_cell[    4991] = 32'h275b0be0;
    ram_cell[    4992] = 32'hcbe18ee9;
    ram_cell[    4993] = 32'h387e2833;
    ram_cell[    4994] = 32'h4f888004;
    ram_cell[    4995] = 32'hbb81f935;
    ram_cell[    4996] = 32'hf476d86d;
    ram_cell[    4997] = 32'ha197d54d;
    ram_cell[    4998] = 32'h1c9e154d;
    ram_cell[    4999] = 32'h9020cede;
    ram_cell[    5000] = 32'h16455019;
    ram_cell[    5001] = 32'hecc763a3;
    ram_cell[    5002] = 32'hb576bc78;
    ram_cell[    5003] = 32'h7ebba805;
    ram_cell[    5004] = 32'h4c56965f;
    ram_cell[    5005] = 32'h536a7114;
    ram_cell[    5006] = 32'hbb85794b;
    ram_cell[    5007] = 32'h7257b5c4;
    ram_cell[    5008] = 32'h4a46c611;
    ram_cell[    5009] = 32'h3cebd57b;
    ram_cell[    5010] = 32'he7b6dd76;
    ram_cell[    5011] = 32'ha6a99f59;
    ram_cell[    5012] = 32'hdd2b487c;
    ram_cell[    5013] = 32'h2f8c0fd5;
    ram_cell[    5014] = 32'hbe55d15f;
    ram_cell[    5015] = 32'hcb338ce6;
    ram_cell[    5016] = 32'hc79780f5;
    ram_cell[    5017] = 32'h98e24c4c;
    ram_cell[    5018] = 32'ha8dfdc85;
    ram_cell[    5019] = 32'hca551981;
    ram_cell[    5020] = 32'h09fb68ec;
    ram_cell[    5021] = 32'hf703f2e4;
    ram_cell[    5022] = 32'h6b5769c7;
    ram_cell[    5023] = 32'hde25a0cb;
    ram_cell[    5024] = 32'h8a5b3ef0;
    ram_cell[    5025] = 32'h17f48db9;
    ram_cell[    5026] = 32'h01fa1f3b;
    ram_cell[    5027] = 32'hc46dc74e;
    ram_cell[    5028] = 32'he5701d12;
    ram_cell[    5029] = 32'hf574093c;
    ram_cell[    5030] = 32'hddd5befc;
    ram_cell[    5031] = 32'h2ad3f07e;
    ram_cell[    5032] = 32'hfabfd0e4;
    ram_cell[    5033] = 32'hbe494425;
    ram_cell[    5034] = 32'hd6e726f1;
    ram_cell[    5035] = 32'h359e9858;
    ram_cell[    5036] = 32'h4dad149c;
    ram_cell[    5037] = 32'h5d4ac70b;
    ram_cell[    5038] = 32'h1167b620;
    ram_cell[    5039] = 32'h661ea60b;
    ram_cell[    5040] = 32'h21f4d37e;
    ram_cell[    5041] = 32'hd17f233c;
    ram_cell[    5042] = 32'h023afd09;
    ram_cell[    5043] = 32'h5aecbb1f;
    ram_cell[    5044] = 32'h2a3fbeea;
    ram_cell[    5045] = 32'h423def9a;
    ram_cell[    5046] = 32'h0872b378;
    ram_cell[    5047] = 32'hf3b5597d;
    ram_cell[    5048] = 32'haa368225;
    ram_cell[    5049] = 32'h921d9b56;
    ram_cell[    5050] = 32'hfdd87321;
    ram_cell[    5051] = 32'h7fdf0cc3;
    ram_cell[    5052] = 32'h3d5fb426;
    ram_cell[    5053] = 32'h24b41e62;
    ram_cell[    5054] = 32'h43b1dcaf;
    ram_cell[    5055] = 32'h030b8d77;
    ram_cell[    5056] = 32'h709b78f5;
    ram_cell[    5057] = 32'hc99e10b1;
    ram_cell[    5058] = 32'h48f8fca4;
    ram_cell[    5059] = 32'h8a048f3f;
    ram_cell[    5060] = 32'hfec47239;
    ram_cell[    5061] = 32'h1e15320f;
    ram_cell[    5062] = 32'hd77d507b;
    ram_cell[    5063] = 32'hbf3279ac;
    ram_cell[    5064] = 32'h220887dd;
    ram_cell[    5065] = 32'hca5b0af2;
    ram_cell[    5066] = 32'h49eb92b2;
    ram_cell[    5067] = 32'h550155ce;
    ram_cell[    5068] = 32'h7817f982;
    ram_cell[    5069] = 32'h1bf09222;
    ram_cell[    5070] = 32'had0213c7;
    ram_cell[    5071] = 32'h97ae4c75;
    ram_cell[    5072] = 32'h24ba98f1;
    ram_cell[    5073] = 32'h3de07552;
    ram_cell[    5074] = 32'hb340cba6;
    ram_cell[    5075] = 32'h7ab5221b;
    ram_cell[    5076] = 32'h0776bf63;
    ram_cell[    5077] = 32'h81b3b46d;
    ram_cell[    5078] = 32'h61a0288b;
    ram_cell[    5079] = 32'h947922f1;
    ram_cell[    5080] = 32'h48e164f3;
    ram_cell[    5081] = 32'hcc8bfe2b;
    ram_cell[    5082] = 32'h2812fea7;
    ram_cell[    5083] = 32'hd4fe67bb;
    ram_cell[    5084] = 32'h21a4a0ca;
    ram_cell[    5085] = 32'hb93aeb08;
    ram_cell[    5086] = 32'hec6032d0;
    ram_cell[    5087] = 32'h706fb04e;
    ram_cell[    5088] = 32'h2f15d798;
    ram_cell[    5089] = 32'h9ecd695d;
    ram_cell[    5090] = 32'h2f829ae1;
    ram_cell[    5091] = 32'h39938f4b;
    ram_cell[    5092] = 32'h06746ad1;
    ram_cell[    5093] = 32'hddb26b61;
    ram_cell[    5094] = 32'h6d4fad88;
    ram_cell[    5095] = 32'hb5a58035;
    ram_cell[    5096] = 32'hf2ac6205;
    ram_cell[    5097] = 32'hde3aae6d;
    ram_cell[    5098] = 32'ha23c83de;
    ram_cell[    5099] = 32'h0b962481;
    ram_cell[    5100] = 32'h2f342099;
    ram_cell[    5101] = 32'h38b5deff;
    ram_cell[    5102] = 32'h48fe9f11;
    ram_cell[    5103] = 32'hbef5bdd0;
    ram_cell[    5104] = 32'h3a4515cc;
    ram_cell[    5105] = 32'h921946b8;
    ram_cell[    5106] = 32'h41f79908;
    ram_cell[    5107] = 32'h12b0efe3;
    ram_cell[    5108] = 32'hb214d804;
    ram_cell[    5109] = 32'h29da67a0;
    ram_cell[    5110] = 32'he85e4e3c;
    ram_cell[    5111] = 32'h8d7ffd07;
    ram_cell[    5112] = 32'h6cf78e8d;
    ram_cell[    5113] = 32'h5bcfb065;
    ram_cell[    5114] = 32'h4a0e1e4c;
    ram_cell[    5115] = 32'h4919d25f;
    ram_cell[    5116] = 32'ha027b551;
    ram_cell[    5117] = 32'hf6a77b95;
    ram_cell[    5118] = 32'h0a8e021f;
    ram_cell[    5119] = 32'h9376e658;
    ram_cell[    5120] = 32'h95b690e7;
    ram_cell[    5121] = 32'h059bee8f;
    ram_cell[    5122] = 32'hbec276b8;
    ram_cell[    5123] = 32'h5c1d7691;
    ram_cell[    5124] = 32'h372a11ac;
    ram_cell[    5125] = 32'hd2f12264;
    ram_cell[    5126] = 32'hfba3c157;
    ram_cell[    5127] = 32'hcc06301a;
    ram_cell[    5128] = 32'hb905fd2b;
    ram_cell[    5129] = 32'hcc3ac199;
    ram_cell[    5130] = 32'he0659d40;
    ram_cell[    5131] = 32'h908ec45f;
    ram_cell[    5132] = 32'h326e19ab;
    ram_cell[    5133] = 32'h49b0c854;
    ram_cell[    5134] = 32'h85a2663f;
    ram_cell[    5135] = 32'h5e032189;
    ram_cell[    5136] = 32'hca8b4fb2;
    ram_cell[    5137] = 32'hcbc71ac0;
    ram_cell[    5138] = 32'h1dc37053;
    ram_cell[    5139] = 32'h706d1757;
    ram_cell[    5140] = 32'hf50229c1;
    ram_cell[    5141] = 32'ha610b5c0;
    ram_cell[    5142] = 32'hc2b0ebf0;
    ram_cell[    5143] = 32'h9e8dc923;
    ram_cell[    5144] = 32'h143b9be6;
    ram_cell[    5145] = 32'ha83a131f;
    ram_cell[    5146] = 32'h328e6d31;
    ram_cell[    5147] = 32'h3cf760c0;
    ram_cell[    5148] = 32'hac47a8a4;
    ram_cell[    5149] = 32'h29eba46a;
    ram_cell[    5150] = 32'hf69fecda;
    ram_cell[    5151] = 32'hc42a9952;
    ram_cell[    5152] = 32'hdf02b1da;
    ram_cell[    5153] = 32'h8faa0d0d;
    ram_cell[    5154] = 32'hade43e26;
    ram_cell[    5155] = 32'h50743658;
    ram_cell[    5156] = 32'hd9354b12;
    ram_cell[    5157] = 32'h8176d571;
    ram_cell[    5158] = 32'ha757b7e7;
    ram_cell[    5159] = 32'h8de1a398;
    ram_cell[    5160] = 32'ha9362655;
    ram_cell[    5161] = 32'h599ffff0;
    ram_cell[    5162] = 32'h4d70ed2b;
    ram_cell[    5163] = 32'he5b5aa84;
    ram_cell[    5164] = 32'h1bb3346d;
    ram_cell[    5165] = 32'hfcff678c;
    ram_cell[    5166] = 32'ha5c64af8;
    ram_cell[    5167] = 32'hb885084e;
    ram_cell[    5168] = 32'h61487a13;
    ram_cell[    5169] = 32'he28a4501;
    ram_cell[    5170] = 32'h255a9ab9;
    ram_cell[    5171] = 32'he40fa6b7;
    ram_cell[    5172] = 32'hf1fdbe24;
    ram_cell[    5173] = 32'hb5c0ba9a;
    ram_cell[    5174] = 32'hf94a295a;
    ram_cell[    5175] = 32'h8ef03fc6;
    ram_cell[    5176] = 32'hb100e04c;
    ram_cell[    5177] = 32'h3ab05384;
    ram_cell[    5178] = 32'h757b940e;
    ram_cell[    5179] = 32'h6b5449e5;
    ram_cell[    5180] = 32'hd077f69f;
    ram_cell[    5181] = 32'h62ab9568;
    ram_cell[    5182] = 32'ha4baf259;
    ram_cell[    5183] = 32'h7cb36cd4;
    ram_cell[    5184] = 32'h7e7e0c6a;
    ram_cell[    5185] = 32'hf0d75cf1;
    ram_cell[    5186] = 32'h52b07d64;
    ram_cell[    5187] = 32'h8e61b7f2;
    ram_cell[    5188] = 32'h81c284e6;
    ram_cell[    5189] = 32'hde8b9c69;
    ram_cell[    5190] = 32'h06ef1701;
    ram_cell[    5191] = 32'hb07b4461;
    ram_cell[    5192] = 32'hff15aebc;
    ram_cell[    5193] = 32'h8c49aad3;
    ram_cell[    5194] = 32'h42598701;
    ram_cell[    5195] = 32'hb2504bb3;
    ram_cell[    5196] = 32'h7fcaca5e;
    ram_cell[    5197] = 32'h9296d98f;
    ram_cell[    5198] = 32'hcfed24a8;
    ram_cell[    5199] = 32'h7f49d978;
    ram_cell[    5200] = 32'hb1abbbcd;
    ram_cell[    5201] = 32'h264c6711;
    ram_cell[    5202] = 32'h5f243b9d;
    ram_cell[    5203] = 32'hde361137;
    ram_cell[    5204] = 32'hb84b7352;
    ram_cell[    5205] = 32'he933df5a;
    ram_cell[    5206] = 32'h4c693a16;
    ram_cell[    5207] = 32'h0d32d136;
    ram_cell[    5208] = 32'h5a5b81e2;
    ram_cell[    5209] = 32'h7b4629fa;
    ram_cell[    5210] = 32'h2951b649;
    ram_cell[    5211] = 32'h82772c1c;
    ram_cell[    5212] = 32'h888320d9;
    ram_cell[    5213] = 32'h2c6bf4aa;
    ram_cell[    5214] = 32'hfca232bf;
    ram_cell[    5215] = 32'h3f79772a;
    ram_cell[    5216] = 32'hadaad469;
    ram_cell[    5217] = 32'h627e6217;
    ram_cell[    5218] = 32'hbc6ab27e;
    ram_cell[    5219] = 32'hee989a80;
    ram_cell[    5220] = 32'h63293f0f;
    ram_cell[    5221] = 32'h70e050cd;
    ram_cell[    5222] = 32'h8052c1c7;
    ram_cell[    5223] = 32'hcfab1f75;
    ram_cell[    5224] = 32'h799fba50;
    ram_cell[    5225] = 32'h3336ba09;
    ram_cell[    5226] = 32'h2edde029;
    ram_cell[    5227] = 32'h10b494ec;
    ram_cell[    5228] = 32'h0328afa4;
    ram_cell[    5229] = 32'ha0cb745e;
    ram_cell[    5230] = 32'hde233a33;
    ram_cell[    5231] = 32'hb826c513;
    ram_cell[    5232] = 32'h6d8fd54b;
    ram_cell[    5233] = 32'hfaf2aefc;
    ram_cell[    5234] = 32'hd56b7d56;
    ram_cell[    5235] = 32'h9b514cf3;
    ram_cell[    5236] = 32'h39a3e1d2;
    ram_cell[    5237] = 32'ha5bbc8f0;
    ram_cell[    5238] = 32'h1e5e3efd;
    ram_cell[    5239] = 32'hba294e24;
    ram_cell[    5240] = 32'hc047e188;
    ram_cell[    5241] = 32'h0eebc478;
    ram_cell[    5242] = 32'h4a33eb90;
    ram_cell[    5243] = 32'h85d66047;
    ram_cell[    5244] = 32'h59ea8145;
    ram_cell[    5245] = 32'h93aa1d95;
    ram_cell[    5246] = 32'hd7f6d5cb;
    ram_cell[    5247] = 32'haaa54305;
    ram_cell[    5248] = 32'h5d4a0df5;
    ram_cell[    5249] = 32'hadcb07af;
    ram_cell[    5250] = 32'h6c475460;
    ram_cell[    5251] = 32'h3aeb22d4;
    ram_cell[    5252] = 32'h4261c55f;
    ram_cell[    5253] = 32'h3561e455;
    ram_cell[    5254] = 32'hc4351d5a;
    ram_cell[    5255] = 32'h91ae2cd2;
    ram_cell[    5256] = 32'he93d9ddf;
    ram_cell[    5257] = 32'h10b213c7;
    ram_cell[    5258] = 32'h7efbf685;
    ram_cell[    5259] = 32'hd4714eca;
    ram_cell[    5260] = 32'hd67964bd;
    ram_cell[    5261] = 32'hf73f358b;
    ram_cell[    5262] = 32'h3c3ecce9;
    ram_cell[    5263] = 32'h26538d49;
    ram_cell[    5264] = 32'h846146a5;
    ram_cell[    5265] = 32'h3e430459;
    ram_cell[    5266] = 32'h58bf6ecd;
    ram_cell[    5267] = 32'h90e62e99;
    ram_cell[    5268] = 32'h7fa6c8d8;
    ram_cell[    5269] = 32'hb5a6f963;
    ram_cell[    5270] = 32'hfbf3ef86;
    ram_cell[    5271] = 32'he137fb11;
    ram_cell[    5272] = 32'h7fb92061;
    ram_cell[    5273] = 32'h8d8de22d;
    ram_cell[    5274] = 32'hd41e4366;
    ram_cell[    5275] = 32'h661ffb38;
    ram_cell[    5276] = 32'hb9170fb4;
    ram_cell[    5277] = 32'h22972d1b;
    ram_cell[    5278] = 32'h4fcf4180;
    ram_cell[    5279] = 32'hcc4e7799;
    ram_cell[    5280] = 32'ha44a14e1;
    ram_cell[    5281] = 32'h6e83056a;
    ram_cell[    5282] = 32'hd0e7b6ba;
    ram_cell[    5283] = 32'h40fbb236;
    ram_cell[    5284] = 32'hbe935b3f;
    ram_cell[    5285] = 32'hdaaaca7a;
    ram_cell[    5286] = 32'hf8c8d1b4;
    ram_cell[    5287] = 32'h805a1202;
    ram_cell[    5288] = 32'hd8f51e6f;
    ram_cell[    5289] = 32'h38f23270;
    ram_cell[    5290] = 32'h5d4ca1c5;
    ram_cell[    5291] = 32'hd4ff9511;
    ram_cell[    5292] = 32'h202d9b7c;
    ram_cell[    5293] = 32'hc76e223b;
    ram_cell[    5294] = 32'hbf727ebf;
    ram_cell[    5295] = 32'h5db1ad7f;
    ram_cell[    5296] = 32'h0080f4f6;
    ram_cell[    5297] = 32'hf1fb4da0;
    ram_cell[    5298] = 32'h111e8642;
    ram_cell[    5299] = 32'hce6921c0;
    ram_cell[    5300] = 32'h5dabef37;
    ram_cell[    5301] = 32'hd06fdfff;
    ram_cell[    5302] = 32'h2ccc3d3a;
    ram_cell[    5303] = 32'h464fa95c;
    ram_cell[    5304] = 32'h1b9c8233;
    ram_cell[    5305] = 32'hbfb64e49;
    ram_cell[    5306] = 32'hc87c5577;
    ram_cell[    5307] = 32'h87e0f3ef;
    ram_cell[    5308] = 32'h8ab5866d;
    ram_cell[    5309] = 32'h1904a00d;
    ram_cell[    5310] = 32'hf6bd3201;
    ram_cell[    5311] = 32'hdc0c490c;
    ram_cell[    5312] = 32'h6925ea85;
    ram_cell[    5313] = 32'h0e4f36d9;
    ram_cell[    5314] = 32'hd89d3bbf;
    ram_cell[    5315] = 32'h5eab83ee;
    ram_cell[    5316] = 32'h7ee3cf92;
    ram_cell[    5317] = 32'h303b9654;
    ram_cell[    5318] = 32'h233bdec0;
    ram_cell[    5319] = 32'h90ee2da1;
    ram_cell[    5320] = 32'h2175ac5b;
    ram_cell[    5321] = 32'ha3def8cf;
    ram_cell[    5322] = 32'hff43fa9c;
    ram_cell[    5323] = 32'hce4ee6f1;
    ram_cell[    5324] = 32'h52353e07;
    ram_cell[    5325] = 32'hc0e966aa;
    ram_cell[    5326] = 32'hcf9c1036;
    ram_cell[    5327] = 32'h783568cc;
    ram_cell[    5328] = 32'ha8eccde0;
    ram_cell[    5329] = 32'h05b1ac04;
    ram_cell[    5330] = 32'h166e7f26;
    ram_cell[    5331] = 32'he72ca566;
    ram_cell[    5332] = 32'h00d32bbe;
    ram_cell[    5333] = 32'h0fea59d6;
    ram_cell[    5334] = 32'h256236d4;
    ram_cell[    5335] = 32'h308e423e;
    ram_cell[    5336] = 32'h1f1bf804;
    ram_cell[    5337] = 32'h74bf3989;
    ram_cell[    5338] = 32'he6e3181b;
    ram_cell[    5339] = 32'h1bc32a5a;
    ram_cell[    5340] = 32'h31bc0910;
    ram_cell[    5341] = 32'h8df2455f;
    ram_cell[    5342] = 32'he0b2ae45;
    ram_cell[    5343] = 32'hf19dd6ec;
    ram_cell[    5344] = 32'h410469a4;
    ram_cell[    5345] = 32'hec6b78f2;
    ram_cell[    5346] = 32'hcf023713;
    ram_cell[    5347] = 32'hfc03f871;
    ram_cell[    5348] = 32'h71b2735d;
    ram_cell[    5349] = 32'hb624aa29;
    ram_cell[    5350] = 32'h8e9b1fc0;
    ram_cell[    5351] = 32'ha1ee5606;
    ram_cell[    5352] = 32'h45ce31aa;
    ram_cell[    5353] = 32'h0fa4a6df;
    ram_cell[    5354] = 32'ha821023e;
    ram_cell[    5355] = 32'h488e96de;
    ram_cell[    5356] = 32'h57d02dc3;
    ram_cell[    5357] = 32'h0ea007d7;
    ram_cell[    5358] = 32'hc0341474;
    ram_cell[    5359] = 32'h4acf6a27;
    ram_cell[    5360] = 32'h5e8f6afd;
    ram_cell[    5361] = 32'h07965276;
    ram_cell[    5362] = 32'hc7a75aa7;
    ram_cell[    5363] = 32'heb7d7bae;
    ram_cell[    5364] = 32'h8401588c;
    ram_cell[    5365] = 32'h12ad6c72;
    ram_cell[    5366] = 32'hc53e55bf;
    ram_cell[    5367] = 32'h4a6889d7;
    ram_cell[    5368] = 32'h17eeb81d;
    ram_cell[    5369] = 32'hd1294e60;
    ram_cell[    5370] = 32'hf7e476ea;
    ram_cell[    5371] = 32'h1c2c16c2;
    ram_cell[    5372] = 32'hb2459535;
    ram_cell[    5373] = 32'hc8c4b1b9;
    ram_cell[    5374] = 32'h443b717f;
    ram_cell[    5375] = 32'hae88eeac;
    ram_cell[    5376] = 32'hd367a94b;
    ram_cell[    5377] = 32'h128ab1bb;
    ram_cell[    5378] = 32'hd7174fbf;
    ram_cell[    5379] = 32'hd3baa489;
    ram_cell[    5380] = 32'h74aa768b;
    ram_cell[    5381] = 32'h2c672716;
    ram_cell[    5382] = 32'hd4004466;
    ram_cell[    5383] = 32'ha645142c;
    ram_cell[    5384] = 32'h251325d9;
    ram_cell[    5385] = 32'h9b03b37a;
    ram_cell[    5386] = 32'hbf83c5b0;
    ram_cell[    5387] = 32'h8505eec3;
    ram_cell[    5388] = 32'h62986752;
    ram_cell[    5389] = 32'h33711332;
    ram_cell[    5390] = 32'hf19ed2d5;
    ram_cell[    5391] = 32'hf9c2c537;
    ram_cell[    5392] = 32'h71fe0337;
    ram_cell[    5393] = 32'h955b2178;
    ram_cell[    5394] = 32'hb4daabd6;
    ram_cell[    5395] = 32'hd3799a5f;
    ram_cell[    5396] = 32'h50ec6116;
    ram_cell[    5397] = 32'hc8cbd5ed;
    ram_cell[    5398] = 32'h8863679a;
    ram_cell[    5399] = 32'h951a72f6;
    ram_cell[    5400] = 32'h8b20a0b1;
    ram_cell[    5401] = 32'h46b4a7d0;
    ram_cell[    5402] = 32'h112e04cc;
    ram_cell[    5403] = 32'h8ea661ed;
    ram_cell[    5404] = 32'h171f983d;
    ram_cell[    5405] = 32'h8e6bf2d5;
    ram_cell[    5406] = 32'h0ed4a55b;
    ram_cell[    5407] = 32'h9795005d;
    ram_cell[    5408] = 32'h8bf1a8c2;
    ram_cell[    5409] = 32'h172407b8;
    ram_cell[    5410] = 32'hf5f1394b;
    ram_cell[    5411] = 32'hc1540901;
    ram_cell[    5412] = 32'h704570f3;
    ram_cell[    5413] = 32'hbc0b81db;
    ram_cell[    5414] = 32'h2ca75564;
    ram_cell[    5415] = 32'h303418e9;
    ram_cell[    5416] = 32'hbf3abd74;
    ram_cell[    5417] = 32'h22f57f4e;
    ram_cell[    5418] = 32'hc67605db;
    ram_cell[    5419] = 32'hbcd0fb71;
    ram_cell[    5420] = 32'hd2b3a397;
    ram_cell[    5421] = 32'he20cdcab;
    ram_cell[    5422] = 32'hd76090cd;
    ram_cell[    5423] = 32'h41626eb4;
    ram_cell[    5424] = 32'h14f3db68;
    ram_cell[    5425] = 32'he6257b18;
    ram_cell[    5426] = 32'h6f69a208;
    ram_cell[    5427] = 32'he2e1e6d1;
    ram_cell[    5428] = 32'h44c38acf;
    ram_cell[    5429] = 32'h3814a59b;
    ram_cell[    5430] = 32'h017b83f0;
    ram_cell[    5431] = 32'h14173207;
    ram_cell[    5432] = 32'h6debaa2c;
    ram_cell[    5433] = 32'h77a01440;
    ram_cell[    5434] = 32'ha2012252;
    ram_cell[    5435] = 32'h9ca7e5fb;
    ram_cell[    5436] = 32'hba977cac;
    ram_cell[    5437] = 32'h11c343d5;
    ram_cell[    5438] = 32'hefe634f7;
    ram_cell[    5439] = 32'h4b03d431;
    ram_cell[    5440] = 32'h1a454d01;
    ram_cell[    5441] = 32'h712544a0;
    ram_cell[    5442] = 32'h7a0781fd;
    ram_cell[    5443] = 32'hc2709c1f;
    ram_cell[    5444] = 32'h04f10dbe;
    ram_cell[    5445] = 32'h3f26f375;
    ram_cell[    5446] = 32'hbaef6a38;
    ram_cell[    5447] = 32'he99a2e6f;
    ram_cell[    5448] = 32'h209bd877;
    ram_cell[    5449] = 32'h5627a62b;
    ram_cell[    5450] = 32'ha522f684;
    ram_cell[    5451] = 32'hc3b81d71;
    ram_cell[    5452] = 32'h8c0fd6e8;
    ram_cell[    5453] = 32'h61d1eb1c;
    ram_cell[    5454] = 32'h18efa72b;
    ram_cell[    5455] = 32'h30a99cd2;
    ram_cell[    5456] = 32'h6697e113;
    ram_cell[    5457] = 32'hf1d3192c;
    ram_cell[    5458] = 32'h555a5971;
    ram_cell[    5459] = 32'h9b1c6e49;
    ram_cell[    5460] = 32'h6e96af83;
    ram_cell[    5461] = 32'h35f7da08;
    ram_cell[    5462] = 32'h042d6f57;
    ram_cell[    5463] = 32'h21363fa9;
    ram_cell[    5464] = 32'h2928ab63;
    ram_cell[    5465] = 32'h44d7c251;
    ram_cell[    5466] = 32'h22c2516c;
    ram_cell[    5467] = 32'hff67b5c6;
    ram_cell[    5468] = 32'h37d67f23;
    ram_cell[    5469] = 32'hdc6f8276;
    ram_cell[    5470] = 32'h71b17932;
    ram_cell[    5471] = 32'h7c758ef7;
    ram_cell[    5472] = 32'h3713ab70;
    ram_cell[    5473] = 32'h667062b6;
    ram_cell[    5474] = 32'h2329c3ca;
    ram_cell[    5475] = 32'h7bed0dc8;
    ram_cell[    5476] = 32'h744a8be7;
    ram_cell[    5477] = 32'h7228ef34;
    ram_cell[    5478] = 32'hbb298765;
    ram_cell[    5479] = 32'h94c88448;
    ram_cell[    5480] = 32'h07800450;
    ram_cell[    5481] = 32'h2c2d279b;
    ram_cell[    5482] = 32'he15c62db;
    ram_cell[    5483] = 32'h838f2b75;
    ram_cell[    5484] = 32'h5f9601dc;
    ram_cell[    5485] = 32'h8442672e;
    ram_cell[    5486] = 32'h1cdae395;
    ram_cell[    5487] = 32'h64dcfd65;
    ram_cell[    5488] = 32'h162a8a12;
    ram_cell[    5489] = 32'hc4460534;
    ram_cell[    5490] = 32'h2ba27d8e;
    ram_cell[    5491] = 32'h75fb70bc;
    ram_cell[    5492] = 32'h767fa1dc;
    ram_cell[    5493] = 32'h091e9e1f;
    ram_cell[    5494] = 32'h5f9023c4;
    ram_cell[    5495] = 32'h1c5b0703;
    ram_cell[    5496] = 32'h4ae04844;
    ram_cell[    5497] = 32'ha92b82dd;
    ram_cell[    5498] = 32'h46174985;
    ram_cell[    5499] = 32'hf9c807e4;
    ram_cell[    5500] = 32'hfb5a479a;
    ram_cell[    5501] = 32'h7996e9fb;
    ram_cell[    5502] = 32'ha66d9c90;
    ram_cell[    5503] = 32'hc72818ec;
    ram_cell[    5504] = 32'h0bf2aeef;
    ram_cell[    5505] = 32'h7bf4e9e2;
    ram_cell[    5506] = 32'ha00b778f;
    ram_cell[    5507] = 32'h74779433;
    ram_cell[    5508] = 32'h379e50d1;
    ram_cell[    5509] = 32'h9c705af3;
    ram_cell[    5510] = 32'h5b63a68d;
    ram_cell[    5511] = 32'h2032ba85;
    ram_cell[    5512] = 32'h9da89788;
    ram_cell[    5513] = 32'h67e61e5f;
    ram_cell[    5514] = 32'h5bdbde6e;
    ram_cell[    5515] = 32'h3d59c657;
    ram_cell[    5516] = 32'hdda545be;
    ram_cell[    5517] = 32'ha2cb47b0;
    ram_cell[    5518] = 32'hb6a974c3;
    ram_cell[    5519] = 32'h63150cfb;
    ram_cell[    5520] = 32'h5f35eb66;
    ram_cell[    5521] = 32'hc5d3231d;
    ram_cell[    5522] = 32'hfac561a7;
    ram_cell[    5523] = 32'h3635e52d;
    ram_cell[    5524] = 32'h2db66d9a;
    ram_cell[    5525] = 32'h9cb5bf05;
    ram_cell[    5526] = 32'hc063a70c;
    ram_cell[    5527] = 32'h3a0562ba;
    ram_cell[    5528] = 32'ha021b018;
    ram_cell[    5529] = 32'h9cf3accb;
    ram_cell[    5530] = 32'hd9a9efb3;
    ram_cell[    5531] = 32'h517c9bd0;
    ram_cell[    5532] = 32'hf9f92204;
    ram_cell[    5533] = 32'heb0a674c;
    ram_cell[    5534] = 32'hd3222a90;
    ram_cell[    5535] = 32'h829a4a85;
    ram_cell[    5536] = 32'h6e28e8cb;
    ram_cell[    5537] = 32'h6e2763fe;
    ram_cell[    5538] = 32'h0a3073ce;
    ram_cell[    5539] = 32'hf016a8d5;
    ram_cell[    5540] = 32'ha729c0f9;
    ram_cell[    5541] = 32'hee67e0af;
    ram_cell[    5542] = 32'ha31c5fb4;
    ram_cell[    5543] = 32'ha4ee17b4;
    ram_cell[    5544] = 32'h9b250a83;
    ram_cell[    5545] = 32'hda971e21;
    ram_cell[    5546] = 32'h02a1b8b1;
    ram_cell[    5547] = 32'hb8a9eed5;
    ram_cell[    5548] = 32'h16a7b480;
    ram_cell[    5549] = 32'ha70960ea;
    ram_cell[    5550] = 32'h3066eefc;
    ram_cell[    5551] = 32'hebbd6ba9;
    ram_cell[    5552] = 32'h8953371c;
    ram_cell[    5553] = 32'hecf5cebd;
    ram_cell[    5554] = 32'h3e2da554;
    ram_cell[    5555] = 32'h315a628e;
    ram_cell[    5556] = 32'h51b285b2;
    ram_cell[    5557] = 32'h64111835;
    ram_cell[    5558] = 32'hb4a93057;
    ram_cell[    5559] = 32'hce3934f5;
    ram_cell[    5560] = 32'ha93c4818;
    ram_cell[    5561] = 32'h22a29816;
    ram_cell[    5562] = 32'hf0fa9e5a;
    ram_cell[    5563] = 32'hf4376448;
    ram_cell[    5564] = 32'he61e49c6;
    ram_cell[    5565] = 32'h5753ffb7;
    ram_cell[    5566] = 32'hd7004f19;
    ram_cell[    5567] = 32'h412bf6cc;
    ram_cell[    5568] = 32'h28d6c1c6;
    ram_cell[    5569] = 32'hc25c9d98;
    ram_cell[    5570] = 32'h16b8a8b1;
    ram_cell[    5571] = 32'h6a75345b;
    ram_cell[    5572] = 32'hc95dac48;
    ram_cell[    5573] = 32'h49d76334;
    ram_cell[    5574] = 32'h26f6d7f8;
    ram_cell[    5575] = 32'hf71a0fdb;
    ram_cell[    5576] = 32'h78adfd1f;
    ram_cell[    5577] = 32'hab102346;
    ram_cell[    5578] = 32'hbb93bb1b;
    ram_cell[    5579] = 32'h4b9110fe;
    ram_cell[    5580] = 32'hb03bd55d;
    ram_cell[    5581] = 32'hc6657680;
    ram_cell[    5582] = 32'ha3ce742c;
    ram_cell[    5583] = 32'h6321c7d6;
    ram_cell[    5584] = 32'h7a81d24a;
    ram_cell[    5585] = 32'h0c935f1c;
    ram_cell[    5586] = 32'he1e576c9;
    ram_cell[    5587] = 32'haa9131d0;
    ram_cell[    5588] = 32'h8978bb41;
    ram_cell[    5589] = 32'hdfa32325;
    ram_cell[    5590] = 32'hff7ee1ac;
    ram_cell[    5591] = 32'h70a72254;
    ram_cell[    5592] = 32'h3797d484;
    ram_cell[    5593] = 32'h9cbca863;
    ram_cell[    5594] = 32'h0c6a1670;
    ram_cell[    5595] = 32'h7c55e457;
    ram_cell[    5596] = 32'hef8ac073;
    ram_cell[    5597] = 32'hc87933e5;
    ram_cell[    5598] = 32'he8be18fe;
    ram_cell[    5599] = 32'hf6cf8d84;
    ram_cell[    5600] = 32'hf4336b1a;
    ram_cell[    5601] = 32'hfb62b2d7;
    ram_cell[    5602] = 32'h08c18b21;
    ram_cell[    5603] = 32'h89cb6cd8;
    ram_cell[    5604] = 32'hf7e869ee;
    ram_cell[    5605] = 32'h6526738f;
    ram_cell[    5606] = 32'h18160afa;
    ram_cell[    5607] = 32'hfb9ba194;
    ram_cell[    5608] = 32'hf856d4af;
    ram_cell[    5609] = 32'hf4e36bda;
    ram_cell[    5610] = 32'he3d98588;
    ram_cell[    5611] = 32'h3d306acb;
    ram_cell[    5612] = 32'haed250ca;
    ram_cell[    5613] = 32'h5b42d3fe;
    ram_cell[    5614] = 32'h949d2984;
    ram_cell[    5615] = 32'ha187b43c;
    ram_cell[    5616] = 32'h99a31e61;
    ram_cell[    5617] = 32'hecd313b4;
    ram_cell[    5618] = 32'h97904f96;
    ram_cell[    5619] = 32'h847c4702;
    ram_cell[    5620] = 32'h601ab413;
    ram_cell[    5621] = 32'hdc393965;
    ram_cell[    5622] = 32'heb7b5195;
    ram_cell[    5623] = 32'ha40715de;
    ram_cell[    5624] = 32'h90dced56;
    ram_cell[    5625] = 32'ha1c0f3bd;
    ram_cell[    5626] = 32'h45075c67;
    ram_cell[    5627] = 32'h8a71c401;
    ram_cell[    5628] = 32'h35285b16;
    ram_cell[    5629] = 32'hbb65dbbe;
    ram_cell[    5630] = 32'h002d5c1f;
    ram_cell[    5631] = 32'hbf834ae0;
    ram_cell[    5632] = 32'hca19f053;
    ram_cell[    5633] = 32'hd33560bf;
    ram_cell[    5634] = 32'hfbbe7873;
    ram_cell[    5635] = 32'h96d77530;
    ram_cell[    5636] = 32'h04d0d111;
    ram_cell[    5637] = 32'h77f99657;
    ram_cell[    5638] = 32'hf7c8f50e;
    ram_cell[    5639] = 32'h8decf076;
    ram_cell[    5640] = 32'h1641f2fc;
    ram_cell[    5641] = 32'h974e168a;
    ram_cell[    5642] = 32'h106d10e1;
    ram_cell[    5643] = 32'h3d9a193f;
    ram_cell[    5644] = 32'h8ae97e88;
    ram_cell[    5645] = 32'h409edfda;
    ram_cell[    5646] = 32'h2d9522f7;
    ram_cell[    5647] = 32'h3d650e9d;
    ram_cell[    5648] = 32'hd434368e;
    ram_cell[    5649] = 32'hea21643d;
    ram_cell[    5650] = 32'h7b6511da;
    ram_cell[    5651] = 32'h4f5b4303;
    ram_cell[    5652] = 32'hc3d12007;
    ram_cell[    5653] = 32'h4cab43a0;
    ram_cell[    5654] = 32'h24118542;
    ram_cell[    5655] = 32'h8fa9a047;
    ram_cell[    5656] = 32'h4b016149;
    ram_cell[    5657] = 32'habf07d94;
    ram_cell[    5658] = 32'h86ffc262;
    ram_cell[    5659] = 32'h27aaf7db;
    ram_cell[    5660] = 32'he12b8ad7;
    ram_cell[    5661] = 32'h5bad3dc6;
    ram_cell[    5662] = 32'h1508b2af;
    ram_cell[    5663] = 32'h08cd8aff;
    ram_cell[    5664] = 32'h02b9edf4;
    ram_cell[    5665] = 32'h7caf7102;
    ram_cell[    5666] = 32'hb4249c08;
    ram_cell[    5667] = 32'h555d156f;
    ram_cell[    5668] = 32'hd047d4ee;
    ram_cell[    5669] = 32'h191be1cc;
    ram_cell[    5670] = 32'hc09371a3;
    ram_cell[    5671] = 32'hbdd6109e;
    ram_cell[    5672] = 32'h11285baf;
    ram_cell[    5673] = 32'h282410cc;
    ram_cell[    5674] = 32'h204532aa;
    ram_cell[    5675] = 32'hcf0ea412;
    ram_cell[    5676] = 32'h9de7b495;
    ram_cell[    5677] = 32'h13fb2684;
    ram_cell[    5678] = 32'hf62f1a1b;
    ram_cell[    5679] = 32'hf958f0c7;
    ram_cell[    5680] = 32'h480206fc;
    ram_cell[    5681] = 32'he1ece3aa;
    ram_cell[    5682] = 32'h73d43824;
    ram_cell[    5683] = 32'h0dc7beb8;
    ram_cell[    5684] = 32'hb53f6a3e;
    ram_cell[    5685] = 32'hd92ccddf;
    ram_cell[    5686] = 32'hd426cdd2;
    ram_cell[    5687] = 32'h953ec5fd;
    ram_cell[    5688] = 32'h5f4b2c49;
    ram_cell[    5689] = 32'hbf96dd64;
    ram_cell[    5690] = 32'hada4e62d;
    ram_cell[    5691] = 32'hef6886d0;
    ram_cell[    5692] = 32'h0ba71e24;
    ram_cell[    5693] = 32'h89c08f82;
    ram_cell[    5694] = 32'hc69cfca1;
    ram_cell[    5695] = 32'h979da5c3;
    ram_cell[    5696] = 32'h3b1e5ba1;
    ram_cell[    5697] = 32'h80e53968;
    ram_cell[    5698] = 32'h8dfcf698;
    ram_cell[    5699] = 32'h02c59efd;
    ram_cell[    5700] = 32'h0b4cc735;
    ram_cell[    5701] = 32'hf4355bdc;
    ram_cell[    5702] = 32'h1d5df8d8;
    ram_cell[    5703] = 32'hb0f42562;
    ram_cell[    5704] = 32'h721dfeca;
    ram_cell[    5705] = 32'h87f51816;
    ram_cell[    5706] = 32'hca15b809;
    ram_cell[    5707] = 32'h9281968b;
    ram_cell[    5708] = 32'hc52019c4;
    ram_cell[    5709] = 32'hb7260e62;
    ram_cell[    5710] = 32'h4e282bb2;
    ram_cell[    5711] = 32'h74c0e7f9;
    ram_cell[    5712] = 32'hef2d0858;
    ram_cell[    5713] = 32'hcfbb815a;
    ram_cell[    5714] = 32'h66849155;
    ram_cell[    5715] = 32'h0dbe65f4;
    ram_cell[    5716] = 32'h85bbb7ac;
    ram_cell[    5717] = 32'h59d94133;
    ram_cell[    5718] = 32'hc15cd203;
    ram_cell[    5719] = 32'h13a00259;
    ram_cell[    5720] = 32'h1cfcc6b9;
    ram_cell[    5721] = 32'h4a3a303d;
    ram_cell[    5722] = 32'h00b612d8;
    ram_cell[    5723] = 32'h5e9c8698;
    ram_cell[    5724] = 32'h3a40ac89;
    ram_cell[    5725] = 32'hfa331a28;
    ram_cell[    5726] = 32'h0291584e;
    ram_cell[    5727] = 32'he1476b38;
    ram_cell[    5728] = 32'h8bf56202;
    ram_cell[    5729] = 32'h89b30893;
    ram_cell[    5730] = 32'h0dfcc4a3;
    ram_cell[    5731] = 32'h07bc7883;
    ram_cell[    5732] = 32'h83a7cdbf;
    ram_cell[    5733] = 32'h03b94976;
    ram_cell[    5734] = 32'h8cd95cd1;
    ram_cell[    5735] = 32'ha45250a9;
    ram_cell[    5736] = 32'hb6e591ac;
    ram_cell[    5737] = 32'h695a79e4;
    ram_cell[    5738] = 32'hce610359;
    ram_cell[    5739] = 32'h7e246cdb;
    ram_cell[    5740] = 32'hdfc8f99c;
    ram_cell[    5741] = 32'he93f5c07;
    ram_cell[    5742] = 32'h9e5e5694;
    ram_cell[    5743] = 32'h4e1686ef;
    ram_cell[    5744] = 32'h8de19dee;
    ram_cell[    5745] = 32'h6454f40a;
    ram_cell[    5746] = 32'h73dd8285;
    ram_cell[    5747] = 32'h6ad46920;
    ram_cell[    5748] = 32'h6ed44d76;
    ram_cell[    5749] = 32'h38c2c9ce;
    ram_cell[    5750] = 32'h7126f0e9;
    ram_cell[    5751] = 32'hff84d5e5;
    ram_cell[    5752] = 32'hdf8c8c10;
    ram_cell[    5753] = 32'h3b8ededf;
    ram_cell[    5754] = 32'hdfb38c44;
    ram_cell[    5755] = 32'h9fa7e398;
    ram_cell[    5756] = 32'hd503aebd;
    ram_cell[    5757] = 32'h2bd773f9;
    ram_cell[    5758] = 32'h0520804c;
    ram_cell[    5759] = 32'he05698d3;
    ram_cell[    5760] = 32'h8c77723b;
    ram_cell[    5761] = 32'he509290c;
    ram_cell[    5762] = 32'h91c98193;
    ram_cell[    5763] = 32'h83a6d53f;
    ram_cell[    5764] = 32'h918829d9;
    ram_cell[    5765] = 32'h75fc4023;
    ram_cell[    5766] = 32'hab503b92;
    ram_cell[    5767] = 32'h39988bf6;
    ram_cell[    5768] = 32'h0a9c9e2c;
    ram_cell[    5769] = 32'h05b746a7;
    ram_cell[    5770] = 32'h17b4e4a1;
    ram_cell[    5771] = 32'hf3611f91;
    ram_cell[    5772] = 32'h5805c0ec;
    ram_cell[    5773] = 32'h2096d514;
    ram_cell[    5774] = 32'hf377ce0e;
    ram_cell[    5775] = 32'hdfd1855e;
    ram_cell[    5776] = 32'hf9307cbc;
    ram_cell[    5777] = 32'h909c28cd;
    ram_cell[    5778] = 32'hd3c5dc0e;
    ram_cell[    5779] = 32'h5e793a24;
    ram_cell[    5780] = 32'hbacf67b3;
    ram_cell[    5781] = 32'h3a2492cd;
    ram_cell[    5782] = 32'hef00a038;
    ram_cell[    5783] = 32'he551148c;
    ram_cell[    5784] = 32'hf44119b9;
    ram_cell[    5785] = 32'h6b359217;
    ram_cell[    5786] = 32'hd7e6e588;
    ram_cell[    5787] = 32'h05743422;
    ram_cell[    5788] = 32'h09f201ab;
    ram_cell[    5789] = 32'hc1341de0;
    ram_cell[    5790] = 32'h7f155145;
    ram_cell[    5791] = 32'h6d53b34e;
    ram_cell[    5792] = 32'h10a1bd28;
    ram_cell[    5793] = 32'hf9e2cc52;
    ram_cell[    5794] = 32'h4c098b20;
    ram_cell[    5795] = 32'he78839a2;
    ram_cell[    5796] = 32'h65a2d0fb;
    ram_cell[    5797] = 32'h25850916;
    ram_cell[    5798] = 32'h78a4e961;
    ram_cell[    5799] = 32'h3bc817ca;
    ram_cell[    5800] = 32'hf1541da0;
    ram_cell[    5801] = 32'h32154208;
    ram_cell[    5802] = 32'hb97b2b42;
    ram_cell[    5803] = 32'h37ca84d3;
    ram_cell[    5804] = 32'h98f8bdfa;
    ram_cell[    5805] = 32'hd1e3a80f;
    ram_cell[    5806] = 32'ha667a3fb;
    ram_cell[    5807] = 32'h89cdda55;
    ram_cell[    5808] = 32'h94bddf14;
    ram_cell[    5809] = 32'h54df9234;
    ram_cell[    5810] = 32'hb2fe226f;
    ram_cell[    5811] = 32'h77f509b7;
    ram_cell[    5812] = 32'h541217bb;
    ram_cell[    5813] = 32'hfd4d5be9;
    ram_cell[    5814] = 32'he8a46b0d;
    ram_cell[    5815] = 32'hfc30f952;
    ram_cell[    5816] = 32'hd9074bbb;
    ram_cell[    5817] = 32'he429cff1;
    ram_cell[    5818] = 32'hb5d2aeee;
    ram_cell[    5819] = 32'h938cfb3c;
    ram_cell[    5820] = 32'h6e647380;
    ram_cell[    5821] = 32'hb6f38891;
    ram_cell[    5822] = 32'hfe02edc4;
    ram_cell[    5823] = 32'h69554900;
    ram_cell[    5824] = 32'h5558ed44;
    ram_cell[    5825] = 32'hadfadad3;
    ram_cell[    5826] = 32'h21d25d22;
    ram_cell[    5827] = 32'h5de447d0;
    ram_cell[    5828] = 32'h1b313370;
    ram_cell[    5829] = 32'h8931d5bf;
    ram_cell[    5830] = 32'h1310b40f;
    ram_cell[    5831] = 32'hce73e67a;
    ram_cell[    5832] = 32'h9f136bd1;
    ram_cell[    5833] = 32'hadde9a27;
    ram_cell[    5834] = 32'h285c6b2b;
    ram_cell[    5835] = 32'h33211c57;
    ram_cell[    5836] = 32'h47b57815;
    ram_cell[    5837] = 32'h1f7deb57;
    ram_cell[    5838] = 32'h3708c60e;
    ram_cell[    5839] = 32'h81958425;
    ram_cell[    5840] = 32'h038efee4;
    ram_cell[    5841] = 32'hf1b916bb;
    ram_cell[    5842] = 32'hcb66b048;
    ram_cell[    5843] = 32'ha2f41d5f;
    ram_cell[    5844] = 32'h392eef47;
    ram_cell[    5845] = 32'hcfdf94e6;
    ram_cell[    5846] = 32'hc01fed6e;
    ram_cell[    5847] = 32'h7848b2eb;
    ram_cell[    5848] = 32'h5d4ba1b9;
    ram_cell[    5849] = 32'ha4bc7a3e;
    ram_cell[    5850] = 32'he3f80d7e;
    ram_cell[    5851] = 32'h1564d0d9;
    ram_cell[    5852] = 32'hfa6b6cb9;
    ram_cell[    5853] = 32'h0c0f2d66;
    ram_cell[    5854] = 32'h74a626e8;
    ram_cell[    5855] = 32'hd4e4bb8b;
    ram_cell[    5856] = 32'h94da14ca;
    ram_cell[    5857] = 32'hd7e39dc2;
    ram_cell[    5858] = 32'h999ca078;
    ram_cell[    5859] = 32'h01a3a84f;
    ram_cell[    5860] = 32'h905bca87;
    ram_cell[    5861] = 32'h834c9f7d;
    ram_cell[    5862] = 32'h358a9e41;
    ram_cell[    5863] = 32'h290f1c65;
    ram_cell[    5864] = 32'h51321f6d;
    ram_cell[    5865] = 32'hef24b5e1;
    ram_cell[    5866] = 32'h98135dd0;
    ram_cell[    5867] = 32'he4ea421a;
    ram_cell[    5868] = 32'h585d6d6b;
    ram_cell[    5869] = 32'haad20ea0;
    ram_cell[    5870] = 32'h6939979b;
    ram_cell[    5871] = 32'he5bd6987;
    ram_cell[    5872] = 32'h1163b028;
    ram_cell[    5873] = 32'h52b8a7f0;
    ram_cell[    5874] = 32'h9e1e1ad9;
    ram_cell[    5875] = 32'hc0d9308f;
    ram_cell[    5876] = 32'hee0467d9;
    ram_cell[    5877] = 32'h30085e34;
    ram_cell[    5878] = 32'hd601c151;
    ram_cell[    5879] = 32'h9e22a156;
    ram_cell[    5880] = 32'h0c0af64a;
    ram_cell[    5881] = 32'h3808ce9a;
    ram_cell[    5882] = 32'h88e6fc9a;
    ram_cell[    5883] = 32'h738d2edc;
    ram_cell[    5884] = 32'hdf81bdb6;
    ram_cell[    5885] = 32'h4b1133ee;
    ram_cell[    5886] = 32'h62bd2227;
    ram_cell[    5887] = 32'h7e4eb9f4;
    ram_cell[    5888] = 32'hacc5cb20;
    ram_cell[    5889] = 32'h37c09d78;
    ram_cell[    5890] = 32'he86f8423;
    ram_cell[    5891] = 32'hf74c024e;
    ram_cell[    5892] = 32'h8da84c8c;
    ram_cell[    5893] = 32'hf7115bc6;
    ram_cell[    5894] = 32'h78f8c84b;
    ram_cell[    5895] = 32'h4e75a875;
    ram_cell[    5896] = 32'hbd668e38;
    ram_cell[    5897] = 32'h1fe6d572;
    ram_cell[    5898] = 32'h97ec0a20;
    ram_cell[    5899] = 32'h36e64fcf;
    ram_cell[    5900] = 32'h0c607f0f;
    ram_cell[    5901] = 32'h14a938c4;
    ram_cell[    5902] = 32'h58237e8e;
    ram_cell[    5903] = 32'h2e60ed11;
    ram_cell[    5904] = 32'hcf78c845;
    ram_cell[    5905] = 32'h8c18ad39;
    ram_cell[    5906] = 32'hf2443291;
    ram_cell[    5907] = 32'h8587f0aa;
    ram_cell[    5908] = 32'h543ad087;
    ram_cell[    5909] = 32'h08c46aae;
    ram_cell[    5910] = 32'hf9d01f2c;
    ram_cell[    5911] = 32'h7aa552e9;
    ram_cell[    5912] = 32'hd7aaf7e1;
    ram_cell[    5913] = 32'h90eaa714;
    ram_cell[    5914] = 32'h0c50e785;
    ram_cell[    5915] = 32'h752df733;
    ram_cell[    5916] = 32'hd57bed10;
    ram_cell[    5917] = 32'h01ba836e;
    ram_cell[    5918] = 32'h0ba22416;
    ram_cell[    5919] = 32'h2cdd22b4;
    ram_cell[    5920] = 32'hc9bc0f19;
    ram_cell[    5921] = 32'h594d896e;
    ram_cell[    5922] = 32'h33342aa9;
    ram_cell[    5923] = 32'h1f9e2596;
    ram_cell[    5924] = 32'h473bc2b2;
    ram_cell[    5925] = 32'h85216522;
    ram_cell[    5926] = 32'hf1ee7649;
    ram_cell[    5927] = 32'h5b6c5e67;
    ram_cell[    5928] = 32'h6e66c5ae;
    ram_cell[    5929] = 32'h52a1b75b;
    ram_cell[    5930] = 32'h3f122bdc;
    ram_cell[    5931] = 32'h2aa10236;
    ram_cell[    5932] = 32'h7d32ac5d;
    ram_cell[    5933] = 32'h957bb4fc;
    ram_cell[    5934] = 32'ha90f3aa2;
    ram_cell[    5935] = 32'h96b6c52e;
    ram_cell[    5936] = 32'h97ceb65b;
    ram_cell[    5937] = 32'h32e6c20d;
    ram_cell[    5938] = 32'hbc73c989;
    ram_cell[    5939] = 32'h300e20e8;
    ram_cell[    5940] = 32'h52177202;
    ram_cell[    5941] = 32'hff4d5d1c;
    ram_cell[    5942] = 32'h13ea563a;
    ram_cell[    5943] = 32'h4750295c;
    ram_cell[    5944] = 32'h1c5f17c6;
    ram_cell[    5945] = 32'h8f850060;
    ram_cell[    5946] = 32'h164287e7;
    ram_cell[    5947] = 32'hab6f0090;
    ram_cell[    5948] = 32'h0c6399df;
    ram_cell[    5949] = 32'hd52079a8;
    ram_cell[    5950] = 32'ha429daa3;
    ram_cell[    5951] = 32'hcd6bea39;
    ram_cell[    5952] = 32'h2c4beef6;
    ram_cell[    5953] = 32'haceee497;
    ram_cell[    5954] = 32'he8eec028;
    ram_cell[    5955] = 32'h49796ff4;
    ram_cell[    5956] = 32'he613bfab;
    ram_cell[    5957] = 32'haac03cf0;
    ram_cell[    5958] = 32'hce5f9938;
    ram_cell[    5959] = 32'h18c8b633;
    ram_cell[    5960] = 32'hc17953bd;
    ram_cell[    5961] = 32'hfcb92d65;
    ram_cell[    5962] = 32'h5c51525d;
    ram_cell[    5963] = 32'h7d6e7e44;
    ram_cell[    5964] = 32'h6a701a46;
    ram_cell[    5965] = 32'h55ceb170;
    ram_cell[    5966] = 32'h70931eb5;
    ram_cell[    5967] = 32'h92acd26f;
    ram_cell[    5968] = 32'h9cbbf8cf;
    ram_cell[    5969] = 32'hc3e95514;
    ram_cell[    5970] = 32'h55ee4265;
    ram_cell[    5971] = 32'h4b1c2e53;
    ram_cell[    5972] = 32'ha834d8ac;
    ram_cell[    5973] = 32'h34df54db;
    ram_cell[    5974] = 32'h59bab907;
    ram_cell[    5975] = 32'he1ba4766;
    ram_cell[    5976] = 32'hdd265dd0;
    ram_cell[    5977] = 32'h9f2975a3;
    ram_cell[    5978] = 32'hf7b8b9b8;
    ram_cell[    5979] = 32'hbbecc9e7;
    ram_cell[    5980] = 32'habc13f8c;
    ram_cell[    5981] = 32'h894bd2a5;
    ram_cell[    5982] = 32'hdbe46bf6;
    ram_cell[    5983] = 32'h63df98ce;
    ram_cell[    5984] = 32'h54d4ce17;
    ram_cell[    5985] = 32'h9eae4e99;
    ram_cell[    5986] = 32'hc353ce0b;
    ram_cell[    5987] = 32'hdb6a9d4b;
    ram_cell[    5988] = 32'h1d8ec52b;
    ram_cell[    5989] = 32'h6381c195;
    ram_cell[    5990] = 32'h1a2bc968;
    ram_cell[    5991] = 32'hd017978e;
    ram_cell[    5992] = 32'h377602f1;
    ram_cell[    5993] = 32'ha552be77;
    ram_cell[    5994] = 32'h970f2a76;
    ram_cell[    5995] = 32'he9f72bbe;
    ram_cell[    5996] = 32'h3b7d5b36;
    ram_cell[    5997] = 32'hcaf5a9fa;
    ram_cell[    5998] = 32'hd112f83b;
    ram_cell[    5999] = 32'h372f19ed;
    ram_cell[    6000] = 32'h023ae2c9;
    ram_cell[    6001] = 32'hea53caf6;
    ram_cell[    6002] = 32'hf3947e4d;
    ram_cell[    6003] = 32'h10b8b72d;
    ram_cell[    6004] = 32'hddaa791d;
    ram_cell[    6005] = 32'h02b43dd9;
    ram_cell[    6006] = 32'hc47b7b02;
    ram_cell[    6007] = 32'ha8d2f3f0;
    ram_cell[    6008] = 32'h6815e5d5;
    ram_cell[    6009] = 32'hf9bebc7e;
    ram_cell[    6010] = 32'h06dc76b6;
    ram_cell[    6011] = 32'hb441f3e6;
    ram_cell[    6012] = 32'h323a1b97;
    ram_cell[    6013] = 32'h86be9b3f;
    ram_cell[    6014] = 32'h289009d4;
    ram_cell[    6015] = 32'h56c2d770;
    ram_cell[    6016] = 32'h95184ac2;
    ram_cell[    6017] = 32'h62a3c45c;
    ram_cell[    6018] = 32'ha9e2e6fb;
    ram_cell[    6019] = 32'hb37d5bf3;
    ram_cell[    6020] = 32'h7bb8a223;
    ram_cell[    6021] = 32'h1d6b85ba;
    ram_cell[    6022] = 32'ha1955897;
    ram_cell[    6023] = 32'h127365e2;
    ram_cell[    6024] = 32'h36d9af96;
    ram_cell[    6025] = 32'h7c642160;
    ram_cell[    6026] = 32'hc47d1075;
    ram_cell[    6027] = 32'he91d61fa;
    ram_cell[    6028] = 32'h0d8c2f3d;
    ram_cell[    6029] = 32'h51de189f;
    ram_cell[    6030] = 32'hda5f4c68;
    ram_cell[    6031] = 32'hba2b39a5;
    ram_cell[    6032] = 32'h5a246554;
    ram_cell[    6033] = 32'h6dd10962;
    ram_cell[    6034] = 32'h035730b4;
    ram_cell[    6035] = 32'h589fde6d;
    ram_cell[    6036] = 32'hfab9930f;
    ram_cell[    6037] = 32'h7a2ffbfe;
    ram_cell[    6038] = 32'h264558b7;
    ram_cell[    6039] = 32'h31d5b7bd;
    ram_cell[    6040] = 32'h70b10189;
    ram_cell[    6041] = 32'ha15869ff;
    ram_cell[    6042] = 32'hf149eb18;
    ram_cell[    6043] = 32'h27234feb;
    ram_cell[    6044] = 32'h2db281cb;
    ram_cell[    6045] = 32'h4520183b;
    ram_cell[    6046] = 32'hd9c47c2c;
    ram_cell[    6047] = 32'h5a8a007c;
    ram_cell[    6048] = 32'h6715a6ea;
    ram_cell[    6049] = 32'hef382493;
    ram_cell[    6050] = 32'h33ff8b41;
    ram_cell[    6051] = 32'hcef36fce;
    ram_cell[    6052] = 32'h14672934;
    ram_cell[    6053] = 32'h20ec8e14;
    ram_cell[    6054] = 32'h51d778ef;
    ram_cell[    6055] = 32'hcbe27d45;
    ram_cell[    6056] = 32'he6b1e98c;
    ram_cell[    6057] = 32'h384ac47b;
    ram_cell[    6058] = 32'h9f5e3163;
    ram_cell[    6059] = 32'hfac9a1fc;
    ram_cell[    6060] = 32'h3391533b;
    ram_cell[    6061] = 32'hc3db6804;
    ram_cell[    6062] = 32'hc5a8f9e0;
    ram_cell[    6063] = 32'h2c8a3895;
    ram_cell[    6064] = 32'h5940e80f;
    ram_cell[    6065] = 32'hfd4002f5;
    ram_cell[    6066] = 32'hf7975644;
    ram_cell[    6067] = 32'h2b043be9;
    ram_cell[    6068] = 32'h3d151523;
    ram_cell[    6069] = 32'h1040c003;
    ram_cell[    6070] = 32'hc036bb0b;
    ram_cell[    6071] = 32'hc4bc054c;
    ram_cell[    6072] = 32'hfe1d55f1;
    ram_cell[    6073] = 32'hb244a7dc;
    ram_cell[    6074] = 32'h5c53c1ae;
    ram_cell[    6075] = 32'hc18ec4da;
    ram_cell[    6076] = 32'h40fced3a;
    ram_cell[    6077] = 32'h6b33c821;
    ram_cell[    6078] = 32'h829201f8;
    ram_cell[    6079] = 32'h63b2aaff;
    ram_cell[    6080] = 32'h7abcace0;
    ram_cell[    6081] = 32'hf5ed4449;
    ram_cell[    6082] = 32'he81c6d6a;
    ram_cell[    6083] = 32'h56763d55;
    ram_cell[    6084] = 32'hfcfa0822;
    ram_cell[    6085] = 32'h2d64f85a;
    ram_cell[    6086] = 32'hd9a84550;
    ram_cell[    6087] = 32'hc908aa14;
    ram_cell[    6088] = 32'hea31774e;
    ram_cell[    6089] = 32'hd9226723;
    ram_cell[    6090] = 32'hf0e56fbc;
    ram_cell[    6091] = 32'h74d82f04;
    ram_cell[    6092] = 32'hd505b899;
    ram_cell[    6093] = 32'hb4218c72;
    ram_cell[    6094] = 32'ha905308d;
    ram_cell[    6095] = 32'h3697f238;
    ram_cell[    6096] = 32'hd97af07b;
    ram_cell[    6097] = 32'hd79e14fe;
    ram_cell[    6098] = 32'hdf0e1b78;
    ram_cell[    6099] = 32'h83f52c50;
    ram_cell[    6100] = 32'h180533a9;
    ram_cell[    6101] = 32'h5f08843b;
    ram_cell[    6102] = 32'hfd660273;
    ram_cell[    6103] = 32'h5b45c6fc;
    ram_cell[    6104] = 32'hb25a77c8;
    ram_cell[    6105] = 32'h73dbb5c7;
    ram_cell[    6106] = 32'h0043349c;
    ram_cell[    6107] = 32'hd288a40d;
    ram_cell[    6108] = 32'h353c9aa4;
    ram_cell[    6109] = 32'h6930df18;
    ram_cell[    6110] = 32'h3cfad756;
    ram_cell[    6111] = 32'h95b392b7;
    ram_cell[    6112] = 32'h8ff735bd;
    ram_cell[    6113] = 32'hb6716ec4;
    ram_cell[    6114] = 32'hc6ca7895;
    ram_cell[    6115] = 32'h31c631e4;
    ram_cell[    6116] = 32'hc1c98d66;
    ram_cell[    6117] = 32'h8fcc7413;
    ram_cell[    6118] = 32'hfba71285;
    ram_cell[    6119] = 32'h9d183f13;
    ram_cell[    6120] = 32'hf799cc8a;
    ram_cell[    6121] = 32'h7fd049bc;
    ram_cell[    6122] = 32'h4fe0891e;
    ram_cell[    6123] = 32'h67f89e72;
    ram_cell[    6124] = 32'h8618b24f;
    ram_cell[    6125] = 32'h17efec26;
    ram_cell[    6126] = 32'h32f749c1;
    ram_cell[    6127] = 32'hdcc3c393;
    ram_cell[    6128] = 32'h9940ab62;
    ram_cell[    6129] = 32'h0d75f12f;
    ram_cell[    6130] = 32'h5ec8ea35;
    ram_cell[    6131] = 32'hb3085be4;
    ram_cell[    6132] = 32'h0662ba76;
    ram_cell[    6133] = 32'h8d77b915;
    ram_cell[    6134] = 32'hcb7c1a0a;
    ram_cell[    6135] = 32'hb2a9cbe1;
    ram_cell[    6136] = 32'h9a5d9ff4;
    ram_cell[    6137] = 32'hf7f6b5e9;
    ram_cell[    6138] = 32'h0563efa6;
    ram_cell[    6139] = 32'hb6d1c0d3;
    ram_cell[    6140] = 32'h0d9f0894;
    ram_cell[    6141] = 32'h3205aa8f;
    ram_cell[    6142] = 32'h66d8536a;
    ram_cell[    6143] = 32'hec423d63;
    ram_cell[    6144] = 32'h2f50ed04;
    ram_cell[    6145] = 32'h1f4cec99;
    ram_cell[    6146] = 32'h8df8156f;
    ram_cell[    6147] = 32'hfc5a4311;
    ram_cell[    6148] = 32'h7b849f67;
    ram_cell[    6149] = 32'hfe7f7544;
    ram_cell[    6150] = 32'ha062e71b;
    ram_cell[    6151] = 32'h95dad7bd;
    ram_cell[    6152] = 32'hdf924935;
    ram_cell[    6153] = 32'h4b28b123;
    ram_cell[    6154] = 32'h79295b5e;
    ram_cell[    6155] = 32'hda490c3a;
    ram_cell[    6156] = 32'h5c2f14af;
    ram_cell[    6157] = 32'he59fb090;
    ram_cell[    6158] = 32'h3e7bdda3;
    ram_cell[    6159] = 32'hc2e22b6a;
    ram_cell[    6160] = 32'he8d6161e;
    ram_cell[    6161] = 32'hb8651a5d;
    ram_cell[    6162] = 32'hcb0e7bea;
    ram_cell[    6163] = 32'heb5ab16f;
    ram_cell[    6164] = 32'h369b194c;
    ram_cell[    6165] = 32'h6674e736;
    ram_cell[    6166] = 32'h304d1395;
    ram_cell[    6167] = 32'hb5d65efc;
    ram_cell[    6168] = 32'hcc5d78ee;
    ram_cell[    6169] = 32'hb8909521;
    ram_cell[    6170] = 32'hd37f59b1;
    ram_cell[    6171] = 32'h820eb2b3;
    ram_cell[    6172] = 32'h3ce93eb4;
    ram_cell[    6173] = 32'h71523c0d;
    ram_cell[    6174] = 32'hd20fbca8;
    ram_cell[    6175] = 32'hcee8d31f;
    ram_cell[    6176] = 32'hbd696456;
    ram_cell[    6177] = 32'h74f5c8d6;
    ram_cell[    6178] = 32'hc2cbfc99;
    ram_cell[    6179] = 32'h562aae00;
    ram_cell[    6180] = 32'h8701fd66;
    ram_cell[    6181] = 32'h950662a6;
    ram_cell[    6182] = 32'h1f37a72d;
    ram_cell[    6183] = 32'h9e2f1184;
    ram_cell[    6184] = 32'hfa153d19;
    ram_cell[    6185] = 32'h7ba6b964;
    ram_cell[    6186] = 32'h61c583aa;
    ram_cell[    6187] = 32'hf483fdf3;
    ram_cell[    6188] = 32'hf20f2013;
    ram_cell[    6189] = 32'h36ee0230;
    ram_cell[    6190] = 32'h83868afa;
    ram_cell[    6191] = 32'he71edecb;
    ram_cell[    6192] = 32'h4c9b637d;
    ram_cell[    6193] = 32'hdf56cd4a;
    ram_cell[    6194] = 32'hbda6d9b9;
    ram_cell[    6195] = 32'h3f2237ec;
    ram_cell[    6196] = 32'hb593a0f8;
    ram_cell[    6197] = 32'hf49676e3;
    ram_cell[    6198] = 32'hca7c7b54;
    ram_cell[    6199] = 32'hf34373b3;
    ram_cell[    6200] = 32'h31f6a5bb;
    ram_cell[    6201] = 32'h133e4153;
    ram_cell[    6202] = 32'h1e6598d5;
    ram_cell[    6203] = 32'h250d1b49;
    ram_cell[    6204] = 32'h1368baf4;
    ram_cell[    6205] = 32'hc69fcd18;
    ram_cell[    6206] = 32'h6032ad96;
    ram_cell[    6207] = 32'hb6d0968d;
    ram_cell[    6208] = 32'h4315cc7f;
    ram_cell[    6209] = 32'hcd056593;
    ram_cell[    6210] = 32'h136bac8c;
    ram_cell[    6211] = 32'h6b5ce56d;
    ram_cell[    6212] = 32'h286020fd;
    ram_cell[    6213] = 32'h99fce3fb;
    ram_cell[    6214] = 32'ha32e419f;
    ram_cell[    6215] = 32'h0dfcb390;
    ram_cell[    6216] = 32'h545ca330;
    ram_cell[    6217] = 32'hba0da431;
    ram_cell[    6218] = 32'h64f5aaef;
    ram_cell[    6219] = 32'hcdc09e58;
    ram_cell[    6220] = 32'h9ac485d4;
    ram_cell[    6221] = 32'hc72d9766;
    ram_cell[    6222] = 32'h82d5392f;
    ram_cell[    6223] = 32'h234ee407;
    ram_cell[    6224] = 32'h7b8db2df;
    ram_cell[    6225] = 32'h8e953f31;
    ram_cell[    6226] = 32'h5f062006;
    ram_cell[    6227] = 32'h243db359;
    ram_cell[    6228] = 32'h5d7edf29;
    ram_cell[    6229] = 32'ha77d8cd3;
    ram_cell[    6230] = 32'h11334a8e;
    ram_cell[    6231] = 32'hef54f423;
    ram_cell[    6232] = 32'h58009363;
    ram_cell[    6233] = 32'h18b50ac9;
    ram_cell[    6234] = 32'h7c69cb13;
    ram_cell[    6235] = 32'h70c6c91a;
    ram_cell[    6236] = 32'ha1902e1f;
    ram_cell[    6237] = 32'h70b5451b;
    ram_cell[    6238] = 32'hed5eab5d;
    ram_cell[    6239] = 32'h9cf68f94;
    ram_cell[    6240] = 32'h7dabce58;
    ram_cell[    6241] = 32'hbc6a761e;
    ram_cell[    6242] = 32'hef240e3e;
    ram_cell[    6243] = 32'h321752b8;
    ram_cell[    6244] = 32'hd94d2bb8;
    ram_cell[    6245] = 32'h5f50e41f;
    ram_cell[    6246] = 32'hc3b55c3a;
    ram_cell[    6247] = 32'h2faf161a;
    ram_cell[    6248] = 32'h00bca2b1;
    ram_cell[    6249] = 32'h4902e1cb;
    ram_cell[    6250] = 32'hbf7a5ccf;
    ram_cell[    6251] = 32'hf61dafd1;
    ram_cell[    6252] = 32'he0a12ebc;
    ram_cell[    6253] = 32'h84a1ebeb;
    ram_cell[    6254] = 32'hb6d65f77;
    ram_cell[    6255] = 32'h4613c80a;
    ram_cell[    6256] = 32'hbcc3886f;
    ram_cell[    6257] = 32'hc6b7be82;
    ram_cell[    6258] = 32'h7c4b58e6;
    ram_cell[    6259] = 32'h7d5c1452;
    ram_cell[    6260] = 32'hec9551e1;
    ram_cell[    6261] = 32'h1ce2a2cb;
    ram_cell[    6262] = 32'hfee71a8b;
    ram_cell[    6263] = 32'h32c6b2de;
    ram_cell[    6264] = 32'haeab7598;
    ram_cell[    6265] = 32'hbcaad34f;
    ram_cell[    6266] = 32'hde571db7;
    ram_cell[    6267] = 32'h00e98057;
    ram_cell[    6268] = 32'haef42863;
    ram_cell[    6269] = 32'h3b1b017f;
    ram_cell[    6270] = 32'h86de8d2c;
    ram_cell[    6271] = 32'h30fcc086;
    ram_cell[    6272] = 32'hc8aa4c85;
    ram_cell[    6273] = 32'h8a37d015;
    ram_cell[    6274] = 32'h1dcba06d;
    ram_cell[    6275] = 32'hcc8cbffd;
    ram_cell[    6276] = 32'h2e416739;
    ram_cell[    6277] = 32'h0dd5a722;
    ram_cell[    6278] = 32'he9e5682f;
    ram_cell[    6279] = 32'hd929e2e3;
    ram_cell[    6280] = 32'h389bb17a;
    ram_cell[    6281] = 32'h3ad888c4;
    ram_cell[    6282] = 32'hc900d634;
    ram_cell[    6283] = 32'hb262312b;
    ram_cell[    6284] = 32'ha2de7187;
    ram_cell[    6285] = 32'h3f9a7f1a;
    ram_cell[    6286] = 32'hbc142c2d;
    ram_cell[    6287] = 32'h69f35955;
    ram_cell[    6288] = 32'h1748b419;
    ram_cell[    6289] = 32'hbb5d3539;
    ram_cell[    6290] = 32'h2074c4a1;
    ram_cell[    6291] = 32'h5cc1c581;
    ram_cell[    6292] = 32'h6258fda3;
    ram_cell[    6293] = 32'hd44fa493;
    ram_cell[    6294] = 32'h6383a140;
    ram_cell[    6295] = 32'h46d93553;
    ram_cell[    6296] = 32'h89805602;
    ram_cell[    6297] = 32'h35a30be7;
    ram_cell[    6298] = 32'h0ec3a620;
    ram_cell[    6299] = 32'h5533fdc9;
    ram_cell[    6300] = 32'h8456ba3b;
    ram_cell[    6301] = 32'hed63398b;
    ram_cell[    6302] = 32'hd2f8383c;
    ram_cell[    6303] = 32'hc666c137;
    ram_cell[    6304] = 32'h4740ab82;
    ram_cell[    6305] = 32'h88941747;
    ram_cell[    6306] = 32'h60e2693d;
    ram_cell[    6307] = 32'h1e7d337b;
    ram_cell[    6308] = 32'h5921894e;
    ram_cell[    6309] = 32'hdfe234b8;
    ram_cell[    6310] = 32'h543ce2cd;
    ram_cell[    6311] = 32'h34803c6c;
    ram_cell[    6312] = 32'h24385635;
    ram_cell[    6313] = 32'h6d151a19;
    ram_cell[    6314] = 32'h59635f9a;
    ram_cell[    6315] = 32'h3525d3e4;
    ram_cell[    6316] = 32'h6607a64c;
    ram_cell[    6317] = 32'h194cce68;
    ram_cell[    6318] = 32'hdc81a37c;
    ram_cell[    6319] = 32'h2101467f;
    ram_cell[    6320] = 32'h7309f27f;
    ram_cell[    6321] = 32'h9c000286;
    ram_cell[    6322] = 32'ha114d5ac;
    ram_cell[    6323] = 32'hc904a1ac;
    ram_cell[    6324] = 32'hf28eeb1d;
    ram_cell[    6325] = 32'h2fde155d;
    ram_cell[    6326] = 32'h85aabb70;
    ram_cell[    6327] = 32'hc5c32ba8;
    ram_cell[    6328] = 32'h9794bc88;
    ram_cell[    6329] = 32'h06f1e83a;
    ram_cell[    6330] = 32'hca27b051;
    ram_cell[    6331] = 32'h5c251885;
    ram_cell[    6332] = 32'he37c9f5f;
    ram_cell[    6333] = 32'h8e9ee756;
    ram_cell[    6334] = 32'h8cf1f21b;
    ram_cell[    6335] = 32'h3ac3bf3c;
    ram_cell[    6336] = 32'h04b7b4e1;
    ram_cell[    6337] = 32'h0378dcab;
    ram_cell[    6338] = 32'h501c5036;
    ram_cell[    6339] = 32'he9a44228;
    ram_cell[    6340] = 32'hc27de831;
    ram_cell[    6341] = 32'h967e3d51;
    ram_cell[    6342] = 32'he32a4a6c;
    ram_cell[    6343] = 32'h8c8deaca;
    ram_cell[    6344] = 32'h1ed86b37;
    ram_cell[    6345] = 32'heb99f142;
    ram_cell[    6346] = 32'hb352a7b8;
    ram_cell[    6347] = 32'h46d336e9;
    ram_cell[    6348] = 32'h58476458;
    ram_cell[    6349] = 32'h2a02d62b;
    ram_cell[    6350] = 32'h724fef89;
    ram_cell[    6351] = 32'h51697589;
    ram_cell[    6352] = 32'hfb0961aa;
    ram_cell[    6353] = 32'h7560b76e;
    ram_cell[    6354] = 32'hda2461e0;
    ram_cell[    6355] = 32'h9beea56f;
    ram_cell[    6356] = 32'h717e2746;
    ram_cell[    6357] = 32'h846d1c2a;
    ram_cell[    6358] = 32'h7d748b58;
    ram_cell[    6359] = 32'h4a0e8180;
    ram_cell[    6360] = 32'hf9d1d449;
    ram_cell[    6361] = 32'h26113ab9;
    ram_cell[    6362] = 32'h7d5fbc4a;
    ram_cell[    6363] = 32'h11e7be49;
    ram_cell[    6364] = 32'h13760009;
    ram_cell[    6365] = 32'hc1141bb2;
    ram_cell[    6366] = 32'hf6594673;
    ram_cell[    6367] = 32'h01fd2c50;
    ram_cell[    6368] = 32'h23f26471;
    ram_cell[    6369] = 32'h9ef7c5f4;
    ram_cell[    6370] = 32'hd8549957;
    ram_cell[    6371] = 32'h30bd98f1;
    ram_cell[    6372] = 32'ha6ca9e9c;
    ram_cell[    6373] = 32'h57b05604;
    ram_cell[    6374] = 32'hc0390a70;
    ram_cell[    6375] = 32'h6a015a57;
    ram_cell[    6376] = 32'hfeffa01a;
    ram_cell[    6377] = 32'h4615cf47;
    ram_cell[    6378] = 32'hd3e7a66f;
    ram_cell[    6379] = 32'h5b6159ec;
    ram_cell[    6380] = 32'h4f440f99;
    ram_cell[    6381] = 32'h3473728d;
    ram_cell[    6382] = 32'h5efc40f4;
    ram_cell[    6383] = 32'h1b688dc9;
    ram_cell[    6384] = 32'h6144f943;
    ram_cell[    6385] = 32'h138cca93;
    ram_cell[    6386] = 32'h8c80d94d;
    ram_cell[    6387] = 32'h73ed1474;
    ram_cell[    6388] = 32'h679c7134;
    ram_cell[    6389] = 32'h11603168;
    ram_cell[    6390] = 32'h777cf8c7;
    ram_cell[    6391] = 32'h8afb2cc0;
    ram_cell[    6392] = 32'hb4af5159;
    ram_cell[    6393] = 32'h9e11d2bb;
    ram_cell[    6394] = 32'hffd2dd21;
    ram_cell[    6395] = 32'h10b95aba;
    ram_cell[    6396] = 32'h260d9425;
    ram_cell[    6397] = 32'h9a27b00a;
    ram_cell[    6398] = 32'hee54b31e;
    ram_cell[    6399] = 32'h5ea482e8;
    ram_cell[    6400] = 32'hb4d8e261;
    ram_cell[    6401] = 32'h91d3f525;
    ram_cell[    6402] = 32'h3180a019;
    ram_cell[    6403] = 32'h46bf015d;
    ram_cell[    6404] = 32'hb9eaffbf;
    ram_cell[    6405] = 32'h74867a3a;
    ram_cell[    6406] = 32'h697c4001;
    ram_cell[    6407] = 32'h39269ff0;
    ram_cell[    6408] = 32'h490bac6c;
    ram_cell[    6409] = 32'h83a886c6;
    ram_cell[    6410] = 32'h7a6a2aa0;
    ram_cell[    6411] = 32'hdee4697a;
    ram_cell[    6412] = 32'h202d8467;
    ram_cell[    6413] = 32'he16a73c9;
    ram_cell[    6414] = 32'h610b0773;
    ram_cell[    6415] = 32'hdf206bef;
    ram_cell[    6416] = 32'hff8133f2;
    ram_cell[    6417] = 32'h62a63bb1;
    ram_cell[    6418] = 32'h09ec9f80;
    ram_cell[    6419] = 32'hcb9ec2f6;
    ram_cell[    6420] = 32'ha2af6809;
    ram_cell[    6421] = 32'h6fe254f4;
    ram_cell[    6422] = 32'h22b85d5c;
    ram_cell[    6423] = 32'h79edc41c;
    ram_cell[    6424] = 32'h8ece7d14;
    ram_cell[    6425] = 32'h464fbbc1;
    ram_cell[    6426] = 32'h235eb8fe;
    ram_cell[    6427] = 32'h314e0455;
    ram_cell[    6428] = 32'h8832b7c3;
    ram_cell[    6429] = 32'h53a6d12b;
    ram_cell[    6430] = 32'hbce0a95c;
    ram_cell[    6431] = 32'h6064db1f;
    ram_cell[    6432] = 32'h67d5f796;
    ram_cell[    6433] = 32'hbd63173c;
    ram_cell[    6434] = 32'h074a2f3e;
    ram_cell[    6435] = 32'h07d60fe5;
    ram_cell[    6436] = 32'h10e124cb;
    ram_cell[    6437] = 32'h40d1e0d2;
    ram_cell[    6438] = 32'h2146e989;
    ram_cell[    6439] = 32'h9d65681a;
    ram_cell[    6440] = 32'h0807f464;
    ram_cell[    6441] = 32'hccd4ff64;
    ram_cell[    6442] = 32'h658d0cf4;
    ram_cell[    6443] = 32'h2d84a978;
    ram_cell[    6444] = 32'h6be8fc47;
    ram_cell[    6445] = 32'h698d36a0;
    ram_cell[    6446] = 32'h566f4cea;
    ram_cell[    6447] = 32'ha9f40cc8;
    ram_cell[    6448] = 32'h5fd1cec2;
    ram_cell[    6449] = 32'h0a79cd42;
    ram_cell[    6450] = 32'h95646c22;
    ram_cell[    6451] = 32'h6d38b0b3;
    ram_cell[    6452] = 32'h03f9046e;
    ram_cell[    6453] = 32'hffa759f7;
    ram_cell[    6454] = 32'h8a4635d7;
    ram_cell[    6455] = 32'h0c0d355c;
    ram_cell[    6456] = 32'hc7310907;
    ram_cell[    6457] = 32'h2f461aaf;
    ram_cell[    6458] = 32'h3a204ccc;
    ram_cell[    6459] = 32'h1e34f076;
    ram_cell[    6460] = 32'h5f1afff6;
    ram_cell[    6461] = 32'h18da8798;
    ram_cell[    6462] = 32'h98f8821c;
    ram_cell[    6463] = 32'h32680705;
    ram_cell[    6464] = 32'ha3626be9;
    ram_cell[    6465] = 32'h0559b019;
    ram_cell[    6466] = 32'h8e41cf46;
    ram_cell[    6467] = 32'h32acfb83;
    ram_cell[    6468] = 32'h3f737700;
    ram_cell[    6469] = 32'h838bc4d3;
    ram_cell[    6470] = 32'heefe02fa;
    ram_cell[    6471] = 32'h5ec94c0a;
    ram_cell[    6472] = 32'hf105cb04;
    ram_cell[    6473] = 32'hed2db70b;
    ram_cell[    6474] = 32'h03af48fb;
    ram_cell[    6475] = 32'hc0f1436d;
    ram_cell[    6476] = 32'h58f4c65a;
    ram_cell[    6477] = 32'he686f568;
    ram_cell[    6478] = 32'haa762ae1;
    ram_cell[    6479] = 32'h05df8fbe;
    ram_cell[    6480] = 32'hc294a378;
    ram_cell[    6481] = 32'h6d113f7c;
    ram_cell[    6482] = 32'h2c79311e;
    ram_cell[    6483] = 32'hea20c335;
    ram_cell[    6484] = 32'h1c6309e7;
    ram_cell[    6485] = 32'h4e04f0d4;
    ram_cell[    6486] = 32'h037f2bf6;
    ram_cell[    6487] = 32'h8364cf55;
    ram_cell[    6488] = 32'h8dffff6a;
    ram_cell[    6489] = 32'h44d3d8f1;
    ram_cell[    6490] = 32'hcf1fcda1;
    ram_cell[    6491] = 32'h680ce19d;
    ram_cell[    6492] = 32'h41f9db91;
    ram_cell[    6493] = 32'h09531250;
    ram_cell[    6494] = 32'h34099eac;
    ram_cell[    6495] = 32'hb0e6b302;
    ram_cell[    6496] = 32'hea589af3;
    ram_cell[    6497] = 32'hc33b9fca;
    ram_cell[    6498] = 32'h23a3bba5;
    ram_cell[    6499] = 32'h5c2d710f;
    ram_cell[    6500] = 32'hf4036bc1;
    ram_cell[    6501] = 32'hc06c5e24;
    ram_cell[    6502] = 32'h0fca6bbd;
    ram_cell[    6503] = 32'h6a789c56;
    ram_cell[    6504] = 32'h890da26b;
    ram_cell[    6505] = 32'h49a9bf1f;
    ram_cell[    6506] = 32'h8f81cd04;
    ram_cell[    6507] = 32'hd1527d0e;
    ram_cell[    6508] = 32'h39bb363e;
    ram_cell[    6509] = 32'heef4c231;
    ram_cell[    6510] = 32'h1d3a860e;
    ram_cell[    6511] = 32'h0d01626f;
    ram_cell[    6512] = 32'h922883f5;
    ram_cell[    6513] = 32'hb011920a;
    ram_cell[    6514] = 32'hf3845bcf;
    ram_cell[    6515] = 32'h392476ff;
    ram_cell[    6516] = 32'ha2aa2319;
    ram_cell[    6517] = 32'haab5b69b;
    ram_cell[    6518] = 32'hfc94f49c;
    ram_cell[    6519] = 32'hbd4a0154;
    ram_cell[    6520] = 32'h3efc6795;
    ram_cell[    6521] = 32'hfb19fc5d;
    ram_cell[    6522] = 32'h90279b24;
    ram_cell[    6523] = 32'h4661809f;
    ram_cell[    6524] = 32'h39454898;
    ram_cell[    6525] = 32'h454cce08;
    ram_cell[    6526] = 32'h309d6ec5;
    ram_cell[    6527] = 32'hfa710891;
    ram_cell[    6528] = 32'ha972cc94;
    ram_cell[    6529] = 32'ha6d81b40;
    ram_cell[    6530] = 32'ha0bb6b04;
    ram_cell[    6531] = 32'h9cf3eddd;
    ram_cell[    6532] = 32'h50c285cb;
    ram_cell[    6533] = 32'h2c9b2139;
    ram_cell[    6534] = 32'h2f6ca947;
    ram_cell[    6535] = 32'h7da4d9a4;
    ram_cell[    6536] = 32'h7ceb0f6d;
    ram_cell[    6537] = 32'h50240f2e;
    ram_cell[    6538] = 32'h6a3796b4;
    ram_cell[    6539] = 32'h7c3ea65f;
    ram_cell[    6540] = 32'he06af3e8;
    ram_cell[    6541] = 32'hcbef88b4;
    ram_cell[    6542] = 32'h9464a8e5;
    ram_cell[    6543] = 32'hc2e2f7d0;
    ram_cell[    6544] = 32'hdef34b2c;
    ram_cell[    6545] = 32'h3c7a36b6;
    ram_cell[    6546] = 32'hd5e50cc5;
    ram_cell[    6547] = 32'h33b2062a;
    ram_cell[    6548] = 32'h0d635d43;
    ram_cell[    6549] = 32'ha0825998;
    ram_cell[    6550] = 32'h17572bee;
    ram_cell[    6551] = 32'h534019ee;
    ram_cell[    6552] = 32'hc5027aa3;
    ram_cell[    6553] = 32'h293240ba;
    ram_cell[    6554] = 32'hfcd35123;
    ram_cell[    6555] = 32'ha362d178;
    ram_cell[    6556] = 32'h412a8296;
    ram_cell[    6557] = 32'hdc1fa420;
    ram_cell[    6558] = 32'hc7849d7f;
    ram_cell[    6559] = 32'h3a1f4247;
    ram_cell[    6560] = 32'hb5e37adb;
    ram_cell[    6561] = 32'hbd41016d;
    ram_cell[    6562] = 32'h032354d0;
    ram_cell[    6563] = 32'hafeec2a4;
    ram_cell[    6564] = 32'hf9647919;
    ram_cell[    6565] = 32'ha8c7b655;
    ram_cell[    6566] = 32'h97656fbe;
    ram_cell[    6567] = 32'ha70b9c49;
    ram_cell[    6568] = 32'hf4402d04;
    ram_cell[    6569] = 32'hb96e1822;
    ram_cell[    6570] = 32'hdcd39bd0;
    ram_cell[    6571] = 32'h848b4a41;
    ram_cell[    6572] = 32'h7ee84c59;
    ram_cell[    6573] = 32'h1613a689;
    ram_cell[    6574] = 32'hd667e224;
    ram_cell[    6575] = 32'h63bc8e41;
    ram_cell[    6576] = 32'h8255a8ba;
    ram_cell[    6577] = 32'h100ae8d8;
    ram_cell[    6578] = 32'h03c0830a;
    ram_cell[    6579] = 32'he768f8b9;
    ram_cell[    6580] = 32'he699d8ae;
    ram_cell[    6581] = 32'h96efe6be;
    ram_cell[    6582] = 32'ha4e7a976;
    ram_cell[    6583] = 32'hf848307a;
    ram_cell[    6584] = 32'h694d46a8;
    ram_cell[    6585] = 32'hed58cafd;
    ram_cell[    6586] = 32'hf9c1ed07;
    ram_cell[    6587] = 32'h8a39658b;
    ram_cell[    6588] = 32'hd985e461;
    ram_cell[    6589] = 32'hfce0d0ed;
    ram_cell[    6590] = 32'h4cd330a3;
    ram_cell[    6591] = 32'hf93c6a21;
    ram_cell[    6592] = 32'h8880ef25;
    ram_cell[    6593] = 32'h19bf664d;
    ram_cell[    6594] = 32'h6dc26ed9;
    ram_cell[    6595] = 32'h2353f8f5;
    ram_cell[    6596] = 32'h5b48b1c6;
    ram_cell[    6597] = 32'h4a861b6e;
    ram_cell[    6598] = 32'he8fb19c3;
    ram_cell[    6599] = 32'h0b9c9235;
    ram_cell[    6600] = 32'h0b2364d8;
    ram_cell[    6601] = 32'h6485d3bd;
    ram_cell[    6602] = 32'hea79f8ae;
    ram_cell[    6603] = 32'h88dde358;
    ram_cell[    6604] = 32'h6211095b;
    ram_cell[    6605] = 32'h74933b5b;
    ram_cell[    6606] = 32'h0dc7b7c2;
    ram_cell[    6607] = 32'h0a0593b2;
    ram_cell[    6608] = 32'h4b4b1484;
    ram_cell[    6609] = 32'h676c8867;
    ram_cell[    6610] = 32'hc0f22b21;
    ram_cell[    6611] = 32'h2c54541d;
    ram_cell[    6612] = 32'hbd097c06;
    ram_cell[    6613] = 32'hfcdbb2c8;
    ram_cell[    6614] = 32'h62e33a11;
    ram_cell[    6615] = 32'hace5effd;
    ram_cell[    6616] = 32'hd1b1e768;
    ram_cell[    6617] = 32'he566a3c7;
    ram_cell[    6618] = 32'h83c12b3f;
    ram_cell[    6619] = 32'hfa37422d;
    ram_cell[    6620] = 32'hec980b95;
    ram_cell[    6621] = 32'h804908d7;
    ram_cell[    6622] = 32'h3b02a79d;
    ram_cell[    6623] = 32'h402694ae;
    ram_cell[    6624] = 32'h93b0b0c8;
    ram_cell[    6625] = 32'hf99b4ad2;
    ram_cell[    6626] = 32'h8d9bd51b;
    ram_cell[    6627] = 32'h0bebeab1;
    ram_cell[    6628] = 32'hbac78011;
    ram_cell[    6629] = 32'h5b4b8e8c;
    ram_cell[    6630] = 32'ha8e0a424;
    ram_cell[    6631] = 32'haece5bbb;
    ram_cell[    6632] = 32'h82df8f8e;
    ram_cell[    6633] = 32'hd1999cf2;
    ram_cell[    6634] = 32'h38812724;
    ram_cell[    6635] = 32'heb4d8730;
    ram_cell[    6636] = 32'h197d2954;
    ram_cell[    6637] = 32'h890502b7;
    ram_cell[    6638] = 32'hdc969a90;
    ram_cell[    6639] = 32'h1321e7ca;
    ram_cell[    6640] = 32'h4edd59a2;
    ram_cell[    6641] = 32'h934f160d;
    ram_cell[    6642] = 32'hfd10a1e5;
    ram_cell[    6643] = 32'hf29ea65b;
    ram_cell[    6644] = 32'he4116b01;
    ram_cell[    6645] = 32'h26a1b2ca;
    ram_cell[    6646] = 32'h077ade5b;
    ram_cell[    6647] = 32'h72c65bb8;
    ram_cell[    6648] = 32'ha2cc2844;
    ram_cell[    6649] = 32'hbeeab91d;
    ram_cell[    6650] = 32'h94d0b1b2;
    ram_cell[    6651] = 32'h34d8aac0;
    ram_cell[    6652] = 32'hdd4d6dcb;
    ram_cell[    6653] = 32'ha1e19654;
    ram_cell[    6654] = 32'h94be888c;
    ram_cell[    6655] = 32'hbe836f7b;
    ram_cell[    6656] = 32'h9e57a791;
    ram_cell[    6657] = 32'h897f418d;
    ram_cell[    6658] = 32'hcd5413f3;
    ram_cell[    6659] = 32'hea850978;
    ram_cell[    6660] = 32'h2a6e4c63;
    ram_cell[    6661] = 32'hb49d3bad;
    ram_cell[    6662] = 32'h65f6237d;
    ram_cell[    6663] = 32'h4c7e0195;
    ram_cell[    6664] = 32'h5cd6c588;
    ram_cell[    6665] = 32'h35259da4;
    ram_cell[    6666] = 32'hac2208e3;
    ram_cell[    6667] = 32'h5c7ea043;
    ram_cell[    6668] = 32'hb5d55150;
    ram_cell[    6669] = 32'hb17bfb3e;
    ram_cell[    6670] = 32'h6993358a;
    ram_cell[    6671] = 32'hde62a3f0;
    ram_cell[    6672] = 32'hff127502;
    ram_cell[    6673] = 32'hd60f8c9b;
    ram_cell[    6674] = 32'hb58cf3c2;
    ram_cell[    6675] = 32'had53aa3e;
    ram_cell[    6676] = 32'h1ce63b29;
    ram_cell[    6677] = 32'he8be89ff;
    ram_cell[    6678] = 32'haeeaa504;
    ram_cell[    6679] = 32'ha2e0f532;
    ram_cell[    6680] = 32'h48244bfb;
    ram_cell[    6681] = 32'h44d406dc;
    ram_cell[    6682] = 32'h290d6469;
    ram_cell[    6683] = 32'h4bc9c609;
    ram_cell[    6684] = 32'h4c79a7cf;
    ram_cell[    6685] = 32'h2bbe0297;
    ram_cell[    6686] = 32'h98be7ea4;
    ram_cell[    6687] = 32'ha8630ecc;
    ram_cell[    6688] = 32'h284c5a7d;
    ram_cell[    6689] = 32'h499132e9;
    ram_cell[    6690] = 32'he99517b7;
    ram_cell[    6691] = 32'h832f1ff7;
    ram_cell[    6692] = 32'he0a3996a;
    ram_cell[    6693] = 32'h609a3f16;
    ram_cell[    6694] = 32'h957bd311;
    ram_cell[    6695] = 32'hfd51eab8;
    ram_cell[    6696] = 32'h56752ac6;
    ram_cell[    6697] = 32'h3d4b6943;
    ram_cell[    6698] = 32'h0d7440bf;
    ram_cell[    6699] = 32'hfadb7090;
    ram_cell[    6700] = 32'h89454c93;
    ram_cell[    6701] = 32'hd2842c64;
    ram_cell[    6702] = 32'h876fb518;
    ram_cell[    6703] = 32'h9b7acab9;
    ram_cell[    6704] = 32'ha0f5c79f;
    ram_cell[    6705] = 32'h98e6b3ec;
    ram_cell[    6706] = 32'h999c91e3;
    ram_cell[    6707] = 32'h88b05886;
    ram_cell[    6708] = 32'h677e8e29;
    ram_cell[    6709] = 32'h5bbf78e6;
    ram_cell[    6710] = 32'hdecec63a;
    ram_cell[    6711] = 32'hb14e9c5f;
    ram_cell[    6712] = 32'hdb200bd8;
    ram_cell[    6713] = 32'h2893f7cd;
    ram_cell[    6714] = 32'hdc9f9d88;
    ram_cell[    6715] = 32'h67c69fb4;
    ram_cell[    6716] = 32'h1405f46f;
    ram_cell[    6717] = 32'hf213c1bd;
    ram_cell[    6718] = 32'h63d18fec;
    ram_cell[    6719] = 32'hd4820c11;
    ram_cell[    6720] = 32'hbfafb214;
    ram_cell[    6721] = 32'h88301316;
    ram_cell[    6722] = 32'h01043d39;
    ram_cell[    6723] = 32'h97fac42c;
    ram_cell[    6724] = 32'h80980a65;
    ram_cell[    6725] = 32'hda6dbd45;
    ram_cell[    6726] = 32'h66b6019a;
    ram_cell[    6727] = 32'h284b1056;
    ram_cell[    6728] = 32'h4f1a13db;
    ram_cell[    6729] = 32'hd3439a49;
    ram_cell[    6730] = 32'h97c8c30d;
    ram_cell[    6731] = 32'h55aa8151;
    ram_cell[    6732] = 32'he159d6d8;
    ram_cell[    6733] = 32'h6e76b3f7;
    ram_cell[    6734] = 32'h1060b472;
    ram_cell[    6735] = 32'hd33e22c0;
    ram_cell[    6736] = 32'hc33ea95f;
    ram_cell[    6737] = 32'h80bd76ea;
    ram_cell[    6738] = 32'hc28087bb;
    ram_cell[    6739] = 32'h8d5f8861;
    ram_cell[    6740] = 32'hacfb6efe;
    ram_cell[    6741] = 32'h99df5261;
    ram_cell[    6742] = 32'h9b960158;
    ram_cell[    6743] = 32'h5776a0ea;
    ram_cell[    6744] = 32'h5487ca6c;
    ram_cell[    6745] = 32'hea826644;
    ram_cell[    6746] = 32'h0835675d;
    ram_cell[    6747] = 32'h3a545a3c;
    ram_cell[    6748] = 32'h2c99d365;
    ram_cell[    6749] = 32'hd718c167;
    ram_cell[    6750] = 32'h5ce95296;
    ram_cell[    6751] = 32'he5895f56;
    ram_cell[    6752] = 32'h6eb3d4c4;
    ram_cell[    6753] = 32'h7c283835;
    ram_cell[    6754] = 32'h99553cc8;
    ram_cell[    6755] = 32'h4a899c82;
    ram_cell[    6756] = 32'h22675e71;
    ram_cell[    6757] = 32'h1dcc8a48;
    ram_cell[    6758] = 32'h136f9e48;
    ram_cell[    6759] = 32'h3167e9ec;
    ram_cell[    6760] = 32'h9a7e3547;
    ram_cell[    6761] = 32'hebda3c3c;
    ram_cell[    6762] = 32'h828ec2f0;
    ram_cell[    6763] = 32'h4a316203;
    ram_cell[    6764] = 32'hf890803f;
    ram_cell[    6765] = 32'h29156226;
    ram_cell[    6766] = 32'h8f0a1854;
    ram_cell[    6767] = 32'h425c7ee4;
    ram_cell[    6768] = 32'h86108250;
    ram_cell[    6769] = 32'h125414ec;
    ram_cell[    6770] = 32'h14ad1990;
    ram_cell[    6771] = 32'h50c7e9cd;
    ram_cell[    6772] = 32'hd9386586;
    ram_cell[    6773] = 32'h4ecb8f86;
    ram_cell[    6774] = 32'hbe6acba5;
    ram_cell[    6775] = 32'h27a51cb6;
    ram_cell[    6776] = 32'he30c744c;
    ram_cell[    6777] = 32'hdff981fb;
    ram_cell[    6778] = 32'h7304a8aa;
    ram_cell[    6779] = 32'h549018ca;
    ram_cell[    6780] = 32'h2f927d37;
    ram_cell[    6781] = 32'h9362cbda;
    ram_cell[    6782] = 32'h610e1a9b;
    ram_cell[    6783] = 32'h3de1c5b9;
    ram_cell[    6784] = 32'h44884111;
    ram_cell[    6785] = 32'h0e977f0c;
    ram_cell[    6786] = 32'h8da519e3;
    ram_cell[    6787] = 32'h4b7d4e03;
    ram_cell[    6788] = 32'h53b266b7;
    ram_cell[    6789] = 32'h2c9882e1;
    ram_cell[    6790] = 32'hc6840766;
    ram_cell[    6791] = 32'h3490a4e2;
    ram_cell[    6792] = 32'hd9820fbb;
    ram_cell[    6793] = 32'hb69b0ecf;
    ram_cell[    6794] = 32'ha377a2b0;
    ram_cell[    6795] = 32'h25ef58d0;
    ram_cell[    6796] = 32'h00cc9aaa;
    ram_cell[    6797] = 32'hecacfcf7;
    ram_cell[    6798] = 32'h1ef71189;
    ram_cell[    6799] = 32'h2185bd5f;
    ram_cell[    6800] = 32'h27631671;
    ram_cell[    6801] = 32'hce120b17;
    ram_cell[    6802] = 32'h3a38160e;
    ram_cell[    6803] = 32'heaa72bdd;
    ram_cell[    6804] = 32'h3a49d894;
    ram_cell[    6805] = 32'h3dbb7287;
    ram_cell[    6806] = 32'hcdbb9a64;
    ram_cell[    6807] = 32'h32054706;
    ram_cell[    6808] = 32'h0c1e8b56;
    ram_cell[    6809] = 32'h55e49687;
    ram_cell[    6810] = 32'h478f41ec;
    ram_cell[    6811] = 32'hd6a98974;
    ram_cell[    6812] = 32'h06d6b7dd;
    ram_cell[    6813] = 32'h4e783925;
    ram_cell[    6814] = 32'hcf21f1bb;
    ram_cell[    6815] = 32'hebe451a8;
    ram_cell[    6816] = 32'he91f808f;
    ram_cell[    6817] = 32'h0c118d12;
    ram_cell[    6818] = 32'h973013a2;
    ram_cell[    6819] = 32'ha5060741;
    ram_cell[    6820] = 32'h5ae99b3c;
    ram_cell[    6821] = 32'h2dba4484;
    ram_cell[    6822] = 32'h0b459fb5;
    ram_cell[    6823] = 32'hc61e13ee;
    ram_cell[    6824] = 32'h5b26d303;
    ram_cell[    6825] = 32'h47e2a626;
    ram_cell[    6826] = 32'h91b6460e;
    ram_cell[    6827] = 32'h85952d1b;
    ram_cell[    6828] = 32'h33bd9fdd;
    ram_cell[    6829] = 32'h655c7ed7;
    ram_cell[    6830] = 32'h25d66437;
    ram_cell[    6831] = 32'h3b8134e4;
    ram_cell[    6832] = 32'h15514380;
    ram_cell[    6833] = 32'h7651b111;
    ram_cell[    6834] = 32'h825b39f9;
    ram_cell[    6835] = 32'h85ab7587;
    ram_cell[    6836] = 32'h0bdbdb21;
    ram_cell[    6837] = 32'hbeefdbe7;
    ram_cell[    6838] = 32'h2eda8a16;
    ram_cell[    6839] = 32'he4b972ac;
    ram_cell[    6840] = 32'he2ff9dd8;
    ram_cell[    6841] = 32'h75191852;
    ram_cell[    6842] = 32'hb2931bae;
    ram_cell[    6843] = 32'hba0a2189;
    ram_cell[    6844] = 32'haf7314b4;
    ram_cell[    6845] = 32'h8008a276;
    ram_cell[    6846] = 32'hf58eb942;
    ram_cell[    6847] = 32'h40db48e3;
    ram_cell[    6848] = 32'h6a1a75f9;
    ram_cell[    6849] = 32'h4cc0d287;
    ram_cell[    6850] = 32'hf7301913;
    ram_cell[    6851] = 32'h9340cdad;
    ram_cell[    6852] = 32'hcf968aa9;
    ram_cell[    6853] = 32'hf707b954;
    ram_cell[    6854] = 32'h87911e86;
    ram_cell[    6855] = 32'hc74433d5;
    ram_cell[    6856] = 32'h05c0d80b;
    ram_cell[    6857] = 32'h38ba09e1;
    ram_cell[    6858] = 32'h269d74cf;
    ram_cell[    6859] = 32'h6a3b4c9e;
    ram_cell[    6860] = 32'hbc1dc098;
    ram_cell[    6861] = 32'h8a6aabbb;
    ram_cell[    6862] = 32'h136762bf;
    ram_cell[    6863] = 32'haa8a9f9c;
    ram_cell[    6864] = 32'h65f87bc4;
    ram_cell[    6865] = 32'h0a07f82c;
    ram_cell[    6866] = 32'hc1e2649e;
    ram_cell[    6867] = 32'h901e82a7;
    ram_cell[    6868] = 32'hffa9509a;
    ram_cell[    6869] = 32'hbfba2c88;
    ram_cell[    6870] = 32'h60980dea;
    ram_cell[    6871] = 32'h102ce960;
    ram_cell[    6872] = 32'h8e0b223a;
    ram_cell[    6873] = 32'h799fd5c8;
    ram_cell[    6874] = 32'h6dd6781f;
    ram_cell[    6875] = 32'hfa15b80e;
    ram_cell[    6876] = 32'hd022dc74;
    ram_cell[    6877] = 32'hd56773cd;
    ram_cell[    6878] = 32'h07de9ec5;
    ram_cell[    6879] = 32'h85702aa0;
    ram_cell[    6880] = 32'h91ceab12;
    ram_cell[    6881] = 32'h75f20f94;
    ram_cell[    6882] = 32'h3108a2e8;
    ram_cell[    6883] = 32'hd5a071af;
    ram_cell[    6884] = 32'hf0a7ca13;
    ram_cell[    6885] = 32'hcbf26060;
    ram_cell[    6886] = 32'ha9cf8a25;
    ram_cell[    6887] = 32'h8324335d;
    ram_cell[    6888] = 32'h3cc5be46;
    ram_cell[    6889] = 32'h73c41caa;
    ram_cell[    6890] = 32'hb8b4fad0;
    ram_cell[    6891] = 32'hd3384916;
    ram_cell[    6892] = 32'had3151ca;
    ram_cell[    6893] = 32'h0f879ce2;
    ram_cell[    6894] = 32'h9711217b;
    ram_cell[    6895] = 32'hd3c72df6;
    ram_cell[    6896] = 32'h1fbd2721;
    ram_cell[    6897] = 32'h9ac01fc0;
    ram_cell[    6898] = 32'hffa11c96;
    ram_cell[    6899] = 32'h51662965;
    ram_cell[    6900] = 32'h68cba8bd;
    ram_cell[    6901] = 32'h510d5d48;
    ram_cell[    6902] = 32'hdf84ed15;
    ram_cell[    6903] = 32'hc0471a0f;
    ram_cell[    6904] = 32'h4ac5ebbb;
    ram_cell[    6905] = 32'he9082247;
    ram_cell[    6906] = 32'h8a909075;
    ram_cell[    6907] = 32'h959a6d9a;
    ram_cell[    6908] = 32'h98003c35;
    ram_cell[    6909] = 32'h90910bd8;
    ram_cell[    6910] = 32'h000f6b32;
    ram_cell[    6911] = 32'hb0af853c;
    ram_cell[    6912] = 32'h1eba7078;
    ram_cell[    6913] = 32'h5b91d5e7;
    ram_cell[    6914] = 32'h9897e59f;
    ram_cell[    6915] = 32'hbabe508f;
    ram_cell[    6916] = 32'h1daee5a8;
    ram_cell[    6917] = 32'hd467188e;
    ram_cell[    6918] = 32'hae54b50f;
    ram_cell[    6919] = 32'h699eac8d;
    ram_cell[    6920] = 32'h9a1987bf;
    ram_cell[    6921] = 32'h26f6969d;
    ram_cell[    6922] = 32'h0eefcb1f;
    ram_cell[    6923] = 32'hcdd02045;
    ram_cell[    6924] = 32'ha7f3dba0;
    ram_cell[    6925] = 32'hade9d7b9;
    ram_cell[    6926] = 32'hf07e6707;
    ram_cell[    6927] = 32'hea10bd9d;
    ram_cell[    6928] = 32'hf4d22e0c;
    ram_cell[    6929] = 32'h3b26e1d9;
    ram_cell[    6930] = 32'ha3b20766;
    ram_cell[    6931] = 32'h11adbcc3;
    ram_cell[    6932] = 32'h8697b720;
    ram_cell[    6933] = 32'h515c3ab4;
    ram_cell[    6934] = 32'h31d9fbce;
    ram_cell[    6935] = 32'h91c86c56;
    ram_cell[    6936] = 32'h08b4635a;
    ram_cell[    6937] = 32'h0d37300a;
    ram_cell[    6938] = 32'hc20de7d7;
    ram_cell[    6939] = 32'h9719d28f;
    ram_cell[    6940] = 32'hf144ee33;
    ram_cell[    6941] = 32'hb34c3aa1;
    ram_cell[    6942] = 32'hfa7e2729;
    ram_cell[    6943] = 32'hcc3431c3;
    ram_cell[    6944] = 32'hbb953115;
    ram_cell[    6945] = 32'h4dbef4ed;
    ram_cell[    6946] = 32'h1ee2ea8a;
    ram_cell[    6947] = 32'hf666b449;
    ram_cell[    6948] = 32'h6b48d12f;
    ram_cell[    6949] = 32'h29109460;
    ram_cell[    6950] = 32'hfc120a5f;
    ram_cell[    6951] = 32'hb4916530;
    ram_cell[    6952] = 32'hde66bf78;
    ram_cell[    6953] = 32'hba8bd4a5;
    ram_cell[    6954] = 32'h163a2746;
    ram_cell[    6955] = 32'hb2dcc605;
    ram_cell[    6956] = 32'h554bde20;
    ram_cell[    6957] = 32'h07c44dec;
    ram_cell[    6958] = 32'h540f9f29;
    ram_cell[    6959] = 32'h6a414065;
    ram_cell[    6960] = 32'h4542890b;
    ram_cell[    6961] = 32'h367f379c;
    ram_cell[    6962] = 32'h977903ff;
    ram_cell[    6963] = 32'h30ae4c45;
    ram_cell[    6964] = 32'h1ec80ca7;
    ram_cell[    6965] = 32'h957d4df6;
    ram_cell[    6966] = 32'hab4e817d;
    ram_cell[    6967] = 32'hb2026b60;
    ram_cell[    6968] = 32'hbbf718e5;
    ram_cell[    6969] = 32'h4ca8e986;
    ram_cell[    6970] = 32'h6810f0f7;
    ram_cell[    6971] = 32'hdfcdf00e;
    ram_cell[    6972] = 32'hd1128708;
    ram_cell[    6973] = 32'h0db59749;
    ram_cell[    6974] = 32'hc6326132;
    ram_cell[    6975] = 32'h99b0bbf9;
    ram_cell[    6976] = 32'hb9fa0066;
    ram_cell[    6977] = 32'h0770738f;
    ram_cell[    6978] = 32'h1a7fd85b;
    ram_cell[    6979] = 32'hdb2a602a;
    ram_cell[    6980] = 32'h9affd985;
    ram_cell[    6981] = 32'h9ac1ee1b;
    ram_cell[    6982] = 32'hbcfc7d6a;
    ram_cell[    6983] = 32'hb549032a;
    ram_cell[    6984] = 32'h9afd62fe;
    ram_cell[    6985] = 32'hb2ccf543;
    ram_cell[    6986] = 32'h17aea225;
    ram_cell[    6987] = 32'h4ce54d9b;
    ram_cell[    6988] = 32'h4dd38db6;
    ram_cell[    6989] = 32'ha667ce39;
    ram_cell[    6990] = 32'h71424624;
    ram_cell[    6991] = 32'h0417c664;
    ram_cell[    6992] = 32'h521cfb36;
    ram_cell[    6993] = 32'h5524ba5f;
    ram_cell[    6994] = 32'h8114869b;
    ram_cell[    6995] = 32'h0bd633d6;
    ram_cell[    6996] = 32'h97b3d408;
    ram_cell[    6997] = 32'h1e6f4cd1;
    ram_cell[    6998] = 32'h978cc485;
    ram_cell[    6999] = 32'h47bf48b2;
    ram_cell[    7000] = 32'h5601691c;
    ram_cell[    7001] = 32'h69f872a8;
    ram_cell[    7002] = 32'hf25dfa56;
    ram_cell[    7003] = 32'h962ccb9d;
    ram_cell[    7004] = 32'h20bf6b39;
    ram_cell[    7005] = 32'h4e83de38;
    ram_cell[    7006] = 32'h99bbeff5;
    ram_cell[    7007] = 32'ha6ca2ef8;
    ram_cell[    7008] = 32'h54a87a82;
    ram_cell[    7009] = 32'h1437daac;
    ram_cell[    7010] = 32'h9ec40744;
    ram_cell[    7011] = 32'h759e6cd8;
    ram_cell[    7012] = 32'h95dbdfb4;
    ram_cell[    7013] = 32'he1230389;
    ram_cell[    7014] = 32'hcb66584a;
    ram_cell[    7015] = 32'h304b563b;
    ram_cell[    7016] = 32'h76291bb3;
    ram_cell[    7017] = 32'h6c9ccea8;
    ram_cell[    7018] = 32'hfadd4ce5;
    ram_cell[    7019] = 32'h0196d6b6;
    ram_cell[    7020] = 32'h4dc6df8e;
    ram_cell[    7021] = 32'h987cd326;
    ram_cell[    7022] = 32'h517a5d65;
    ram_cell[    7023] = 32'h8c187bc3;
    ram_cell[    7024] = 32'h2dfdd50b;
    ram_cell[    7025] = 32'h4b5863f7;
    ram_cell[    7026] = 32'h80824b8c;
    ram_cell[    7027] = 32'h4a5645b9;
    ram_cell[    7028] = 32'h05626048;
    ram_cell[    7029] = 32'h897517ce;
    ram_cell[    7030] = 32'hec65a948;
    ram_cell[    7031] = 32'h0a91e8ef;
    ram_cell[    7032] = 32'hd092c639;
    ram_cell[    7033] = 32'h0c98b0a3;
    ram_cell[    7034] = 32'h0eae3f50;
    ram_cell[    7035] = 32'h00404566;
    ram_cell[    7036] = 32'h64c554b4;
    ram_cell[    7037] = 32'h4e6e4ef9;
    ram_cell[    7038] = 32'hdc34ba04;
    ram_cell[    7039] = 32'h2c74c666;
    ram_cell[    7040] = 32'hda056c55;
    ram_cell[    7041] = 32'h974ff310;
    ram_cell[    7042] = 32'h58b41490;
    ram_cell[    7043] = 32'h9b60ad10;
    ram_cell[    7044] = 32'h866a325a;
    ram_cell[    7045] = 32'h1c2d6465;
    ram_cell[    7046] = 32'hfdd573ab;
    ram_cell[    7047] = 32'hdeabb4df;
    ram_cell[    7048] = 32'hb0dac42c;
    ram_cell[    7049] = 32'hea5eb616;
    ram_cell[    7050] = 32'h1c2b3c95;
    ram_cell[    7051] = 32'h3c381c61;
    ram_cell[    7052] = 32'h6eac54f1;
    ram_cell[    7053] = 32'hb5c72509;
    ram_cell[    7054] = 32'h49fb1200;
    ram_cell[    7055] = 32'h37fb28e5;
    ram_cell[    7056] = 32'h57c3c1e4;
    ram_cell[    7057] = 32'h6ce57919;
    ram_cell[    7058] = 32'h2c769a40;
    ram_cell[    7059] = 32'hf048e2cb;
    ram_cell[    7060] = 32'h29666ab2;
    ram_cell[    7061] = 32'h05472dd1;
    ram_cell[    7062] = 32'hecdabfd1;
    ram_cell[    7063] = 32'hd951f46e;
    ram_cell[    7064] = 32'h408cb64e;
    ram_cell[    7065] = 32'h1cb7ad90;
    ram_cell[    7066] = 32'h2038bf08;
    ram_cell[    7067] = 32'h44518317;
    ram_cell[    7068] = 32'h7b2458c9;
    ram_cell[    7069] = 32'h73ac2412;
    ram_cell[    7070] = 32'h8f3a3e50;
    ram_cell[    7071] = 32'h0cfdfe67;
    ram_cell[    7072] = 32'h31a8fa55;
    ram_cell[    7073] = 32'hac93e010;
    ram_cell[    7074] = 32'hdb57aec7;
    ram_cell[    7075] = 32'hda329320;
    ram_cell[    7076] = 32'h4d78f645;
    ram_cell[    7077] = 32'hc9ac430d;
    ram_cell[    7078] = 32'h708e3394;
    ram_cell[    7079] = 32'h21b8803c;
    ram_cell[    7080] = 32'h1dfd80e6;
    ram_cell[    7081] = 32'hb942c0e3;
    ram_cell[    7082] = 32'h033dea1b;
    ram_cell[    7083] = 32'h924d8693;
    ram_cell[    7084] = 32'he7b9bcd3;
    ram_cell[    7085] = 32'h2c067c14;
    ram_cell[    7086] = 32'h04fe1066;
    ram_cell[    7087] = 32'h049b6e09;
    ram_cell[    7088] = 32'h71e4e267;
    ram_cell[    7089] = 32'h1049e999;
    ram_cell[    7090] = 32'h51bd63b0;
    ram_cell[    7091] = 32'h761d5bc2;
    ram_cell[    7092] = 32'h2dee8c2b;
    ram_cell[    7093] = 32'h3be3dd33;
    ram_cell[    7094] = 32'h74b75ad8;
    ram_cell[    7095] = 32'h8ac7fa35;
    ram_cell[    7096] = 32'he83b0acd;
    ram_cell[    7097] = 32'hf195fefd;
    ram_cell[    7098] = 32'h6e525642;
    ram_cell[    7099] = 32'h120afe55;
    ram_cell[    7100] = 32'h0b4a3833;
    ram_cell[    7101] = 32'hb7995ad1;
    ram_cell[    7102] = 32'hac7c8398;
    ram_cell[    7103] = 32'h9eb0b6e5;
    ram_cell[    7104] = 32'hfacdfde5;
    ram_cell[    7105] = 32'h67d60a94;
    ram_cell[    7106] = 32'h2e5501a8;
    ram_cell[    7107] = 32'hff4d167f;
    ram_cell[    7108] = 32'h688cbfec;
    ram_cell[    7109] = 32'hf08cfd03;
    ram_cell[    7110] = 32'ha23fc407;
    ram_cell[    7111] = 32'h2d8d0c94;
    ram_cell[    7112] = 32'ha3d5fe8c;
    ram_cell[    7113] = 32'hb9f99eab;
    ram_cell[    7114] = 32'hc645cf46;
    ram_cell[    7115] = 32'h2adadb65;
    ram_cell[    7116] = 32'h83dd0d1b;
    ram_cell[    7117] = 32'h77e5c5dc;
    ram_cell[    7118] = 32'h1fc5647f;
    ram_cell[    7119] = 32'h7b1f9b47;
    ram_cell[    7120] = 32'h4d7e4468;
    ram_cell[    7121] = 32'h222d3e4e;
    ram_cell[    7122] = 32'h4e18e13e;
    ram_cell[    7123] = 32'ha9e9baca;
    ram_cell[    7124] = 32'hf7070d40;
    ram_cell[    7125] = 32'h711b5655;
    ram_cell[    7126] = 32'h3002a07d;
    ram_cell[    7127] = 32'h06b10da3;
    ram_cell[    7128] = 32'hde0cdaa1;
    ram_cell[    7129] = 32'h4f492a76;
    ram_cell[    7130] = 32'h5c0046a8;
    ram_cell[    7131] = 32'h99d4ea5e;
    ram_cell[    7132] = 32'h98f73df5;
    ram_cell[    7133] = 32'h57dbba33;
    ram_cell[    7134] = 32'h309abc7a;
    ram_cell[    7135] = 32'hc3b43cc6;
    ram_cell[    7136] = 32'h2b7ad447;
    ram_cell[    7137] = 32'h602af3bf;
    ram_cell[    7138] = 32'h943ef146;
    ram_cell[    7139] = 32'h9023ee04;
    ram_cell[    7140] = 32'h1c83b684;
    ram_cell[    7141] = 32'h58ab29d5;
    ram_cell[    7142] = 32'hf681be7d;
    ram_cell[    7143] = 32'h18d0ce05;
    ram_cell[    7144] = 32'hdcfe4488;
    ram_cell[    7145] = 32'h52b8a4bd;
    ram_cell[    7146] = 32'h239896e9;
    ram_cell[    7147] = 32'h7d675e49;
    ram_cell[    7148] = 32'hb66b8e63;
    ram_cell[    7149] = 32'hd0c5d0e6;
    ram_cell[    7150] = 32'hc30d4f20;
    ram_cell[    7151] = 32'hf462a509;
    ram_cell[    7152] = 32'hf6fb015f;
    ram_cell[    7153] = 32'h7250120f;
    ram_cell[    7154] = 32'h9ce4866c;
    ram_cell[    7155] = 32'h14de4079;
    ram_cell[    7156] = 32'hb5f7cc2f;
    ram_cell[    7157] = 32'h9c55edfb;
    ram_cell[    7158] = 32'hc034174d;
    ram_cell[    7159] = 32'h608786b2;
    ram_cell[    7160] = 32'h2569de9a;
    ram_cell[    7161] = 32'h7e65ba48;
    ram_cell[    7162] = 32'he50c2bde;
    ram_cell[    7163] = 32'h47a08d55;
    ram_cell[    7164] = 32'hbcb65ac2;
    ram_cell[    7165] = 32'h2f970bdd;
    ram_cell[    7166] = 32'h767bebbe;
    ram_cell[    7167] = 32'h3f99ea6f;
    ram_cell[    7168] = 32'hdc0e987c;
    ram_cell[    7169] = 32'haaded663;
    ram_cell[    7170] = 32'h540862a2;
    ram_cell[    7171] = 32'h6a3b284a;
    ram_cell[    7172] = 32'h5829529c;
    ram_cell[    7173] = 32'hf80a9f0a;
    ram_cell[    7174] = 32'h8ab08add;
    ram_cell[    7175] = 32'h4e44ff3f;
    ram_cell[    7176] = 32'h8b2384ae;
    ram_cell[    7177] = 32'h86d14b4c;
    ram_cell[    7178] = 32'ha629cbe3;
    ram_cell[    7179] = 32'h758750e7;
    ram_cell[    7180] = 32'h21c013b2;
    ram_cell[    7181] = 32'h1b9903cc;
    ram_cell[    7182] = 32'h216e14bb;
    ram_cell[    7183] = 32'h362514f5;
    ram_cell[    7184] = 32'h6f307227;
    ram_cell[    7185] = 32'hc278b490;
    ram_cell[    7186] = 32'hbb73d3ef;
    ram_cell[    7187] = 32'hc4ac48f6;
    ram_cell[    7188] = 32'ha140d5b8;
    ram_cell[    7189] = 32'h35ed6d63;
    ram_cell[    7190] = 32'h9b66b189;
    ram_cell[    7191] = 32'h10472832;
    ram_cell[    7192] = 32'hbb26c0bb;
    ram_cell[    7193] = 32'h5a95798f;
    ram_cell[    7194] = 32'hd456e967;
    ram_cell[    7195] = 32'he4b34dbe;
    ram_cell[    7196] = 32'h4eb2c557;
    ram_cell[    7197] = 32'ha88ad122;
    ram_cell[    7198] = 32'h72970164;
    ram_cell[    7199] = 32'h5095a2b3;
    ram_cell[    7200] = 32'ha49d66ac;
    ram_cell[    7201] = 32'ha9675f0d;
    ram_cell[    7202] = 32'h17bd52bd;
    ram_cell[    7203] = 32'hac954c68;
    ram_cell[    7204] = 32'h64eb0be4;
    ram_cell[    7205] = 32'hc23d55e1;
    ram_cell[    7206] = 32'hdfd25364;
    ram_cell[    7207] = 32'hac6f0665;
    ram_cell[    7208] = 32'hdfefdf4f;
    ram_cell[    7209] = 32'hc8ccb50d;
    ram_cell[    7210] = 32'h1fff3d38;
    ram_cell[    7211] = 32'hb880152a;
    ram_cell[    7212] = 32'hc2110e99;
    ram_cell[    7213] = 32'hdeb05b72;
    ram_cell[    7214] = 32'ha19f0663;
    ram_cell[    7215] = 32'hde044b70;
    ram_cell[    7216] = 32'h7754e610;
    ram_cell[    7217] = 32'h2af801a7;
    ram_cell[    7218] = 32'h2d2166b6;
    ram_cell[    7219] = 32'h9ef0a9de;
    ram_cell[    7220] = 32'h2eab8708;
    ram_cell[    7221] = 32'h5060f7a2;
    ram_cell[    7222] = 32'h80875b91;
    ram_cell[    7223] = 32'h3e9c2672;
    ram_cell[    7224] = 32'hc55a7d15;
    ram_cell[    7225] = 32'hc4fb5f6a;
    ram_cell[    7226] = 32'h16f8a482;
    ram_cell[    7227] = 32'h51b8ab07;
    ram_cell[    7228] = 32'h8162e5f7;
    ram_cell[    7229] = 32'h9ff169a9;
    ram_cell[    7230] = 32'h293d45d5;
    ram_cell[    7231] = 32'hdf5d4ab9;
    ram_cell[    7232] = 32'h1e1cdd26;
    ram_cell[    7233] = 32'h6bdf1d86;
    ram_cell[    7234] = 32'hdf2a6769;
    ram_cell[    7235] = 32'h12399af7;
    ram_cell[    7236] = 32'h76c5f498;
    ram_cell[    7237] = 32'h6459bf84;
    ram_cell[    7238] = 32'h6bd735ab;
    ram_cell[    7239] = 32'h90b05177;
    ram_cell[    7240] = 32'hc0581f04;
    ram_cell[    7241] = 32'h49c01197;
    ram_cell[    7242] = 32'h0fb71894;
    ram_cell[    7243] = 32'h2c209888;
    ram_cell[    7244] = 32'hed0169b8;
    ram_cell[    7245] = 32'hf4f06949;
    ram_cell[    7246] = 32'h70a2a822;
    ram_cell[    7247] = 32'hc07b9547;
    ram_cell[    7248] = 32'h0a00bd43;
    ram_cell[    7249] = 32'hb6a8c8dd;
    ram_cell[    7250] = 32'hc2861e91;
    ram_cell[    7251] = 32'ha8e9e540;
    ram_cell[    7252] = 32'he60debff;
    ram_cell[    7253] = 32'h430352ea;
    ram_cell[    7254] = 32'h65df6dcc;
    ram_cell[    7255] = 32'h199cd133;
    ram_cell[    7256] = 32'hf4be5763;
    ram_cell[    7257] = 32'h21926612;
    ram_cell[    7258] = 32'h062e5a31;
    ram_cell[    7259] = 32'hf887acc9;
    ram_cell[    7260] = 32'hbddb3bbc;
    ram_cell[    7261] = 32'h544572d6;
    ram_cell[    7262] = 32'h9ae2a004;
    ram_cell[    7263] = 32'h89a97c4e;
    ram_cell[    7264] = 32'he7310fac;
    ram_cell[    7265] = 32'h91bc33b1;
    ram_cell[    7266] = 32'hedf27944;
    ram_cell[    7267] = 32'h051e161f;
    ram_cell[    7268] = 32'hed88a2ec;
    ram_cell[    7269] = 32'hb93bf975;
    ram_cell[    7270] = 32'h11e4aaf5;
    ram_cell[    7271] = 32'hf177c6ad;
    ram_cell[    7272] = 32'h8fe0018d;
    ram_cell[    7273] = 32'h7341c85e;
    ram_cell[    7274] = 32'h2bad6095;
    ram_cell[    7275] = 32'haf1701df;
    ram_cell[    7276] = 32'h3a3503ff;
    ram_cell[    7277] = 32'h4cec7d6b;
    ram_cell[    7278] = 32'hc92728c8;
    ram_cell[    7279] = 32'hc87c8996;
    ram_cell[    7280] = 32'he168ac97;
    ram_cell[    7281] = 32'hfd150304;
    ram_cell[    7282] = 32'h33b6abd5;
    ram_cell[    7283] = 32'h16b55b7d;
    ram_cell[    7284] = 32'haa7fedd7;
    ram_cell[    7285] = 32'h8825281f;
    ram_cell[    7286] = 32'h48e8eae0;
    ram_cell[    7287] = 32'h01f2329b;
    ram_cell[    7288] = 32'h4ecc7685;
    ram_cell[    7289] = 32'h123fc765;
    ram_cell[    7290] = 32'h19dd3797;
    ram_cell[    7291] = 32'hb393142f;
    ram_cell[    7292] = 32'hea191a39;
    ram_cell[    7293] = 32'h04f5eca7;
    ram_cell[    7294] = 32'hff2e2313;
    ram_cell[    7295] = 32'h94b1baba;
    ram_cell[    7296] = 32'he484cb93;
    ram_cell[    7297] = 32'h10bd09d9;
    ram_cell[    7298] = 32'hefd0e0d4;
    ram_cell[    7299] = 32'h49820ef7;
    ram_cell[    7300] = 32'h8b686a20;
    ram_cell[    7301] = 32'h470a60ba;
    ram_cell[    7302] = 32'h83fd9781;
    ram_cell[    7303] = 32'h42b2743b;
    ram_cell[    7304] = 32'h3dce05cd;
    ram_cell[    7305] = 32'hf63b6cfa;
    ram_cell[    7306] = 32'hb7b850a4;
    ram_cell[    7307] = 32'h21f03d34;
    ram_cell[    7308] = 32'he64bc443;
    ram_cell[    7309] = 32'hf11aa445;
    ram_cell[    7310] = 32'h3d9aa21e;
    ram_cell[    7311] = 32'h9e1bfc40;
    ram_cell[    7312] = 32'h403834c7;
    ram_cell[    7313] = 32'hd9b7437d;
    ram_cell[    7314] = 32'hca38b34b;
    ram_cell[    7315] = 32'h12bace65;
    ram_cell[    7316] = 32'h9529cbc2;
    ram_cell[    7317] = 32'hf67df1d9;
    ram_cell[    7318] = 32'h3fbc536c;
    ram_cell[    7319] = 32'h1ef034a2;
    ram_cell[    7320] = 32'h76632b40;
    ram_cell[    7321] = 32'hf4149ca5;
    ram_cell[    7322] = 32'h43b2e784;
    ram_cell[    7323] = 32'h108052c8;
    ram_cell[    7324] = 32'h08322cac;
    ram_cell[    7325] = 32'h30af519e;
    ram_cell[    7326] = 32'h9ad08565;
    ram_cell[    7327] = 32'h8bb5d05c;
    ram_cell[    7328] = 32'h68a6c37c;
    ram_cell[    7329] = 32'hb0b49de0;
    ram_cell[    7330] = 32'h6ff11aa2;
    ram_cell[    7331] = 32'hc1202f55;
    ram_cell[    7332] = 32'h178f9130;
    ram_cell[    7333] = 32'h9688b30e;
    ram_cell[    7334] = 32'h1f4ae3b4;
    ram_cell[    7335] = 32'hbdf1e0af;
    ram_cell[    7336] = 32'hc5458068;
    ram_cell[    7337] = 32'hc638a7e4;
    ram_cell[    7338] = 32'h02b79fdd;
    ram_cell[    7339] = 32'h141ce6d6;
    ram_cell[    7340] = 32'he9aa7d07;
    ram_cell[    7341] = 32'hb2a993c2;
    ram_cell[    7342] = 32'he73d1f07;
    ram_cell[    7343] = 32'h52bb8706;
    ram_cell[    7344] = 32'h2164291f;
    ram_cell[    7345] = 32'h2c85f70c;
    ram_cell[    7346] = 32'hee405014;
    ram_cell[    7347] = 32'h9a5cc376;
    ram_cell[    7348] = 32'h2cd8b654;
    ram_cell[    7349] = 32'h465a08bd;
    ram_cell[    7350] = 32'h0db9b772;
    ram_cell[    7351] = 32'h8ac2b39f;
    ram_cell[    7352] = 32'h6c0eceec;
    ram_cell[    7353] = 32'h98e182b2;
    ram_cell[    7354] = 32'hc5618372;
    ram_cell[    7355] = 32'hb5edb836;
    ram_cell[    7356] = 32'h200539c7;
    ram_cell[    7357] = 32'h2c9cae0d;
    ram_cell[    7358] = 32'ha6ea862e;
    ram_cell[    7359] = 32'h4a0bf1cf;
    ram_cell[    7360] = 32'hdb08f8ac;
    ram_cell[    7361] = 32'h2a0ea413;
    ram_cell[    7362] = 32'h85d93a5c;
    ram_cell[    7363] = 32'h63544e83;
    ram_cell[    7364] = 32'h4ced7dd1;
    ram_cell[    7365] = 32'h90b87ea6;
    ram_cell[    7366] = 32'hb0f4e68f;
    ram_cell[    7367] = 32'h9101ac51;
    ram_cell[    7368] = 32'ha3204fd7;
    ram_cell[    7369] = 32'h2b4e71cb;
    ram_cell[    7370] = 32'hfa0ea07f;
    ram_cell[    7371] = 32'h557ffd26;
    ram_cell[    7372] = 32'hf53742cc;
    ram_cell[    7373] = 32'hb91ee0ec;
    ram_cell[    7374] = 32'h5517db86;
    ram_cell[    7375] = 32'h0d6ab9af;
    ram_cell[    7376] = 32'h7506ded1;
    ram_cell[    7377] = 32'h0675a4fc;
    ram_cell[    7378] = 32'he2e182bc;
    ram_cell[    7379] = 32'h1ab3ed4b;
    ram_cell[    7380] = 32'h92d2ebee;
    ram_cell[    7381] = 32'h21c74f13;
    ram_cell[    7382] = 32'he0959a7c;
    ram_cell[    7383] = 32'hcc2a5a47;
    ram_cell[    7384] = 32'h85419d13;
    ram_cell[    7385] = 32'hcb0ac9ba;
    ram_cell[    7386] = 32'hf07c9ca7;
    ram_cell[    7387] = 32'h9e624703;
    ram_cell[    7388] = 32'h004f5c16;
    ram_cell[    7389] = 32'h2ca62e20;
    ram_cell[    7390] = 32'hcff92975;
    ram_cell[    7391] = 32'h370484d0;
    ram_cell[    7392] = 32'hf560fe0d;
    ram_cell[    7393] = 32'hd0175e99;
    ram_cell[    7394] = 32'hc261d5fc;
    ram_cell[    7395] = 32'hb3f42b9c;
    ram_cell[    7396] = 32'h50e9e785;
    ram_cell[    7397] = 32'hbbd80a4a;
    ram_cell[    7398] = 32'hc3864b35;
    ram_cell[    7399] = 32'h81b254f7;
    ram_cell[    7400] = 32'h24bc0fb4;
    ram_cell[    7401] = 32'hefa3d457;
    ram_cell[    7402] = 32'hb4d0c091;
    ram_cell[    7403] = 32'hcf03738a;
    ram_cell[    7404] = 32'h7364f59a;
    ram_cell[    7405] = 32'h2928d9a2;
    ram_cell[    7406] = 32'h991fddcc;
    ram_cell[    7407] = 32'hf4165f9b;
    ram_cell[    7408] = 32'hc55ac2e5;
    ram_cell[    7409] = 32'h4cacdbfc;
    ram_cell[    7410] = 32'h6c3e6fd2;
    ram_cell[    7411] = 32'hf701abef;
    ram_cell[    7412] = 32'he11c2c27;
    ram_cell[    7413] = 32'h70de27ae;
    ram_cell[    7414] = 32'hd6a4c894;
    ram_cell[    7415] = 32'hae85c4fe;
    ram_cell[    7416] = 32'hfb2a5c4e;
    ram_cell[    7417] = 32'h169a5f0f;
    ram_cell[    7418] = 32'h19873abd;
    ram_cell[    7419] = 32'h0453e8cd;
    ram_cell[    7420] = 32'h5fa64de8;
    ram_cell[    7421] = 32'h53472e99;
    ram_cell[    7422] = 32'hbc752f5c;
    ram_cell[    7423] = 32'h45d771f8;
    ram_cell[    7424] = 32'hf71e5705;
    ram_cell[    7425] = 32'h353641a9;
    ram_cell[    7426] = 32'h284beaff;
    ram_cell[    7427] = 32'h294b8d5e;
    ram_cell[    7428] = 32'h92c1a497;
    ram_cell[    7429] = 32'h51de7941;
    ram_cell[    7430] = 32'h133fa891;
    ram_cell[    7431] = 32'h0b85e7e2;
    ram_cell[    7432] = 32'hc9004c88;
    ram_cell[    7433] = 32'h2fcc2299;
    ram_cell[    7434] = 32'h57ebfb02;
    ram_cell[    7435] = 32'hd68d5d31;
    ram_cell[    7436] = 32'h11ed4d33;
    ram_cell[    7437] = 32'hd476afab;
    ram_cell[    7438] = 32'h7bbc77e1;
    ram_cell[    7439] = 32'h0cb3aeff;
    ram_cell[    7440] = 32'h2160df56;
    ram_cell[    7441] = 32'h7e340b9e;
    ram_cell[    7442] = 32'hebf22b51;
    ram_cell[    7443] = 32'h139c9cf2;
    ram_cell[    7444] = 32'h9fb47f4a;
    ram_cell[    7445] = 32'hcb42fc97;
    ram_cell[    7446] = 32'h28ea307f;
    ram_cell[    7447] = 32'ha124ce5f;
    ram_cell[    7448] = 32'h157287ce;
    ram_cell[    7449] = 32'hff0498b1;
    ram_cell[    7450] = 32'hae237020;
    ram_cell[    7451] = 32'hfab37edf;
    ram_cell[    7452] = 32'h8e911914;
    ram_cell[    7453] = 32'h8679658e;
    ram_cell[    7454] = 32'h862e75e0;
    ram_cell[    7455] = 32'h1e7b0fd8;
    ram_cell[    7456] = 32'h02607345;
    ram_cell[    7457] = 32'h2b3f7cc9;
    ram_cell[    7458] = 32'h8be1ee2e;
    ram_cell[    7459] = 32'h317823ed;
    ram_cell[    7460] = 32'haa0fb31d;
    ram_cell[    7461] = 32'hddedc611;
    ram_cell[    7462] = 32'h2b2bebee;
    ram_cell[    7463] = 32'h364bb37a;
    ram_cell[    7464] = 32'hf4f1b4b5;
    ram_cell[    7465] = 32'h6798ebc8;
    ram_cell[    7466] = 32'h74d4702a;
    ram_cell[    7467] = 32'h9b3cfa77;
    ram_cell[    7468] = 32'h1a01f665;
    ram_cell[    7469] = 32'h4f7078f0;
    ram_cell[    7470] = 32'h64d568b1;
    ram_cell[    7471] = 32'h772c5883;
    ram_cell[    7472] = 32'hecff1eab;
    ram_cell[    7473] = 32'h9525602e;
    ram_cell[    7474] = 32'h85bbbbad;
    ram_cell[    7475] = 32'hb73be7f7;
    ram_cell[    7476] = 32'hab81d9da;
    ram_cell[    7477] = 32'h33551c86;
    ram_cell[    7478] = 32'h67bed366;
    ram_cell[    7479] = 32'h05edf894;
    ram_cell[    7480] = 32'he235622c;
    ram_cell[    7481] = 32'h1e85d807;
    ram_cell[    7482] = 32'h169b8eee;
    ram_cell[    7483] = 32'haf189b28;
    ram_cell[    7484] = 32'hf1780ab3;
    ram_cell[    7485] = 32'h9997df3b;
    ram_cell[    7486] = 32'hcce2048a;
    ram_cell[    7487] = 32'h1453f4d5;
    ram_cell[    7488] = 32'h00c1b24a;
    ram_cell[    7489] = 32'h81c4bde6;
    ram_cell[    7490] = 32'h3c4cc424;
    ram_cell[    7491] = 32'hbb64e44f;
    ram_cell[    7492] = 32'h036f4482;
    ram_cell[    7493] = 32'h180f9b84;
    ram_cell[    7494] = 32'h8111ce07;
    ram_cell[    7495] = 32'h21bd42e1;
    ram_cell[    7496] = 32'h481b7590;
    ram_cell[    7497] = 32'h2ee60135;
    ram_cell[    7498] = 32'ha57d59ae;
    ram_cell[    7499] = 32'hd4f9dbcc;
    ram_cell[    7500] = 32'h4d42fbb9;
    ram_cell[    7501] = 32'h6dd417d5;
    ram_cell[    7502] = 32'h8b69f7c7;
    ram_cell[    7503] = 32'he5f028d4;
    ram_cell[    7504] = 32'h9c9aa33d;
    ram_cell[    7505] = 32'hf7747417;
    ram_cell[    7506] = 32'haa03d795;
    ram_cell[    7507] = 32'he13823e3;
    ram_cell[    7508] = 32'h5af05089;
    ram_cell[    7509] = 32'he5d3e14b;
    ram_cell[    7510] = 32'h146028ee;
    ram_cell[    7511] = 32'haf8cc5a7;
    ram_cell[    7512] = 32'hb273104c;
    ram_cell[    7513] = 32'h65910cf1;
    ram_cell[    7514] = 32'hc5955c02;
    ram_cell[    7515] = 32'h8314484d;
    ram_cell[    7516] = 32'h3868ba2a;
    ram_cell[    7517] = 32'h4288d16a;
    ram_cell[    7518] = 32'hd57699e3;
    ram_cell[    7519] = 32'h4652b518;
    ram_cell[    7520] = 32'h33c7d6b6;
    ram_cell[    7521] = 32'h107ef983;
    ram_cell[    7522] = 32'hf3646ebd;
    ram_cell[    7523] = 32'hf2704536;
    ram_cell[    7524] = 32'h3cc9f75d;
    ram_cell[    7525] = 32'h12e90629;
    ram_cell[    7526] = 32'hdc0dc485;
    ram_cell[    7527] = 32'h231b7785;
    ram_cell[    7528] = 32'h170aa62d;
    ram_cell[    7529] = 32'he2bf1be0;
    ram_cell[    7530] = 32'hb4d7a861;
    ram_cell[    7531] = 32'h75365138;
    ram_cell[    7532] = 32'h28a2c446;
    ram_cell[    7533] = 32'h6d220681;
    ram_cell[    7534] = 32'h9f806f5d;
    ram_cell[    7535] = 32'hbb08fa59;
    ram_cell[    7536] = 32'h2af8bedb;
    ram_cell[    7537] = 32'h2f330eb8;
    ram_cell[    7538] = 32'h288e1b60;
    ram_cell[    7539] = 32'h19df1226;
    ram_cell[    7540] = 32'hb1d341d5;
    ram_cell[    7541] = 32'h35835e82;
    ram_cell[    7542] = 32'h6ca1acf0;
    ram_cell[    7543] = 32'h8d97d211;
    ram_cell[    7544] = 32'h06b7191a;
    ram_cell[    7545] = 32'hac04aabf;
    ram_cell[    7546] = 32'h331df86f;
    ram_cell[    7547] = 32'h0e049e02;
    ram_cell[    7548] = 32'h8a36d0ef;
    ram_cell[    7549] = 32'hc4e2579d;
    ram_cell[    7550] = 32'h5f6c59fd;
    ram_cell[    7551] = 32'h8187a764;
    ram_cell[    7552] = 32'h526e73f1;
    ram_cell[    7553] = 32'hbc28f32a;
    ram_cell[    7554] = 32'h6db667e9;
    ram_cell[    7555] = 32'h74009e61;
    ram_cell[    7556] = 32'h491f004c;
    ram_cell[    7557] = 32'h0c423d9b;
    ram_cell[    7558] = 32'hce8b2a06;
    ram_cell[    7559] = 32'h3506b1e4;
    ram_cell[    7560] = 32'he4600c60;
    ram_cell[    7561] = 32'h3e38d9d6;
    ram_cell[    7562] = 32'h51711279;
    ram_cell[    7563] = 32'h6232ad92;
    ram_cell[    7564] = 32'hb5879652;
    ram_cell[    7565] = 32'hd7978ae2;
    ram_cell[    7566] = 32'h7d9d674e;
    ram_cell[    7567] = 32'hb5c2ce4c;
    ram_cell[    7568] = 32'h3be44295;
    ram_cell[    7569] = 32'h3e28ee25;
    ram_cell[    7570] = 32'h0719805d;
    ram_cell[    7571] = 32'h70ae56b7;
    ram_cell[    7572] = 32'h8162c470;
    ram_cell[    7573] = 32'hc7d1b76f;
    ram_cell[    7574] = 32'hef805a76;
    ram_cell[    7575] = 32'hb129edb6;
    ram_cell[    7576] = 32'h7bc01074;
    ram_cell[    7577] = 32'h682ded68;
    ram_cell[    7578] = 32'haed73cba;
    ram_cell[    7579] = 32'h4c2a0412;
    ram_cell[    7580] = 32'h7c08d54b;
    ram_cell[    7581] = 32'h57847e75;
    ram_cell[    7582] = 32'hd3ca6b91;
    ram_cell[    7583] = 32'h76de13fb;
    ram_cell[    7584] = 32'h30b6496b;
    ram_cell[    7585] = 32'he359ea35;
    ram_cell[    7586] = 32'ha96e1d4a;
    ram_cell[    7587] = 32'hf272620b;
    ram_cell[    7588] = 32'h6ec19b07;
    ram_cell[    7589] = 32'hbda6a2cb;
    ram_cell[    7590] = 32'h0e6d3a71;
    ram_cell[    7591] = 32'h527823c5;
    ram_cell[    7592] = 32'hd493a811;
    ram_cell[    7593] = 32'h7530fcf8;
    ram_cell[    7594] = 32'h4890ad76;
    ram_cell[    7595] = 32'h3ae3eba8;
    ram_cell[    7596] = 32'h7ba7a9c4;
    ram_cell[    7597] = 32'ha9eb9f94;
    ram_cell[    7598] = 32'h3ae633e7;
    ram_cell[    7599] = 32'hc4f32ee8;
    ram_cell[    7600] = 32'h30a0ae0c;
    ram_cell[    7601] = 32'hefa81828;
    ram_cell[    7602] = 32'hde779544;
    ram_cell[    7603] = 32'hd6b11c8d;
    ram_cell[    7604] = 32'h3b212606;
    ram_cell[    7605] = 32'h0bcb6a52;
    ram_cell[    7606] = 32'h7f94a76f;
    ram_cell[    7607] = 32'hfce7eccc;
    ram_cell[    7608] = 32'hd9ea50dc;
    ram_cell[    7609] = 32'hcb78bcc3;
    ram_cell[    7610] = 32'hfb17138d;
    ram_cell[    7611] = 32'h3f85d974;
    ram_cell[    7612] = 32'h371c76b1;
    ram_cell[    7613] = 32'h93f79739;
    ram_cell[    7614] = 32'h8d37b006;
    ram_cell[    7615] = 32'he45230ff;
    ram_cell[    7616] = 32'h75fc4326;
    ram_cell[    7617] = 32'h7a4ad0f0;
    ram_cell[    7618] = 32'h4c28d27c;
    ram_cell[    7619] = 32'hf8d8f4f1;
    ram_cell[    7620] = 32'he8982982;
    ram_cell[    7621] = 32'h33f94694;
    ram_cell[    7622] = 32'h731d7066;
    ram_cell[    7623] = 32'h8fcdaa0a;
    ram_cell[    7624] = 32'hce97cd9f;
    ram_cell[    7625] = 32'hb40866c6;
    ram_cell[    7626] = 32'h40d76de8;
    ram_cell[    7627] = 32'h9b94c6eb;
    ram_cell[    7628] = 32'h70553914;
    ram_cell[    7629] = 32'hcaa1b3e0;
    ram_cell[    7630] = 32'h36850432;
    ram_cell[    7631] = 32'h7621019f;
    ram_cell[    7632] = 32'ha718976f;
    ram_cell[    7633] = 32'h3a619310;
    ram_cell[    7634] = 32'hffc6a44c;
    ram_cell[    7635] = 32'h5c6508ec;
    ram_cell[    7636] = 32'h6a0c7869;
    ram_cell[    7637] = 32'h5d581fa6;
    ram_cell[    7638] = 32'hf352b1a9;
    ram_cell[    7639] = 32'hadedce70;
    ram_cell[    7640] = 32'h8aa35e21;
    ram_cell[    7641] = 32'h10e973d7;
    ram_cell[    7642] = 32'h5b33cb1b;
    ram_cell[    7643] = 32'h69686ab6;
    ram_cell[    7644] = 32'h95e38e43;
    ram_cell[    7645] = 32'ha41b7e89;
    ram_cell[    7646] = 32'hcc1ff9a1;
    ram_cell[    7647] = 32'h6826da90;
    ram_cell[    7648] = 32'hf90aab5c;
    ram_cell[    7649] = 32'habdf5e2a;
    ram_cell[    7650] = 32'hdddb4740;
    ram_cell[    7651] = 32'h2126c869;
    ram_cell[    7652] = 32'hfb572b1b;
    ram_cell[    7653] = 32'had5b46e6;
    ram_cell[    7654] = 32'h1f04f609;
    ram_cell[    7655] = 32'h96fcfb3c;
    ram_cell[    7656] = 32'hf59db185;
    ram_cell[    7657] = 32'hbbce30d8;
    ram_cell[    7658] = 32'h8ed24509;
    ram_cell[    7659] = 32'h527a4cfb;
    ram_cell[    7660] = 32'hd7ba8231;
    ram_cell[    7661] = 32'h3a18720b;
    ram_cell[    7662] = 32'h96e33bc3;
    ram_cell[    7663] = 32'ha5d66835;
    ram_cell[    7664] = 32'hf1302e47;
    ram_cell[    7665] = 32'hdcb8d647;
    ram_cell[    7666] = 32'h7e19bc0c;
    ram_cell[    7667] = 32'h0463f870;
    ram_cell[    7668] = 32'hbdbc2c15;
    ram_cell[    7669] = 32'ha46b00ed;
    ram_cell[    7670] = 32'hd0507dd9;
    ram_cell[    7671] = 32'h1192eb3e;
    ram_cell[    7672] = 32'hb72b8f75;
    ram_cell[    7673] = 32'h7b3d062c;
    ram_cell[    7674] = 32'h1f31a0c1;
    ram_cell[    7675] = 32'h8c47f6c3;
    ram_cell[    7676] = 32'he91e880b;
    ram_cell[    7677] = 32'hd63084ad;
    ram_cell[    7678] = 32'hd8b1f6f7;
    ram_cell[    7679] = 32'h0b060a2c;
    ram_cell[    7680] = 32'hb04f0c7d;
    ram_cell[    7681] = 32'h5c57017f;
    ram_cell[    7682] = 32'hb7faec68;
    ram_cell[    7683] = 32'h04d075f8;
    ram_cell[    7684] = 32'h7fcf7e63;
    ram_cell[    7685] = 32'he3fa9c9d;
    ram_cell[    7686] = 32'h52c65915;
    ram_cell[    7687] = 32'hd6e30b90;
    ram_cell[    7688] = 32'hb99b371a;
    ram_cell[    7689] = 32'h24517ee5;
    ram_cell[    7690] = 32'h60e1bdf0;
    ram_cell[    7691] = 32'h0af8c107;
    ram_cell[    7692] = 32'h289b16e6;
    ram_cell[    7693] = 32'ha46369f7;
    ram_cell[    7694] = 32'h28e51626;
    ram_cell[    7695] = 32'h4b96be18;
    ram_cell[    7696] = 32'h7d57a6aa;
    ram_cell[    7697] = 32'hd079a5ff;
    ram_cell[    7698] = 32'h9d6e977f;
    ram_cell[    7699] = 32'ha312a06d;
    ram_cell[    7700] = 32'hc4d41a7b;
    ram_cell[    7701] = 32'hec7a6834;
    ram_cell[    7702] = 32'hc59b1b24;
    ram_cell[    7703] = 32'h404c2472;
    ram_cell[    7704] = 32'h3701d98a;
    ram_cell[    7705] = 32'h57cbd848;
    ram_cell[    7706] = 32'h994e45e3;
    ram_cell[    7707] = 32'h317eb7e3;
    ram_cell[    7708] = 32'h418c941b;
    ram_cell[    7709] = 32'ha4bc35ea;
    ram_cell[    7710] = 32'h616a1f4e;
    ram_cell[    7711] = 32'h44e77432;
    ram_cell[    7712] = 32'h5efd9ec3;
    ram_cell[    7713] = 32'h09364fbe;
    ram_cell[    7714] = 32'hfb1a9eaa;
    ram_cell[    7715] = 32'h4bf1e076;
    ram_cell[    7716] = 32'h4e97681c;
    ram_cell[    7717] = 32'h663161f9;
    ram_cell[    7718] = 32'h823b61e8;
    ram_cell[    7719] = 32'h5cbb7647;
    ram_cell[    7720] = 32'h38643be1;
    ram_cell[    7721] = 32'hb85f6939;
    ram_cell[    7722] = 32'h60fc27f6;
    ram_cell[    7723] = 32'h07f04f2b;
    ram_cell[    7724] = 32'hc4f4c8f6;
    ram_cell[    7725] = 32'h55e6e7ba;
    ram_cell[    7726] = 32'h59feeadb;
    ram_cell[    7727] = 32'hf3f24e04;
    ram_cell[    7728] = 32'he3926be8;
    ram_cell[    7729] = 32'he865a899;
    ram_cell[    7730] = 32'h2c83b70a;
    ram_cell[    7731] = 32'h410e56fe;
    ram_cell[    7732] = 32'hc3debf91;
    ram_cell[    7733] = 32'h6f8567d8;
    ram_cell[    7734] = 32'h9bc018ff;
    ram_cell[    7735] = 32'h4f04eabd;
    ram_cell[    7736] = 32'h21c1ea45;
    ram_cell[    7737] = 32'hc5739f66;
    ram_cell[    7738] = 32'hfb639cbe;
    ram_cell[    7739] = 32'h4d8352a5;
    ram_cell[    7740] = 32'h2b2458d9;
    ram_cell[    7741] = 32'h9f3b9d41;
    ram_cell[    7742] = 32'hf700e0f3;
    ram_cell[    7743] = 32'hc3c317c1;
    ram_cell[    7744] = 32'h10298f68;
    ram_cell[    7745] = 32'h1d694ac0;
    ram_cell[    7746] = 32'h392134a5;
    ram_cell[    7747] = 32'hdd4d4541;
    ram_cell[    7748] = 32'h2b4ebf5d;
    ram_cell[    7749] = 32'h05f22e66;
    ram_cell[    7750] = 32'h192791ea;
    ram_cell[    7751] = 32'had399993;
    ram_cell[    7752] = 32'hb5516c05;
    ram_cell[    7753] = 32'h96d9d920;
    ram_cell[    7754] = 32'h314fd2e6;
    ram_cell[    7755] = 32'h95fd8dc7;
    ram_cell[    7756] = 32'ha7469166;
    ram_cell[    7757] = 32'h0f7b5175;
    ram_cell[    7758] = 32'heb0d7130;
    ram_cell[    7759] = 32'h1536283d;
    ram_cell[    7760] = 32'hd00cfd78;
    ram_cell[    7761] = 32'hdc735b52;
    ram_cell[    7762] = 32'ha034e55e;
    ram_cell[    7763] = 32'h3f6e5f28;
    ram_cell[    7764] = 32'h9da60e95;
    ram_cell[    7765] = 32'h2b78a400;
    ram_cell[    7766] = 32'h1d4f51c4;
    ram_cell[    7767] = 32'hf56c5608;
    ram_cell[    7768] = 32'hb76b4b38;
    ram_cell[    7769] = 32'h319d191e;
    ram_cell[    7770] = 32'h8ba2cb42;
    ram_cell[    7771] = 32'hf397462f;
    ram_cell[    7772] = 32'hae45f8d4;
    ram_cell[    7773] = 32'h4866f340;
    ram_cell[    7774] = 32'h7a1a2aab;
    ram_cell[    7775] = 32'h1fc45e3b;
    ram_cell[    7776] = 32'ha06fc16f;
    ram_cell[    7777] = 32'h47b6fac7;
    ram_cell[    7778] = 32'hbd5a9d93;
    ram_cell[    7779] = 32'h09a2a425;
    ram_cell[    7780] = 32'h0f988e28;
    ram_cell[    7781] = 32'hf61c17c1;
    ram_cell[    7782] = 32'hd3778549;
    ram_cell[    7783] = 32'h679d83e0;
    ram_cell[    7784] = 32'h3818b95d;
    ram_cell[    7785] = 32'h6ca35e01;
    ram_cell[    7786] = 32'h0f9be021;
    ram_cell[    7787] = 32'h22a87d45;
    ram_cell[    7788] = 32'hadaf39c2;
    ram_cell[    7789] = 32'h7bca118e;
    ram_cell[    7790] = 32'h6f96da88;
    ram_cell[    7791] = 32'haceaa2d4;
    ram_cell[    7792] = 32'hc5c92a55;
    ram_cell[    7793] = 32'h0932cd80;
    ram_cell[    7794] = 32'h45deee18;
    ram_cell[    7795] = 32'h13412b49;
    ram_cell[    7796] = 32'hca46227d;
    ram_cell[    7797] = 32'he8d3481b;
    ram_cell[    7798] = 32'h0074a9ba;
    ram_cell[    7799] = 32'h89963e14;
    ram_cell[    7800] = 32'he7664d39;
    ram_cell[    7801] = 32'h8c06e963;
    ram_cell[    7802] = 32'hd1a80527;
    ram_cell[    7803] = 32'h2f36ca54;
    ram_cell[    7804] = 32'he3965c1d;
    ram_cell[    7805] = 32'h1ddb33af;
    ram_cell[    7806] = 32'hc89b715d;
    ram_cell[    7807] = 32'hb329af0a;
    ram_cell[    7808] = 32'h8fcdbd1f;
    ram_cell[    7809] = 32'h09fb5e7d;
    ram_cell[    7810] = 32'hf688fd1e;
    ram_cell[    7811] = 32'h7f2cf878;
    ram_cell[    7812] = 32'h5b598a8f;
    ram_cell[    7813] = 32'ha6f4ebb5;
    ram_cell[    7814] = 32'h4198cb54;
    ram_cell[    7815] = 32'he6fd0981;
    ram_cell[    7816] = 32'h4573aa3e;
    ram_cell[    7817] = 32'hd6cbafac;
    ram_cell[    7818] = 32'hecaf7d83;
    ram_cell[    7819] = 32'h15d8f522;
    ram_cell[    7820] = 32'h2301a9d6;
    ram_cell[    7821] = 32'h39c69293;
    ram_cell[    7822] = 32'h313eacbb;
    ram_cell[    7823] = 32'h90bbf184;
    ram_cell[    7824] = 32'h23bc82b8;
    ram_cell[    7825] = 32'hbd68aea1;
    ram_cell[    7826] = 32'h2a2f7cde;
    ram_cell[    7827] = 32'hc278e986;
    ram_cell[    7828] = 32'h66c80fa2;
    ram_cell[    7829] = 32'h4285a48d;
    ram_cell[    7830] = 32'hdcfb98ed;
    ram_cell[    7831] = 32'hddf2c090;
    ram_cell[    7832] = 32'h51aa808a;
    ram_cell[    7833] = 32'ha1c68d54;
    ram_cell[    7834] = 32'hf712fee1;
    ram_cell[    7835] = 32'hb0280d6c;
    ram_cell[    7836] = 32'haf09bea3;
    ram_cell[    7837] = 32'h60987581;
    ram_cell[    7838] = 32'hecf66fa3;
    ram_cell[    7839] = 32'hc51a60c3;
    ram_cell[    7840] = 32'hbd55e748;
    ram_cell[    7841] = 32'h6c5f9321;
    ram_cell[    7842] = 32'h11fc1871;
    ram_cell[    7843] = 32'hf452fec2;
    ram_cell[    7844] = 32'h4474d9f7;
    ram_cell[    7845] = 32'h6655d066;
    ram_cell[    7846] = 32'h09357821;
    ram_cell[    7847] = 32'ha40a6aeb;
    ram_cell[    7848] = 32'h7155e83d;
    ram_cell[    7849] = 32'heddb65b2;
    ram_cell[    7850] = 32'hde105844;
    ram_cell[    7851] = 32'hb0f36c93;
    ram_cell[    7852] = 32'hdf5160d2;
    ram_cell[    7853] = 32'h9f96bf04;
    ram_cell[    7854] = 32'h5de8445d;
    ram_cell[    7855] = 32'hc74b1192;
    ram_cell[    7856] = 32'hcfeed935;
    ram_cell[    7857] = 32'h9a1d1ed9;
    ram_cell[    7858] = 32'hff2134b4;
    ram_cell[    7859] = 32'h2d02a76e;
    ram_cell[    7860] = 32'h84eed0ff;
    ram_cell[    7861] = 32'h94041498;
    ram_cell[    7862] = 32'hb251ba9d;
    ram_cell[    7863] = 32'h09fa599f;
    ram_cell[    7864] = 32'h8dd952d0;
    ram_cell[    7865] = 32'ha3d95f26;
    ram_cell[    7866] = 32'hff347737;
    ram_cell[    7867] = 32'h65f49670;
    ram_cell[    7868] = 32'h5987c304;
    ram_cell[    7869] = 32'he21c39bd;
    ram_cell[    7870] = 32'hfa539689;
    ram_cell[    7871] = 32'ha8bd7ce2;
    ram_cell[    7872] = 32'hf7f3dbf0;
    ram_cell[    7873] = 32'hc245e519;
    ram_cell[    7874] = 32'h0e946b54;
    ram_cell[    7875] = 32'h45b20427;
    ram_cell[    7876] = 32'h9eddf3c7;
    ram_cell[    7877] = 32'h47739357;
    ram_cell[    7878] = 32'haad6551b;
    ram_cell[    7879] = 32'h1fbed466;
    ram_cell[    7880] = 32'h03c37fe9;
    ram_cell[    7881] = 32'ha0bd8b7e;
    ram_cell[    7882] = 32'h6e611b8d;
    ram_cell[    7883] = 32'h353cc19b;
    ram_cell[    7884] = 32'h6bd000ed;
    ram_cell[    7885] = 32'h12b60d7a;
    ram_cell[    7886] = 32'hce01786c;
    ram_cell[    7887] = 32'hfefad19a;
    ram_cell[    7888] = 32'h7ec507b3;
    ram_cell[    7889] = 32'h2074c333;
    ram_cell[    7890] = 32'h5078a088;
    ram_cell[    7891] = 32'h071a2115;
    ram_cell[    7892] = 32'h7b39056d;
    ram_cell[    7893] = 32'h727c9871;
    ram_cell[    7894] = 32'h7298d5c0;
    ram_cell[    7895] = 32'ha5078c65;
    ram_cell[    7896] = 32'h4aa7e9ba;
    ram_cell[    7897] = 32'h410b73a8;
    ram_cell[    7898] = 32'h94287ac3;
    ram_cell[    7899] = 32'hb5bd793b;
    ram_cell[    7900] = 32'h9254884f;
    ram_cell[    7901] = 32'h63f10e49;
    ram_cell[    7902] = 32'he71e3111;
    ram_cell[    7903] = 32'h7f8d748b;
    ram_cell[    7904] = 32'h526f8341;
    ram_cell[    7905] = 32'h8cb6c6aa;
    ram_cell[    7906] = 32'h8e17b795;
    ram_cell[    7907] = 32'ha512ae41;
    ram_cell[    7908] = 32'h577f872e;
    ram_cell[    7909] = 32'h75b9f6f9;
    ram_cell[    7910] = 32'h64a042f1;
    ram_cell[    7911] = 32'he038c665;
    ram_cell[    7912] = 32'hdb139ec3;
    ram_cell[    7913] = 32'h5b91e812;
    ram_cell[    7914] = 32'h63ce21dc;
    ram_cell[    7915] = 32'h4a92ef93;
    ram_cell[    7916] = 32'h67a7a4ec;
    ram_cell[    7917] = 32'haf854005;
    ram_cell[    7918] = 32'h59a8d239;
    ram_cell[    7919] = 32'hb34225e7;
    ram_cell[    7920] = 32'h917d008f;
    ram_cell[    7921] = 32'h231ed4b4;
    ram_cell[    7922] = 32'h98d31186;
    ram_cell[    7923] = 32'h0442a4f9;
    ram_cell[    7924] = 32'hf32de4f9;
    ram_cell[    7925] = 32'h26b8387a;
    ram_cell[    7926] = 32'h99b3aa99;
    ram_cell[    7927] = 32'hdee6c24c;
    ram_cell[    7928] = 32'h996d21c2;
    ram_cell[    7929] = 32'hc0c91f65;
    ram_cell[    7930] = 32'h92132a7d;
    ram_cell[    7931] = 32'hebcba37d;
    ram_cell[    7932] = 32'h796ee7c2;
    ram_cell[    7933] = 32'ha86e853e;
    ram_cell[    7934] = 32'h0979b48a;
    ram_cell[    7935] = 32'hf4a45324;
    ram_cell[    7936] = 32'h5ede4804;
    ram_cell[    7937] = 32'h5c52b46b;
    ram_cell[    7938] = 32'h8d74559a;
    ram_cell[    7939] = 32'hdc15154d;
    ram_cell[    7940] = 32'hb6bb15f1;
    ram_cell[    7941] = 32'h24331cef;
    ram_cell[    7942] = 32'h71839c43;
    ram_cell[    7943] = 32'hd0dc7635;
    ram_cell[    7944] = 32'hb12b1fe1;
    ram_cell[    7945] = 32'hcdff25bc;
    ram_cell[    7946] = 32'h14d822c2;
    ram_cell[    7947] = 32'h7d09a555;
    ram_cell[    7948] = 32'h6389599d;
    ram_cell[    7949] = 32'h9091160f;
    ram_cell[    7950] = 32'h7276928f;
    ram_cell[    7951] = 32'hf706408a;
    ram_cell[    7952] = 32'h912903f5;
    ram_cell[    7953] = 32'hf7f61362;
    ram_cell[    7954] = 32'h855b037b;
    ram_cell[    7955] = 32'h89e4b889;
    ram_cell[    7956] = 32'habe8bd3c;
    ram_cell[    7957] = 32'hfabcb9ad;
    ram_cell[    7958] = 32'h891bd481;
    ram_cell[    7959] = 32'h3f4aa1e9;
    ram_cell[    7960] = 32'h5f4e6883;
    ram_cell[    7961] = 32'h077537bb;
    ram_cell[    7962] = 32'he3d0dfb8;
    ram_cell[    7963] = 32'hbfd2dd60;
    ram_cell[    7964] = 32'h3e0425b3;
    ram_cell[    7965] = 32'hf8a8bbd7;
    ram_cell[    7966] = 32'hcab2236b;
    ram_cell[    7967] = 32'hd06f42c9;
    ram_cell[    7968] = 32'h7c59db8e;
    ram_cell[    7969] = 32'h6d21b35f;
    ram_cell[    7970] = 32'h382a03e4;
    ram_cell[    7971] = 32'h71166083;
    ram_cell[    7972] = 32'h01468096;
    ram_cell[    7973] = 32'h6e5415bd;
    ram_cell[    7974] = 32'h7249bee0;
    ram_cell[    7975] = 32'hb95721e5;
    ram_cell[    7976] = 32'hbfdf9166;
    ram_cell[    7977] = 32'h0c1bee72;
    ram_cell[    7978] = 32'h65b2d70e;
    ram_cell[    7979] = 32'h40a138be;
    ram_cell[    7980] = 32'he5938aa3;
    ram_cell[    7981] = 32'h5b8f2206;
    ram_cell[    7982] = 32'h52f55733;
    ram_cell[    7983] = 32'hd7d207f6;
    ram_cell[    7984] = 32'h9e3cf115;
    ram_cell[    7985] = 32'hb8406251;
    ram_cell[    7986] = 32'h75d2e1ba;
    ram_cell[    7987] = 32'h5f6ff0bd;
    ram_cell[    7988] = 32'h701a1583;
    ram_cell[    7989] = 32'h9c78f88a;
    ram_cell[    7990] = 32'h942d0e28;
    ram_cell[    7991] = 32'hbb32959b;
    ram_cell[    7992] = 32'h8fe77edd;
    ram_cell[    7993] = 32'h81abcf07;
    ram_cell[    7994] = 32'hc0ee6ee4;
    ram_cell[    7995] = 32'h5e2f5097;
    ram_cell[    7996] = 32'h331d1576;
    ram_cell[    7997] = 32'h8de8b83e;
    ram_cell[    7998] = 32'hce5bfcb3;
    ram_cell[    7999] = 32'hc0a43b41;
    ram_cell[    8000] = 32'hdfeb81c5;
    ram_cell[    8001] = 32'ha9f52725;
    ram_cell[    8002] = 32'h82899956;
    ram_cell[    8003] = 32'h11f938c1;
    ram_cell[    8004] = 32'hb828881e;
    ram_cell[    8005] = 32'h88b130a8;
    ram_cell[    8006] = 32'h51adc3cd;
    ram_cell[    8007] = 32'h75146ece;
    ram_cell[    8008] = 32'ha4b588cb;
    ram_cell[    8009] = 32'h6b3359fd;
    ram_cell[    8010] = 32'h47604b9f;
    ram_cell[    8011] = 32'h023410f3;
    ram_cell[    8012] = 32'ha4807d5b;
    ram_cell[    8013] = 32'h78e4617c;
    ram_cell[    8014] = 32'he7f504cb;
    ram_cell[    8015] = 32'h5249ba94;
    ram_cell[    8016] = 32'h6142a9c7;
    ram_cell[    8017] = 32'ha85e4422;
    ram_cell[    8018] = 32'h91d32c41;
    ram_cell[    8019] = 32'h85274c5a;
    ram_cell[    8020] = 32'hf0faf7e5;
    ram_cell[    8021] = 32'hcf87d04b;
    ram_cell[    8022] = 32'h1447bfe8;
    ram_cell[    8023] = 32'h9fc06f31;
    ram_cell[    8024] = 32'h71a3556d;
    ram_cell[    8025] = 32'h24799bdf;
    ram_cell[    8026] = 32'h3afbb530;
    ram_cell[    8027] = 32'h0bf5753b;
    ram_cell[    8028] = 32'hce6e92ed;
    ram_cell[    8029] = 32'he8c6301a;
    ram_cell[    8030] = 32'h060838f2;
    ram_cell[    8031] = 32'h60b6ed94;
    ram_cell[    8032] = 32'ha13b52b5;
    ram_cell[    8033] = 32'h7200f896;
    ram_cell[    8034] = 32'h0e7307bb;
    ram_cell[    8035] = 32'h42d9f8ce;
    ram_cell[    8036] = 32'h00e0763b;
    ram_cell[    8037] = 32'h7c78766b;
    ram_cell[    8038] = 32'h3a031654;
    ram_cell[    8039] = 32'haedca5f1;
    ram_cell[    8040] = 32'hd1407ba5;
    ram_cell[    8041] = 32'h7cf532ee;
    ram_cell[    8042] = 32'h371f4acc;
    ram_cell[    8043] = 32'h6ea5a54c;
    ram_cell[    8044] = 32'h1d438781;
    ram_cell[    8045] = 32'hafb38a49;
    ram_cell[    8046] = 32'he5ae678d;
    ram_cell[    8047] = 32'h158d5a85;
    ram_cell[    8048] = 32'hfe62ceaf;
    ram_cell[    8049] = 32'he233d655;
    ram_cell[    8050] = 32'h15d22122;
    ram_cell[    8051] = 32'hc70e8d04;
    ram_cell[    8052] = 32'h3fb61e4c;
    ram_cell[    8053] = 32'h3ab1cff6;
    ram_cell[    8054] = 32'ha62e6e2b;
    ram_cell[    8055] = 32'ha8bcfe91;
    ram_cell[    8056] = 32'h755c3f12;
    ram_cell[    8057] = 32'h4e1c1a72;
    ram_cell[    8058] = 32'h22ef2f19;
    ram_cell[    8059] = 32'hc7a22404;
    ram_cell[    8060] = 32'h825120e7;
    ram_cell[    8061] = 32'h8c805e1e;
    ram_cell[    8062] = 32'h60b182e4;
    ram_cell[    8063] = 32'h078d8fdb;
    ram_cell[    8064] = 32'hf9490fea;
    ram_cell[    8065] = 32'hd72bc262;
    ram_cell[    8066] = 32'he8624d75;
    ram_cell[    8067] = 32'h743b76f9;
    ram_cell[    8068] = 32'haea3900f;
    ram_cell[    8069] = 32'ha7b5444d;
    ram_cell[    8070] = 32'hc66df259;
    ram_cell[    8071] = 32'hc25ca2cd;
    ram_cell[    8072] = 32'hba05196c;
    ram_cell[    8073] = 32'h0f3ac521;
    ram_cell[    8074] = 32'h8b29db04;
    ram_cell[    8075] = 32'h7fe12bf1;
    ram_cell[    8076] = 32'ha27235b3;
    ram_cell[    8077] = 32'h2f12cb5c;
    ram_cell[    8078] = 32'hce02eb9a;
    ram_cell[    8079] = 32'hc3f2ed79;
    ram_cell[    8080] = 32'h531fdd0e;
    ram_cell[    8081] = 32'h8e277f26;
    ram_cell[    8082] = 32'h19cebf61;
    ram_cell[    8083] = 32'h95679e6a;
    ram_cell[    8084] = 32'h48ee3243;
    ram_cell[    8085] = 32'h95c19a14;
    ram_cell[    8086] = 32'hc6bb98d5;
    ram_cell[    8087] = 32'h63dcef0e;
    ram_cell[    8088] = 32'h553ca023;
    ram_cell[    8089] = 32'he2b2587b;
    ram_cell[    8090] = 32'h6ae1ef84;
    ram_cell[    8091] = 32'ha68f5f41;
    ram_cell[    8092] = 32'hae688745;
    ram_cell[    8093] = 32'h96699cfe;
    ram_cell[    8094] = 32'h7f0ebd66;
    ram_cell[    8095] = 32'h2c075495;
    ram_cell[    8096] = 32'heb30b065;
    ram_cell[    8097] = 32'h8a9384fd;
    ram_cell[    8098] = 32'h10cd32b2;
    ram_cell[    8099] = 32'h53455234;
    ram_cell[    8100] = 32'hacecfee8;
    ram_cell[    8101] = 32'h72ae850e;
    ram_cell[    8102] = 32'h0395ecd5;
    ram_cell[    8103] = 32'h965afaff;
    ram_cell[    8104] = 32'h3089127c;
    ram_cell[    8105] = 32'hba4f7f80;
    ram_cell[    8106] = 32'h35ff5fca;
    ram_cell[    8107] = 32'h51b9baff;
    ram_cell[    8108] = 32'h215c1c2b;
    ram_cell[    8109] = 32'hcac6d072;
    ram_cell[    8110] = 32'h8f3b24b9;
    ram_cell[    8111] = 32'h1463520b;
    ram_cell[    8112] = 32'h47939cf7;
    ram_cell[    8113] = 32'hd74fe78a;
    ram_cell[    8114] = 32'h09e98ce5;
    ram_cell[    8115] = 32'h8737aaf9;
    ram_cell[    8116] = 32'h62852a64;
    ram_cell[    8117] = 32'hdd983bf4;
    ram_cell[    8118] = 32'h22811085;
    ram_cell[    8119] = 32'h9eb665b0;
    ram_cell[    8120] = 32'hdfec9775;
    ram_cell[    8121] = 32'hafa41a2a;
    ram_cell[    8122] = 32'h811ceb67;
    ram_cell[    8123] = 32'h8896c3fc;
    ram_cell[    8124] = 32'he3f92ef9;
    ram_cell[    8125] = 32'hc03abb19;
    ram_cell[    8126] = 32'h688b4ced;
    ram_cell[    8127] = 32'hf920bae3;
    ram_cell[    8128] = 32'hceb1792d;
    ram_cell[    8129] = 32'h52e5c8db;
    ram_cell[    8130] = 32'hce1a6066;
    ram_cell[    8131] = 32'ha4b67801;
    ram_cell[    8132] = 32'h10e1f7b8;
    ram_cell[    8133] = 32'h02f6cb62;
    ram_cell[    8134] = 32'h6cbd3e6f;
    ram_cell[    8135] = 32'hce6dd1a3;
    ram_cell[    8136] = 32'h65d8b470;
    ram_cell[    8137] = 32'h7371b797;
    ram_cell[    8138] = 32'hcc040f10;
    ram_cell[    8139] = 32'h290173fb;
    ram_cell[    8140] = 32'hcc307682;
    ram_cell[    8141] = 32'h934ec4f3;
    ram_cell[    8142] = 32'hfc393ce0;
    ram_cell[    8143] = 32'h1c984314;
    ram_cell[    8144] = 32'h91e5515e;
    ram_cell[    8145] = 32'hfd16cdb6;
    ram_cell[    8146] = 32'h6f384f69;
    ram_cell[    8147] = 32'h8750f773;
    ram_cell[    8148] = 32'h14a8aef4;
    ram_cell[    8149] = 32'h8d4eda5a;
    ram_cell[    8150] = 32'ha07b9a82;
    ram_cell[    8151] = 32'h0757a809;
    ram_cell[    8152] = 32'haaec06bd;
    ram_cell[    8153] = 32'h08abfac9;
    ram_cell[    8154] = 32'h60f5f5f4;
    ram_cell[    8155] = 32'hca954bcf;
    ram_cell[    8156] = 32'hd49ced3d;
    ram_cell[    8157] = 32'h84acb023;
    ram_cell[    8158] = 32'h6db64988;
    ram_cell[    8159] = 32'h41a5ffd6;
    ram_cell[    8160] = 32'h05123adb;
    ram_cell[    8161] = 32'hd5a1e1fe;
    ram_cell[    8162] = 32'ha0b37738;
    ram_cell[    8163] = 32'h27e2b1b0;
    ram_cell[    8164] = 32'h75347e1b;
    ram_cell[    8165] = 32'h1bbe3cbf;
    ram_cell[    8166] = 32'h11f09099;
    ram_cell[    8167] = 32'hc121d013;
    ram_cell[    8168] = 32'hc37bf927;
    ram_cell[    8169] = 32'h4fb5a839;
    ram_cell[    8170] = 32'he2b8bced;
    ram_cell[    8171] = 32'h7c524497;
    ram_cell[    8172] = 32'h98909f5b;
    ram_cell[    8173] = 32'h94dab86f;
    ram_cell[    8174] = 32'h1ad842a3;
    ram_cell[    8175] = 32'h554aef45;
    ram_cell[    8176] = 32'hfa1d7a35;
    ram_cell[    8177] = 32'heed85f85;
    ram_cell[    8178] = 32'hd01cbefb;
    ram_cell[    8179] = 32'h689d4b4b;
    ram_cell[    8180] = 32'hec444b1f;
    ram_cell[    8181] = 32'hfaba9450;
    ram_cell[    8182] = 32'h9b33da70;
    ram_cell[    8183] = 32'h2868245b;
    ram_cell[    8184] = 32'h875d8576;
    ram_cell[    8185] = 32'h0f082ef0;
    ram_cell[    8186] = 32'h7d93a17b;
    ram_cell[    8187] = 32'hf2f8dced;
    ram_cell[    8188] = 32'hdc53ae62;
    ram_cell[    8189] = 32'h48cbf396;
    ram_cell[    8190] = 32'h023fcf97;
    ram_cell[    8191] = 32'h83e02403;
    // src matrix B
    ram_cell[    8192] = 32'h4533b3f1;
    ram_cell[    8193] = 32'hafa1f175;
    ram_cell[    8194] = 32'h6cd093f7;
    ram_cell[    8195] = 32'h963df274;
    ram_cell[    8196] = 32'h73f4202a;
    ram_cell[    8197] = 32'he5ad84c9;
    ram_cell[    8198] = 32'h30980e5f;
    ram_cell[    8199] = 32'h53bf94e0;
    ram_cell[    8200] = 32'h9b1661d0;
    ram_cell[    8201] = 32'h51e254bb;
    ram_cell[    8202] = 32'h3d6fcf24;
    ram_cell[    8203] = 32'h4ff37567;
    ram_cell[    8204] = 32'hc4366e3a;
    ram_cell[    8205] = 32'hc5949eac;
    ram_cell[    8206] = 32'h9bb26286;
    ram_cell[    8207] = 32'h91d46be7;
    ram_cell[    8208] = 32'h19eb775e;
    ram_cell[    8209] = 32'h7f13c412;
    ram_cell[    8210] = 32'h05e0b612;
    ram_cell[    8211] = 32'h9e8c31a8;
    ram_cell[    8212] = 32'h1a8bcc91;
    ram_cell[    8213] = 32'h0ade918f;
    ram_cell[    8214] = 32'h18ae1a14;
    ram_cell[    8215] = 32'hbeff31dd;
    ram_cell[    8216] = 32'h5a28e30f;
    ram_cell[    8217] = 32'h0e5c0e29;
    ram_cell[    8218] = 32'ha7dd4213;
    ram_cell[    8219] = 32'hcaed517f;
    ram_cell[    8220] = 32'h399fdab3;
    ram_cell[    8221] = 32'h9c929e50;
    ram_cell[    8222] = 32'h53dd4a76;
    ram_cell[    8223] = 32'h9af528b2;
    ram_cell[    8224] = 32'h86bfe83f;
    ram_cell[    8225] = 32'heb6cea0f;
    ram_cell[    8226] = 32'h3212a3d7;
    ram_cell[    8227] = 32'h0da6ac81;
    ram_cell[    8228] = 32'ha8bb900c;
    ram_cell[    8229] = 32'hca632073;
    ram_cell[    8230] = 32'heece2afc;
    ram_cell[    8231] = 32'h34bf0db1;
    ram_cell[    8232] = 32'hcfd439a4;
    ram_cell[    8233] = 32'h4d6a8d78;
    ram_cell[    8234] = 32'h25f07bce;
    ram_cell[    8235] = 32'h0064accb;
    ram_cell[    8236] = 32'h3b6d4704;
    ram_cell[    8237] = 32'hda3e4064;
    ram_cell[    8238] = 32'h2fe01a4b;
    ram_cell[    8239] = 32'h73b37c98;
    ram_cell[    8240] = 32'h08e6bb45;
    ram_cell[    8241] = 32'ha7d50171;
    ram_cell[    8242] = 32'h22e51088;
    ram_cell[    8243] = 32'h54bfd177;
    ram_cell[    8244] = 32'hc117cae0;
    ram_cell[    8245] = 32'h94f36f66;
    ram_cell[    8246] = 32'h381f1eb6;
    ram_cell[    8247] = 32'hc5949639;
    ram_cell[    8248] = 32'h036ad693;
    ram_cell[    8249] = 32'hacd83f40;
    ram_cell[    8250] = 32'h610f053e;
    ram_cell[    8251] = 32'h125c3aa6;
    ram_cell[    8252] = 32'haeafdbaf;
    ram_cell[    8253] = 32'hb1011d36;
    ram_cell[    8254] = 32'h6bb68e60;
    ram_cell[    8255] = 32'h0096600d;
    ram_cell[    8256] = 32'h7cef7ace;
    ram_cell[    8257] = 32'he8546ad4;
    ram_cell[    8258] = 32'h8722edc3;
    ram_cell[    8259] = 32'h579948fc;
    ram_cell[    8260] = 32'heff358ab;
    ram_cell[    8261] = 32'h225a61f0;
    ram_cell[    8262] = 32'h8fc7378f;
    ram_cell[    8263] = 32'hdcf4f73d;
    ram_cell[    8264] = 32'h12ec7aa3;
    ram_cell[    8265] = 32'hd010e67c;
    ram_cell[    8266] = 32'h4e4ce195;
    ram_cell[    8267] = 32'h328c85d1;
    ram_cell[    8268] = 32'h7ca6e23f;
    ram_cell[    8269] = 32'hcf57d26a;
    ram_cell[    8270] = 32'h5960373d;
    ram_cell[    8271] = 32'h601d1329;
    ram_cell[    8272] = 32'he70129a1;
    ram_cell[    8273] = 32'h2bbd7fcd;
    ram_cell[    8274] = 32'h7da3fffd;
    ram_cell[    8275] = 32'h158f4f1e;
    ram_cell[    8276] = 32'h5be3e728;
    ram_cell[    8277] = 32'h67714918;
    ram_cell[    8278] = 32'hfc6d0006;
    ram_cell[    8279] = 32'h330bd807;
    ram_cell[    8280] = 32'hac5044f3;
    ram_cell[    8281] = 32'h6fd7ac14;
    ram_cell[    8282] = 32'h0fec2e3f;
    ram_cell[    8283] = 32'h9e804d7b;
    ram_cell[    8284] = 32'h58dbe270;
    ram_cell[    8285] = 32'hd5d4c3b7;
    ram_cell[    8286] = 32'hc947e635;
    ram_cell[    8287] = 32'h4147037e;
    ram_cell[    8288] = 32'h93bc771b;
    ram_cell[    8289] = 32'h35b85ad9;
    ram_cell[    8290] = 32'h7528267b;
    ram_cell[    8291] = 32'hfe14cc4e;
    ram_cell[    8292] = 32'hfcf67194;
    ram_cell[    8293] = 32'h58f6c716;
    ram_cell[    8294] = 32'h8da80c0e;
    ram_cell[    8295] = 32'h126c34de;
    ram_cell[    8296] = 32'h5770b133;
    ram_cell[    8297] = 32'h886bfc61;
    ram_cell[    8298] = 32'h10c6b087;
    ram_cell[    8299] = 32'h7f3e75b9;
    ram_cell[    8300] = 32'h9f0e5ccf;
    ram_cell[    8301] = 32'hdc2306f8;
    ram_cell[    8302] = 32'h51271822;
    ram_cell[    8303] = 32'h219cecc7;
    ram_cell[    8304] = 32'hdb56c47a;
    ram_cell[    8305] = 32'h7840cc09;
    ram_cell[    8306] = 32'hd3cc8681;
    ram_cell[    8307] = 32'hba54cb3b;
    ram_cell[    8308] = 32'h248e41a0;
    ram_cell[    8309] = 32'h7ef8d3f5;
    ram_cell[    8310] = 32'hf90318b0;
    ram_cell[    8311] = 32'h39767b17;
    ram_cell[    8312] = 32'h651f387f;
    ram_cell[    8313] = 32'h0ddd499c;
    ram_cell[    8314] = 32'h67ee8a7b;
    ram_cell[    8315] = 32'hb1758bbe;
    ram_cell[    8316] = 32'h6630949a;
    ram_cell[    8317] = 32'h81322c60;
    ram_cell[    8318] = 32'hdba4ac57;
    ram_cell[    8319] = 32'ha82fa4e4;
    ram_cell[    8320] = 32'h33f273bd;
    ram_cell[    8321] = 32'h34883587;
    ram_cell[    8322] = 32'h41ad29a4;
    ram_cell[    8323] = 32'hc9f81822;
    ram_cell[    8324] = 32'h2bdcf83c;
    ram_cell[    8325] = 32'h18f7c998;
    ram_cell[    8326] = 32'hb0cc9c68;
    ram_cell[    8327] = 32'hc403f8bd;
    ram_cell[    8328] = 32'hbeed325b;
    ram_cell[    8329] = 32'h22d30884;
    ram_cell[    8330] = 32'h58322204;
    ram_cell[    8331] = 32'h873ebc13;
    ram_cell[    8332] = 32'h68cb66fc;
    ram_cell[    8333] = 32'h9f4f01aa;
    ram_cell[    8334] = 32'h14b51c1c;
    ram_cell[    8335] = 32'h26d89f77;
    ram_cell[    8336] = 32'h2150a451;
    ram_cell[    8337] = 32'h7aac6207;
    ram_cell[    8338] = 32'hfad4ec25;
    ram_cell[    8339] = 32'h17303176;
    ram_cell[    8340] = 32'h3fe87f10;
    ram_cell[    8341] = 32'h7446759c;
    ram_cell[    8342] = 32'h46a92eb5;
    ram_cell[    8343] = 32'he2c894ee;
    ram_cell[    8344] = 32'he38dec57;
    ram_cell[    8345] = 32'h68b280a8;
    ram_cell[    8346] = 32'hac98db49;
    ram_cell[    8347] = 32'hc1965b64;
    ram_cell[    8348] = 32'hc259c42e;
    ram_cell[    8349] = 32'hcc7a9a94;
    ram_cell[    8350] = 32'h55c1c771;
    ram_cell[    8351] = 32'h7c49832b;
    ram_cell[    8352] = 32'ha7e91842;
    ram_cell[    8353] = 32'heed1ef56;
    ram_cell[    8354] = 32'hf6003978;
    ram_cell[    8355] = 32'h0673290a;
    ram_cell[    8356] = 32'hc7d90ea2;
    ram_cell[    8357] = 32'hf4a0b3c4;
    ram_cell[    8358] = 32'hbd70c81e;
    ram_cell[    8359] = 32'hdd2d7a80;
    ram_cell[    8360] = 32'hbdbf0bf5;
    ram_cell[    8361] = 32'he7b8b2d0;
    ram_cell[    8362] = 32'h201bd509;
    ram_cell[    8363] = 32'h539eead4;
    ram_cell[    8364] = 32'hb6260b54;
    ram_cell[    8365] = 32'hdb3c6b85;
    ram_cell[    8366] = 32'he7513ee8;
    ram_cell[    8367] = 32'h28b4d614;
    ram_cell[    8368] = 32'h6f53d6c1;
    ram_cell[    8369] = 32'hdca2670c;
    ram_cell[    8370] = 32'h15e7feee;
    ram_cell[    8371] = 32'hacc01ddf;
    ram_cell[    8372] = 32'h7cd59b2e;
    ram_cell[    8373] = 32'hf13a548f;
    ram_cell[    8374] = 32'h23d8547c;
    ram_cell[    8375] = 32'h2a6467e5;
    ram_cell[    8376] = 32'h689f0d7d;
    ram_cell[    8377] = 32'h84253f47;
    ram_cell[    8378] = 32'h5fb361fe;
    ram_cell[    8379] = 32'h479e20fc;
    ram_cell[    8380] = 32'hafc40571;
    ram_cell[    8381] = 32'hdfe0f867;
    ram_cell[    8382] = 32'h3ac74dd5;
    ram_cell[    8383] = 32'h4ca9203b;
    ram_cell[    8384] = 32'h37b0cf5c;
    ram_cell[    8385] = 32'had48b98c;
    ram_cell[    8386] = 32'h6c793a45;
    ram_cell[    8387] = 32'ha5e26781;
    ram_cell[    8388] = 32'h26661870;
    ram_cell[    8389] = 32'h156b654f;
    ram_cell[    8390] = 32'hc00bb0d1;
    ram_cell[    8391] = 32'h9dd920e0;
    ram_cell[    8392] = 32'h2af01dcb;
    ram_cell[    8393] = 32'h68f770eb;
    ram_cell[    8394] = 32'h307d452a;
    ram_cell[    8395] = 32'h1e1da0b5;
    ram_cell[    8396] = 32'hc6a85803;
    ram_cell[    8397] = 32'h8ff01d93;
    ram_cell[    8398] = 32'h2795ccc8;
    ram_cell[    8399] = 32'h289ca158;
    ram_cell[    8400] = 32'h0c9b7fb1;
    ram_cell[    8401] = 32'hb3f35e38;
    ram_cell[    8402] = 32'h7281f896;
    ram_cell[    8403] = 32'hcd3ae90b;
    ram_cell[    8404] = 32'ha7fbbc75;
    ram_cell[    8405] = 32'h8d1f292f;
    ram_cell[    8406] = 32'hc1f5560f;
    ram_cell[    8407] = 32'h09a122ec;
    ram_cell[    8408] = 32'hbfd49ea6;
    ram_cell[    8409] = 32'h562f9a2f;
    ram_cell[    8410] = 32'hfcabb9e0;
    ram_cell[    8411] = 32'hc993290d;
    ram_cell[    8412] = 32'hf06ac0b3;
    ram_cell[    8413] = 32'h769932e5;
    ram_cell[    8414] = 32'h52a291e2;
    ram_cell[    8415] = 32'he27cd41d;
    ram_cell[    8416] = 32'h84175538;
    ram_cell[    8417] = 32'h853e7bf4;
    ram_cell[    8418] = 32'h36f8241c;
    ram_cell[    8419] = 32'h631b3f01;
    ram_cell[    8420] = 32'hfefe9c62;
    ram_cell[    8421] = 32'h438dc9de;
    ram_cell[    8422] = 32'h89c980ee;
    ram_cell[    8423] = 32'hce9a9e42;
    ram_cell[    8424] = 32'hc947155e;
    ram_cell[    8425] = 32'h51373d91;
    ram_cell[    8426] = 32'hc2e801d3;
    ram_cell[    8427] = 32'h6cfee8e4;
    ram_cell[    8428] = 32'h2b088b33;
    ram_cell[    8429] = 32'h353f9f72;
    ram_cell[    8430] = 32'h891bf6bb;
    ram_cell[    8431] = 32'h3d829264;
    ram_cell[    8432] = 32'h87c7745e;
    ram_cell[    8433] = 32'h068bab66;
    ram_cell[    8434] = 32'h97804bc0;
    ram_cell[    8435] = 32'hc80d08ed;
    ram_cell[    8436] = 32'h9a29c7de;
    ram_cell[    8437] = 32'h7837bcc7;
    ram_cell[    8438] = 32'hffdfd074;
    ram_cell[    8439] = 32'h271aaf13;
    ram_cell[    8440] = 32'hcf866035;
    ram_cell[    8441] = 32'h6361020e;
    ram_cell[    8442] = 32'hce19e735;
    ram_cell[    8443] = 32'h0621d326;
    ram_cell[    8444] = 32'h47c2d41a;
    ram_cell[    8445] = 32'h9eac7d44;
    ram_cell[    8446] = 32'hfeb5dde6;
    ram_cell[    8447] = 32'h99846a79;
    ram_cell[    8448] = 32'hc73272e8;
    ram_cell[    8449] = 32'h6b364341;
    ram_cell[    8450] = 32'hb25b1fc7;
    ram_cell[    8451] = 32'hd19a3df6;
    ram_cell[    8452] = 32'hb16daeef;
    ram_cell[    8453] = 32'h10c53e65;
    ram_cell[    8454] = 32'h36023a07;
    ram_cell[    8455] = 32'he5952afc;
    ram_cell[    8456] = 32'h3525b7ff;
    ram_cell[    8457] = 32'h948e52a3;
    ram_cell[    8458] = 32'hd2380e25;
    ram_cell[    8459] = 32'h802a19b8;
    ram_cell[    8460] = 32'hf85320a8;
    ram_cell[    8461] = 32'hf61bfafb;
    ram_cell[    8462] = 32'h2e10506d;
    ram_cell[    8463] = 32'hc652d3ec;
    ram_cell[    8464] = 32'h02409971;
    ram_cell[    8465] = 32'h0b95abb0;
    ram_cell[    8466] = 32'h5786c36b;
    ram_cell[    8467] = 32'h58d20e6f;
    ram_cell[    8468] = 32'h113ded13;
    ram_cell[    8469] = 32'he52e8bf0;
    ram_cell[    8470] = 32'h09d9fd75;
    ram_cell[    8471] = 32'h9f377867;
    ram_cell[    8472] = 32'h79ac999a;
    ram_cell[    8473] = 32'h9f551d43;
    ram_cell[    8474] = 32'h548bc324;
    ram_cell[    8475] = 32'h492d62a2;
    ram_cell[    8476] = 32'h32d3c8c0;
    ram_cell[    8477] = 32'h425202d7;
    ram_cell[    8478] = 32'h3ea10fac;
    ram_cell[    8479] = 32'hcd361bda;
    ram_cell[    8480] = 32'hc62cb6b7;
    ram_cell[    8481] = 32'hff9b9c06;
    ram_cell[    8482] = 32'habaaca2b;
    ram_cell[    8483] = 32'h2365adb2;
    ram_cell[    8484] = 32'he090aef6;
    ram_cell[    8485] = 32'hcff89d42;
    ram_cell[    8486] = 32'he4ff0d73;
    ram_cell[    8487] = 32'hfa8c4015;
    ram_cell[    8488] = 32'h391a1b61;
    ram_cell[    8489] = 32'h5c75c57e;
    ram_cell[    8490] = 32'h68d51c47;
    ram_cell[    8491] = 32'h4112070f;
    ram_cell[    8492] = 32'h1b7be611;
    ram_cell[    8493] = 32'h5c151956;
    ram_cell[    8494] = 32'h00f65bdf;
    ram_cell[    8495] = 32'h31178bb5;
    ram_cell[    8496] = 32'h942a0fd3;
    ram_cell[    8497] = 32'h52d8b993;
    ram_cell[    8498] = 32'h94b2e66a;
    ram_cell[    8499] = 32'h03228d2a;
    ram_cell[    8500] = 32'h54a2c900;
    ram_cell[    8501] = 32'hf0304d20;
    ram_cell[    8502] = 32'h4319cf2f;
    ram_cell[    8503] = 32'h38ad0f26;
    ram_cell[    8504] = 32'h67ab1a8d;
    ram_cell[    8505] = 32'hd1dd3835;
    ram_cell[    8506] = 32'h92af68d6;
    ram_cell[    8507] = 32'h444a041f;
    ram_cell[    8508] = 32'h061dd52a;
    ram_cell[    8509] = 32'hdaed2eb5;
    ram_cell[    8510] = 32'hb0aea765;
    ram_cell[    8511] = 32'hb1f41b2e;
    ram_cell[    8512] = 32'h9690ffb2;
    ram_cell[    8513] = 32'h6f6dd7d6;
    ram_cell[    8514] = 32'hc6b4beda;
    ram_cell[    8515] = 32'h27579639;
    ram_cell[    8516] = 32'hfe1f18fc;
    ram_cell[    8517] = 32'hdc25c39d;
    ram_cell[    8518] = 32'h2890ba26;
    ram_cell[    8519] = 32'h6ff624bc;
    ram_cell[    8520] = 32'h97ecb022;
    ram_cell[    8521] = 32'h4f3bbc8c;
    ram_cell[    8522] = 32'h59e219f4;
    ram_cell[    8523] = 32'hc2a59125;
    ram_cell[    8524] = 32'h5e0c1cf2;
    ram_cell[    8525] = 32'hc00c7853;
    ram_cell[    8526] = 32'hcd42fc0d;
    ram_cell[    8527] = 32'h87e12aab;
    ram_cell[    8528] = 32'h4c7a0c4a;
    ram_cell[    8529] = 32'ha32f44ff;
    ram_cell[    8530] = 32'h6d8946fa;
    ram_cell[    8531] = 32'h62364043;
    ram_cell[    8532] = 32'hef5b51e9;
    ram_cell[    8533] = 32'h9e8ee2a0;
    ram_cell[    8534] = 32'h49d5337d;
    ram_cell[    8535] = 32'h582f24c6;
    ram_cell[    8536] = 32'hd4536155;
    ram_cell[    8537] = 32'h744039e3;
    ram_cell[    8538] = 32'ha3c6277b;
    ram_cell[    8539] = 32'ha615c3d9;
    ram_cell[    8540] = 32'hf3f774ca;
    ram_cell[    8541] = 32'h87b91903;
    ram_cell[    8542] = 32'h307e0549;
    ram_cell[    8543] = 32'h35327645;
    ram_cell[    8544] = 32'haa1b34e7;
    ram_cell[    8545] = 32'hdf79fc98;
    ram_cell[    8546] = 32'h76a6042c;
    ram_cell[    8547] = 32'h243f59d3;
    ram_cell[    8548] = 32'h41cca482;
    ram_cell[    8549] = 32'hff350efa;
    ram_cell[    8550] = 32'h3a9efcf3;
    ram_cell[    8551] = 32'h7ebec397;
    ram_cell[    8552] = 32'ha330bc9a;
    ram_cell[    8553] = 32'h6c0cb809;
    ram_cell[    8554] = 32'hb867aae7;
    ram_cell[    8555] = 32'hcae7118f;
    ram_cell[    8556] = 32'h407b56e1;
    ram_cell[    8557] = 32'h609c7918;
    ram_cell[    8558] = 32'hcceaaeb4;
    ram_cell[    8559] = 32'h7ad6f681;
    ram_cell[    8560] = 32'hdfad3163;
    ram_cell[    8561] = 32'h32359458;
    ram_cell[    8562] = 32'hdbf7cb50;
    ram_cell[    8563] = 32'hc78b10bb;
    ram_cell[    8564] = 32'h2d0b0391;
    ram_cell[    8565] = 32'h936e4ebd;
    ram_cell[    8566] = 32'h71f0ae54;
    ram_cell[    8567] = 32'h36f09c53;
    ram_cell[    8568] = 32'h7bef8653;
    ram_cell[    8569] = 32'h2ac2bac8;
    ram_cell[    8570] = 32'h02a48b93;
    ram_cell[    8571] = 32'he667dda8;
    ram_cell[    8572] = 32'h45294838;
    ram_cell[    8573] = 32'ha6c6bbc0;
    ram_cell[    8574] = 32'hb47fc34d;
    ram_cell[    8575] = 32'h98e8a72a;
    ram_cell[    8576] = 32'hd7bcf3ab;
    ram_cell[    8577] = 32'hd41eb595;
    ram_cell[    8578] = 32'h70c148a9;
    ram_cell[    8579] = 32'h2bfd5d4d;
    ram_cell[    8580] = 32'h7d82216b;
    ram_cell[    8581] = 32'h858c3b40;
    ram_cell[    8582] = 32'h0e1635db;
    ram_cell[    8583] = 32'hb3d6d9e8;
    ram_cell[    8584] = 32'hea8f68e6;
    ram_cell[    8585] = 32'h57844121;
    ram_cell[    8586] = 32'h26a357e1;
    ram_cell[    8587] = 32'h7be487c5;
    ram_cell[    8588] = 32'hae5460a8;
    ram_cell[    8589] = 32'h81973367;
    ram_cell[    8590] = 32'h9230159a;
    ram_cell[    8591] = 32'h7bde2343;
    ram_cell[    8592] = 32'h776a9cce;
    ram_cell[    8593] = 32'h2cbd594f;
    ram_cell[    8594] = 32'h3fdf5dd8;
    ram_cell[    8595] = 32'h36b7df46;
    ram_cell[    8596] = 32'h195cf330;
    ram_cell[    8597] = 32'hd11a1059;
    ram_cell[    8598] = 32'hef93d42e;
    ram_cell[    8599] = 32'h70da745e;
    ram_cell[    8600] = 32'hdb7b9bef;
    ram_cell[    8601] = 32'ha4f93d21;
    ram_cell[    8602] = 32'hcee924ce;
    ram_cell[    8603] = 32'h67bbbe40;
    ram_cell[    8604] = 32'h8ecb803c;
    ram_cell[    8605] = 32'h875151d0;
    ram_cell[    8606] = 32'h1d0dba1a;
    ram_cell[    8607] = 32'h6bcacd1b;
    ram_cell[    8608] = 32'hc1ee25a9;
    ram_cell[    8609] = 32'hd472506c;
    ram_cell[    8610] = 32'hbbb0a1b5;
    ram_cell[    8611] = 32'hf4d22e14;
    ram_cell[    8612] = 32'hf5621d07;
    ram_cell[    8613] = 32'h7444bb14;
    ram_cell[    8614] = 32'h9c326ef1;
    ram_cell[    8615] = 32'hc1377826;
    ram_cell[    8616] = 32'hd5173dd2;
    ram_cell[    8617] = 32'h244f5ca1;
    ram_cell[    8618] = 32'haefe0578;
    ram_cell[    8619] = 32'h4ff873d6;
    ram_cell[    8620] = 32'h8db15dda;
    ram_cell[    8621] = 32'hdf6f6dce;
    ram_cell[    8622] = 32'he47136ff;
    ram_cell[    8623] = 32'h9ce21d03;
    ram_cell[    8624] = 32'h8c8d1d67;
    ram_cell[    8625] = 32'hd02eaee6;
    ram_cell[    8626] = 32'h72480c72;
    ram_cell[    8627] = 32'h93e2a33f;
    ram_cell[    8628] = 32'h997b54d2;
    ram_cell[    8629] = 32'h3cc9a784;
    ram_cell[    8630] = 32'hde95bcaf;
    ram_cell[    8631] = 32'ha135d1c5;
    ram_cell[    8632] = 32'h64b09528;
    ram_cell[    8633] = 32'h75ff3486;
    ram_cell[    8634] = 32'he276ea7c;
    ram_cell[    8635] = 32'h0d253c36;
    ram_cell[    8636] = 32'h59116806;
    ram_cell[    8637] = 32'h7f7e58e6;
    ram_cell[    8638] = 32'hc81d2ee3;
    ram_cell[    8639] = 32'hd210edb7;
    ram_cell[    8640] = 32'h26f065e9;
    ram_cell[    8641] = 32'he9da3b72;
    ram_cell[    8642] = 32'hacd83a1f;
    ram_cell[    8643] = 32'hf54ecdfa;
    ram_cell[    8644] = 32'h4622f601;
    ram_cell[    8645] = 32'hbb1e039d;
    ram_cell[    8646] = 32'hebe6b72a;
    ram_cell[    8647] = 32'h0bb421b8;
    ram_cell[    8648] = 32'h220dacfe;
    ram_cell[    8649] = 32'hc5f667fa;
    ram_cell[    8650] = 32'h2b5ed5eb;
    ram_cell[    8651] = 32'h2a119342;
    ram_cell[    8652] = 32'h234fceb3;
    ram_cell[    8653] = 32'h3eb32836;
    ram_cell[    8654] = 32'h3cb04215;
    ram_cell[    8655] = 32'ha38cc512;
    ram_cell[    8656] = 32'h3dbe52d8;
    ram_cell[    8657] = 32'h942c6c26;
    ram_cell[    8658] = 32'hb5840fb6;
    ram_cell[    8659] = 32'hbdf36e93;
    ram_cell[    8660] = 32'hb28b883d;
    ram_cell[    8661] = 32'h4c795343;
    ram_cell[    8662] = 32'h94e94764;
    ram_cell[    8663] = 32'hbfdb0630;
    ram_cell[    8664] = 32'h337a7795;
    ram_cell[    8665] = 32'h98952259;
    ram_cell[    8666] = 32'hb8b40d43;
    ram_cell[    8667] = 32'h59837abc;
    ram_cell[    8668] = 32'h0d42312d;
    ram_cell[    8669] = 32'h52eb114e;
    ram_cell[    8670] = 32'h20b00d29;
    ram_cell[    8671] = 32'h9b9efa69;
    ram_cell[    8672] = 32'h31715746;
    ram_cell[    8673] = 32'ha0dd8e98;
    ram_cell[    8674] = 32'h5661ff70;
    ram_cell[    8675] = 32'h3816f5c7;
    ram_cell[    8676] = 32'hd7f78275;
    ram_cell[    8677] = 32'h40eac424;
    ram_cell[    8678] = 32'h2543ded6;
    ram_cell[    8679] = 32'h95cf6c19;
    ram_cell[    8680] = 32'h67698709;
    ram_cell[    8681] = 32'hb62a0951;
    ram_cell[    8682] = 32'h9783dac7;
    ram_cell[    8683] = 32'h83eb32cc;
    ram_cell[    8684] = 32'h59c6149c;
    ram_cell[    8685] = 32'h958be7c5;
    ram_cell[    8686] = 32'hdd969fb3;
    ram_cell[    8687] = 32'h2c74a942;
    ram_cell[    8688] = 32'ha757bd43;
    ram_cell[    8689] = 32'h6f354e0b;
    ram_cell[    8690] = 32'hf2c43d20;
    ram_cell[    8691] = 32'h9194f53b;
    ram_cell[    8692] = 32'hee339c74;
    ram_cell[    8693] = 32'hf08f7c9d;
    ram_cell[    8694] = 32'he1b7d8f0;
    ram_cell[    8695] = 32'hebba30a6;
    ram_cell[    8696] = 32'h738ebcf6;
    ram_cell[    8697] = 32'hd9c0615b;
    ram_cell[    8698] = 32'h50aad7d5;
    ram_cell[    8699] = 32'hdc11f40f;
    ram_cell[    8700] = 32'h20615c2a;
    ram_cell[    8701] = 32'he2f0e34e;
    ram_cell[    8702] = 32'h1c9e87c5;
    ram_cell[    8703] = 32'h1aed9063;
    ram_cell[    8704] = 32'h6fc38c54;
    ram_cell[    8705] = 32'h42460870;
    ram_cell[    8706] = 32'h0382c3e0;
    ram_cell[    8707] = 32'h93e05218;
    ram_cell[    8708] = 32'hf6640731;
    ram_cell[    8709] = 32'hb634539c;
    ram_cell[    8710] = 32'h8c3f81d8;
    ram_cell[    8711] = 32'hf7814913;
    ram_cell[    8712] = 32'hac7683af;
    ram_cell[    8713] = 32'hcc35b1f2;
    ram_cell[    8714] = 32'h6c5c776f;
    ram_cell[    8715] = 32'h53a8910c;
    ram_cell[    8716] = 32'h1d5c3f19;
    ram_cell[    8717] = 32'hd7b98154;
    ram_cell[    8718] = 32'hcf0d2c53;
    ram_cell[    8719] = 32'h84e83c8b;
    ram_cell[    8720] = 32'hbd31e3f9;
    ram_cell[    8721] = 32'hfb5d1578;
    ram_cell[    8722] = 32'h619a6a78;
    ram_cell[    8723] = 32'h4ee836cf;
    ram_cell[    8724] = 32'heef55ed4;
    ram_cell[    8725] = 32'h3fcdf8eb;
    ram_cell[    8726] = 32'hc1217bed;
    ram_cell[    8727] = 32'h5fe3cd49;
    ram_cell[    8728] = 32'hdd6eb99c;
    ram_cell[    8729] = 32'h242054a0;
    ram_cell[    8730] = 32'h512b57e4;
    ram_cell[    8731] = 32'h887a6621;
    ram_cell[    8732] = 32'h304a05b6;
    ram_cell[    8733] = 32'hfd839d11;
    ram_cell[    8734] = 32'h6b499c24;
    ram_cell[    8735] = 32'h2591f383;
    ram_cell[    8736] = 32'h48069aa7;
    ram_cell[    8737] = 32'hbb5ff0b2;
    ram_cell[    8738] = 32'hbbb682d5;
    ram_cell[    8739] = 32'h855c1562;
    ram_cell[    8740] = 32'hbceb8e01;
    ram_cell[    8741] = 32'ha0e94b1a;
    ram_cell[    8742] = 32'hfa9b3af1;
    ram_cell[    8743] = 32'he181b9d6;
    ram_cell[    8744] = 32'h94183726;
    ram_cell[    8745] = 32'hf34e3e97;
    ram_cell[    8746] = 32'haa3eac03;
    ram_cell[    8747] = 32'hb72758c1;
    ram_cell[    8748] = 32'hf9c82122;
    ram_cell[    8749] = 32'h5f2e5b27;
    ram_cell[    8750] = 32'h8c2ae0f0;
    ram_cell[    8751] = 32'hd10e9521;
    ram_cell[    8752] = 32'h710c619a;
    ram_cell[    8753] = 32'hb241269e;
    ram_cell[    8754] = 32'h83fd2e33;
    ram_cell[    8755] = 32'h99149985;
    ram_cell[    8756] = 32'h2a12648a;
    ram_cell[    8757] = 32'haa74b6d2;
    ram_cell[    8758] = 32'hc1a09ff7;
    ram_cell[    8759] = 32'h92182c8f;
    ram_cell[    8760] = 32'h06732d8b;
    ram_cell[    8761] = 32'h3dde5ca4;
    ram_cell[    8762] = 32'h6876b2c0;
    ram_cell[    8763] = 32'hc2ad4b4d;
    ram_cell[    8764] = 32'haaff1893;
    ram_cell[    8765] = 32'hc7812b62;
    ram_cell[    8766] = 32'h49d2ce3d;
    ram_cell[    8767] = 32'hd68d66db;
    ram_cell[    8768] = 32'h03a864e1;
    ram_cell[    8769] = 32'hcc862915;
    ram_cell[    8770] = 32'h34924f1b;
    ram_cell[    8771] = 32'h8e328812;
    ram_cell[    8772] = 32'h04a0ad18;
    ram_cell[    8773] = 32'h6569d527;
    ram_cell[    8774] = 32'h986c5180;
    ram_cell[    8775] = 32'ha657902c;
    ram_cell[    8776] = 32'hd15ad950;
    ram_cell[    8777] = 32'h73f760bf;
    ram_cell[    8778] = 32'h8b0f4a32;
    ram_cell[    8779] = 32'h2d6ac392;
    ram_cell[    8780] = 32'h14111a56;
    ram_cell[    8781] = 32'h1023b337;
    ram_cell[    8782] = 32'h2e11e727;
    ram_cell[    8783] = 32'ha5d2b0dd;
    ram_cell[    8784] = 32'h3adb063f;
    ram_cell[    8785] = 32'hdda78c32;
    ram_cell[    8786] = 32'h32ce89f3;
    ram_cell[    8787] = 32'hb2eb6a4a;
    ram_cell[    8788] = 32'h54719db8;
    ram_cell[    8789] = 32'h9ca3b31c;
    ram_cell[    8790] = 32'hf7cebef2;
    ram_cell[    8791] = 32'ha0eea849;
    ram_cell[    8792] = 32'hf9ad1eee;
    ram_cell[    8793] = 32'hac11b350;
    ram_cell[    8794] = 32'hdc69e838;
    ram_cell[    8795] = 32'h51997ce0;
    ram_cell[    8796] = 32'h0504efdd;
    ram_cell[    8797] = 32'h48b71ae2;
    ram_cell[    8798] = 32'hb5c37480;
    ram_cell[    8799] = 32'ha792998e;
    ram_cell[    8800] = 32'h4bed1c11;
    ram_cell[    8801] = 32'h089920dd;
    ram_cell[    8802] = 32'h1094606a;
    ram_cell[    8803] = 32'hecba4116;
    ram_cell[    8804] = 32'habaedb97;
    ram_cell[    8805] = 32'h00ccad59;
    ram_cell[    8806] = 32'hcef4fd20;
    ram_cell[    8807] = 32'h8526428c;
    ram_cell[    8808] = 32'hcb03025b;
    ram_cell[    8809] = 32'h062c1ccb;
    ram_cell[    8810] = 32'h3b9541c1;
    ram_cell[    8811] = 32'hd53a315e;
    ram_cell[    8812] = 32'heba2258c;
    ram_cell[    8813] = 32'h3bf27899;
    ram_cell[    8814] = 32'h913cb17d;
    ram_cell[    8815] = 32'h42ffb206;
    ram_cell[    8816] = 32'hd2b2834b;
    ram_cell[    8817] = 32'hbb4a5e6b;
    ram_cell[    8818] = 32'hd4c9518a;
    ram_cell[    8819] = 32'h96924a86;
    ram_cell[    8820] = 32'hf84de274;
    ram_cell[    8821] = 32'hb02ba707;
    ram_cell[    8822] = 32'hd89f6b62;
    ram_cell[    8823] = 32'ha49dda63;
    ram_cell[    8824] = 32'h50660749;
    ram_cell[    8825] = 32'hc940fe0a;
    ram_cell[    8826] = 32'h6d40c974;
    ram_cell[    8827] = 32'h80b4e2ab;
    ram_cell[    8828] = 32'h9551f1dc;
    ram_cell[    8829] = 32'hd327b115;
    ram_cell[    8830] = 32'ha1565390;
    ram_cell[    8831] = 32'hb99e4a02;
    ram_cell[    8832] = 32'hb14bd8d7;
    ram_cell[    8833] = 32'h609e67a3;
    ram_cell[    8834] = 32'hb41d495e;
    ram_cell[    8835] = 32'h4305dd23;
    ram_cell[    8836] = 32'h8298951f;
    ram_cell[    8837] = 32'h57bb3e42;
    ram_cell[    8838] = 32'h5ac46a3e;
    ram_cell[    8839] = 32'h0dd9eaca;
    ram_cell[    8840] = 32'haea35b23;
    ram_cell[    8841] = 32'h6bdd1fd5;
    ram_cell[    8842] = 32'h7539d3a6;
    ram_cell[    8843] = 32'hb2b40aba;
    ram_cell[    8844] = 32'h2f9ece2f;
    ram_cell[    8845] = 32'h9c42bd1c;
    ram_cell[    8846] = 32'hb4e5a3ba;
    ram_cell[    8847] = 32'ha1851f78;
    ram_cell[    8848] = 32'h52265a40;
    ram_cell[    8849] = 32'h15fc0e39;
    ram_cell[    8850] = 32'hddf5c989;
    ram_cell[    8851] = 32'h325e8289;
    ram_cell[    8852] = 32'h09a543e5;
    ram_cell[    8853] = 32'h1d9313e3;
    ram_cell[    8854] = 32'h8f471ba9;
    ram_cell[    8855] = 32'hc0410c03;
    ram_cell[    8856] = 32'h06306325;
    ram_cell[    8857] = 32'hb8b56968;
    ram_cell[    8858] = 32'he19623a5;
    ram_cell[    8859] = 32'hafe0ebdd;
    ram_cell[    8860] = 32'h78ab9166;
    ram_cell[    8861] = 32'head18568;
    ram_cell[    8862] = 32'h2977eac4;
    ram_cell[    8863] = 32'h45d3f32d;
    ram_cell[    8864] = 32'h1a28396e;
    ram_cell[    8865] = 32'h0ad8fc69;
    ram_cell[    8866] = 32'ha4e27aad;
    ram_cell[    8867] = 32'hca1759a6;
    ram_cell[    8868] = 32'h0a833c47;
    ram_cell[    8869] = 32'hd1614a72;
    ram_cell[    8870] = 32'h5396aa59;
    ram_cell[    8871] = 32'hb20f167e;
    ram_cell[    8872] = 32'hd0fecf1d;
    ram_cell[    8873] = 32'h48e9124c;
    ram_cell[    8874] = 32'hc3a210fa;
    ram_cell[    8875] = 32'h3bd91052;
    ram_cell[    8876] = 32'h72b6b30f;
    ram_cell[    8877] = 32'h0d2a8b16;
    ram_cell[    8878] = 32'hf08700a1;
    ram_cell[    8879] = 32'h2f4395ce;
    ram_cell[    8880] = 32'he722da12;
    ram_cell[    8881] = 32'h1d660eb4;
    ram_cell[    8882] = 32'h8ea0ba06;
    ram_cell[    8883] = 32'hf10690ba;
    ram_cell[    8884] = 32'h7bef09ce;
    ram_cell[    8885] = 32'h8dafc693;
    ram_cell[    8886] = 32'hb4291c93;
    ram_cell[    8887] = 32'h859c0b81;
    ram_cell[    8888] = 32'h53d61ce0;
    ram_cell[    8889] = 32'he111f7f8;
    ram_cell[    8890] = 32'h9c7f2671;
    ram_cell[    8891] = 32'h1e574b2f;
    ram_cell[    8892] = 32'h62da7dc6;
    ram_cell[    8893] = 32'h296e2a25;
    ram_cell[    8894] = 32'h0ec02736;
    ram_cell[    8895] = 32'h654f9275;
    ram_cell[    8896] = 32'h711391b3;
    ram_cell[    8897] = 32'h5fad9016;
    ram_cell[    8898] = 32'h61048911;
    ram_cell[    8899] = 32'hbcfdbea7;
    ram_cell[    8900] = 32'h5b923e4e;
    ram_cell[    8901] = 32'h04764b03;
    ram_cell[    8902] = 32'h301f7f3c;
    ram_cell[    8903] = 32'h08cfee8c;
    ram_cell[    8904] = 32'h0a6d2080;
    ram_cell[    8905] = 32'h825275c1;
    ram_cell[    8906] = 32'hdd8c2a1d;
    ram_cell[    8907] = 32'hb061d48a;
    ram_cell[    8908] = 32'hcdeae728;
    ram_cell[    8909] = 32'ha070e5ed;
    ram_cell[    8910] = 32'hcf25daaf;
    ram_cell[    8911] = 32'h8454d7d1;
    ram_cell[    8912] = 32'hb221ae5d;
    ram_cell[    8913] = 32'hc8b2619e;
    ram_cell[    8914] = 32'h0bcdf762;
    ram_cell[    8915] = 32'he0e6e256;
    ram_cell[    8916] = 32'hf9811af4;
    ram_cell[    8917] = 32'h03de296b;
    ram_cell[    8918] = 32'h826ddc0a;
    ram_cell[    8919] = 32'he0c425a8;
    ram_cell[    8920] = 32'hf626cc99;
    ram_cell[    8921] = 32'hc0d1f68f;
    ram_cell[    8922] = 32'h42d0f50d;
    ram_cell[    8923] = 32'h168482b5;
    ram_cell[    8924] = 32'h018a7c0c;
    ram_cell[    8925] = 32'hc728d91f;
    ram_cell[    8926] = 32'h44205a13;
    ram_cell[    8927] = 32'h1c85795a;
    ram_cell[    8928] = 32'hbc9d15da;
    ram_cell[    8929] = 32'h17922f02;
    ram_cell[    8930] = 32'ha9175d2d;
    ram_cell[    8931] = 32'hd99c057f;
    ram_cell[    8932] = 32'h47f7d903;
    ram_cell[    8933] = 32'h501334b3;
    ram_cell[    8934] = 32'hd78d9ad4;
    ram_cell[    8935] = 32'h80a6a39c;
    ram_cell[    8936] = 32'hcc0d2002;
    ram_cell[    8937] = 32'h13df93a2;
    ram_cell[    8938] = 32'h6d3a13a6;
    ram_cell[    8939] = 32'hb02db78b;
    ram_cell[    8940] = 32'h1864b8aa;
    ram_cell[    8941] = 32'he927c2dd;
    ram_cell[    8942] = 32'hc8893f05;
    ram_cell[    8943] = 32'ha9153099;
    ram_cell[    8944] = 32'hef800e72;
    ram_cell[    8945] = 32'h5b83df90;
    ram_cell[    8946] = 32'hc74e93aa;
    ram_cell[    8947] = 32'hfba09980;
    ram_cell[    8948] = 32'h049b2c4a;
    ram_cell[    8949] = 32'hf4be0e81;
    ram_cell[    8950] = 32'h0b9322d5;
    ram_cell[    8951] = 32'h9ddd4592;
    ram_cell[    8952] = 32'ha4c6b029;
    ram_cell[    8953] = 32'h3f1fd8c3;
    ram_cell[    8954] = 32'h035267c7;
    ram_cell[    8955] = 32'h2701d024;
    ram_cell[    8956] = 32'he9c8b179;
    ram_cell[    8957] = 32'h1c342b44;
    ram_cell[    8958] = 32'h0804f98b;
    ram_cell[    8959] = 32'h02641a89;
    ram_cell[    8960] = 32'hc31457ed;
    ram_cell[    8961] = 32'hfc4b2676;
    ram_cell[    8962] = 32'h3ef3d51a;
    ram_cell[    8963] = 32'hbe42ffe2;
    ram_cell[    8964] = 32'h523086ad;
    ram_cell[    8965] = 32'h91d25fa0;
    ram_cell[    8966] = 32'hf50f12fe;
    ram_cell[    8967] = 32'h10a25180;
    ram_cell[    8968] = 32'h55f6d859;
    ram_cell[    8969] = 32'hff52038c;
    ram_cell[    8970] = 32'hff374762;
    ram_cell[    8971] = 32'h250d909c;
    ram_cell[    8972] = 32'ha132d8b2;
    ram_cell[    8973] = 32'h984bc4fa;
    ram_cell[    8974] = 32'h7fa64cbe;
    ram_cell[    8975] = 32'hbea4b898;
    ram_cell[    8976] = 32'h7a980e18;
    ram_cell[    8977] = 32'h8cd45efb;
    ram_cell[    8978] = 32'h88d0e0ec;
    ram_cell[    8979] = 32'h368991f4;
    ram_cell[    8980] = 32'h0b12b959;
    ram_cell[    8981] = 32'h55abe22e;
    ram_cell[    8982] = 32'heb927a3f;
    ram_cell[    8983] = 32'hb59b7dfe;
    ram_cell[    8984] = 32'h79630d3d;
    ram_cell[    8985] = 32'h3cf4cbdf;
    ram_cell[    8986] = 32'hb85ebc20;
    ram_cell[    8987] = 32'h7e5e0f6a;
    ram_cell[    8988] = 32'hc214d90c;
    ram_cell[    8989] = 32'ha046110d;
    ram_cell[    8990] = 32'h703a4d1f;
    ram_cell[    8991] = 32'h96758c3d;
    ram_cell[    8992] = 32'h9620ccd8;
    ram_cell[    8993] = 32'h2e0a0350;
    ram_cell[    8994] = 32'hbbbf9fef;
    ram_cell[    8995] = 32'hf97dc63f;
    ram_cell[    8996] = 32'h5de6041c;
    ram_cell[    8997] = 32'hf5e836f2;
    ram_cell[    8998] = 32'h9511cd78;
    ram_cell[    8999] = 32'hd5d7c6ab;
    ram_cell[    9000] = 32'hbf1357f9;
    ram_cell[    9001] = 32'hc4d523a2;
    ram_cell[    9002] = 32'habcbaffc;
    ram_cell[    9003] = 32'h7a541bd5;
    ram_cell[    9004] = 32'h5183e038;
    ram_cell[    9005] = 32'h0c712c93;
    ram_cell[    9006] = 32'hd3c1aae4;
    ram_cell[    9007] = 32'h65543b28;
    ram_cell[    9008] = 32'ha1c2363c;
    ram_cell[    9009] = 32'h6b07cc3f;
    ram_cell[    9010] = 32'h560d585c;
    ram_cell[    9011] = 32'h983023cc;
    ram_cell[    9012] = 32'h7d0bf001;
    ram_cell[    9013] = 32'h977777f4;
    ram_cell[    9014] = 32'hc51b18a3;
    ram_cell[    9015] = 32'h57673e1e;
    ram_cell[    9016] = 32'h6622ae0c;
    ram_cell[    9017] = 32'h4d688750;
    ram_cell[    9018] = 32'h94eee536;
    ram_cell[    9019] = 32'h8368315a;
    ram_cell[    9020] = 32'h347b0672;
    ram_cell[    9021] = 32'h96c41ceb;
    ram_cell[    9022] = 32'h502d70da;
    ram_cell[    9023] = 32'h35dfeeea;
    ram_cell[    9024] = 32'h2179353f;
    ram_cell[    9025] = 32'h8175837a;
    ram_cell[    9026] = 32'h89baffd7;
    ram_cell[    9027] = 32'h1e20e102;
    ram_cell[    9028] = 32'h16d58f52;
    ram_cell[    9029] = 32'h5b5cc794;
    ram_cell[    9030] = 32'h2b0c33a5;
    ram_cell[    9031] = 32'h22fe4a26;
    ram_cell[    9032] = 32'hf2ce22ae;
    ram_cell[    9033] = 32'h4bdae0cf;
    ram_cell[    9034] = 32'hf9e61108;
    ram_cell[    9035] = 32'hbf3cd391;
    ram_cell[    9036] = 32'h57bb6557;
    ram_cell[    9037] = 32'h18345ddd;
    ram_cell[    9038] = 32'ha3d886b5;
    ram_cell[    9039] = 32'h252eec56;
    ram_cell[    9040] = 32'hbb05a5b3;
    ram_cell[    9041] = 32'h06790270;
    ram_cell[    9042] = 32'hd4d1436e;
    ram_cell[    9043] = 32'h4fd7bbb7;
    ram_cell[    9044] = 32'h33496c06;
    ram_cell[    9045] = 32'he645d60c;
    ram_cell[    9046] = 32'h3ecbeddc;
    ram_cell[    9047] = 32'h84afa67f;
    ram_cell[    9048] = 32'hfdc9abad;
    ram_cell[    9049] = 32'h7f92c374;
    ram_cell[    9050] = 32'h835e90e6;
    ram_cell[    9051] = 32'h62c051b3;
    ram_cell[    9052] = 32'hf6c79102;
    ram_cell[    9053] = 32'hbc7d5ed1;
    ram_cell[    9054] = 32'had0bfedf;
    ram_cell[    9055] = 32'h917765ce;
    ram_cell[    9056] = 32'h4f35eeb9;
    ram_cell[    9057] = 32'h506ff082;
    ram_cell[    9058] = 32'h17afa341;
    ram_cell[    9059] = 32'h39669c2b;
    ram_cell[    9060] = 32'hbd550985;
    ram_cell[    9061] = 32'h683d2efc;
    ram_cell[    9062] = 32'h1c41f120;
    ram_cell[    9063] = 32'hbe68e5ac;
    ram_cell[    9064] = 32'hd6cb6d9a;
    ram_cell[    9065] = 32'h0b0f0820;
    ram_cell[    9066] = 32'h319559be;
    ram_cell[    9067] = 32'hc64f085b;
    ram_cell[    9068] = 32'h48199349;
    ram_cell[    9069] = 32'h802af053;
    ram_cell[    9070] = 32'he62da27e;
    ram_cell[    9071] = 32'he4c4cf6b;
    ram_cell[    9072] = 32'h31159d67;
    ram_cell[    9073] = 32'h1342f189;
    ram_cell[    9074] = 32'hba86eb1d;
    ram_cell[    9075] = 32'h88e05d59;
    ram_cell[    9076] = 32'h8075e485;
    ram_cell[    9077] = 32'h7fdcacea;
    ram_cell[    9078] = 32'hc79e2e0f;
    ram_cell[    9079] = 32'hf1458770;
    ram_cell[    9080] = 32'hf3753c66;
    ram_cell[    9081] = 32'hfcce842c;
    ram_cell[    9082] = 32'h7c1e8aa7;
    ram_cell[    9083] = 32'h1e1871e4;
    ram_cell[    9084] = 32'h8510cdc3;
    ram_cell[    9085] = 32'h596abd3e;
    ram_cell[    9086] = 32'h5e16615a;
    ram_cell[    9087] = 32'he567c0c1;
    ram_cell[    9088] = 32'h8540dbc6;
    ram_cell[    9089] = 32'hadfd356d;
    ram_cell[    9090] = 32'h6013b990;
    ram_cell[    9091] = 32'hb355a902;
    ram_cell[    9092] = 32'hd9b60014;
    ram_cell[    9093] = 32'h30c94ff5;
    ram_cell[    9094] = 32'ha01e44eb;
    ram_cell[    9095] = 32'h4c0ace72;
    ram_cell[    9096] = 32'h98dee830;
    ram_cell[    9097] = 32'h4c829ccb;
    ram_cell[    9098] = 32'hf43f5ae0;
    ram_cell[    9099] = 32'hc6a79e6b;
    ram_cell[    9100] = 32'h5d445033;
    ram_cell[    9101] = 32'ha83722bb;
    ram_cell[    9102] = 32'h06887363;
    ram_cell[    9103] = 32'h7a11f4c7;
    ram_cell[    9104] = 32'ha2ff7bf5;
    ram_cell[    9105] = 32'hc2eebcdd;
    ram_cell[    9106] = 32'hf5742d18;
    ram_cell[    9107] = 32'h65233faa;
    ram_cell[    9108] = 32'hc38ce60f;
    ram_cell[    9109] = 32'h11eb84ba;
    ram_cell[    9110] = 32'hef57e233;
    ram_cell[    9111] = 32'hf2ba6ac1;
    ram_cell[    9112] = 32'he17df433;
    ram_cell[    9113] = 32'h6e93a946;
    ram_cell[    9114] = 32'hffd83f8f;
    ram_cell[    9115] = 32'h11b8c3c6;
    ram_cell[    9116] = 32'h7995e57c;
    ram_cell[    9117] = 32'h171fd110;
    ram_cell[    9118] = 32'h2db936db;
    ram_cell[    9119] = 32'h5151c08b;
    ram_cell[    9120] = 32'h79d8a5cf;
    ram_cell[    9121] = 32'hdc918af8;
    ram_cell[    9122] = 32'hdd9b1302;
    ram_cell[    9123] = 32'hf61a9ad1;
    ram_cell[    9124] = 32'h9c0cbf4e;
    ram_cell[    9125] = 32'h2a69047c;
    ram_cell[    9126] = 32'h4a2ca965;
    ram_cell[    9127] = 32'he8ae1744;
    ram_cell[    9128] = 32'hdc5ac06a;
    ram_cell[    9129] = 32'h4531345b;
    ram_cell[    9130] = 32'h78d6349a;
    ram_cell[    9131] = 32'h28b157ed;
    ram_cell[    9132] = 32'ha48a2cc6;
    ram_cell[    9133] = 32'hb1adaed5;
    ram_cell[    9134] = 32'h3c9b9d49;
    ram_cell[    9135] = 32'h8d5ab01b;
    ram_cell[    9136] = 32'hc5279652;
    ram_cell[    9137] = 32'h67bda411;
    ram_cell[    9138] = 32'h4c1f026e;
    ram_cell[    9139] = 32'h04e8a32c;
    ram_cell[    9140] = 32'h16a8c4ee;
    ram_cell[    9141] = 32'h0e26a329;
    ram_cell[    9142] = 32'he3b4553e;
    ram_cell[    9143] = 32'h9e37d071;
    ram_cell[    9144] = 32'hd982886b;
    ram_cell[    9145] = 32'h75d46de6;
    ram_cell[    9146] = 32'h9a4732f7;
    ram_cell[    9147] = 32'hb6562410;
    ram_cell[    9148] = 32'h3d2bb34d;
    ram_cell[    9149] = 32'h8ef63531;
    ram_cell[    9150] = 32'h36c65ffb;
    ram_cell[    9151] = 32'h35220b92;
    ram_cell[    9152] = 32'hf7b80691;
    ram_cell[    9153] = 32'h68824931;
    ram_cell[    9154] = 32'hd11e4f77;
    ram_cell[    9155] = 32'h8f245e0a;
    ram_cell[    9156] = 32'h252203d5;
    ram_cell[    9157] = 32'h81d58ce8;
    ram_cell[    9158] = 32'h8552bcf6;
    ram_cell[    9159] = 32'hd5ca72ff;
    ram_cell[    9160] = 32'hda06d8cd;
    ram_cell[    9161] = 32'hbb03ba01;
    ram_cell[    9162] = 32'h278d32ac;
    ram_cell[    9163] = 32'h4cc6d33f;
    ram_cell[    9164] = 32'h4e47a07d;
    ram_cell[    9165] = 32'h9f85b162;
    ram_cell[    9166] = 32'ha8dd3f63;
    ram_cell[    9167] = 32'h667ce0f6;
    ram_cell[    9168] = 32'h3957f08c;
    ram_cell[    9169] = 32'h3ce5eaed;
    ram_cell[    9170] = 32'hed54eed3;
    ram_cell[    9171] = 32'h3e2c938a;
    ram_cell[    9172] = 32'h7e1ac45a;
    ram_cell[    9173] = 32'h74c17037;
    ram_cell[    9174] = 32'hb7ee829f;
    ram_cell[    9175] = 32'hd3fdf52f;
    ram_cell[    9176] = 32'h790623e7;
    ram_cell[    9177] = 32'he187d9c9;
    ram_cell[    9178] = 32'h7a7b3fc9;
    ram_cell[    9179] = 32'h9684ea1d;
    ram_cell[    9180] = 32'h84142e0f;
    ram_cell[    9181] = 32'h79b45265;
    ram_cell[    9182] = 32'h5558b6b3;
    ram_cell[    9183] = 32'h9830ac79;
    ram_cell[    9184] = 32'h0ec090bb;
    ram_cell[    9185] = 32'h4640d3c0;
    ram_cell[    9186] = 32'h92103b4d;
    ram_cell[    9187] = 32'h2fb95d58;
    ram_cell[    9188] = 32'h38fc6295;
    ram_cell[    9189] = 32'hfbede302;
    ram_cell[    9190] = 32'h4f8974a6;
    ram_cell[    9191] = 32'h1ec68682;
    ram_cell[    9192] = 32'h1d136961;
    ram_cell[    9193] = 32'h071acbae;
    ram_cell[    9194] = 32'h92ecc878;
    ram_cell[    9195] = 32'hea6ca74c;
    ram_cell[    9196] = 32'hb84b6ee1;
    ram_cell[    9197] = 32'h5ad7b9e3;
    ram_cell[    9198] = 32'ha2c3ad3a;
    ram_cell[    9199] = 32'hd3b7d231;
    ram_cell[    9200] = 32'h35318822;
    ram_cell[    9201] = 32'h82dac3e8;
    ram_cell[    9202] = 32'had332063;
    ram_cell[    9203] = 32'h2caacff9;
    ram_cell[    9204] = 32'h4e1be4bb;
    ram_cell[    9205] = 32'h9d1a1337;
    ram_cell[    9206] = 32'h4c972f44;
    ram_cell[    9207] = 32'h6f0d6e64;
    ram_cell[    9208] = 32'hfb5f6d2b;
    ram_cell[    9209] = 32'h99e752d1;
    ram_cell[    9210] = 32'hf280f47c;
    ram_cell[    9211] = 32'hd3388b67;
    ram_cell[    9212] = 32'h29ad9325;
    ram_cell[    9213] = 32'h44e6adaf;
    ram_cell[    9214] = 32'hc2c2ab19;
    ram_cell[    9215] = 32'hea77ff52;
    ram_cell[    9216] = 32'h5b7d0dda;
    ram_cell[    9217] = 32'h2ebb2cda;
    ram_cell[    9218] = 32'hca5bac42;
    ram_cell[    9219] = 32'h75adb702;
    ram_cell[    9220] = 32'hc7c75622;
    ram_cell[    9221] = 32'hf564b1a0;
    ram_cell[    9222] = 32'h66b5db78;
    ram_cell[    9223] = 32'h8ec502be;
    ram_cell[    9224] = 32'h2faaa4ef;
    ram_cell[    9225] = 32'h1c36e0ae;
    ram_cell[    9226] = 32'h96a81a9a;
    ram_cell[    9227] = 32'h432722f0;
    ram_cell[    9228] = 32'h6e197e55;
    ram_cell[    9229] = 32'hd7a92b88;
    ram_cell[    9230] = 32'h397a56d0;
    ram_cell[    9231] = 32'hb66238b4;
    ram_cell[    9232] = 32'h358d5b56;
    ram_cell[    9233] = 32'h46dc237e;
    ram_cell[    9234] = 32'hbdf119e9;
    ram_cell[    9235] = 32'h73570b78;
    ram_cell[    9236] = 32'h5b62ff23;
    ram_cell[    9237] = 32'h22d1caec;
    ram_cell[    9238] = 32'h42325058;
    ram_cell[    9239] = 32'h127695c4;
    ram_cell[    9240] = 32'hd878498e;
    ram_cell[    9241] = 32'hce33b626;
    ram_cell[    9242] = 32'h2b500a6d;
    ram_cell[    9243] = 32'h92150794;
    ram_cell[    9244] = 32'h2c73b9de;
    ram_cell[    9245] = 32'h2de786d3;
    ram_cell[    9246] = 32'h0a98cdd1;
    ram_cell[    9247] = 32'h0d353215;
    ram_cell[    9248] = 32'h0fceeeb2;
    ram_cell[    9249] = 32'h864d7441;
    ram_cell[    9250] = 32'h170b433e;
    ram_cell[    9251] = 32'h305c6902;
    ram_cell[    9252] = 32'h709c1c88;
    ram_cell[    9253] = 32'hc9f94d30;
    ram_cell[    9254] = 32'h9c8861d2;
    ram_cell[    9255] = 32'he6c5cd8c;
    ram_cell[    9256] = 32'he9412ec1;
    ram_cell[    9257] = 32'hd4f615e1;
    ram_cell[    9258] = 32'h671b3a8b;
    ram_cell[    9259] = 32'h7308b185;
    ram_cell[    9260] = 32'h343001ec;
    ram_cell[    9261] = 32'hfd2e826f;
    ram_cell[    9262] = 32'h1e64c9b4;
    ram_cell[    9263] = 32'h833d3882;
    ram_cell[    9264] = 32'h2bf21a39;
    ram_cell[    9265] = 32'h8a049e16;
    ram_cell[    9266] = 32'he2abc2e3;
    ram_cell[    9267] = 32'h0dcd4131;
    ram_cell[    9268] = 32'hc7f82cd4;
    ram_cell[    9269] = 32'h7e2b9b95;
    ram_cell[    9270] = 32'h894d0957;
    ram_cell[    9271] = 32'he2ff90b9;
    ram_cell[    9272] = 32'h0c0c1813;
    ram_cell[    9273] = 32'h2d420878;
    ram_cell[    9274] = 32'h955356cc;
    ram_cell[    9275] = 32'hae3ebb5e;
    ram_cell[    9276] = 32'h394b859f;
    ram_cell[    9277] = 32'hb30be03a;
    ram_cell[    9278] = 32'h5bbfec89;
    ram_cell[    9279] = 32'hb053cd04;
    ram_cell[    9280] = 32'h3e1e0525;
    ram_cell[    9281] = 32'h5923d362;
    ram_cell[    9282] = 32'h8f639954;
    ram_cell[    9283] = 32'h4945fbf6;
    ram_cell[    9284] = 32'h765b9f80;
    ram_cell[    9285] = 32'h7a8f21a3;
    ram_cell[    9286] = 32'hab05bb20;
    ram_cell[    9287] = 32'h1848622c;
    ram_cell[    9288] = 32'hc4ba4f67;
    ram_cell[    9289] = 32'he33e0e95;
    ram_cell[    9290] = 32'h865be841;
    ram_cell[    9291] = 32'h0d39c343;
    ram_cell[    9292] = 32'h63e886f1;
    ram_cell[    9293] = 32'h5b6b7cd3;
    ram_cell[    9294] = 32'h2113f042;
    ram_cell[    9295] = 32'h16bc7190;
    ram_cell[    9296] = 32'h96494293;
    ram_cell[    9297] = 32'h502a09a1;
    ram_cell[    9298] = 32'h33c2ddb4;
    ram_cell[    9299] = 32'h1a9b50d0;
    ram_cell[    9300] = 32'he38246bf;
    ram_cell[    9301] = 32'hb8d2020e;
    ram_cell[    9302] = 32'h71a84ebb;
    ram_cell[    9303] = 32'h2499cb23;
    ram_cell[    9304] = 32'h86428da3;
    ram_cell[    9305] = 32'hcf5fc279;
    ram_cell[    9306] = 32'h3b32d562;
    ram_cell[    9307] = 32'hb77c2497;
    ram_cell[    9308] = 32'hf106036c;
    ram_cell[    9309] = 32'h95d1cb9f;
    ram_cell[    9310] = 32'he1d5b8a8;
    ram_cell[    9311] = 32'h30fdc12d;
    ram_cell[    9312] = 32'hf3f524ae;
    ram_cell[    9313] = 32'h28dfd0c4;
    ram_cell[    9314] = 32'h72daef2e;
    ram_cell[    9315] = 32'h4637e652;
    ram_cell[    9316] = 32'hea8742b8;
    ram_cell[    9317] = 32'hd3f58f03;
    ram_cell[    9318] = 32'h4f643b29;
    ram_cell[    9319] = 32'hb1e01560;
    ram_cell[    9320] = 32'h328217d4;
    ram_cell[    9321] = 32'h99ac56d1;
    ram_cell[    9322] = 32'hc201e751;
    ram_cell[    9323] = 32'h979f274c;
    ram_cell[    9324] = 32'hfe3c484f;
    ram_cell[    9325] = 32'h510136bf;
    ram_cell[    9326] = 32'h7291caa5;
    ram_cell[    9327] = 32'hbc1d5a28;
    ram_cell[    9328] = 32'h77234a42;
    ram_cell[    9329] = 32'hc45ec71e;
    ram_cell[    9330] = 32'h9cbe52e9;
    ram_cell[    9331] = 32'hdbb61aa6;
    ram_cell[    9332] = 32'h73b43fb3;
    ram_cell[    9333] = 32'hcff7bb24;
    ram_cell[    9334] = 32'hb42e5c50;
    ram_cell[    9335] = 32'h89298e18;
    ram_cell[    9336] = 32'h072b1d0b;
    ram_cell[    9337] = 32'hbeb509d8;
    ram_cell[    9338] = 32'hd0fbc2ea;
    ram_cell[    9339] = 32'h657eedaa;
    ram_cell[    9340] = 32'hee7ad48f;
    ram_cell[    9341] = 32'h86337569;
    ram_cell[    9342] = 32'hbd8668df;
    ram_cell[    9343] = 32'he4ef2977;
    ram_cell[    9344] = 32'h5151a07b;
    ram_cell[    9345] = 32'h99fd425a;
    ram_cell[    9346] = 32'h31305b8f;
    ram_cell[    9347] = 32'he07a5485;
    ram_cell[    9348] = 32'h095a3781;
    ram_cell[    9349] = 32'h74a8ba09;
    ram_cell[    9350] = 32'h5a784f8f;
    ram_cell[    9351] = 32'h9bd2065a;
    ram_cell[    9352] = 32'h0c0d24e2;
    ram_cell[    9353] = 32'hf27caccf;
    ram_cell[    9354] = 32'hfd21b315;
    ram_cell[    9355] = 32'hb65dec41;
    ram_cell[    9356] = 32'h3f063a71;
    ram_cell[    9357] = 32'h52f80139;
    ram_cell[    9358] = 32'hb9f8d4ac;
    ram_cell[    9359] = 32'h5da01736;
    ram_cell[    9360] = 32'hd4154761;
    ram_cell[    9361] = 32'h86a46e55;
    ram_cell[    9362] = 32'h490f5779;
    ram_cell[    9363] = 32'h9bb66867;
    ram_cell[    9364] = 32'h66c4f9ce;
    ram_cell[    9365] = 32'h7d222d03;
    ram_cell[    9366] = 32'h1ef432c9;
    ram_cell[    9367] = 32'hab3f33e7;
    ram_cell[    9368] = 32'h483eb666;
    ram_cell[    9369] = 32'h855c722b;
    ram_cell[    9370] = 32'hd153be93;
    ram_cell[    9371] = 32'h67814306;
    ram_cell[    9372] = 32'h71277c59;
    ram_cell[    9373] = 32'h07508b18;
    ram_cell[    9374] = 32'hc76c1e85;
    ram_cell[    9375] = 32'hd8bc8047;
    ram_cell[    9376] = 32'h863de662;
    ram_cell[    9377] = 32'he4cc6448;
    ram_cell[    9378] = 32'ha741598d;
    ram_cell[    9379] = 32'hf23148cf;
    ram_cell[    9380] = 32'h84c0c3de;
    ram_cell[    9381] = 32'hd8ff408c;
    ram_cell[    9382] = 32'h0202966f;
    ram_cell[    9383] = 32'h875e690c;
    ram_cell[    9384] = 32'h6eb95b51;
    ram_cell[    9385] = 32'h0a5a75ad;
    ram_cell[    9386] = 32'hbe0dcbc3;
    ram_cell[    9387] = 32'h4cd2dc7f;
    ram_cell[    9388] = 32'h9aafd6a0;
    ram_cell[    9389] = 32'hbdf58f86;
    ram_cell[    9390] = 32'h9179d427;
    ram_cell[    9391] = 32'he5db0abf;
    ram_cell[    9392] = 32'haeb3ff36;
    ram_cell[    9393] = 32'h5b103520;
    ram_cell[    9394] = 32'h86b87563;
    ram_cell[    9395] = 32'h6641b25b;
    ram_cell[    9396] = 32'h9ef15600;
    ram_cell[    9397] = 32'hfd422307;
    ram_cell[    9398] = 32'h0bb1d7e0;
    ram_cell[    9399] = 32'h95783729;
    ram_cell[    9400] = 32'hc24cf78c;
    ram_cell[    9401] = 32'h3dabafb5;
    ram_cell[    9402] = 32'h22a88827;
    ram_cell[    9403] = 32'h8baf6e91;
    ram_cell[    9404] = 32'h4946eed9;
    ram_cell[    9405] = 32'h2c3516d1;
    ram_cell[    9406] = 32'h4f9f5653;
    ram_cell[    9407] = 32'h0acec099;
    ram_cell[    9408] = 32'h6e8b835c;
    ram_cell[    9409] = 32'h4e3a2392;
    ram_cell[    9410] = 32'h0c69137c;
    ram_cell[    9411] = 32'h902b043a;
    ram_cell[    9412] = 32'hbbf62fd7;
    ram_cell[    9413] = 32'h71aff6e2;
    ram_cell[    9414] = 32'h1581b66a;
    ram_cell[    9415] = 32'h09291301;
    ram_cell[    9416] = 32'hb3ee37d5;
    ram_cell[    9417] = 32'h600c7e97;
    ram_cell[    9418] = 32'h08ce155e;
    ram_cell[    9419] = 32'hb48fb6f3;
    ram_cell[    9420] = 32'h3d36f12e;
    ram_cell[    9421] = 32'hecc44e77;
    ram_cell[    9422] = 32'h6ec841b3;
    ram_cell[    9423] = 32'hac1ee442;
    ram_cell[    9424] = 32'hb8cbcd6b;
    ram_cell[    9425] = 32'hb0d2abc9;
    ram_cell[    9426] = 32'h3942a964;
    ram_cell[    9427] = 32'h616c7e6a;
    ram_cell[    9428] = 32'hdddeea3a;
    ram_cell[    9429] = 32'h3999de52;
    ram_cell[    9430] = 32'ha90755fa;
    ram_cell[    9431] = 32'ha5f3740d;
    ram_cell[    9432] = 32'hfc87e2fc;
    ram_cell[    9433] = 32'hea7fffcd;
    ram_cell[    9434] = 32'h24e62e9c;
    ram_cell[    9435] = 32'h2f7e0e35;
    ram_cell[    9436] = 32'h9d4adb1b;
    ram_cell[    9437] = 32'h3f34a9fa;
    ram_cell[    9438] = 32'h67477611;
    ram_cell[    9439] = 32'he3a03c62;
    ram_cell[    9440] = 32'h2222b3de;
    ram_cell[    9441] = 32'hf8a341d5;
    ram_cell[    9442] = 32'he6e444c9;
    ram_cell[    9443] = 32'hb239e4c3;
    ram_cell[    9444] = 32'hdb34702a;
    ram_cell[    9445] = 32'hffbfc9b7;
    ram_cell[    9446] = 32'hd1df4fe5;
    ram_cell[    9447] = 32'h68e77b77;
    ram_cell[    9448] = 32'h84db56da;
    ram_cell[    9449] = 32'h764daea5;
    ram_cell[    9450] = 32'hc81a0452;
    ram_cell[    9451] = 32'h9c11c849;
    ram_cell[    9452] = 32'hf68418b8;
    ram_cell[    9453] = 32'h504335d4;
    ram_cell[    9454] = 32'he4f23073;
    ram_cell[    9455] = 32'h4421ea0d;
    ram_cell[    9456] = 32'h0d6f20c0;
    ram_cell[    9457] = 32'h143aebad;
    ram_cell[    9458] = 32'hf56c63f2;
    ram_cell[    9459] = 32'h5d5a7b18;
    ram_cell[    9460] = 32'h70391de2;
    ram_cell[    9461] = 32'h511f1fa6;
    ram_cell[    9462] = 32'h7e0a59dc;
    ram_cell[    9463] = 32'h6189232c;
    ram_cell[    9464] = 32'he5a91c58;
    ram_cell[    9465] = 32'h687ed99e;
    ram_cell[    9466] = 32'h7396da17;
    ram_cell[    9467] = 32'hecffe90d;
    ram_cell[    9468] = 32'h7e3fbf50;
    ram_cell[    9469] = 32'h9287912b;
    ram_cell[    9470] = 32'hdf7851fe;
    ram_cell[    9471] = 32'ha47ae04b;
    ram_cell[    9472] = 32'h407b36ba;
    ram_cell[    9473] = 32'h6d21198b;
    ram_cell[    9474] = 32'h1bda5ccd;
    ram_cell[    9475] = 32'h33930f2a;
    ram_cell[    9476] = 32'h5be3510b;
    ram_cell[    9477] = 32'h1ef74d5c;
    ram_cell[    9478] = 32'h0035d73a;
    ram_cell[    9479] = 32'h3ed920da;
    ram_cell[    9480] = 32'h2e2246ee;
    ram_cell[    9481] = 32'hc7fb26a2;
    ram_cell[    9482] = 32'h8e8706d7;
    ram_cell[    9483] = 32'h363afb52;
    ram_cell[    9484] = 32'h5bb15e13;
    ram_cell[    9485] = 32'h115c308e;
    ram_cell[    9486] = 32'h79a2f29a;
    ram_cell[    9487] = 32'h6a470544;
    ram_cell[    9488] = 32'hd85d2965;
    ram_cell[    9489] = 32'h298341ef;
    ram_cell[    9490] = 32'h5070d0dd;
    ram_cell[    9491] = 32'hd4d9b51f;
    ram_cell[    9492] = 32'ha1a93e18;
    ram_cell[    9493] = 32'h993ab696;
    ram_cell[    9494] = 32'h53d78c29;
    ram_cell[    9495] = 32'ha0c69ef2;
    ram_cell[    9496] = 32'h50577e79;
    ram_cell[    9497] = 32'h6e7cccd5;
    ram_cell[    9498] = 32'h380881a8;
    ram_cell[    9499] = 32'hb8f08c9f;
    ram_cell[    9500] = 32'hed00f536;
    ram_cell[    9501] = 32'hb7562ca2;
    ram_cell[    9502] = 32'hd3b3ad59;
    ram_cell[    9503] = 32'he9e47100;
    ram_cell[    9504] = 32'hce92ea49;
    ram_cell[    9505] = 32'h41c7feff;
    ram_cell[    9506] = 32'h8242fa77;
    ram_cell[    9507] = 32'h4fb8b9e6;
    ram_cell[    9508] = 32'ha12dcb18;
    ram_cell[    9509] = 32'had18fc2f;
    ram_cell[    9510] = 32'h48c123df;
    ram_cell[    9511] = 32'hd4c78c15;
    ram_cell[    9512] = 32'h6a16fb8e;
    ram_cell[    9513] = 32'h76dedd3a;
    ram_cell[    9514] = 32'h6c568971;
    ram_cell[    9515] = 32'hd1dabe68;
    ram_cell[    9516] = 32'h8f378e6a;
    ram_cell[    9517] = 32'hfcb0c917;
    ram_cell[    9518] = 32'h5cd37db1;
    ram_cell[    9519] = 32'hea50b203;
    ram_cell[    9520] = 32'he8c039d8;
    ram_cell[    9521] = 32'h41ae0dbb;
    ram_cell[    9522] = 32'hb05aa2f6;
    ram_cell[    9523] = 32'h2fe0f413;
    ram_cell[    9524] = 32'h973c2ff6;
    ram_cell[    9525] = 32'heeed52ef;
    ram_cell[    9526] = 32'hd6efbe83;
    ram_cell[    9527] = 32'h747b3caf;
    ram_cell[    9528] = 32'h3a164071;
    ram_cell[    9529] = 32'h0d5ac027;
    ram_cell[    9530] = 32'h961beba9;
    ram_cell[    9531] = 32'h8497433a;
    ram_cell[    9532] = 32'h4c24e9ad;
    ram_cell[    9533] = 32'hf9162e1c;
    ram_cell[    9534] = 32'h14ef0277;
    ram_cell[    9535] = 32'hd50476a1;
    ram_cell[    9536] = 32'hc1d4d54e;
    ram_cell[    9537] = 32'h589ecfab;
    ram_cell[    9538] = 32'hbb31f2bc;
    ram_cell[    9539] = 32'h8aae19b3;
    ram_cell[    9540] = 32'hc95a5d0f;
    ram_cell[    9541] = 32'h418e7c00;
    ram_cell[    9542] = 32'h07996c84;
    ram_cell[    9543] = 32'h4b4f3ae1;
    ram_cell[    9544] = 32'he25de0ab;
    ram_cell[    9545] = 32'h545f4e2f;
    ram_cell[    9546] = 32'hed5357bb;
    ram_cell[    9547] = 32'h7a17ee65;
    ram_cell[    9548] = 32'h10d6fc89;
    ram_cell[    9549] = 32'h03557f72;
    ram_cell[    9550] = 32'h77c313dc;
    ram_cell[    9551] = 32'h63f4b099;
    ram_cell[    9552] = 32'h5ad721a9;
    ram_cell[    9553] = 32'hbdae7a27;
    ram_cell[    9554] = 32'h5fde9422;
    ram_cell[    9555] = 32'he6070a93;
    ram_cell[    9556] = 32'habcdde5e;
    ram_cell[    9557] = 32'h49184812;
    ram_cell[    9558] = 32'h701e8a67;
    ram_cell[    9559] = 32'hb3a1cbdd;
    ram_cell[    9560] = 32'h11bbc543;
    ram_cell[    9561] = 32'h9ff7b19f;
    ram_cell[    9562] = 32'h45beedac;
    ram_cell[    9563] = 32'h5c7ecd25;
    ram_cell[    9564] = 32'h07062646;
    ram_cell[    9565] = 32'he5cee665;
    ram_cell[    9566] = 32'heb6fba30;
    ram_cell[    9567] = 32'hcc64fffb;
    ram_cell[    9568] = 32'hb2fa17ec;
    ram_cell[    9569] = 32'h9fd69080;
    ram_cell[    9570] = 32'h76d1a36f;
    ram_cell[    9571] = 32'h56216888;
    ram_cell[    9572] = 32'h4c6bf10d;
    ram_cell[    9573] = 32'hf37e6568;
    ram_cell[    9574] = 32'ha906e328;
    ram_cell[    9575] = 32'h29567c18;
    ram_cell[    9576] = 32'h0de4fbc0;
    ram_cell[    9577] = 32'h061e1685;
    ram_cell[    9578] = 32'h7fa111fe;
    ram_cell[    9579] = 32'he29845d2;
    ram_cell[    9580] = 32'h95fc0b43;
    ram_cell[    9581] = 32'h774eab16;
    ram_cell[    9582] = 32'hfc6ad5fa;
    ram_cell[    9583] = 32'h8ea611c5;
    ram_cell[    9584] = 32'h3af70228;
    ram_cell[    9585] = 32'hde967823;
    ram_cell[    9586] = 32'h08d1a341;
    ram_cell[    9587] = 32'hbd339074;
    ram_cell[    9588] = 32'he41ab909;
    ram_cell[    9589] = 32'h85d16229;
    ram_cell[    9590] = 32'h576b98f7;
    ram_cell[    9591] = 32'h3bf467a6;
    ram_cell[    9592] = 32'h79d086e2;
    ram_cell[    9593] = 32'hedcf0fa5;
    ram_cell[    9594] = 32'h492e4141;
    ram_cell[    9595] = 32'h1170e5ed;
    ram_cell[    9596] = 32'hcef35481;
    ram_cell[    9597] = 32'ha1e512a4;
    ram_cell[    9598] = 32'hac5a77d4;
    ram_cell[    9599] = 32'h84859f6b;
    ram_cell[    9600] = 32'h5d6a8295;
    ram_cell[    9601] = 32'hc292cdb1;
    ram_cell[    9602] = 32'h1931cd2f;
    ram_cell[    9603] = 32'ha33fa979;
    ram_cell[    9604] = 32'h2d89aba9;
    ram_cell[    9605] = 32'ha4d4f790;
    ram_cell[    9606] = 32'h86f894e1;
    ram_cell[    9607] = 32'h51c36143;
    ram_cell[    9608] = 32'hb2f1147d;
    ram_cell[    9609] = 32'h810699db;
    ram_cell[    9610] = 32'hfb3874ea;
    ram_cell[    9611] = 32'h93505fe2;
    ram_cell[    9612] = 32'h947b9672;
    ram_cell[    9613] = 32'h8725b479;
    ram_cell[    9614] = 32'ha846dc00;
    ram_cell[    9615] = 32'h9716bf63;
    ram_cell[    9616] = 32'h723e520f;
    ram_cell[    9617] = 32'hc14ef397;
    ram_cell[    9618] = 32'h45a1b237;
    ram_cell[    9619] = 32'h06cd2bf3;
    ram_cell[    9620] = 32'h61962cd5;
    ram_cell[    9621] = 32'h0f5ef939;
    ram_cell[    9622] = 32'h93f7b721;
    ram_cell[    9623] = 32'h7a8ffc26;
    ram_cell[    9624] = 32'h62d360fc;
    ram_cell[    9625] = 32'hc00799e1;
    ram_cell[    9626] = 32'h5f61017a;
    ram_cell[    9627] = 32'h086e05e8;
    ram_cell[    9628] = 32'h99cf4728;
    ram_cell[    9629] = 32'hb8b499e5;
    ram_cell[    9630] = 32'he132f2e0;
    ram_cell[    9631] = 32'h541733f9;
    ram_cell[    9632] = 32'h0e2b7b9e;
    ram_cell[    9633] = 32'h9a1c46e2;
    ram_cell[    9634] = 32'h7f39963a;
    ram_cell[    9635] = 32'h25005dfe;
    ram_cell[    9636] = 32'h28a4eeb2;
    ram_cell[    9637] = 32'h18d4b2fc;
    ram_cell[    9638] = 32'h5e1a92a3;
    ram_cell[    9639] = 32'hcf267339;
    ram_cell[    9640] = 32'h349dec3c;
    ram_cell[    9641] = 32'h3ef23f8f;
    ram_cell[    9642] = 32'hba798146;
    ram_cell[    9643] = 32'h9a34af8a;
    ram_cell[    9644] = 32'hce24a656;
    ram_cell[    9645] = 32'h6cb7ca30;
    ram_cell[    9646] = 32'h5a2b3973;
    ram_cell[    9647] = 32'ha0b3582c;
    ram_cell[    9648] = 32'hc8ae88e4;
    ram_cell[    9649] = 32'h815d532d;
    ram_cell[    9650] = 32'hff8dc587;
    ram_cell[    9651] = 32'h40eb40b0;
    ram_cell[    9652] = 32'heb41e2d1;
    ram_cell[    9653] = 32'hab2314ab;
    ram_cell[    9654] = 32'h2e11d09e;
    ram_cell[    9655] = 32'h2db17095;
    ram_cell[    9656] = 32'h40324aa6;
    ram_cell[    9657] = 32'h3e1b9e9b;
    ram_cell[    9658] = 32'h0e0f5ce5;
    ram_cell[    9659] = 32'h5cc6eb75;
    ram_cell[    9660] = 32'hee4a8d67;
    ram_cell[    9661] = 32'h43d42c09;
    ram_cell[    9662] = 32'hac1e15f6;
    ram_cell[    9663] = 32'h8fa40548;
    ram_cell[    9664] = 32'h702b2656;
    ram_cell[    9665] = 32'h49e6afb8;
    ram_cell[    9666] = 32'h785da952;
    ram_cell[    9667] = 32'h89552e6f;
    ram_cell[    9668] = 32'hef21b603;
    ram_cell[    9669] = 32'hab745c73;
    ram_cell[    9670] = 32'h96d9698a;
    ram_cell[    9671] = 32'hd79a04e6;
    ram_cell[    9672] = 32'h0e36b079;
    ram_cell[    9673] = 32'h1a5f8140;
    ram_cell[    9674] = 32'h8cc20d9c;
    ram_cell[    9675] = 32'h8161fdb4;
    ram_cell[    9676] = 32'ha4b9ec6b;
    ram_cell[    9677] = 32'hdecea77a;
    ram_cell[    9678] = 32'h56fc1f09;
    ram_cell[    9679] = 32'h9790524f;
    ram_cell[    9680] = 32'h0d7a105c;
    ram_cell[    9681] = 32'h130fa6ba;
    ram_cell[    9682] = 32'hee7770e6;
    ram_cell[    9683] = 32'hb230e6d5;
    ram_cell[    9684] = 32'hb83c955b;
    ram_cell[    9685] = 32'hb0e23709;
    ram_cell[    9686] = 32'h581e0b53;
    ram_cell[    9687] = 32'h49e3123c;
    ram_cell[    9688] = 32'h1cac4f03;
    ram_cell[    9689] = 32'h27e9a664;
    ram_cell[    9690] = 32'h681a9903;
    ram_cell[    9691] = 32'hb8c34048;
    ram_cell[    9692] = 32'h6345b717;
    ram_cell[    9693] = 32'ha97d726c;
    ram_cell[    9694] = 32'h33ed00e6;
    ram_cell[    9695] = 32'habc1093d;
    ram_cell[    9696] = 32'h666be322;
    ram_cell[    9697] = 32'h9098826e;
    ram_cell[    9698] = 32'h9a727f0a;
    ram_cell[    9699] = 32'h549c9ddb;
    ram_cell[    9700] = 32'h7d5716fe;
    ram_cell[    9701] = 32'h037a2f36;
    ram_cell[    9702] = 32'hfd1f1cd3;
    ram_cell[    9703] = 32'h7ab2d339;
    ram_cell[    9704] = 32'hf5e24825;
    ram_cell[    9705] = 32'h13ade343;
    ram_cell[    9706] = 32'hec963af4;
    ram_cell[    9707] = 32'h4273f472;
    ram_cell[    9708] = 32'h87b6508f;
    ram_cell[    9709] = 32'hca8d8217;
    ram_cell[    9710] = 32'h73c6a7ba;
    ram_cell[    9711] = 32'h161f240b;
    ram_cell[    9712] = 32'h4f94cfdf;
    ram_cell[    9713] = 32'h1c438787;
    ram_cell[    9714] = 32'h37f05438;
    ram_cell[    9715] = 32'h70140357;
    ram_cell[    9716] = 32'h407faf33;
    ram_cell[    9717] = 32'hf2bf6fc6;
    ram_cell[    9718] = 32'hba5d3fdf;
    ram_cell[    9719] = 32'h82c6ac15;
    ram_cell[    9720] = 32'h90b18eb8;
    ram_cell[    9721] = 32'h26ad7a02;
    ram_cell[    9722] = 32'hdcc0c2ff;
    ram_cell[    9723] = 32'hd73dadfa;
    ram_cell[    9724] = 32'h369a3354;
    ram_cell[    9725] = 32'he088bae5;
    ram_cell[    9726] = 32'h0d31530e;
    ram_cell[    9727] = 32'h3df00342;
    ram_cell[    9728] = 32'h94ae4be1;
    ram_cell[    9729] = 32'h59eeec54;
    ram_cell[    9730] = 32'h558a02ce;
    ram_cell[    9731] = 32'h14769483;
    ram_cell[    9732] = 32'h7789b636;
    ram_cell[    9733] = 32'ha1ce8057;
    ram_cell[    9734] = 32'h2a33cf08;
    ram_cell[    9735] = 32'hfcff5332;
    ram_cell[    9736] = 32'h77924583;
    ram_cell[    9737] = 32'h666be019;
    ram_cell[    9738] = 32'h1dfaa32f;
    ram_cell[    9739] = 32'h42b3bcad;
    ram_cell[    9740] = 32'hedf7818e;
    ram_cell[    9741] = 32'h316357c4;
    ram_cell[    9742] = 32'h037dfc52;
    ram_cell[    9743] = 32'hbbcdb996;
    ram_cell[    9744] = 32'h8d5bbba3;
    ram_cell[    9745] = 32'h4cd2a028;
    ram_cell[    9746] = 32'hbad8b520;
    ram_cell[    9747] = 32'hdfa41c87;
    ram_cell[    9748] = 32'h8fcb0685;
    ram_cell[    9749] = 32'hc131182a;
    ram_cell[    9750] = 32'hf12eea56;
    ram_cell[    9751] = 32'hea5156a9;
    ram_cell[    9752] = 32'h1e3adb34;
    ram_cell[    9753] = 32'h7568cacc;
    ram_cell[    9754] = 32'h0c04559c;
    ram_cell[    9755] = 32'h2b732b79;
    ram_cell[    9756] = 32'hc11aa0f8;
    ram_cell[    9757] = 32'heaa7601c;
    ram_cell[    9758] = 32'h34ec0eaa;
    ram_cell[    9759] = 32'hd0b30775;
    ram_cell[    9760] = 32'h8bb9b9c4;
    ram_cell[    9761] = 32'hf000d18d;
    ram_cell[    9762] = 32'h4ebe2e57;
    ram_cell[    9763] = 32'ha2b7f40f;
    ram_cell[    9764] = 32'hdaa48aaa;
    ram_cell[    9765] = 32'ha874f987;
    ram_cell[    9766] = 32'h48ef8eed;
    ram_cell[    9767] = 32'h6dfaaaf8;
    ram_cell[    9768] = 32'h9ac9b758;
    ram_cell[    9769] = 32'h3767841f;
    ram_cell[    9770] = 32'h6c2638b5;
    ram_cell[    9771] = 32'hf3196dce;
    ram_cell[    9772] = 32'h62eb81fd;
    ram_cell[    9773] = 32'h745217a7;
    ram_cell[    9774] = 32'he25efcbd;
    ram_cell[    9775] = 32'h5966fd09;
    ram_cell[    9776] = 32'h33fbf698;
    ram_cell[    9777] = 32'h24197ee8;
    ram_cell[    9778] = 32'h8f9abd10;
    ram_cell[    9779] = 32'h9e114054;
    ram_cell[    9780] = 32'h6502e89e;
    ram_cell[    9781] = 32'ha68d6f03;
    ram_cell[    9782] = 32'h8f48b668;
    ram_cell[    9783] = 32'h4b60ff7f;
    ram_cell[    9784] = 32'h7fa56ad5;
    ram_cell[    9785] = 32'hc9070e79;
    ram_cell[    9786] = 32'hfd060b90;
    ram_cell[    9787] = 32'h002aa0b1;
    ram_cell[    9788] = 32'h333e4e99;
    ram_cell[    9789] = 32'hb9ec45ce;
    ram_cell[    9790] = 32'hbf098b63;
    ram_cell[    9791] = 32'hba9d58f2;
    ram_cell[    9792] = 32'h48b21d45;
    ram_cell[    9793] = 32'h56affca2;
    ram_cell[    9794] = 32'h88a1818e;
    ram_cell[    9795] = 32'h9ce2b17f;
    ram_cell[    9796] = 32'hd3398f69;
    ram_cell[    9797] = 32'h37678aa9;
    ram_cell[    9798] = 32'h74f62b50;
    ram_cell[    9799] = 32'hefd4be8a;
    ram_cell[    9800] = 32'hedccaed9;
    ram_cell[    9801] = 32'h16dd9b7f;
    ram_cell[    9802] = 32'h64e32a33;
    ram_cell[    9803] = 32'ha31437ce;
    ram_cell[    9804] = 32'h69b82f6b;
    ram_cell[    9805] = 32'h10d74572;
    ram_cell[    9806] = 32'hd8acee20;
    ram_cell[    9807] = 32'h12d0918b;
    ram_cell[    9808] = 32'hd78688f0;
    ram_cell[    9809] = 32'hd96366b4;
    ram_cell[    9810] = 32'h410c012d;
    ram_cell[    9811] = 32'h56f0edd0;
    ram_cell[    9812] = 32'h81bfd788;
    ram_cell[    9813] = 32'h10a2e637;
    ram_cell[    9814] = 32'hadca0a58;
    ram_cell[    9815] = 32'h135c8b77;
    ram_cell[    9816] = 32'h588c0848;
    ram_cell[    9817] = 32'h81f87b2d;
    ram_cell[    9818] = 32'hf48dd05f;
    ram_cell[    9819] = 32'hf8326222;
    ram_cell[    9820] = 32'h4784d076;
    ram_cell[    9821] = 32'hd5494af3;
    ram_cell[    9822] = 32'h395f8c73;
    ram_cell[    9823] = 32'he0c0b3a8;
    ram_cell[    9824] = 32'hcd8c69cc;
    ram_cell[    9825] = 32'h773ce949;
    ram_cell[    9826] = 32'h6815eae1;
    ram_cell[    9827] = 32'h9894fbf4;
    ram_cell[    9828] = 32'h1de6741b;
    ram_cell[    9829] = 32'h6e162a49;
    ram_cell[    9830] = 32'h3921e178;
    ram_cell[    9831] = 32'h158c3430;
    ram_cell[    9832] = 32'h866c471f;
    ram_cell[    9833] = 32'h07ce72bf;
    ram_cell[    9834] = 32'h23799eb4;
    ram_cell[    9835] = 32'h93772282;
    ram_cell[    9836] = 32'h6df1c98f;
    ram_cell[    9837] = 32'h3c5a81c4;
    ram_cell[    9838] = 32'he64d4596;
    ram_cell[    9839] = 32'h4cc985ca;
    ram_cell[    9840] = 32'hdba1ea15;
    ram_cell[    9841] = 32'hdb9881ae;
    ram_cell[    9842] = 32'h72168d68;
    ram_cell[    9843] = 32'h4b3f5a89;
    ram_cell[    9844] = 32'hfec67072;
    ram_cell[    9845] = 32'h9b723b03;
    ram_cell[    9846] = 32'h64beba31;
    ram_cell[    9847] = 32'h65751648;
    ram_cell[    9848] = 32'h7a9ab5ad;
    ram_cell[    9849] = 32'hf046d1c0;
    ram_cell[    9850] = 32'h2f7dfd58;
    ram_cell[    9851] = 32'h62ad5f5d;
    ram_cell[    9852] = 32'h33a67986;
    ram_cell[    9853] = 32'he6876089;
    ram_cell[    9854] = 32'h806b385a;
    ram_cell[    9855] = 32'h7a891da3;
    ram_cell[    9856] = 32'hdbb8a6db;
    ram_cell[    9857] = 32'hce7f5ef2;
    ram_cell[    9858] = 32'h322073f1;
    ram_cell[    9859] = 32'h4c724008;
    ram_cell[    9860] = 32'h42bda9e0;
    ram_cell[    9861] = 32'h8229d5f1;
    ram_cell[    9862] = 32'h358b6732;
    ram_cell[    9863] = 32'ha1f511f7;
    ram_cell[    9864] = 32'h50be582e;
    ram_cell[    9865] = 32'h7dedfbb4;
    ram_cell[    9866] = 32'he0ddd20c;
    ram_cell[    9867] = 32'ha8587b36;
    ram_cell[    9868] = 32'ha59a7e1c;
    ram_cell[    9869] = 32'hb5aae576;
    ram_cell[    9870] = 32'h55834b0e;
    ram_cell[    9871] = 32'h5d4cde18;
    ram_cell[    9872] = 32'hb587c7fd;
    ram_cell[    9873] = 32'h515d2231;
    ram_cell[    9874] = 32'h942ccb87;
    ram_cell[    9875] = 32'hc12d5550;
    ram_cell[    9876] = 32'hd3498d2e;
    ram_cell[    9877] = 32'h95fde0c6;
    ram_cell[    9878] = 32'heac7b532;
    ram_cell[    9879] = 32'h5421b466;
    ram_cell[    9880] = 32'he3979fc9;
    ram_cell[    9881] = 32'hcda3ff2e;
    ram_cell[    9882] = 32'h0a889cad;
    ram_cell[    9883] = 32'h6dbe9a10;
    ram_cell[    9884] = 32'hb6e721b3;
    ram_cell[    9885] = 32'ha2f35cba;
    ram_cell[    9886] = 32'h72ae4800;
    ram_cell[    9887] = 32'hb84a0c05;
    ram_cell[    9888] = 32'hdea69a3d;
    ram_cell[    9889] = 32'hebe521d1;
    ram_cell[    9890] = 32'hf871db4d;
    ram_cell[    9891] = 32'h968a454b;
    ram_cell[    9892] = 32'h00713caf;
    ram_cell[    9893] = 32'h294c5a5a;
    ram_cell[    9894] = 32'hc1f7f32e;
    ram_cell[    9895] = 32'hcacc1982;
    ram_cell[    9896] = 32'hf6c4615b;
    ram_cell[    9897] = 32'h95264bb5;
    ram_cell[    9898] = 32'h39f37efc;
    ram_cell[    9899] = 32'h2b2b8449;
    ram_cell[    9900] = 32'h1af436e4;
    ram_cell[    9901] = 32'h481dd2bc;
    ram_cell[    9902] = 32'ha78d0aef;
    ram_cell[    9903] = 32'h48deedc0;
    ram_cell[    9904] = 32'he768e433;
    ram_cell[    9905] = 32'hfc491fdf;
    ram_cell[    9906] = 32'hd7591ce7;
    ram_cell[    9907] = 32'hc6a0818f;
    ram_cell[    9908] = 32'h3622e006;
    ram_cell[    9909] = 32'hf63e78b2;
    ram_cell[    9910] = 32'h750645a1;
    ram_cell[    9911] = 32'hb8bed53e;
    ram_cell[    9912] = 32'hd733db1b;
    ram_cell[    9913] = 32'h97759161;
    ram_cell[    9914] = 32'hfea18f07;
    ram_cell[    9915] = 32'h9faf4d19;
    ram_cell[    9916] = 32'h7bd30305;
    ram_cell[    9917] = 32'h9c7c901e;
    ram_cell[    9918] = 32'h3e1bb336;
    ram_cell[    9919] = 32'hb2c7a2e3;
    ram_cell[    9920] = 32'h27ba7df9;
    ram_cell[    9921] = 32'h1e10f76c;
    ram_cell[    9922] = 32'h3fe931e2;
    ram_cell[    9923] = 32'h0ce7c346;
    ram_cell[    9924] = 32'h22f8359b;
    ram_cell[    9925] = 32'hc65f2dc1;
    ram_cell[    9926] = 32'ha6322eca;
    ram_cell[    9927] = 32'h82bcaa91;
    ram_cell[    9928] = 32'hf6807149;
    ram_cell[    9929] = 32'hc8b9b212;
    ram_cell[    9930] = 32'h42d79f37;
    ram_cell[    9931] = 32'h75cbfc3e;
    ram_cell[    9932] = 32'h152daff2;
    ram_cell[    9933] = 32'h34cd9f9e;
    ram_cell[    9934] = 32'hcfe2ffe5;
    ram_cell[    9935] = 32'h4b329d21;
    ram_cell[    9936] = 32'h8b88022b;
    ram_cell[    9937] = 32'h9e4192c9;
    ram_cell[    9938] = 32'h4e46471a;
    ram_cell[    9939] = 32'hb5ba0f84;
    ram_cell[    9940] = 32'h6edf82a9;
    ram_cell[    9941] = 32'hb293cff2;
    ram_cell[    9942] = 32'h648fc80e;
    ram_cell[    9943] = 32'h3b6dfca7;
    ram_cell[    9944] = 32'h3d7d45c3;
    ram_cell[    9945] = 32'h40964358;
    ram_cell[    9946] = 32'h8f37c3dd;
    ram_cell[    9947] = 32'h12007866;
    ram_cell[    9948] = 32'h924525ca;
    ram_cell[    9949] = 32'hcc5eff60;
    ram_cell[    9950] = 32'had35d692;
    ram_cell[    9951] = 32'hd52811d7;
    ram_cell[    9952] = 32'h17f446e8;
    ram_cell[    9953] = 32'h9bc3d263;
    ram_cell[    9954] = 32'h96ad99d3;
    ram_cell[    9955] = 32'h57e7c460;
    ram_cell[    9956] = 32'h67def303;
    ram_cell[    9957] = 32'h2399e22c;
    ram_cell[    9958] = 32'hf7738115;
    ram_cell[    9959] = 32'h46826dfc;
    ram_cell[    9960] = 32'hccd4fb97;
    ram_cell[    9961] = 32'hfa34def3;
    ram_cell[    9962] = 32'h91fab340;
    ram_cell[    9963] = 32'h9fece138;
    ram_cell[    9964] = 32'h077304ff;
    ram_cell[    9965] = 32'h0988c2fc;
    ram_cell[    9966] = 32'h28caa7d6;
    ram_cell[    9967] = 32'hb490cbe2;
    ram_cell[    9968] = 32'h9d129805;
    ram_cell[    9969] = 32'h284cf3a7;
    ram_cell[    9970] = 32'h32541687;
    ram_cell[    9971] = 32'h2546b1cc;
    ram_cell[    9972] = 32'hfe6173ef;
    ram_cell[    9973] = 32'h7e7ce638;
    ram_cell[    9974] = 32'h2bac0246;
    ram_cell[    9975] = 32'hbaedd34f;
    ram_cell[    9976] = 32'h30b248e2;
    ram_cell[    9977] = 32'h607bfa5f;
    ram_cell[    9978] = 32'h04bf5dad;
    ram_cell[    9979] = 32'h140277f3;
    ram_cell[    9980] = 32'h9219a8d0;
    ram_cell[    9981] = 32'hf89627d7;
    ram_cell[    9982] = 32'h25361244;
    ram_cell[    9983] = 32'h3afda4b2;
    ram_cell[    9984] = 32'h4ede0edb;
    ram_cell[    9985] = 32'hb51d5d3e;
    ram_cell[    9986] = 32'h84ef7d80;
    ram_cell[    9987] = 32'h783e8288;
    ram_cell[    9988] = 32'hc75d7afd;
    ram_cell[    9989] = 32'h5d439c65;
    ram_cell[    9990] = 32'h3e6d30ca;
    ram_cell[    9991] = 32'h1550c172;
    ram_cell[    9992] = 32'h1d5a670e;
    ram_cell[    9993] = 32'h6e20032e;
    ram_cell[    9994] = 32'h21a92f45;
    ram_cell[    9995] = 32'h9f123cc5;
    ram_cell[    9996] = 32'h7efa915d;
    ram_cell[    9997] = 32'hd07ede0b;
    ram_cell[    9998] = 32'hd593eeec;
    ram_cell[    9999] = 32'h0ae5e5c6;
    ram_cell[   10000] = 32'hfdf001e5;
    ram_cell[   10001] = 32'h2656f640;
    ram_cell[   10002] = 32'h98c43aae;
    ram_cell[   10003] = 32'h2d7cd2a1;
    ram_cell[   10004] = 32'hb8ca71ab;
    ram_cell[   10005] = 32'h661af9ae;
    ram_cell[   10006] = 32'h15a77d9b;
    ram_cell[   10007] = 32'h39683a30;
    ram_cell[   10008] = 32'hdfcff3a5;
    ram_cell[   10009] = 32'hc7b6012d;
    ram_cell[   10010] = 32'h4e3e1a77;
    ram_cell[   10011] = 32'hd21e2df1;
    ram_cell[   10012] = 32'hcaa06446;
    ram_cell[   10013] = 32'hd4c6004f;
    ram_cell[   10014] = 32'h1600c849;
    ram_cell[   10015] = 32'hbd298d0a;
    ram_cell[   10016] = 32'hc68fe5f0;
    ram_cell[   10017] = 32'hc020a7a0;
    ram_cell[   10018] = 32'h55709b32;
    ram_cell[   10019] = 32'hf252ae26;
    ram_cell[   10020] = 32'h7e84fb1a;
    ram_cell[   10021] = 32'h194810d3;
    ram_cell[   10022] = 32'h80d9b60a;
    ram_cell[   10023] = 32'hcce1be41;
    ram_cell[   10024] = 32'h7efb5f39;
    ram_cell[   10025] = 32'h24068e5f;
    ram_cell[   10026] = 32'he7e2f640;
    ram_cell[   10027] = 32'h403c73b5;
    ram_cell[   10028] = 32'h25f6d8de;
    ram_cell[   10029] = 32'h773aa6b6;
    ram_cell[   10030] = 32'h49a51de2;
    ram_cell[   10031] = 32'hb84e3a28;
    ram_cell[   10032] = 32'hea0741ff;
    ram_cell[   10033] = 32'h8a1b03ab;
    ram_cell[   10034] = 32'heb9ab4f6;
    ram_cell[   10035] = 32'h68467a83;
    ram_cell[   10036] = 32'h9fd28515;
    ram_cell[   10037] = 32'h5a2f46fe;
    ram_cell[   10038] = 32'h60d02ee9;
    ram_cell[   10039] = 32'h4b6e4d25;
    ram_cell[   10040] = 32'h97e0dd72;
    ram_cell[   10041] = 32'h1ae9b5aa;
    ram_cell[   10042] = 32'hd968b50d;
    ram_cell[   10043] = 32'hd34cebb4;
    ram_cell[   10044] = 32'hccfc451b;
    ram_cell[   10045] = 32'h427cd1ff;
    ram_cell[   10046] = 32'h26e8d717;
    ram_cell[   10047] = 32'h3d08f397;
    ram_cell[   10048] = 32'hc7748d8f;
    ram_cell[   10049] = 32'h4307e9cf;
    ram_cell[   10050] = 32'h11b88ada;
    ram_cell[   10051] = 32'h4d679d18;
    ram_cell[   10052] = 32'h9e269668;
    ram_cell[   10053] = 32'h0a41a5c9;
    ram_cell[   10054] = 32'h447c62ac;
    ram_cell[   10055] = 32'h7fb08806;
    ram_cell[   10056] = 32'h5a081494;
    ram_cell[   10057] = 32'h887981d0;
    ram_cell[   10058] = 32'hdf7d34e8;
    ram_cell[   10059] = 32'h05bfced1;
    ram_cell[   10060] = 32'h786fde7d;
    ram_cell[   10061] = 32'h30993b4a;
    ram_cell[   10062] = 32'hc043267e;
    ram_cell[   10063] = 32'h2bc0ffb0;
    ram_cell[   10064] = 32'h242f976d;
    ram_cell[   10065] = 32'h93890e9c;
    ram_cell[   10066] = 32'h09c661ea;
    ram_cell[   10067] = 32'h7a391787;
    ram_cell[   10068] = 32'h3a3962a6;
    ram_cell[   10069] = 32'hf6cdf4a3;
    ram_cell[   10070] = 32'hd605b5bd;
    ram_cell[   10071] = 32'hf0856343;
    ram_cell[   10072] = 32'ha045a272;
    ram_cell[   10073] = 32'h7a816c05;
    ram_cell[   10074] = 32'ha74fa02b;
    ram_cell[   10075] = 32'hf0f7f9de;
    ram_cell[   10076] = 32'h63498438;
    ram_cell[   10077] = 32'h50abbd0b;
    ram_cell[   10078] = 32'h04763f79;
    ram_cell[   10079] = 32'hfb97666d;
    ram_cell[   10080] = 32'h64ac74be;
    ram_cell[   10081] = 32'h00560576;
    ram_cell[   10082] = 32'hf5d2f229;
    ram_cell[   10083] = 32'hc23b498b;
    ram_cell[   10084] = 32'h52b8adf0;
    ram_cell[   10085] = 32'h0f0e478b;
    ram_cell[   10086] = 32'hf3d80bb9;
    ram_cell[   10087] = 32'ha1361846;
    ram_cell[   10088] = 32'hb0ebcc3e;
    ram_cell[   10089] = 32'hd8bfb0bb;
    ram_cell[   10090] = 32'h4fa4a55b;
    ram_cell[   10091] = 32'h45841621;
    ram_cell[   10092] = 32'h0ef7fecb;
    ram_cell[   10093] = 32'h61f031fc;
    ram_cell[   10094] = 32'hfd0752ac;
    ram_cell[   10095] = 32'hd7778cbd;
    ram_cell[   10096] = 32'h4e3d9bcb;
    ram_cell[   10097] = 32'h6d40e109;
    ram_cell[   10098] = 32'h75795edd;
    ram_cell[   10099] = 32'h49699765;
    ram_cell[   10100] = 32'h0003fbbb;
    ram_cell[   10101] = 32'h80116dbb;
    ram_cell[   10102] = 32'h9bcb7962;
    ram_cell[   10103] = 32'hf55a00ee;
    ram_cell[   10104] = 32'h44153614;
    ram_cell[   10105] = 32'h37eee76a;
    ram_cell[   10106] = 32'hd0f76a91;
    ram_cell[   10107] = 32'h2d651523;
    ram_cell[   10108] = 32'h4e57a5f1;
    ram_cell[   10109] = 32'h16b2d10f;
    ram_cell[   10110] = 32'h69799104;
    ram_cell[   10111] = 32'hdb1911b6;
    ram_cell[   10112] = 32'h87117f27;
    ram_cell[   10113] = 32'h7b96379e;
    ram_cell[   10114] = 32'h30e691ca;
    ram_cell[   10115] = 32'h050929f6;
    ram_cell[   10116] = 32'h8b4f2289;
    ram_cell[   10117] = 32'h0d2ef9ff;
    ram_cell[   10118] = 32'hb663d620;
    ram_cell[   10119] = 32'h6771689a;
    ram_cell[   10120] = 32'ha7864d33;
    ram_cell[   10121] = 32'hf47281e2;
    ram_cell[   10122] = 32'ha71a1d05;
    ram_cell[   10123] = 32'hef618af5;
    ram_cell[   10124] = 32'hfc237c37;
    ram_cell[   10125] = 32'hf172e060;
    ram_cell[   10126] = 32'hae6ae314;
    ram_cell[   10127] = 32'h09fd3a10;
    ram_cell[   10128] = 32'h6f572cce;
    ram_cell[   10129] = 32'hbc0e52bf;
    ram_cell[   10130] = 32'h9cfbed2b;
    ram_cell[   10131] = 32'hee86bcf1;
    ram_cell[   10132] = 32'h165f123a;
    ram_cell[   10133] = 32'h9f8edcc1;
    ram_cell[   10134] = 32'hcbbb3406;
    ram_cell[   10135] = 32'hb0609269;
    ram_cell[   10136] = 32'hb56b155d;
    ram_cell[   10137] = 32'hc1313474;
    ram_cell[   10138] = 32'h8230cb74;
    ram_cell[   10139] = 32'h8f2c45e8;
    ram_cell[   10140] = 32'h8321e847;
    ram_cell[   10141] = 32'hefe16bfa;
    ram_cell[   10142] = 32'h12a53077;
    ram_cell[   10143] = 32'h255e5564;
    ram_cell[   10144] = 32'h86c72cbd;
    ram_cell[   10145] = 32'h535f0218;
    ram_cell[   10146] = 32'he0cef8ae;
    ram_cell[   10147] = 32'h29ad2e94;
    ram_cell[   10148] = 32'h01f44be1;
    ram_cell[   10149] = 32'ha9e060e1;
    ram_cell[   10150] = 32'h0408540c;
    ram_cell[   10151] = 32'h61634f1f;
    ram_cell[   10152] = 32'h71c3d743;
    ram_cell[   10153] = 32'h6bd19b3a;
    ram_cell[   10154] = 32'hb4de80d7;
    ram_cell[   10155] = 32'h439c7402;
    ram_cell[   10156] = 32'h75efaee7;
    ram_cell[   10157] = 32'hffa268b0;
    ram_cell[   10158] = 32'had0f6664;
    ram_cell[   10159] = 32'hf53e6da9;
    ram_cell[   10160] = 32'h5648c1ca;
    ram_cell[   10161] = 32'he73a99bb;
    ram_cell[   10162] = 32'h7d9121aa;
    ram_cell[   10163] = 32'h0cc89d6b;
    ram_cell[   10164] = 32'hf210b99e;
    ram_cell[   10165] = 32'h0901669d;
    ram_cell[   10166] = 32'h9daa3b41;
    ram_cell[   10167] = 32'h740042e1;
    ram_cell[   10168] = 32'he24aff73;
    ram_cell[   10169] = 32'h8410869d;
    ram_cell[   10170] = 32'hde7520f1;
    ram_cell[   10171] = 32'hde37beef;
    ram_cell[   10172] = 32'h89cd732a;
    ram_cell[   10173] = 32'h9ad8a88f;
    ram_cell[   10174] = 32'h90812133;
    ram_cell[   10175] = 32'hecfb02b2;
    ram_cell[   10176] = 32'h677383fe;
    ram_cell[   10177] = 32'heb9b0e92;
    ram_cell[   10178] = 32'h984afd01;
    ram_cell[   10179] = 32'hc5678b1f;
    ram_cell[   10180] = 32'hba3b108a;
    ram_cell[   10181] = 32'h96fca7fd;
    ram_cell[   10182] = 32'h75e515f6;
    ram_cell[   10183] = 32'heaf63332;
    ram_cell[   10184] = 32'hc7eefde8;
    ram_cell[   10185] = 32'hbe1527fd;
    ram_cell[   10186] = 32'h6c5c0ce6;
    ram_cell[   10187] = 32'h0f221fde;
    ram_cell[   10188] = 32'h052dcd8c;
    ram_cell[   10189] = 32'h061089e7;
    ram_cell[   10190] = 32'h928e5ad2;
    ram_cell[   10191] = 32'h1018c1bb;
    ram_cell[   10192] = 32'h9d782569;
    ram_cell[   10193] = 32'h140d4e2e;
    ram_cell[   10194] = 32'hf705a3a3;
    ram_cell[   10195] = 32'hc2a0f6b9;
    ram_cell[   10196] = 32'hf2c557e1;
    ram_cell[   10197] = 32'h4131f5aa;
    ram_cell[   10198] = 32'hb0c33f4d;
    ram_cell[   10199] = 32'h595a3123;
    ram_cell[   10200] = 32'h62a5779a;
    ram_cell[   10201] = 32'h50311f8f;
    ram_cell[   10202] = 32'h9d6b86b8;
    ram_cell[   10203] = 32'hbc2820d0;
    ram_cell[   10204] = 32'h1053d2c7;
    ram_cell[   10205] = 32'hdffff776;
    ram_cell[   10206] = 32'hd81ecc6b;
    ram_cell[   10207] = 32'hc9607367;
    ram_cell[   10208] = 32'h546aa972;
    ram_cell[   10209] = 32'he99b35d5;
    ram_cell[   10210] = 32'h900f23c2;
    ram_cell[   10211] = 32'h6d7076e9;
    ram_cell[   10212] = 32'haaa9f5d1;
    ram_cell[   10213] = 32'he21ed30c;
    ram_cell[   10214] = 32'h86d5738d;
    ram_cell[   10215] = 32'he9717ea1;
    ram_cell[   10216] = 32'h852117cc;
    ram_cell[   10217] = 32'h64ee050b;
    ram_cell[   10218] = 32'hf9c28adb;
    ram_cell[   10219] = 32'hb58e8ee2;
    ram_cell[   10220] = 32'h68ab901d;
    ram_cell[   10221] = 32'h26221667;
    ram_cell[   10222] = 32'h82317f44;
    ram_cell[   10223] = 32'ha20a8968;
    ram_cell[   10224] = 32'h4b453f23;
    ram_cell[   10225] = 32'ha8add019;
    ram_cell[   10226] = 32'h7917b8c5;
    ram_cell[   10227] = 32'h6f7f7b9a;
    ram_cell[   10228] = 32'h95b20d5b;
    ram_cell[   10229] = 32'h7c528189;
    ram_cell[   10230] = 32'h028f78ed;
    ram_cell[   10231] = 32'h20c09dd6;
    ram_cell[   10232] = 32'h9d35895b;
    ram_cell[   10233] = 32'h57b04f2d;
    ram_cell[   10234] = 32'h376e9f87;
    ram_cell[   10235] = 32'hebfc614f;
    ram_cell[   10236] = 32'hf6afb068;
    ram_cell[   10237] = 32'h5f03aebf;
    ram_cell[   10238] = 32'hf358a1d9;
    ram_cell[   10239] = 32'h6cfd1ddb;
    ram_cell[   10240] = 32'ha41301db;
    ram_cell[   10241] = 32'h919696d3;
    ram_cell[   10242] = 32'hcb88b7f2;
    ram_cell[   10243] = 32'h4a3adc8b;
    ram_cell[   10244] = 32'hbf46dfbc;
    ram_cell[   10245] = 32'haf2e58c3;
    ram_cell[   10246] = 32'ha6a3aa6c;
    ram_cell[   10247] = 32'hbad2b940;
    ram_cell[   10248] = 32'hea1ba4cd;
    ram_cell[   10249] = 32'h2bb7ef2e;
    ram_cell[   10250] = 32'hee1d2fb2;
    ram_cell[   10251] = 32'hef29bc0f;
    ram_cell[   10252] = 32'h66307a1a;
    ram_cell[   10253] = 32'h184eacfc;
    ram_cell[   10254] = 32'h179a8736;
    ram_cell[   10255] = 32'he39ff642;
    ram_cell[   10256] = 32'h78cccca0;
    ram_cell[   10257] = 32'h75370f50;
    ram_cell[   10258] = 32'hbcfe0003;
    ram_cell[   10259] = 32'h8601fd07;
    ram_cell[   10260] = 32'h552a5b9a;
    ram_cell[   10261] = 32'h3e4d543c;
    ram_cell[   10262] = 32'h90316826;
    ram_cell[   10263] = 32'hcabefa22;
    ram_cell[   10264] = 32'hd3b24d3a;
    ram_cell[   10265] = 32'h4fc3a1fc;
    ram_cell[   10266] = 32'h15fb2f29;
    ram_cell[   10267] = 32'hdfcbd9b5;
    ram_cell[   10268] = 32'h0edd05f2;
    ram_cell[   10269] = 32'h07f5c85d;
    ram_cell[   10270] = 32'hcc8360a0;
    ram_cell[   10271] = 32'h88d8055f;
    ram_cell[   10272] = 32'h06462e53;
    ram_cell[   10273] = 32'hc4c9e4f0;
    ram_cell[   10274] = 32'he97822f5;
    ram_cell[   10275] = 32'hea3bf54e;
    ram_cell[   10276] = 32'hf9351c9d;
    ram_cell[   10277] = 32'h90ac1157;
    ram_cell[   10278] = 32'h5d173d5c;
    ram_cell[   10279] = 32'h17ed7ca3;
    ram_cell[   10280] = 32'hef74b287;
    ram_cell[   10281] = 32'hcb2326e4;
    ram_cell[   10282] = 32'hcda107b5;
    ram_cell[   10283] = 32'h94fed6ee;
    ram_cell[   10284] = 32'h7f239e45;
    ram_cell[   10285] = 32'h8df35465;
    ram_cell[   10286] = 32'h37c53892;
    ram_cell[   10287] = 32'h60784e3d;
    ram_cell[   10288] = 32'h3cc4b041;
    ram_cell[   10289] = 32'haef635ae;
    ram_cell[   10290] = 32'h8a14d3cb;
    ram_cell[   10291] = 32'he0e2bfc9;
    ram_cell[   10292] = 32'h4ed6c1b2;
    ram_cell[   10293] = 32'h95ab0ac7;
    ram_cell[   10294] = 32'h91475284;
    ram_cell[   10295] = 32'h5e4c4ab4;
    ram_cell[   10296] = 32'ha0067f95;
    ram_cell[   10297] = 32'h8c1fdd16;
    ram_cell[   10298] = 32'h379f69ec;
    ram_cell[   10299] = 32'hd249808e;
    ram_cell[   10300] = 32'h96933450;
    ram_cell[   10301] = 32'hc34b0c0c;
    ram_cell[   10302] = 32'hfc152553;
    ram_cell[   10303] = 32'h574ec973;
    ram_cell[   10304] = 32'hef7b9bab;
    ram_cell[   10305] = 32'h724bce89;
    ram_cell[   10306] = 32'h13683c49;
    ram_cell[   10307] = 32'hd2b0cbee;
    ram_cell[   10308] = 32'h76d3a953;
    ram_cell[   10309] = 32'he073f254;
    ram_cell[   10310] = 32'h086b271f;
    ram_cell[   10311] = 32'h3ab30c74;
    ram_cell[   10312] = 32'h75afbca7;
    ram_cell[   10313] = 32'hcbfebfe1;
    ram_cell[   10314] = 32'hba9efe6d;
    ram_cell[   10315] = 32'h734da9f8;
    ram_cell[   10316] = 32'h51ab4ec7;
    ram_cell[   10317] = 32'hdfd69579;
    ram_cell[   10318] = 32'h002fa56a;
    ram_cell[   10319] = 32'h9287cef4;
    ram_cell[   10320] = 32'h3a9660c2;
    ram_cell[   10321] = 32'h87bd24bb;
    ram_cell[   10322] = 32'h22a24d66;
    ram_cell[   10323] = 32'h83ab9e1a;
    ram_cell[   10324] = 32'h7173a1b9;
    ram_cell[   10325] = 32'h169984fc;
    ram_cell[   10326] = 32'hb4aa2309;
    ram_cell[   10327] = 32'hfc0f0bf0;
    ram_cell[   10328] = 32'hb8f67348;
    ram_cell[   10329] = 32'hbe6d9470;
    ram_cell[   10330] = 32'h614cd1e9;
    ram_cell[   10331] = 32'h32d8e2c5;
    ram_cell[   10332] = 32'h5e481ff9;
    ram_cell[   10333] = 32'h7973b8b5;
    ram_cell[   10334] = 32'h094fc563;
    ram_cell[   10335] = 32'h0f97d404;
    ram_cell[   10336] = 32'h09845e77;
    ram_cell[   10337] = 32'h90d72835;
    ram_cell[   10338] = 32'had097072;
    ram_cell[   10339] = 32'h86bdb09f;
    ram_cell[   10340] = 32'hc203b2ee;
    ram_cell[   10341] = 32'h6061c27d;
    ram_cell[   10342] = 32'h0a3693ad;
    ram_cell[   10343] = 32'h9f32d23a;
    ram_cell[   10344] = 32'h4101fc1c;
    ram_cell[   10345] = 32'h2ad658a1;
    ram_cell[   10346] = 32'h9fe0bbdf;
    ram_cell[   10347] = 32'h2e482d46;
    ram_cell[   10348] = 32'h4ab7c9e4;
    ram_cell[   10349] = 32'hfd43b63a;
    ram_cell[   10350] = 32'h2cd753c6;
    ram_cell[   10351] = 32'h49181510;
    ram_cell[   10352] = 32'hf6300c1e;
    ram_cell[   10353] = 32'h3c3d4a8f;
    ram_cell[   10354] = 32'h71a87519;
    ram_cell[   10355] = 32'hdbed2cf2;
    ram_cell[   10356] = 32'hae859aea;
    ram_cell[   10357] = 32'hc12702d3;
    ram_cell[   10358] = 32'hd8c3647f;
    ram_cell[   10359] = 32'hfe0a5372;
    ram_cell[   10360] = 32'h63e2d9cc;
    ram_cell[   10361] = 32'h0c085768;
    ram_cell[   10362] = 32'hab52148d;
    ram_cell[   10363] = 32'hadd1b665;
    ram_cell[   10364] = 32'hb6d5a986;
    ram_cell[   10365] = 32'h4da1773a;
    ram_cell[   10366] = 32'h773012c6;
    ram_cell[   10367] = 32'ha1ce27c8;
    ram_cell[   10368] = 32'hc81197d4;
    ram_cell[   10369] = 32'h98023977;
    ram_cell[   10370] = 32'ha08f11d9;
    ram_cell[   10371] = 32'ha01d10ef;
    ram_cell[   10372] = 32'h6ba98f96;
    ram_cell[   10373] = 32'h96ad52dd;
    ram_cell[   10374] = 32'h01ebeb5e;
    ram_cell[   10375] = 32'h129becc4;
    ram_cell[   10376] = 32'h600bb7ea;
    ram_cell[   10377] = 32'h38e65423;
    ram_cell[   10378] = 32'h11ab16ba;
    ram_cell[   10379] = 32'h183d84a7;
    ram_cell[   10380] = 32'h07e6de5c;
    ram_cell[   10381] = 32'h5bf58004;
    ram_cell[   10382] = 32'h86ef1877;
    ram_cell[   10383] = 32'h1e9c03fe;
    ram_cell[   10384] = 32'h441de94a;
    ram_cell[   10385] = 32'ha151ed1f;
    ram_cell[   10386] = 32'h7bc2d542;
    ram_cell[   10387] = 32'h7255f0f5;
    ram_cell[   10388] = 32'h4eb99dd8;
    ram_cell[   10389] = 32'hff21f4d4;
    ram_cell[   10390] = 32'h1e0e37c3;
    ram_cell[   10391] = 32'h67503fb2;
    ram_cell[   10392] = 32'he919415d;
    ram_cell[   10393] = 32'h29825e57;
    ram_cell[   10394] = 32'h6d23d7e8;
    ram_cell[   10395] = 32'hb8730eac;
    ram_cell[   10396] = 32'h57507ee6;
    ram_cell[   10397] = 32'h60d47e16;
    ram_cell[   10398] = 32'h012d3fa7;
    ram_cell[   10399] = 32'ha9ffe361;
    ram_cell[   10400] = 32'h478ca932;
    ram_cell[   10401] = 32'hdcf6cb2d;
    ram_cell[   10402] = 32'h3569ad8f;
    ram_cell[   10403] = 32'h5086fb3b;
    ram_cell[   10404] = 32'haaadc921;
    ram_cell[   10405] = 32'h77650cf3;
    ram_cell[   10406] = 32'hcffc50d0;
    ram_cell[   10407] = 32'he5cdf1dc;
    ram_cell[   10408] = 32'h7834985d;
    ram_cell[   10409] = 32'h2b0366c7;
    ram_cell[   10410] = 32'h6c021f76;
    ram_cell[   10411] = 32'h0c001174;
    ram_cell[   10412] = 32'ha56c5597;
    ram_cell[   10413] = 32'h009ec06d;
    ram_cell[   10414] = 32'h4da1bf98;
    ram_cell[   10415] = 32'h6addd92b;
    ram_cell[   10416] = 32'h4d2e5d73;
    ram_cell[   10417] = 32'h43801d7e;
    ram_cell[   10418] = 32'h7bda35e8;
    ram_cell[   10419] = 32'h49ec0628;
    ram_cell[   10420] = 32'hf6507788;
    ram_cell[   10421] = 32'h48f3bfb7;
    ram_cell[   10422] = 32'h3751594d;
    ram_cell[   10423] = 32'h39069fc8;
    ram_cell[   10424] = 32'h6b57d333;
    ram_cell[   10425] = 32'h345ff5b2;
    ram_cell[   10426] = 32'hfb57abb8;
    ram_cell[   10427] = 32'h7803e861;
    ram_cell[   10428] = 32'hef534821;
    ram_cell[   10429] = 32'hf07beaf8;
    ram_cell[   10430] = 32'ha980423f;
    ram_cell[   10431] = 32'hf298c6e3;
    ram_cell[   10432] = 32'ha1c749c6;
    ram_cell[   10433] = 32'h0020ef58;
    ram_cell[   10434] = 32'hf1512be9;
    ram_cell[   10435] = 32'h3dc6574e;
    ram_cell[   10436] = 32'hcd134629;
    ram_cell[   10437] = 32'hef980ece;
    ram_cell[   10438] = 32'h90382f8d;
    ram_cell[   10439] = 32'h937baa3a;
    ram_cell[   10440] = 32'h935c2dbb;
    ram_cell[   10441] = 32'h56848535;
    ram_cell[   10442] = 32'h62ad94dc;
    ram_cell[   10443] = 32'h764fe7b6;
    ram_cell[   10444] = 32'hbc41d6c1;
    ram_cell[   10445] = 32'h8236877d;
    ram_cell[   10446] = 32'h78a8ec07;
    ram_cell[   10447] = 32'hd4767ec0;
    ram_cell[   10448] = 32'h3d495983;
    ram_cell[   10449] = 32'h2c4c59d3;
    ram_cell[   10450] = 32'h0732449e;
    ram_cell[   10451] = 32'h76dce183;
    ram_cell[   10452] = 32'h049c8c7c;
    ram_cell[   10453] = 32'hc9039be4;
    ram_cell[   10454] = 32'hb1adcaf9;
    ram_cell[   10455] = 32'h035d2c5e;
    ram_cell[   10456] = 32'h689b2116;
    ram_cell[   10457] = 32'h31509053;
    ram_cell[   10458] = 32'h4b0c1358;
    ram_cell[   10459] = 32'hbf07cfdd;
    ram_cell[   10460] = 32'h1fe8f3c6;
    ram_cell[   10461] = 32'h435535a5;
    ram_cell[   10462] = 32'h01dd3191;
    ram_cell[   10463] = 32'h6ba63f8f;
    ram_cell[   10464] = 32'hf5448a82;
    ram_cell[   10465] = 32'h2b4558e9;
    ram_cell[   10466] = 32'h9cdbc0db;
    ram_cell[   10467] = 32'h55b44c5e;
    ram_cell[   10468] = 32'h81e40346;
    ram_cell[   10469] = 32'h19130fa5;
    ram_cell[   10470] = 32'h26bdb830;
    ram_cell[   10471] = 32'hd4e78d46;
    ram_cell[   10472] = 32'h300a779c;
    ram_cell[   10473] = 32'h1d4a3c0b;
    ram_cell[   10474] = 32'hf95c4344;
    ram_cell[   10475] = 32'h04aa2296;
    ram_cell[   10476] = 32'hd6f16a43;
    ram_cell[   10477] = 32'hf8d53244;
    ram_cell[   10478] = 32'hd4f1de80;
    ram_cell[   10479] = 32'h0250f016;
    ram_cell[   10480] = 32'h2c709228;
    ram_cell[   10481] = 32'h50fcca1e;
    ram_cell[   10482] = 32'h1202dd40;
    ram_cell[   10483] = 32'he647e0a1;
    ram_cell[   10484] = 32'h2f97f75b;
    ram_cell[   10485] = 32'h3856386a;
    ram_cell[   10486] = 32'h2cc3c249;
    ram_cell[   10487] = 32'h86b2ef4b;
    ram_cell[   10488] = 32'h4701ccbb;
    ram_cell[   10489] = 32'hc234114f;
    ram_cell[   10490] = 32'h0fd1d374;
    ram_cell[   10491] = 32'h432cfec5;
    ram_cell[   10492] = 32'h2bd22c7c;
    ram_cell[   10493] = 32'h72ad84f4;
    ram_cell[   10494] = 32'h3ecfbe1b;
    ram_cell[   10495] = 32'h77c8d48a;
    ram_cell[   10496] = 32'hf61b6f15;
    ram_cell[   10497] = 32'h6b51c933;
    ram_cell[   10498] = 32'hc898dfb3;
    ram_cell[   10499] = 32'h038a9b20;
    ram_cell[   10500] = 32'hbb62b2ba;
    ram_cell[   10501] = 32'h0a0d2585;
    ram_cell[   10502] = 32'had719efc;
    ram_cell[   10503] = 32'h7a883d71;
    ram_cell[   10504] = 32'hed3ba2a1;
    ram_cell[   10505] = 32'hcb6cb76e;
    ram_cell[   10506] = 32'hfb62c713;
    ram_cell[   10507] = 32'h9afd69d3;
    ram_cell[   10508] = 32'hb38e20c7;
    ram_cell[   10509] = 32'h9422e2ee;
    ram_cell[   10510] = 32'hf3140cff;
    ram_cell[   10511] = 32'ha0617927;
    ram_cell[   10512] = 32'h76d3b5c7;
    ram_cell[   10513] = 32'hc6a0da65;
    ram_cell[   10514] = 32'ha1376959;
    ram_cell[   10515] = 32'hd783f95d;
    ram_cell[   10516] = 32'h374fb5ff;
    ram_cell[   10517] = 32'h950d404b;
    ram_cell[   10518] = 32'h5f2b8683;
    ram_cell[   10519] = 32'hbf5c720a;
    ram_cell[   10520] = 32'h019393e5;
    ram_cell[   10521] = 32'he5a30b08;
    ram_cell[   10522] = 32'h4aebf25d;
    ram_cell[   10523] = 32'h7db627dd;
    ram_cell[   10524] = 32'hec3df82b;
    ram_cell[   10525] = 32'hab991b51;
    ram_cell[   10526] = 32'h6e621149;
    ram_cell[   10527] = 32'hb7cd8313;
    ram_cell[   10528] = 32'h6d9b1439;
    ram_cell[   10529] = 32'h9960a5a5;
    ram_cell[   10530] = 32'hab3fce30;
    ram_cell[   10531] = 32'h4b5bed2f;
    ram_cell[   10532] = 32'h96398efe;
    ram_cell[   10533] = 32'hc5e04c78;
    ram_cell[   10534] = 32'h31b95084;
    ram_cell[   10535] = 32'h16ee6511;
    ram_cell[   10536] = 32'h7a68e32e;
    ram_cell[   10537] = 32'h7ae4014d;
    ram_cell[   10538] = 32'h17b94ecb;
    ram_cell[   10539] = 32'h6974ae29;
    ram_cell[   10540] = 32'hb7e272cf;
    ram_cell[   10541] = 32'h24e941b0;
    ram_cell[   10542] = 32'h51a8c69e;
    ram_cell[   10543] = 32'h83ce04de;
    ram_cell[   10544] = 32'h46a81dbc;
    ram_cell[   10545] = 32'hfa4a3df0;
    ram_cell[   10546] = 32'heda89f58;
    ram_cell[   10547] = 32'h8ea07aae;
    ram_cell[   10548] = 32'heb84f9b6;
    ram_cell[   10549] = 32'h0ee5f3af;
    ram_cell[   10550] = 32'hbf5677ac;
    ram_cell[   10551] = 32'h421986c6;
    ram_cell[   10552] = 32'h3aedeeec;
    ram_cell[   10553] = 32'he1e3c7fc;
    ram_cell[   10554] = 32'ha53a405e;
    ram_cell[   10555] = 32'hd78375a7;
    ram_cell[   10556] = 32'hfc026327;
    ram_cell[   10557] = 32'h85fa6765;
    ram_cell[   10558] = 32'h24627e3f;
    ram_cell[   10559] = 32'h2fcfd799;
    ram_cell[   10560] = 32'h89082d06;
    ram_cell[   10561] = 32'h49f79a71;
    ram_cell[   10562] = 32'h62949ebb;
    ram_cell[   10563] = 32'hc1d85558;
    ram_cell[   10564] = 32'hfd826f87;
    ram_cell[   10565] = 32'h7390ff7b;
    ram_cell[   10566] = 32'h0af89f24;
    ram_cell[   10567] = 32'ha21d3b8b;
    ram_cell[   10568] = 32'hfe6a037e;
    ram_cell[   10569] = 32'hc3212d67;
    ram_cell[   10570] = 32'h8a6d4268;
    ram_cell[   10571] = 32'h420c92f0;
    ram_cell[   10572] = 32'hd801a705;
    ram_cell[   10573] = 32'hf29d7b29;
    ram_cell[   10574] = 32'h1bc13e5d;
    ram_cell[   10575] = 32'h0c678e39;
    ram_cell[   10576] = 32'h93f641a8;
    ram_cell[   10577] = 32'h221c5b7c;
    ram_cell[   10578] = 32'h69078201;
    ram_cell[   10579] = 32'hc56c735b;
    ram_cell[   10580] = 32'h779307f7;
    ram_cell[   10581] = 32'h879bd21b;
    ram_cell[   10582] = 32'h55101e2e;
    ram_cell[   10583] = 32'h8a8b92e3;
    ram_cell[   10584] = 32'h36fdde3a;
    ram_cell[   10585] = 32'h9f6a7334;
    ram_cell[   10586] = 32'ha44219a4;
    ram_cell[   10587] = 32'h564fef39;
    ram_cell[   10588] = 32'ha99387be;
    ram_cell[   10589] = 32'h48dfb1c6;
    ram_cell[   10590] = 32'h9bfea407;
    ram_cell[   10591] = 32'hc3100b53;
    ram_cell[   10592] = 32'h4c7f9186;
    ram_cell[   10593] = 32'h0d0f711d;
    ram_cell[   10594] = 32'hb33631f7;
    ram_cell[   10595] = 32'h59e5338b;
    ram_cell[   10596] = 32'heddbc5ee;
    ram_cell[   10597] = 32'h4d740eb6;
    ram_cell[   10598] = 32'he862cafa;
    ram_cell[   10599] = 32'h2abcf44b;
    ram_cell[   10600] = 32'he184cfad;
    ram_cell[   10601] = 32'h7ddd322c;
    ram_cell[   10602] = 32'h7989d31e;
    ram_cell[   10603] = 32'hbc9dfb8b;
    ram_cell[   10604] = 32'h42b6bc94;
    ram_cell[   10605] = 32'hcf254518;
    ram_cell[   10606] = 32'h6a6e69be;
    ram_cell[   10607] = 32'hab6b9da3;
    ram_cell[   10608] = 32'h15660aef;
    ram_cell[   10609] = 32'h640f89e2;
    ram_cell[   10610] = 32'hbb4954e3;
    ram_cell[   10611] = 32'h332623c7;
    ram_cell[   10612] = 32'he4c2a838;
    ram_cell[   10613] = 32'ha4323b34;
    ram_cell[   10614] = 32'hb4dfcf2e;
    ram_cell[   10615] = 32'hde875c24;
    ram_cell[   10616] = 32'h8170f36b;
    ram_cell[   10617] = 32'h70cb6fe4;
    ram_cell[   10618] = 32'h4e6fecd6;
    ram_cell[   10619] = 32'h4f3040ec;
    ram_cell[   10620] = 32'h2aac98f0;
    ram_cell[   10621] = 32'hd965ecc6;
    ram_cell[   10622] = 32'hb4cb4b29;
    ram_cell[   10623] = 32'h754c6d2a;
    ram_cell[   10624] = 32'hf99814f4;
    ram_cell[   10625] = 32'h49203ac9;
    ram_cell[   10626] = 32'h11625220;
    ram_cell[   10627] = 32'hfe318b99;
    ram_cell[   10628] = 32'h58ecdd8e;
    ram_cell[   10629] = 32'heaf8ddcd;
    ram_cell[   10630] = 32'h2d3cf5a9;
    ram_cell[   10631] = 32'h5b06160f;
    ram_cell[   10632] = 32'hf8117846;
    ram_cell[   10633] = 32'h90162ae8;
    ram_cell[   10634] = 32'h2bdcc60a;
    ram_cell[   10635] = 32'h99c998c5;
    ram_cell[   10636] = 32'h1a3f412a;
    ram_cell[   10637] = 32'h299ffe17;
    ram_cell[   10638] = 32'h10f07635;
    ram_cell[   10639] = 32'h09ded08f;
    ram_cell[   10640] = 32'hfdb684f6;
    ram_cell[   10641] = 32'h862c5279;
    ram_cell[   10642] = 32'hfd657c33;
    ram_cell[   10643] = 32'h14bc0260;
    ram_cell[   10644] = 32'hb02823ae;
    ram_cell[   10645] = 32'h3ce5e61c;
    ram_cell[   10646] = 32'h5f1053f0;
    ram_cell[   10647] = 32'h22f90670;
    ram_cell[   10648] = 32'h02f21251;
    ram_cell[   10649] = 32'ha371b5af;
    ram_cell[   10650] = 32'hf2b25a22;
    ram_cell[   10651] = 32'h51d45ccb;
    ram_cell[   10652] = 32'h50a3a906;
    ram_cell[   10653] = 32'h152fc3fe;
    ram_cell[   10654] = 32'hcd88dcf7;
    ram_cell[   10655] = 32'heb0362f0;
    ram_cell[   10656] = 32'hed682668;
    ram_cell[   10657] = 32'hbbbd662c;
    ram_cell[   10658] = 32'h9554121b;
    ram_cell[   10659] = 32'h01da2cbe;
    ram_cell[   10660] = 32'h499e2f40;
    ram_cell[   10661] = 32'h9a6ebf6c;
    ram_cell[   10662] = 32'h9ce77c3e;
    ram_cell[   10663] = 32'h9e33347b;
    ram_cell[   10664] = 32'ha36de8ee;
    ram_cell[   10665] = 32'h45db469b;
    ram_cell[   10666] = 32'h5807172f;
    ram_cell[   10667] = 32'h07f09764;
    ram_cell[   10668] = 32'h9c948b9f;
    ram_cell[   10669] = 32'h1238bbf8;
    ram_cell[   10670] = 32'h2f5b93db;
    ram_cell[   10671] = 32'hb962615b;
    ram_cell[   10672] = 32'h05c9e530;
    ram_cell[   10673] = 32'h13810a9d;
    ram_cell[   10674] = 32'h2330f093;
    ram_cell[   10675] = 32'hd03b220f;
    ram_cell[   10676] = 32'h533e1db5;
    ram_cell[   10677] = 32'h73fe2972;
    ram_cell[   10678] = 32'h294f31b5;
    ram_cell[   10679] = 32'hb8518782;
    ram_cell[   10680] = 32'h3a39a27e;
    ram_cell[   10681] = 32'h0c0a5974;
    ram_cell[   10682] = 32'h468b6965;
    ram_cell[   10683] = 32'hb2b6479a;
    ram_cell[   10684] = 32'hd56697c5;
    ram_cell[   10685] = 32'ha25e9a43;
    ram_cell[   10686] = 32'h330d371e;
    ram_cell[   10687] = 32'hed63e014;
    ram_cell[   10688] = 32'hfeb22a09;
    ram_cell[   10689] = 32'h82d59606;
    ram_cell[   10690] = 32'hd5296514;
    ram_cell[   10691] = 32'h2d3e51fb;
    ram_cell[   10692] = 32'h83447576;
    ram_cell[   10693] = 32'h19874fb6;
    ram_cell[   10694] = 32'hc2db852e;
    ram_cell[   10695] = 32'h8444b957;
    ram_cell[   10696] = 32'h73031e6d;
    ram_cell[   10697] = 32'ha0dfa837;
    ram_cell[   10698] = 32'h08bb5894;
    ram_cell[   10699] = 32'hf04dd593;
    ram_cell[   10700] = 32'h4677c297;
    ram_cell[   10701] = 32'hc1c724be;
    ram_cell[   10702] = 32'h1cf314f9;
    ram_cell[   10703] = 32'h35d796d1;
    ram_cell[   10704] = 32'ha76acdf2;
    ram_cell[   10705] = 32'h881b8e5b;
    ram_cell[   10706] = 32'he119b474;
    ram_cell[   10707] = 32'ha9311678;
    ram_cell[   10708] = 32'ha7adc22e;
    ram_cell[   10709] = 32'hb14bc494;
    ram_cell[   10710] = 32'h0e4edd0f;
    ram_cell[   10711] = 32'h0fa82173;
    ram_cell[   10712] = 32'hb0154eb0;
    ram_cell[   10713] = 32'h6635433e;
    ram_cell[   10714] = 32'hddac1a81;
    ram_cell[   10715] = 32'ha10df639;
    ram_cell[   10716] = 32'hceb13948;
    ram_cell[   10717] = 32'hf50bdfa7;
    ram_cell[   10718] = 32'h35297c0a;
    ram_cell[   10719] = 32'ha8dedf01;
    ram_cell[   10720] = 32'ha9db1e25;
    ram_cell[   10721] = 32'h51ee3962;
    ram_cell[   10722] = 32'hb163349f;
    ram_cell[   10723] = 32'ha575021b;
    ram_cell[   10724] = 32'h788e10ae;
    ram_cell[   10725] = 32'h5036a86b;
    ram_cell[   10726] = 32'h4e163001;
    ram_cell[   10727] = 32'h7e20572c;
    ram_cell[   10728] = 32'h81a5de2b;
    ram_cell[   10729] = 32'hd8dbdb03;
    ram_cell[   10730] = 32'hc4e51bf6;
    ram_cell[   10731] = 32'hec0dc40d;
    ram_cell[   10732] = 32'h41c4918d;
    ram_cell[   10733] = 32'h3595cc7c;
    ram_cell[   10734] = 32'h153bd50a;
    ram_cell[   10735] = 32'hc611a860;
    ram_cell[   10736] = 32'hba511a7b;
    ram_cell[   10737] = 32'hb2176bfe;
    ram_cell[   10738] = 32'h58e6d718;
    ram_cell[   10739] = 32'h0950ee57;
    ram_cell[   10740] = 32'h46828c1a;
    ram_cell[   10741] = 32'h0a96b7cd;
    ram_cell[   10742] = 32'h2f1a8e3a;
    ram_cell[   10743] = 32'hdef8580c;
    ram_cell[   10744] = 32'h22bcb925;
    ram_cell[   10745] = 32'he5aa40b5;
    ram_cell[   10746] = 32'h4797efcd;
    ram_cell[   10747] = 32'hbc959edf;
    ram_cell[   10748] = 32'hc902392f;
    ram_cell[   10749] = 32'h305756c5;
    ram_cell[   10750] = 32'h8dd04bc2;
    ram_cell[   10751] = 32'h81ee339e;
    ram_cell[   10752] = 32'he93a11ec;
    ram_cell[   10753] = 32'h089f41a9;
    ram_cell[   10754] = 32'h170a7c27;
    ram_cell[   10755] = 32'h60b03657;
    ram_cell[   10756] = 32'hc96a5a07;
    ram_cell[   10757] = 32'hedc9792e;
    ram_cell[   10758] = 32'h170c4524;
    ram_cell[   10759] = 32'h554df0b4;
    ram_cell[   10760] = 32'hbf54ef4d;
    ram_cell[   10761] = 32'h327db181;
    ram_cell[   10762] = 32'hcca3ae32;
    ram_cell[   10763] = 32'hf4bd52e1;
    ram_cell[   10764] = 32'h7b381d31;
    ram_cell[   10765] = 32'h008d1931;
    ram_cell[   10766] = 32'h9e1f4925;
    ram_cell[   10767] = 32'h41f79e00;
    ram_cell[   10768] = 32'hdf2097f2;
    ram_cell[   10769] = 32'h0fc820da;
    ram_cell[   10770] = 32'hd92fe1ff;
    ram_cell[   10771] = 32'h323231df;
    ram_cell[   10772] = 32'h4b06b165;
    ram_cell[   10773] = 32'hcc62b928;
    ram_cell[   10774] = 32'hf610abd1;
    ram_cell[   10775] = 32'he55d2fab;
    ram_cell[   10776] = 32'hafaa7eb8;
    ram_cell[   10777] = 32'h0cbf30ec;
    ram_cell[   10778] = 32'h19187337;
    ram_cell[   10779] = 32'h0d9583f4;
    ram_cell[   10780] = 32'h7558cd8d;
    ram_cell[   10781] = 32'hbf35d49f;
    ram_cell[   10782] = 32'h6da6fd41;
    ram_cell[   10783] = 32'h5ce9ba57;
    ram_cell[   10784] = 32'h413b5618;
    ram_cell[   10785] = 32'hcb9f2e26;
    ram_cell[   10786] = 32'haa7b525c;
    ram_cell[   10787] = 32'hccf23dbe;
    ram_cell[   10788] = 32'h1725ae41;
    ram_cell[   10789] = 32'he2c327be;
    ram_cell[   10790] = 32'hed368e30;
    ram_cell[   10791] = 32'h17b98bb1;
    ram_cell[   10792] = 32'h762c3a05;
    ram_cell[   10793] = 32'hbd097c4c;
    ram_cell[   10794] = 32'h53223a32;
    ram_cell[   10795] = 32'h7e92ab3e;
    ram_cell[   10796] = 32'h60001596;
    ram_cell[   10797] = 32'hfa6d6e93;
    ram_cell[   10798] = 32'he9d93909;
    ram_cell[   10799] = 32'hafc3ac60;
    ram_cell[   10800] = 32'h895f2e9b;
    ram_cell[   10801] = 32'h8a2c1312;
    ram_cell[   10802] = 32'hc6fa0ca5;
    ram_cell[   10803] = 32'hdd6e2269;
    ram_cell[   10804] = 32'h7adc9579;
    ram_cell[   10805] = 32'he53a2248;
    ram_cell[   10806] = 32'h04440663;
    ram_cell[   10807] = 32'he3aec96f;
    ram_cell[   10808] = 32'hdf0f52ab;
    ram_cell[   10809] = 32'ha78f906f;
    ram_cell[   10810] = 32'hab9da2b6;
    ram_cell[   10811] = 32'h51f59c0d;
    ram_cell[   10812] = 32'hf1e14fd8;
    ram_cell[   10813] = 32'hcfce29dd;
    ram_cell[   10814] = 32'hdace3de9;
    ram_cell[   10815] = 32'h2e990b5b;
    ram_cell[   10816] = 32'hd837107e;
    ram_cell[   10817] = 32'hfb905e66;
    ram_cell[   10818] = 32'h278e7974;
    ram_cell[   10819] = 32'h46f767a5;
    ram_cell[   10820] = 32'h065f6860;
    ram_cell[   10821] = 32'h3680003b;
    ram_cell[   10822] = 32'h5f5b9181;
    ram_cell[   10823] = 32'h71c96e1b;
    ram_cell[   10824] = 32'hb2d3b53b;
    ram_cell[   10825] = 32'hc2f2375d;
    ram_cell[   10826] = 32'h1951de36;
    ram_cell[   10827] = 32'h3832adf7;
    ram_cell[   10828] = 32'h855f1522;
    ram_cell[   10829] = 32'h7a333078;
    ram_cell[   10830] = 32'h8c5f7a7c;
    ram_cell[   10831] = 32'h57ed5d16;
    ram_cell[   10832] = 32'hbae41879;
    ram_cell[   10833] = 32'h0d39b442;
    ram_cell[   10834] = 32'h4045dc07;
    ram_cell[   10835] = 32'haef800cd;
    ram_cell[   10836] = 32'hd02c9605;
    ram_cell[   10837] = 32'hcff84811;
    ram_cell[   10838] = 32'h65bc56e8;
    ram_cell[   10839] = 32'h58a26416;
    ram_cell[   10840] = 32'h58cfa4bd;
    ram_cell[   10841] = 32'hdcc05f30;
    ram_cell[   10842] = 32'haf1b12fe;
    ram_cell[   10843] = 32'hf77ba205;
    ram_cell[   10844] = 32'h697a80f7;
    ram_cell[   10845] = 32'h8f54be5d;
    ram_cell[   10846] = 32'h1a260cd3;
    ram_cell[   10847] = 32'h3cf0e9f3;
    ram_cell[   10848] = 32'hb0cea261;
    ram_cell[   10849] = 32'h6eed8d0e;
    ram_cell[   10850] = 32'haf8b312b;
    ram_cell[   10851] = 32'h8fe65669;
    ram_cell[   10852] = 32'h5e1ce929;
    ram_cell[   10853] = 32'h6e8dee5d;
    ram_cell[   10854] = 32'hc7dc3de3;
    ram_cell[   10855] = 32'h1611a2ff;
    ram_cell[   10856] = 32'h08bf8029;
    ram_cell[   10857] = 32'h06afbe40;
    ram_cell[   10858] = 32'h9a7a3aab;
    ram_cell[   10859] = 32'h7cd4843a;
    ram_cell[   10860] = 32'hf472ba3b;
    ram_cell[   10861] = 32'h972db61d;
    ram_cell[   10862] = 32'h914cb93d;
    ram_cell[   10863] = 32'h0c42d0ec;
    ram_cell[   10864] = 32'h15a1bc25;
    ram_cell[   10865] = 32'h7084dc8b;
    ram_cell[   10866] = 32'h248013d6;
    ram_cell[   10867] = 32'h72032d52;
    ram_cell[   10868] = 32'h011ffbb4;
    ram_cell[   10869] = 32'h30ef1877;
    ram_cell[   10870] = 32'hc94c2c25;
    ram_cell[   10871] = 32'hda7594d9;
    ram_cell[   10872] = 32'h4aad9341;
    ram_cell[   10873] = 32'hb0883bdc;
    ram_cell[   10874] = 32'h6e6aee2a;
    ram_cell[   10875] = 32'h3b125fa7;
    ram_cell[   10876] = 32'h3ce13018;
    ram_cell[   10877] = 32'h1d8dcd4f;
    ram_cell[   10878] = 32'heb9912a0;
    ram_cell[   10879] = 32'hb4053c4f;
    ram_cell[   10880] = 32'h40def8c7;
    ram_cell[   10881] = 32'h9ea62910;
    ram_cell[   10882] = 32'h4383ed4c;
    ram_cell[   10883] = 32'h8eb6e935;
    ram_cell[   10884] = 32'hd2d31cfa;
    ram_cell[   10885] = 32'h0746cc06;
    ram_cell[   10886] = 32'h2fd7d1db;
    ram_cell[   10887] = 32'h7e03da71;
    ram_cell[   10888] = 32'h59cd06c8;
    ram_cell[   10889] = 32'hccbdfc9b;
    ram_cell[   10890] = 32'h86c23378;
    ram_cell[   10891] = 32'h5e982b0b;
    ram_cell[   10892] = 32'h033b3540;
    ram_cell[   10893] = 32'h278940d0;
    ram_cell[   10894] = 32'h7d6d9b0e;
    ram_cell[   10895] = 32'ha0e4e502;
    ram_cell[   10896] = 32'h11994451;
    ram_cell[   10897] = 32'h49aa65df;
    ram_cell[   10898] = 32'h42cb726b;
    ram_cell[   10899] = 32'hbba84817;
    ram_cell[   10900] = 32'hcd1e4348;
    ram_cell[   10901] = 32'h470c4242;
    ram_cell[   10902] = 32'heecdcabb;
    ram_cell[   10903] = 32'hbf58d145;
    ram_cell[   10904] = 32'hfbf2da86;
    ram_cell[   10905] = 32'h20c8ef67;
    ram_cell[   10906] = 32'hbb372756;
    ram_cell[   10907] = 32'h31fdfb12;
    ram_cell[   10908] = 32'h7c918b18;
    ram_cell[   10909] = 32'hce09a860;
    ram_cell[   10910] = 32'h7991bced;
    ram_cell[   10911] = 32'h25d67d82;
    ram_cell[   10912] = 32'hf9110ab5;
    ram_cell[   10913] = 32'hc3e5558e;
    ram_cell[   10914] = 32'h4120dd02;
    ram_cell[   10915] = 32'hf86a87db;
    ram_cell[   10916] = 32'hc2f6bd83;
    ram_cell[   10917] = 32'hd65fbf33;
    ram_cell[   10918] = 32'heebfb010;
    ram_cell[   10919] = 32'h990f015e;
    ram_cell[   10920] = 32'h2fe07a2c;
    ram_cell[   10921] = 32'h00dbd1df;
    ram_cell[   10922] = 32'h589005fe;
    ram_cell[   10923] = 32'he485a032;
    ram_cell[   10924] = 32'hb218cd98;
    ram_cell[   10925] = 32'h20264bbc;
    ram_cell[   10926] = 32'h5a37f77c;
    ram_cell[   10927] = 32'h081a4330;
    ram_cell[   10928] = 32'hc7072325;
    ram_cell[   10929] = 32'h77472eb0;
    ram_cell[   10930] = 32'hf2e7bf66;
    ram_cell[   10931] = 32'h877416ec;
    ram_cell[   10932] = 32'h7f4d6b8a;
    ram_cell[   10933] = 32'h7287cf8e;
    ram_cell[   10934] = 32'h91462ffc;
    ram_cell[   10935] = 32'ha92f6ee6;
    ram_cell[   10936] = 32'h474c59c2;
    ram_cell[   10937] = 32'hcba8a302;
    ram_cell[   10938] = 32'h0e1ae045;
    ram_cell[   10939] = 32'h70b4a393;
    ram_cell[   10940] = 32'h797bd9dd;
    ram_cell[   10941] = 32'hcde1d676;
    ram_cell[   10942] = 32'hc1dd9649;
    ram_cell[   10943] = 32'hdab74089;
    ram_cell[   10944] = 32'h1432936b;
    ram_cell[   10945] = 32'h51228e3d;
    ram_cell[   10946] = 32'h70a6b83a;
    ram_cell[   10947] = 32'hf4eea56c;
    ram_cell[   10948] = 32'h5b0c924b;
    ram_cell[   10949] = 32'h73c5f750;
    ram_cell[   10950] = 32'h520fe6e6;
    ram_cell[   10951] = 32'h3d6549de;
    ram_cell[   10952] = 32'h75083624;
    ram_cell[   10953] = 32'hdc4501a0;
    ram_cell[   10954] = 32'h67f54161;
    ram_cell[   10955] = 32'hb74b3fd7;
    ram_cell[   10956] = 32'h1902928f;
    ram_cell[   10957] = 32'h8cfd4993;
    ram_cell[   10958] = 32'h90f28170;
    ram_cell[   10959] = 32'ha44c10c8;
    ram_cell[   10960] = 32'h42f481d7;
    ram_cell[   10961] = 32'h8cbda308;
    ram_cell[   10962] = 32'h377c9de2;
    ram_cell[   10963] = 32'h2df7c36e;
    ram_cell[   10964] = 32'h4a770b83;
    ram_cell[   10965] = 32'h4bf4899f;
    ram_cell[   10966] = 32'hcd8d160c;
    ram_cell[   10967] = 32'h6846a3bf;
    ram_cell[   10968] = 32'h8125dd6a;
    ram_cell[   10969] = 32'h02931297;
    ram_cell[   10970] = 32'hec2c86d7;
    ram_cell[   10971] = 32'hdcd4c00d;
    ram_cell[   10972] = 32'hbf385972;
    ram_cell[   10973] = 32'hb81e061e;
    ram_cell[   10974] = 32'h4e1a99d9;
    ram_cell[   10975] = 32'h82dd4e1d;
    ram_cell[   10976] = 32'h6bc36550;
    ram_cell[   10977] = 32'h21fe5f32;
    ram_cell[   10978] = 32'h4ad07546;
    ram_cell[   10979] = 32'h3c74654f;
    ram_cell[   10980] = 32'h7efe143e;
    ram_cell[   10981] = 32'h803da5a3;
    ram_cell[   10982] = 32'h8bdf048d;
    ram_cell[   10983] = 32'h1c4693ae;
    ram_cell[   10984] = 32'hfa79c954;
    ram_cell[   10985] = 32'h40b982ed;
    ram_cell[   10986] = 32'h36021656;
    ram_cell[   10987] = 32'ha1e227f3;
    ram_cell[   10988] = 32'h4589dba9;
    ram_cell[   10989] = 32'h2f892158;
    ram_cell[   10990] = 32'h5c1c8392;
    ram_cell[   10991] = 32'hd070692c;
    ram_cell[   10992] = 32'h65642bfd;
    ram_cell[   10993] = 32'h2ea36e7a;
    ram_cell[   10994] = 32'hc3d7e0db;
    ram_cell[   10995] = 32'h4f2c97c8;
    ram_cell[   10996] = 32'hc52c51ba;
    ram_cell[   10997] = 32'h85aeba8d;
    ram_cell[   10998] = 32'h4b74d266;
    ram_cell[   10999] = 32'h3ceb6960;
    ram_cell[   11000] = 32'h196e6896;
    ram_cell[   11001] = 32'h1818b2ee;
    ram_cell[   11002] = 32'h9d1398a0;
    ram_cell[   11003] = 32'had3e9c40;
    ram_cell[   11004] = 32'hf0cee14a;
    ram_cell[   11005] = 32'hbf45205f;
    ram_cell[   11006] = 32'hed995a7e;
    ram_cell[   11007] = 32'h2d49fa17;
    ram_cell[   11008] = 32'h43b98db7;
    ram_cell[   11009] = 32'h36db01ac;
    ram_cell[   11010] = 32'h065b9fb9;
    ram_cell[   11011] = 32'h67318f35;
    ram_cell[   11012] = 32'hb64c84f7;
    ram_cell[   11013] = 32'h0071a8ef;
    ram_cell[   11014] = 32'hcc50d719;
    ram_cell[   11015] = 32'hf9992761;
    ram_cell[   11016] = 32'he499e2e0;
    ram_cell[   11017] = 32'h66dac089;
    ram_cell[   11018] = 32'h51884172;
    ram_cell[   11019] = 32'h8209f0e0;
    ram_cell[   11020] = 32'h5b8bb291;
    ram_cell[   11021] = 32'hb5a81e86;
    ram_cell[   11022] = 32'he51208ed;
    ram_cell[   11023] = 32'h23563f97;
    ram_cell[   11024] = 32'h2cca6b53;
    ram_cell[   11025] = 32'h6c057d6c;
    ram_cell[   11026] = 32'h91ae64cf;
    ram_cell[   11027] = 32'h68b5cbad;
    ram_cell[   11028] = 32'hf4601c29;
    ram_cell[   11029] = 32'h8d56259b;
    ram_cell[   11030] = 32'he38f0a7c;
    ram_cell[   11031] = 32'habd0cb34;
    ram_cell[   11032] = 32'he2c8d975;
    ram_cell[   11033] = 32'h62f7ff4c;
    ram_cell[   11034] = 32'h1017aa68;
    ram_cell[   11035] = 32'hb06eb1d8;
    ram_cell[   11036] = 32'h7dee2508;
    ram_cell[   11037] = 32'ha53c23c0;
    ram_cell[   11038] = 32'h27ab11fb;
    ram_cell[   11039] = 32'hcbbbd9e6;
    ram_cell[   11040] = 32'hf18c5d16;
    ram_cell[   11041] = 32'h7bab7e51;
    ram_cell[   11042] = 32'hc86c04fb;
    ram_cell[   11043] = 32'head3a94c;
    ram_cell[   11044] = 32'hf91f06e2;
    ram_cell[   11045] = 32'he552181c;
    ram_cell[   11046] = 32'h6706394f;
    ram_cell[   11047] = 32'h7e9d3d54;
    ram_cell[   11048] = 32'h68292bb3;
    ram_cell[   11049] = 32'hba9d2330;
    ram_cell[   11050] = 32'hcf85ab3e;
    ram_cell[   11051] = 32'hbfa052b4;
    ram_cell[   11052] = 32'hfae7b9ef;
    ram_cell[   11053] = 32'hd3b789d2;
    ram_cell[   11054] = 32'hc83d74af;
    ram_cell[   11055] = 32'h22f307b7;
    ram_cell[   11056] = 32'h09d5e7dc;
    ram_cell[   11057] = 32'ha0277182;
    ram_cell[   11058] = 32'hf9ff6d0f;
    ram_cell[   11059] = 32'h7ab337f9;
    ram_cell[   11060] = 32'h63c42bd9;
    ram_cell[   11061] = 32'h8d3c7a0c;
    ram_cell[   11062] = 32'hf23cdf77;
    ram_cell[   11063] = 32'he3529e34;
    ram_cell[   11064] = 32'h3fa9688c;
    ram_cell[   11065] = 32'h495804f0;
    ram_cell[   11066] = 32'h4ae79ea6;
    ram_cell[   11067] = 32'hee016989;
    ram_cell[   11068] = 32'h95cc1553;
    ram_cell[   11069] = 32'h15426e3c;
    ram_cell[   11070] = 32'h9d1a0151;
    ram_cell[   11071] = 32'h67be7910;
    ram_cell[   11072] = 32'ha69fde6f;
    ram_cell[   11073] = 32'h5e1846eb;
    ram_cell[   11074] = 32'h9a65a7a3;
    ram_cell[   11075] = 32'h006e8812;
    ram_cell[   11076] = 32'he5e0dfcd;
    ram_cell[   11077] = 32'h9f25b21d;
    ram_cell[   11078] = 32'h5bc3ed4e;
    ram_cell[   11079] = 32'hf29b71be;
    ram_cell[   11080] = 32'hc9741881;
    ram_cell[   11081] = 32'h101a0317;
    ram_cell[   11082] = 32'hf20b5d8a;
    ram_cell[   11083] = 32'hbebf2751;
    ram_cell[   11084] = 32'h3971e0bf;
    ram_cell[   11085] = 32'hcfeb08c4;
    ram_cell[   11086] = 32'h9b869dfb;
    ram_cell[   11087] = 32'hba448b49;
    ram_cell[   11088] = 32'he8bfbc2d;
    ram_cell[   11089] = 32'h067e1c52;
    ram_cell[   11090] = 32'h48a94061;
    ram_cell[   11091] = 32'h1d3d6c18;
    ram_cell[   11092] = 32'h91c06d1b;
    ram_cell[   11093] = 32'h67fb0aeb;
    ram_cell[   11094] = 32'hc9ac87b1;
    ram_cell[   11095] = 32'h52c69dbe;
    ram_cell[   11096] = 32'hd9f1cac0;
    ram_cell[   11097] = 32'hbc55833d;
    ram_cell[   11098] = 32'h985c3a0f;
    ram_cell[   11099] = 32'h6b677dcc;
    ram_cell[   11100] = 32'h4c7525ab;
    ram_cell[   11101] = 32'hd6cd08a2;
    ram_cell[   11102] = 32'h1e66066f;
    ram_cell[   11103] = 32'hbe700b8b;
    ram_cell[   11104] = 32'h8a8ccece;
    ram_cell[   11105] = 32'h50dbf9d2;
    ram_cell[   11106] = 32'h36b03ae9;
    ram_cell[   11107] = 32'h12fce86d;
    ram_cell[   11108] = 32'h2298668b;
    ram_cell[   11109] = 32'h464b800a;
    ram_cell[   11110] = 32'h4f1001a0;
    ram_cell[   11111] = 32'h03efda7a;
    ram_cell[   11112] = 32'h14d07e0d;
    ram_cell[   11113] = 32'h856de055;
    ram_cell[   11114] = 32'h58fae31e;
    ram_cell[   11115] = 32'h965f6fbe;
    ram_cell[   11116] = 32'h714b78d4;
    ram_cell[   11117] = 32'hce79762f;
    ram_cell[   11118] = 32'h49b089f3;
    ram_cell[   11119] = 32'h7ef839ec;
    ram_cell[   11120] = 32'h99f8d24f;
    ram_cell[   11121] = 32'h7a2f9c77;
    ram_cell[   11122] = 32'h98718c8d;
    ram_cell[   11123] = 32'h5d7984b9;
    ram_cell[   11124] = 32'hb45c60cb;
    ram_cell[   11125] = 32'h78ee2a8c;
    ram_cell[   11126] = 32'h64d9d926;
    ram_cell[   11127] = 32'h2f4f3249;
    ram_cell[   11128] = 32'h5a34ad6c;
    ram_cell[   11129] = 32'h9fbc7690;
    ram_cell[   11130] = 32'h08e9f540;
    ram_cell[   11131] = 32'h958b8fc5;
    ram_cell[   11132] = 32'hc9647999;
    ram_cell[   11133] = 32'hc52e64d6;
    ram_cell[   11134] = 32'hbe11f9b3;
    ram_cell[   11135] = 32'h3d663853;
    ram_cell[   11136] = 32'hf1da7380;
    ram_cell[   11137] = 32'h7a30e7ab;
    ram_cell[   11138] = 32'h86884d8e;
    ram_cell[   11139] = 32'hd3bf0430;
    ram_cell[   11140] = 32'h2a11f0b9;
    ram_cell[   11141] = 32'hc283356b;
    ram_cell[   11142] = 32'hbb1103dd;
    ram_cell[   11143] = 32'he7eaabca;
    ram_cell[   11144] = 32'h902fcab6;
    ram_cell[   11145] = 32'h7e49ae48;
    ram_cell[   11146] = 32'h1273e8b4;
    ram_cell[   11147] = 32'hd0ec07f6;
    ram_cell[   11148] = 32'hae29c9cf;
    ram_cell[   11149] = 32'hc9294273;
    ram_cell[   11150] = 32'h841fde67;
    ram_cell[   11151] = 32'hd1ad9dfb;
    ram_cell[   11152] = 32'h01a1bd37;
    ram_cell[   11153] = 32'hb58fecb0;
    ram_cell[   11154] = 32'hba29579d;
    ram_cell[   11155] = 32'h8a845ecb;
    ram_cell[   11156] = 32'h73d55d18;
    ram_cell[   11157] = 32'h5c6beb83;
    ram_cell[   11158] = 32'h1264c107;
    ram_cell[   11159] = 32'h3be274c1;
    ram_cell[   11160] = 32'h14d055f2;
    ram_cell[   11161] = 32'h4d38db72;
    ram_cell[   11162] = 32'h391e429d;
    ram_cell[   11163] = 32'hc7adc4ee;
    ram_cell[   11164] = 32'hff1072ed;
    ram_cell[   11165] = 32'hd99c4f88;
    ram_cell[   11166] = 32'hf945612b;
    ram_cell[   11167] = 32'h06a98fe5;
    ram_cell[   11168] = 32'hc6b8e30d;
    ram_cell[   11169] = 32'h7e0ecb72;
    ram_cell[   11170] = 32'hc501c0db;
    ram_cell[   11171] = 32'h54a40968;
    ram_cell[   11172] = 32'h5132148a;
    ram_cell[   11173] = 32'ha77ffb23;
    ram_cell[   11174] = 32'h3e53a3ca;
    ram_cell[   11175] = 32'hbea9418b;
    ram_cell[   11176] = 32'hc774bd96;
    ram_cell[   11177] = 32'h07d8d1db;
    ram_cell[   11178] = 32'he9e8b46b;
    ram_cell[   11179] = 32'h70022039;
    ram_cell[   11180] = 32'h551bbe71;
    ram_cell[   11181] = 32'h40d42548;
    ram_cell[   11182] = 32'hba6817f1;
    ram_cell[   11183] = 32'ha07babb3;
    ram_cell[   11184] = 32'h32bf3bc0;
    ram_cell[   11185] = 32'hd8a04153;
    ram_cell[   11186] = 32'h2cf9684b;
    ram_cell[   11187] = 32'hdda43be5;
    ram_cell[   11188] = 32'ha46d4ba7;
    ram_cell[   11189] = 32'hcc838bfa;
    ram_cell[   11190] = 32'h25867ef2;
    ram_cell[   11191] = 32'h0269bb6b;
    ram_cell[   11192] = 32'hc98f109b;
    ram_cell[   11193] = 32'h5ed48094;
    ram_cell[   11194] = 32'h88688620;
    ram_cell[   11195] = 32'haf7ac925;
    ram_cell[   11196] = 32'h1fadabae;
    ram_cell[   11197] = 32'h1584c9e6;
    ram_cell[   11198] = 32'h9d9afe4a;
    ram_cell[   11199] = 32'h3680c6ec;
    ram_cell[   11200] = 32'h67ec994e;
    ram_cell[   11201] = 32'h4f5a0521;
    ram_cell[   11202] = 32'h5615ef5c;
    ram_cell[   11203] = 32'hdf9fe85c;
    ram_cell[   11204] = 32'hc146fc58;
    ram_cell[   11205] = 32'h2b162731;
    ram_cell[   11206] = 32'h55ac0f7a;
    ram_cell[   11207] = 32'h3eebf321;
    ram_cell[   11208] = 32'h9ee764d0;
    ram_cell[   11209] = 32'h1d6e49d1;
    ram_cell[   11210] = 32'hef190f77;
    ram_cell[   11211] = 32'hf89afbdd;
    ram_cell[   11212] = 32'h35d7428c;
    ram_cell[   11213] = 32'h74f7b5b8;
    ram_cell[   11214] = 32'hb0b55537;
    ram_cell[   11215] = 32'h07581b64;
    ram_cell[   11216] = 32'h62964b53;
    ram_cell[   11217] = 32'hdae9a7e6;
    ram_cell[   11218] = 32'hb7f27b7d;
    ram_cell[   11219] = 32'h72bacb8d;
    ram_cell[   11220] = 32'h75aa269a;
    ram_cell[   11221] = 32'h6079afbe;
    ram_cell[   11222] = 32'h3dba8d36;
    ram_cell[   11223] = 32'h6993d508;
    ram_cell[   11224] = 32'hec77286a;
    ram_cell[   11225] = 32'h8f6ac62d;
    ram_cell[   11226] = 32'h14986df0;
    ram_cell[   11227] = 32'ha52e7270;
    ram_cell[   11228] = 32'h84cfea23;
    ram_cell[   11229] = 32'h693504a2;
    ram_cell[   11230] = 32'ha2cb2014;
    ram_cell[   11231] = 32'h9c5d32e7;
    ram_cell[   11232] = 32'hf06c40c4;
    ram_cell[   11233] = 32'h1fc939ae;
    ram_cell[   11234] = 32'h871a975b;
    ram_cell[   11235] = 32'hd9d95636;
    ram_cell[   11236] = 32'h6bfbf4e0;
    ram_cell[   11237] = 32'h500e56ea;
    ram_cell[   11238] = 32'hce7b41c8;
    ram_cell[   11239] = 32'h075090a9;
    ram_cell[   11240] = 32'hef4d197f;
    ram_cell[   11241] = 32'h043c913b;
    ram_cell[   11242] = 32'h6710b908;
    ram_cell[   11243] = 32'ha8b73835;
    ram_cell[   11244] = 32'hef85b1e5;
    ram_cell[   11245] = 32'h858e22a5;
    ram_cell[   11246] = 32'h2978ce07;
    ram_cell[   11247] = 32'he4b1fd29;
    ram_cell[   11248] = 32'h457d5002;
    ram_cell[   11249] = 32'h079771cb;
    ram_cell[   11250] = 32'ha9472068;
    ram_cell[   11251] = 32'h7a7e77a7;
    ram_cell[   11252] = 32'h3c70813b;
    ram_cell[   11253] = 32'h06a94e94;
    ram_cell[   11254] = 32'h672dc07d;
    ram_cell[   11255] = 32'h41ab625f;
    ram_cell[   11256] = 32'h33944e48;
    ram_cell[   11257] = 32'h7526a57d;
    ram_cell[   11258] = 32'h74d4c4da;
    ram_cell[   11259] = 32'heeca68b1;
    ram_cell[   11260] = 32'h8bfe9ccb;
    ram_cell[   11261] = 32'h17b3cbd5;
    ram_cell[   11262] = 32'hc8604a69;
    ram_cell[   11263] = 32'hd536b911;
    ram_cell[   11264] = 32'h12f909bb;
    ram_cell[   11265] = 32'h4191b866;
    ram_cell[   11266] = 32'h8872a905;
    ram_cell[   11267] = 32'hef0d6ae9;
    ram_cell[   11268] = 32'hfd0840a6;
    ram_cell[   11269] = 32'h9f633a26;
    ram_cell[   11270] = 32'h485d2573;
    ram_cell[   11271] = 32'h86f19ca0;
    ram_cell[   11272] = 32'ha559a30e;
    ram_cell[   11273] = 32'hf64088e2;
    ram_cell[   11274] = 32'h3f474d85;
    ram_cell[   11275] = 32'h51b0e4b4;
    ram_cell[   11276] = 32'h8b245a17;
    ram_cell[   11277] = 32'hf0a47d8d;
    ram_cell[   11278] = 32'h3e90069d;
    ram_cell[   11279] = 32'h2e341415;
    ram_cell[   11280] = 32'h3f4d4487;
    ram_cell[   11281] = 32'h7ae2d85c;
    ram_cell[   11282] = 32'h03cd3200;
    ram_cell[   11283] = 32'h023a8232;
    ram_cell[   11284] = 32'ha99bdeb8;
    ram_cell[   11285] = 32'h553fa9c9;
    ram_cell[   11286] = 32'h521ed91f;
    ram_cell[   11287] = 32'hf6ded80a;
    ram_cell[   11288] = 32'h1db3ea4c;
    ram_cell[   11289] = 32'hed8713db;
    ram_cell[   11290] = 32'h1702c950;
    ram_cell[   11291] = 32'h0584a201;
    ram_cell[   11292] = 32'h0a315c6d;
    ram_cell[   11293] = 32'h5bf676f1;
    ram_cell[   11294] = 32'h1579774b;
    ram_cell[   11295] = 32'hd80b3d6b;
    ram_cell[   11296] = 32'h831dd8f4;
    ram_cell[   11297] = 32'h8af2ab48;
    ram_cell[   11298] = 32'h9fd6a8ba;
    ram_cell[   11299] = 32'he407a01f;
    ram_cell[   11300] = 32'hfdf4e1f8;
    ram_cell[   11301] = 32'h4c932bd4;
    ram_cell[   11302] = 32'h298963a9;
    ram_cell[   11303] = 32'hc984edab;
    ram_cell[   11304] = 32'h054c5cf1;
    ram_cell[   11305] = 32'hd4d844e3;
    ram_cell[   11306] = 32'hc8c0202e;
    ram_cell[   11307] = 32'h05a8faea;
    ram_cell[   11308] = 32'h7cbfd883;
    ram_cell[   11309] = 32'hcc637d7e;
    ram_cell[   11310] = 32'h9695b011;
    ram_cell[   11311] = 32'h550538c6;
    ram_cell[   11312] = 32'hc7f4c021;
    ram_cell[   11313] = 32'h44a6a043;
    ram_cell[   11314] = 32'h9b8178b3;
    ram_cell[   11315] = 32'h11936ee6;
    ram_cell[   11316] = 32'h125ff14b;
    ram_cell[   11317] = 32'hf50af3e4;
    ram_cell[   11318] = 32'h49ad51d3;
    ram_cell[   11319] = 32'h8b272857;
    ram_cell[   11320] = 32'he1788a13;
    ram_cell[   11321] = 32'h4971d8cc;
    ram_cell[   11322] = 32'h8a8f22aa;
    ram_cell[   11323] = 32'h6922f091;
    ram_cell[   11324] = 32'h90667a95;
    ram_cell[   11325] = 32'h78f2aecd;
    ram_cell[   11326] = 32'hdb3d8e70;
    ram_cell[   11327] = 32'h5ec61075;
    ram_cell[   11328] = 32'hf3a6c0a8;
    ram_cell[   11329] = 32'h892d9a3e;
    ram_cell[   11330] = 32'h90e25b76;
    ram_cell[   11331] = 32'h25c915e3;
    ram_cell[   11332] = 32'h80b1ae72;
    ram_cell[   11333] = 32'h278583f7;
    ram_cell[   11334] = 32'hbe07915c;
    ram_cell[   11335] = 32'h441dbca7;
    ram_cell[   11336] = 32'h92ac504e;
    ram_cell[   11337] = 32'h997b3ba1;
    ram_cell[   11338] = 32'h9c8293b9;
    ram_cell[   11339] = 32'h1eb9ff4a;
    ram_cell[   11340] = 32'h863a39e6;
    ram_cell[   11341] = 32'h0420eb86;
    ram_cell[   11342] = 32'h491fe2d5;
    ram_cell[   11343] = 32'hffae3828;
    ram_cell[   11344] = 32'hd4e0dc08;
    ram_cell[   11345] = 32'hc8cd94bd;
    ram_cell[   11346] = 32'hf16a387d;
    ram_cell[   11347] = 32'h36a0eb61;
    ram_cell[   11348] = 32'h73f7d940;
    ram_cell[   11349] = 32'h301a9b09;
    ram_cell[   11350] = 32'h88b82296;
    ram_cell[   11351] = 32'h89440314;
    ram_cell[   11352] = 32'hdec3b64b;
    ram_cell[   11353] = 32'he525301b;
    ram_cell[   11354] = 32'he5522452;
    ram_cell[   11355] = 32'h01a1fc29;
    ram_cell[   11356] = 32'h95407c14;
    ram_cell[   11357] = 32'h5de70d3e;
    ram_cell[   11358] = 32'ha22fcf2f;
    ram_cell[   11359] = 32'hb8e3e034;
    ram_cell[   11360] = 32'h27be0e32;
    ram_cell[   11361] = 32'h9c4d3dcd;
    ram_cell[   11362] = 32'h7a841ad0;
    ram_cell[   11363] = 32'h7a52acce;
    ram_cell[   11364] = 32'hf681e236;
    ram_cell[   11365] = 32'h22db941b;
    ram_cell[   11366] = 32'h8321f735;
    ram_cell[   11367] = 32'h7f53dddf;
    ram_cell[   11368] = 32'ha52289f3;
    ram_cell[   11369] = 32'he7fa4833;
    ram_cell[   11370] = 32'h958058a5;
    ram_cell[   11371] = 32'h151a1d4e;
    ram_cell[   11372] = 32'hd548afbf;
    ram_cell[   11373] = 32'h887a572d;
    ram_cell[   11374] = 32'h4587848a;
    ram_cell[   11375] = 32'h14afee9b;
    ram_cell[   11376] = 32'he53d0712;
    ram_cell[   11377] = 32'hcf330138;
    ram_cell[   11378] = 32'h4af95d81;
    ram_cell[   11379] = 32'h6aaed525;
    ram_cell[   11380] = 32'h887a4f7f;
    ram_cell[   11381] = 32'h985a1b2f;
    ram_cell[   11382] = 32'hdb819487;
    ram_cell[   11383] = 32'h837a7020;
    ram_cell[   11384] = 32'h52a16ddb;
    ram_cell[   11385] = 32'h761cc6e1;
    ram_cell[   11386] = 32'h08c60a42;
    ram_cell[   11387] = 32'hd2fd5108;
    ram_cell[   11388] = 32'h1f702c01;
    ram_cell[   11389] = 32'h5105ca54;
    ram_cell[   11390] = 32'h2f579cc4;
    ram_cell[   11391] = 32'hce489b6c;
    ram_cell[   11392] = 32'h6ef92dca;
    ram_cell[   11393] = 32'h32652b9a;
    ram_cell[   11394] = 32'h9e29926c;
    ram_cell[   11395] = 32'h206b7dba;
    ram_cell[   11396] = 32'h6036c92d;
    ram_cell[   11397] = 32'hb2beded5;
    ram_cell[   11398] = 32'h10d5c3e8;
    ram_cell[   11399] = 32'h5eb8a7fc;
    ram_cell[   11400] = 32'hb0e84850;
    ram_cell[   11401] = 32'h66be08a9;
    ram_cell[   11402] = 32'h10bd5769;
    ram_cell[   11403] = 32'hac3197f9;
    ram_cell[   11404] = 32'h2316f7d5;
    ram_cell[   11405] = 32'hd82ae707;
    ram_cell[   11406] = 32'hd45591f5;
    ram_cell[   11407] = 32'h93d4723e;
    ram_cell[   11408] = 32'hd77912ac;
    ram_cell[   11409] = 32'hc155d6ba;
    ram_cell[   11410] = 32'h1fcdb962;
    ram_cell[   11411] = 32'h805415e8;
    ram_cell[   11412] = 32'hd6aad0fb;
    ram_cell[   11413] = 32'hc0c6d4be;
    ram_cell[   11414] = 32'h8f1b695c;
    ram_cell[   11415] = 32'h3420de36;
    ram_cell[   11416] = 32'h0e958365;
    ram_cell[   11417] = 32'h85f66a17;
    ram_cell[   11418] = 32'h2c52fdbc;
    ram_cell[   11419] = 32'hf728da39;
    ram_cell[   11420] = 32'h550a29b1;
    ram_cell[   11421] = 32'hf4f7682b;
    ram_cell[   11422] = 32'he993b1cc;
    ram_cell[   11423] = 32'ha0a67aac;
    ram_cell[   11424] = 32'hc8e4b76f;
    ram_cell[   11425] = 32'h1bd8ae96;
    ram_cell[   11426] = 32'hf0022f2f;
    ram_cell[   11427] = 32'h8da99c5f;
    ram_cell[   11428] = 32'hbc6a6db6;
    ram_cell[   11429] = 32'h60b49bd2;
    ram_cell[   11430] = 32'hecbd0290;
    ram_cell[   11431] = 32'hca51ab1b;
    ram_cell[   11432] = 32'h44a9e8fc;
    ram_cell[   11433] = 32'h2dc229c8;
    ram_cell[   11434] = 32'h3e3d936a;
    ram_cell[   11435] = 32'h4b1b38d6;
    ram_cell[   11436] = 32'h2f3d0c37;
    ram_cell[   11437] = 32'h278bb7e2;
    ram_cell[   11438] = 32'heb272f8f;
    ram_cell[   11439] = 32'h8b35593b;
    ram_cell[   11440] = 32'hf5e9c30d;
    ram_cell[   11441] = 32'h7dc8576e;
    ram_cell[   11442] = 32'ha36b6c7b;
    ram_cell[   11443] = 32'h315fb766;
    ram_cell[   11444] = 32'h65633dd4;
    ram_cell[   11445] = 32'h49575a31;
    ram_cell[   11446] = 32'h5aa20a32;
    ram_cell[   11447] = 32'ha336e79d;
    ram_cell[   11448] = 32'hc7363c92;
    ram_cell[   11449] = 32'ha7e3fa4b;
    ram_cell[   11450] = 32'h42654d5e;
    ram_cell[   11451] = 32'h8e93fe85;
    ram_cell[   11452] = 32'hbce680c2;
    ram_cell[   11453] = 32'h1307d70f;
    ram_cell[   11454] = 32'h556b63a1;
    ram_cell[   11455] = 32'ha6a9e6f3;
    ram_cell[   11456] = 32'he13c52c8;
    ram_cell[   11457] = 32'h2d9134a8;
    ram_cell[   11458] = 32'h41a96f55;
    ram_cell[   11459] = 32'hc52eb355;
    ram_cell[   11460] = 32'h31c84ccf;
    ram_cell[   11461] = 32'heb82ff02;
    ram_cell[   11462] = 32'hac8b2dea;
    ram_cell[   11463] = 32'hfe58340e;
    ram_cell[   11464] = 32'hf71d03e2;
    ram_cell[   11465] = 32'h67fe2769;
    ram_cell[   11466] = 32'h4751189f;
    ram_cell[   11467] = 32'h5be81ccc;
    ram_cell[   11468] = 32'h00cd4440;
    ram_cell[   11469] = 32'h5dbbe995;
    ram_cell[   11470] = 32'ha2c16010;
    ram_cell[   11471] = 32'h2c2ef2cf;
    ram_cell[   11472] = 32'h3ac523dc;
    ram_cell[   11473] = 32'hcc07d712;
    ram_cell[   11474] = 32'h6bfdede4;
    ram_cell[   11475] = 32'hc9c28458;
    ram_cell[   11476] = 32'hcb90f632;
    ram_cell[   11477] = 32'hddbcd296;
    ram_cell[   11478] = 32'h93f8b2d9;
    ram_cell[   11479] = 32'h0e4d9227;
    ram_cell[   11480] = 32'h07d2619b;
    ram_cell[   11481] = 32'hd1dd3a21;
    ram_cell[   11482] = 32'hfb4d0f25;
    ram_cell[   11483] = 32'h9b60fe4a;
    ram_cell[   11484] = 32'h0ecfd01b;
    ram_cell[   11485] = 32'hf80612c4;
    ram_cell[   11486] = 32'h0a2b3b2a;
    ram_cell[   11487] = 32'h7362e720;
    ram_cell[   11488] = 32'hf928c348;
    ram_cell[   11489] = 32'ha632286e;
    ram_cell[   11490] = 32'hb4bfd39f;
    ram_cell[   11491] = 32'hd202b583;
    ram_cell[   11492] = 32'hf4f30cfc;
    ram_cell[   11493] = 32'h43f77913;
    ram_cell[   11494] = 32'h09536e59;
    ram_cell[   11495] = 32'h07ae4e15;
    ram_cell[   11496] = 32'h44500b70;
    ram_cell[   11497] = 32'h9b3cff67;
    ram_cell[   11498] = 32'hca0c964b;
    ram_cell[   11499] = 32'h2f067584;
    ram_cell[   11500] = 32'h95d6c31d;
    ram_cell[   11501] = 32'hdbfb0e73;
    ram_cell[   11502] = 32'h35e4afe4;
    ram_cell[   11503] = 32'ha78876ba;
    ram_cell[   11504] = 32'h81ee52d3;
    ram_cell[   11505] = 32'he23ecad1;
    ram_cell[   11506] = 32'hed3c2fc7;
    ram_cell[   11507] = 32'h89bd7dca;
    ram_cell[   11508] = 32'h8c325c0c;
    ram_cell[   11509] = 32'h2ab1e3c4;
    ram_cell[   11510] = 32'h1bd2ac5a;
    ram_cell[   11511] = 32'hbd58e3ef;
    ram_cell[   11512] = 32'h2744df41;
    ram_cell[   11513] = 32'h61774e71;
    ram_cell[   11514] = 32'he5928ac8;
    ram_cell[   11515] = 32'hc3968603;
    ram_cell[   11516] = 32'h8ab1954a;
    ram_cell[   11517] = 32'hbc1bc111;
    ram_cell[   11518] = 32'h9473e412;
    ram_cell[   11519] = 32'hf52e5d02;
    ram_cell[   11520] = 32'h63bd7387;
    ram_cell[   11521] = 32'hd98d2a96;
    ram_cell[   11522] = 32'h21607eb3;
    ram_cell[   11523] = 32'h04e2243a;
    ram_cell[   11524] = 32'h3d4f1183;
    ram_cell[   11525] = 32'he9989d54;
    ram_cell[   11526] = 32'h7f7eb0fc;
    ram_cell[   11527] = 32'hfdcab085;
    ram_cell[   11528] = 32'h53b33772;
    ram_cell[   11529] = 32'h2c4ad1fc;
    ram_cell[   11530] = 32'h007e6d4b;
    ram_cell[   11531] = 32'hb9f35f7d;
    ram_cell[   11532] = 32'hbb4735c1;
    ram_cell[   11533] = 32'h15d2db5d;
    ram_cell[   11534] = 32'h7f613a3f;
    ram_cell[   11535] = 32'h3ed0c208;
    ram_cell[   11536] = 32'hfe5462d1;
    ram_cell[   11537] = 32'h5bfdfebb;
    ram_cell[   11538] = 32'h628af41d;
    ram_cell[   11539] = 32'h93ba2d1d;
    ram_cell[   11540] = 32'ha21b5111;
    ram_cell[   11541] = 32'h544e2f74;
    ram_cell[   11542] = 32'h255feb91;
    ram_cell[   11543] = 32'h87553932;
    ram_cell[   11544] = 32'h49ac4a23;
    ram_cell[   11545] = 32'h87b056aa;
    ram_cell[   11546] = 32'h675aa9cb;
    ram_cell[   11547] = 32'hd86c165a;
    ram_cell[   11548] = 32'h1bb5c1fb;
    ram_cell[   11549] = 32'h2f32e921;
    ram_cell[   11550] = 32'he8011d66;
    ram_cell[   11551] = 32'h6d05bb27;
    ram_cell[   11552] = 32'h07580be4;
    ram_cell[   11553] = 32'h5c57c38f;
    ram_cell[   11554] = 32'hbe6b08db;
    ram_cell[   11555] = 32'h7ab2aae6;
    ram_cell[   11556] = 32'haede5694;
    ram_cell[   11557] = 32'ha38b4c58;
    ram_cell[   11558] = 32'h039c3c8e;
    ram_cell[   11559] = 32'hb92f5eca;
    ram_cell[   11560] = 32'h6a2ed7a2;
    ram_cell[   11561] = 32'hff09840e;
    ram_cell[   11562] = 32'h9ca88f3b;
    ram_cell[   11563] = 32'h6353ed3b;
    ram_cell[   11564] = 32'h076dd1cc;
    ram_cell[   11565] = 32'h87ae60e9;
    ram_cell[   11566] = 32'hc376f18b;
    ram_cell[   11567] = 32'heb9f7cc2;
    ram_cell[   11568] = 32'hb6cb3af1;
    ram_cell[   11569] = 32'h7bf25d1e;
    ram_cell[   11570] = 32'h082704f3;
    ram_cell[   11571] = 32'h36ee9aa6;
    ram_cell[   11572] = 32'h9faaabcb;
    ram_cell[   11573] = 32'h53b75abe;
    ram_cell[   11574] = 32'h842f605a;
    ram_cell[   11575] = 32'h21173ac2;
    ram_cell[   11576] = 32'h1d3e9ea9;
    ram_cell[   11577] = 32'hf1f96877;
    ram_cell[   11578] = 32'h5f43b415;
    ram_cell[   11579] = 32'hf3fad886;
    ram_cell[   11580] = 32'h9449f908;
    ram_cell[   11581] = 32'h161394c6;
    ram_cell[   11582] = 32'h1d35c685;
    ram_cell[   11583] = 32'he2922b4c;
    ram_cell[   11584] = 32'h2563a336;
    ram_cell[   11585] = 32'h35cf45b0;
    ram_cell[   11586] = 32'h11e4702a;
    ram_cell[   11587] = 32'h56194156;
    ram_cell[   11588] = 32'h61928cdd;
    ram_cell[   11589] = 32'h7d36f0ef;
    ram_cell[   11590] = 32'h8697c573;
    ram_cell[   11591] = 32'hd3b618b9;
    ram_cell[   11592] = 32'h49b6e950;
    ram_cell[   11593] = 32'h1710fb76;
    ram_cell[   11594] = 32'h8c4421c5;
    ram_cell[   11595] = 32'hda46a216;
    ram_cell[   11596] = 32'h3447ce41;
    ram_cell[   11597] = 32'h8b0a14e4;
    ram_cell[   11598] = 32'hb6123dc6;
    ram_cell[   11599] = 32'h114d3ba8;
    ram_cell[   11600] = 32'h3ce3b944;
    ram_cell[   11601] = 32'h0dab312e;
    ram_cell[   11602] = 32'h588aa05a;
    ram_cell[   11603] = 32'hd0bc8786;
    ram_cell[   11604] = 32'h684001cf;
    ram_cell[   11605] = 32'hffc5fb90;
    ram_cell[   11606] = 32'hb2fe84a8;
    ram_cell[   11607] = 32'ha036291a;
    ram_cell[   11608] = 32'hebd13593;
    ram_cell[   11609] = 32'h69da1906;
    ram_cell[   11610] = 32'h39655bce;
    ram_cell[   11611] = 32'h88435654;
    ram_cell[   11612] = 32'h99d3564e;
    ram_cell[   11613] = 32'h26d75bb2;
    ram_cell[   11614] = 32'h2ce0afef;
    ram_cell[   11615] = 32'h9055e3af;
    ram_cell[   11616] = 32'hed299348;
    ram_cell[   11617] = 32'h022302c4;
    ram_cell[   11618] = 32'hea5342f4;
    ram_cell[   11619] = 32'h4450e2b5;
    ram_cell[   11620] = 32'h0e3ea1f6;
    ram_cell[   11621] = 32'hcac97b7e;
    ram_cell[   11622] = 32'h9c4d53d7;
    ram_cell[   11623] = 32'h0e1a2a73;
    ram_cell[   11624] = 32'h63250e05;
    ram_cell[   11625] = 32'hd649c14d;
    ram_cell[   11626] = 32'hedd990f5;
    ram_cell[   11627] = 32'hec791d50;
    ram_cell[   11628] = 32'he2c4e9d6;
    ram_cell[   11629] = 32'h966a8bdc;
    ram_cell[   11630] = 32'hefadacc5;
    ram_cell[   11631] = 32'h33730be6;
    ram_cell[   11632] = 32'h9d8963e2;
    ram_cell[   11633] = 32'h399e1158;
    ram_cell[   11634] = 32'h4441fe86;
    ram_cell[   11635] = 32'he221a3da;
    ram_cell[   11636] = 32'h63ea1c92;
    ram_cell[   11637] = 32'he3e3ee31;
    ram_cell[   11638] = 32'h9f6df09c;
    ram_cell[   11639] = 32'h88269c1a;
    ram_cell[   11640] = 32'h70fe04e6;
    ram_cell[   11641] = 32'h6904c996;
    ram_cell[   11642] = 32'h2242ff2d;
    ram_cell[   11643] = 32'h4adb08cb;
    ram_cell[   11644] = 32'h605b23a8;
    ram_cell[   11645] = 32'hf9f240e0;
    ram_cell[   11646] = 32'hbd0ebfc3;
    ram_cell[   11647] = 32'h40242fa1;
    ram_cell[   11648] = 32'h1d2f8e34;
    ram_cell[   11649] = 32'h112c840b;
    ram_cell[   11650] = 32'h3cf4332a;
    ram_cell[   11651] = 32'h672a6d3f;
    ram_cell[   11652] = 32'hf8c2874b;
    ram_cell[   11653] = 32'h50e2212e;
    ram_cell[   11654] = 32'h3d207c47;
    ram_cell[   11655] = 32'h170779c1;
    ram_cell[   11656] = 32'hddb151ae;
    ram_cell[   11657] = 32'h63f36fb0;
    ram_cell[   11658] = 32'h056618c1;
    ram_cell[   11659] = 32'h361ce35e;
    ram_cell[   11660] = 32'h5563c400;
    ram_cell[   11661] = 32'h8a922ee8;
    ram_cell[   11662] = 32'h9865bd48;
    ram_cell[   11663] = 32'hfc486573;
    ram_cell[   11664] = 32'h462ce9ff;
    ram_cell[   11665] = 32'h66611b96;
    ram_cell[   11666] = 32'h175e8bc0;
    ram_cell[   11667] = 32'ha7a593c4;
    ram_cell[   11668] = 32'h9014a1c8;
    ram_cell[   11669] = 32'h5db9cb71;
    ram_cell[   11670] = 32'h485d1211;
    ram_cell[   11671] = 32'h649f9a55;
    ram_cell[   11672] = 32'h4b2e1f7e;
    ram_cell[   11673] = 32'h7a58119e;
    ram_cell[   11674] = 32'h297a3f81;
    ram_cell[   11675] = 32'hf1ddc4c3;
    ram_cell[   11676] = 32'hff646847;
    ram_cell[   11677] = 32'h0c779f22;
    ram_cell[   11678] = 32'h84d3ee16;
    ram_cell[   11679] = 32'hcc06435a;
    ram_cell[   11680] = 32'h21ed97f5;
    ram_cell[   11681] = 32'hef428b22;
    ram_cell[   11682] = 32'hb639e7db;
    ram_cell[   11683] = 32'hd3b43231;
    ram_cell[   11684] = 32'he43aaf44;
    ram_cell[   11685] = 32'h275acdaa;
    ram_cell[   11686] = 32'h630a2bf3;
    ram_cell[   11687] = 32'hcc6a9554;
    ram_cell[   11688] = 32'h19c6a470;
    ram_cell[   11689] = 32'h5bea1b2b;
    ram_cell[   11690] = 32'ha6cb5f98;
    ram_cell[   11691] = 32'hc37cd5af;
    ram_cell[   11692] = 32'h8d3fce8d;
    ram_cell[   11693] = 32'h47a7fae9;
    ram_cell[   11694] = 32'hcfd719c2;
    ram_cell[   11695] = 32'h0b43fd37;
    ram_cell[   11696] = 32'h10412e03;
    ram_cell[   11697] = 32'hbaed4f92;
    ram_cell[   11698] = 32'h961bac08;
    ram_cell[   11699] = 32'h78d3b7b6;
    ram_cell[   11700] = 32'hfe33a7c9;
    ram_cell[   11701] = 32'h8cadfb67;
    ram_cell[   11702] = 32'hfa1ca433;
    ram_cell[   11703] = 32'h38b9f16a;
    ram_cell[   11704] = 32'h00da3677;
    ram_cell[   11705] = 32'h496742be;
    ram_cell[   11706] = 32'h7401df0c;
    ram_cell[   11707] = 32'h6699029b;
    ram_cell[   11708] = 32'h70359ae0;
    ram_cell[   11709] = 32'hd5f6c72d;
    ram_cell[   11710] = 32'hd4fb1402;
    ram_cell[   11711] = 32'he317e8bc;
    ram_cell[   11712] = 32'hd284f54a;
    ram_cell[   11713] = 32'h2467ebcd;
    ram_cell[   11714] = 32'h44857a0a;
    ram_cell[   11715] = 32'hd401626d;
    ram_cell[   11716] = 32'ha0a69d21;
    ram_cell[   11717] = 32'he05f5279;
    ram_cell[   11718] = 32'h5670cc5a;
    ram_cell[   11719] = 32'h73b6c08f;
    ram_cell[   11720] = 32'hae81a9d5;
    ram_cell[   11721] = 32'hae6096aa;
    ram_cell[   11722] = 32'h9110ae62;
    ram_cell[   11723] = 32'h4065411d;
    ram_cell[   11724] = 32'h12e9fb3c;
    ram_cell[   11725] = 32'h9fd443aa;
    ram_cell[   11726] = 32'h22ea5033;
    ram_cell[   11727] = 32'hcd50848d;
    ram_cell[   11728] = 32'h3324c3c1;
    ram_cell[   11729] = 32'h5fb21531;
    ram_cell[   11730] = 32'hcf8b72f6;
    ram_cell[   11731] = 32'h59802beb;
    ram_cell[   11732] = 32'hfe3b7225;
    ram_cell[   11733] = 32'h7c2e318d;
    ram_cell[   11734] = 32'h21d4b962;
    ram_cell[   11735] = 32'h53a1078d;
    ram_cell[   11736] = 32'hf539c565;
    ram_cell[   11737] = 32'ha8bae9e1;
    ram_cell[   11738] = 32'hb268a36d;
    ram_cell[   11739] = 32'h10fe2d6a;
    ram_cell[   11740] = 32'h476ddde4;
    ram_cell[   11741] = 32'heeeb91c0;
    ram_cell[   11742] = 32'h5c2a9d5b;
    ram_cell[   11743] = 32'h4f800413;
    ram_cell[   11744] = 32'h2c4d04b3;
    ram_cell[   11745] = 32'h4052f533;
    ram_cell[   11746] = 32'h5acb1485;
    ram_cell[   11747] = 32'hdfaf69b8;
    ram_cell[   11748] = 32'hc985417a;
    ram_cell[   11749] = 32'h54a3b585;
    ram_cell[   11750] = 32'h43468b05;
    ram_cell[   11751] = 32'hb69cdd47;
    ram_cell[   11752] = 32'hf87eb42e;
    ram_cell[   11753] = 32'hd56d011f;
    ram_cell[   11754] = 32'h7bfc5261;
    ram_cell[   11755] = 32'hede29dd7;
    ram_cell[   11756] = 32'hdc0b4fce;
    ram_cell[   11757] = 32'h77bc95ea;
    ram_cell[   11758] = 32'h6c882361;
    ram_cell[   11759] = 32'he6bf55e5;
    ram_cell[   11760] = 32'h8df87e02;
    ram_cell[   11761] = 32'h824e7973;
    ram_cell[   11762] = 32'h2013860e;
    ram_cell[   11763] = 32'hec3331ad;
    ram_cell[   11764] = 32'he02aec0d;
    ram_cell[   11765] = 32'hcd0846a5;
    ram_cell[   11766] = 32'h45e7911a;
    ram_cell[   11767] = 32'hfb02cd0c;
    ram_cell[   11768] = 32'hc5ee4a5e;
    ram_cell[   11769] = 32'h16ece1dd;
    ram_cell[   11770] = 32'h35f2689e;
    ram_cell[   11771] = 32'h54758019;
    ram_cell[   11772] = 32'h74bada56;
    ram_cell[   11773] = 32'h67553010;
    ram_cell[   11774] = 32'h55108e64;
    ram_cell[   11775] = 32'hee4487e5;
    ram_cell[   11776] = 32'h2812c9e5;
    ram_cell[   11777] = 32'hf369274a;
    ram_cell[   11778] = 32'hf659a5c3;
    ram_cell[   11779] = 32'heb581270;
    ram_cell[   11780] = 32'h1ac2275f;
    ram_cell[   11781] = 32'h7fd1cd46;
    ram_cell[   11782] = 32'h46c6cb9f;
    ram_cell[   11783] = 32'h13439d74;
    ram_cell[   11784] = 32'h15b0c938;
    ram_cell[   11785] = 32'hea82fecb;
    ram_cell[   11786] = 32'h3fc22116;
    ram_cell[   11787] = 32'h45171dd9;
    ram_cell[   11788] = 32'h598e4ab0;
    ram_cell[   11789] = 32'h9104805a;
    ram_cell[   11790] = 32'h3e4a968d;
    ram_cell[   11791] = 32'h82e31c84;
    ram_cell[   11792] = 32'hd0800e71;
    ram_cell[   11793] = 32'hdaf380f2;
    ram_cell[   11794] = 32'hd28bb3b3;
    ram_cell[   11795] = 32'h6e88543f;
    ram_cell[   11796] = 32'heea8b700;
    ram_cell[   11797] = 32'h3526911b;
    ram_cell[   11798] = 32'h55658267;
    ram_cell[   11799] = 32'hff18e5ad;
    ram_cell[   11800] = 32'ha8a8a5c8;
    ram_cell[   11801] = 32'h6f6c1248;
    ram_cell[   11802] = 32'h4025aa02;
    ram_cell[   11803] = 32'hce9fae35;
    ram_cell[   11804] = 32'hde9a1cf1;
    ram_cell[   11805] = 32'ha2359126;
    ram_cell[   11806] = 32'hfeb5f0ec;
    ram_cell[   11807] = 32'h45a8a381;
    ram_cell[   11808] = 32'h059547bc;
    ram_cell[   11809] = 32'hc1e4dbac;
    ram_cell[   11810] = 32'h12288815;
    ram_cell[   11811] = 32'h99c77bc9;
    ram_cell[   11812] = 32'h5e531c3a;
    ram_cell[   11813] = 32'hbf57aac1;
    ram_cell[   11814] = 32'h6eb91477;
    ram_cell[   11815] = 32'h0fdf77a4;
    ram_cell[   11816] = 32'hdf4900e2;
    ram_cell[   11817] = 32'hf3ff03a0;
    ram_cell[   11818] = 32'h75a08c8a;
    ram_cell[   11819] = 32'he087f8c6;
    ram_cell[   11820] = 32'h1c45f4b0;
    ram_cell[   11821] = 32'hbf872a62;
    ram_cell[   11822] = 32'h15dd52fe;
    ram_cell[   11823] = 32'h319ed77d;
    ram_cell[   11824] = 32'h4dac0920;
    ram_cell[   11825] = 32'hfd80c8ab;
    ram_cell[   11826] = 32'ha270815a;
    ram_cell[   11827] = 32'hf8e2500a;
    ram_cell[   11828] = 32'hafecea98;
    ram_cell[   11829] = 32'h40c0b8f9;
    ram_cell[   11830] = 32'hb0bf1ec7;
    ram_cell[   11831] = 32'hc812b92d;
    ram_cell[   11832] = 32'h689c9404;
    ram_cell[   11833] = 32'hf2bc379c;
    ram_cell[   11834] = 32'h8beb8206;
    ram_cell[   11835] = 32'h0c07aaa1;
    ram_cell[   11836] = 32'h90fcdbc5;
    ram_cell[   11837] = 32'h25af0ff2;
    ram_cell[   11838] = 32'h96120ccf;
    ram_cell[   11839] = 32'hdacb4fe9;
    ram_cell[   11840] = 32'h50c8020f;
    ram_cell[   11841] = 32'h8505a0d8;
    ram_cell[   11842] = 32'hb1f15bdf;
    ram_cell[   11843] = 32'h65b7d94c;
    ram_cell[   11844] = 32'hf80c7dad;
    ram_cell[   11845] = 32'he5cfb5e9;
    ram_cell[   11846] = 32'hfc92a54f;
    ram_cell[   11847] = 32'h7328d476;
    ram_cell[   11848] = 32'he5373139;
    ram_cell[   11849] = 32'h9bb4539e;
    ram_cell[   11850] = 32'h8e80e962;
    ram_cell[   11851] = 32'hc9489353;
    ram_cell[   11852] = 32'hd9c66a5a;
    ram_cell[   11853] = 32'h62f3169f;
    ram_cell[   11854] = 32'hece16969;
    ram_cell[   11855] = 32'h2db28e47;
    ram_cell[   11856] = 32'h7c684551;
    ram_cell[   11857] = 32'h0aedac88;
    ram_cell[   11858] = 32'h3809983e;
    ram_cell[   11859] = 32'he153800c;
    ram_cell[   11860] = 32'h41d8f1dc;
    ram_cell[   11861] = 32'h94167f8b;
    ram_cell[   11862] = 32'h42e134a3;
    ram_cell[   11863] = 32'h895b91fa;
    ram_cell[   11864] = 32'h82da972e;
    ram_cell[   11865] = 32'he796d988;
    ram_cell[   11866] = 32'h8a613bf9;
    ram_cell[   11867] = 32'h3d9912e6;
    ram_cell[   11868] = 32'h561f0896;
    ram_cell[   11869] = 32'h358392c5;
    ram_cell[   11870] = 32'h665e67e7;
    ram_cell[   11871] = 32'hef716bae;
    ram_cell[   11872] = 32'h50b709ce;
    ram_cell[   11873] = 32'h6c6ccfba;
    ram_cell[   11874] = 32'h149d17cb;
    ram_cell[   11875] = 32'h6d2e4e31;
    ram_cell[   11876] = 32'h8cdea6a4;
    ram_cell[   11877] = 32'hf0034b2e;
    ram_cell[   11878] = 32'hfc2a3b1b;
    ram_cell[   11879] = 32'h725b926c;
    ram_cell[   11880] = 32'h18202c73;
    ram_cell[   11881] = 32'h937184a4;
    ram_cell[   11882] = 32'h22936c30;
    ram_cell[   11883] = 32'hb938b2c4;
    ram_cell[   11884] = 32'hd9d59c0d;
    ram_cell[   11885] = 32'h77804b81;
    ram_cell[   11886] = 32'ha01c7545;
    ram_cell[   11887] = 32'h764acbbb;
    ram_cell[   11888] = 32'h6655b773;
    ram_cell[   11889] = 32'hb3e5b834;
    ram_cell[   11890] = 32'h826a5e8e;
    ram_cell[   11891] = 32'h91fcc97b;
    ram_cell[   11892] = 32'hdaea0c47;
    ram_cell[   11893] = 32'h09cf12ef;
    ram_cell[   11894] = 32'hac91df54;
    ram_cell[   11895] = 32'h6003d972;
    ram_cell[   11896] = 32'hd8471974;
    ram_cell[   11897] = 32'h6b78f50c;
    ram_cell[   11898] = 32'h874040fd;
    ram_cell[   11899] = 32'h904b5f6c;
    ram_cell[   11900] = 32'hc5020e4d;
    ram_cell[   11901] = 32'h4553926e;
    ram_cell[   11902] = 32'hc826324e;
    ram_cell[   11903] = 32'h13c920e2;
    ram_cell[   11904] = 32'he389c40d;
    ram_cell[   11905] = 32'h384379db;
    ram_cell[   11906] = 32'h4d2be73d;
    ram_cell[   11907] = 32'hb2eab55f;
    ram_cell[   11908] = 32'h6a26e94d;
    ram_cell[   11909] = 32'h21dbdcb1;
    ram_cell[   11910] = 32'h3cd56f80;
    ram_cell[   11911] = 32'h5d3cb61b;
    ram_cell[   11912] = 32'h50a54f1a;
    ram_cell[   11913] = 32'hd93e51ea;
    ram_cell[   11914] = 32'h7831c14a;
    ram_cell[   11915] = 32'hc85990d9;
    ram_cell[   11916] = 32'he113f0d5;
    ram_cell[   11917] = 32'h8f612643;
    ram_cell[   11918] = 32'hb67511ea;
    ram_cell[   11919] = 32'hcf1913ed;
    ram_cell[   11920] = 32'h07013456;
    ram_cell[   11921] = 32'hc423e114;
    ram_cell[   11922] = 32'h5189383d;
    ram_cell[   11923] = 32'h2d674e4f;
    ram_cell[   11924] = 32'he279ac02;
    ram_cell[   11925] = 32'h3954191e;
    ram_cell[   11926] = 32'hc9fa7f8c;
    ram_cell[   11927] = 32'hae3121b7;
    ram_cell[   11928] = 32'h0d466382;
    ram_cell[   11929] = 32'h3ebef890;
    ram_cell[   11930] = 32'hc6797856;
    ram_cell[   11931] = 32'h8bdf039e;
    ram_cell[   11932] = 32'hb31b6539;
    ram_cell[   11933] = 32'h9fdba663;
    ram_cell[   11934] = 32'ha3d6063a;
    ram_cell[   11935] = 32'hbbbb58af;
    ram_cell[   11936] = 32'h60281bd2;
    ram_cell[   11937] = 32'h2730041b;
    ram_cell[   11938] = 32'h2302f6eb;
    ram_cell[   11939] = 32'hb23ccb17;
    ram_cell[   11940] = 32'h1facf677;
    ram_cell[   11941] = 32'h2ce47919;
    ram_cell[   11942] = 32'h26415420;
    ram_cell[   11943] = 32'h4601c56a;
    ram_cell[   11944] = 32'ha70526e5;
    ram_cell[   11945] = 32'hd5e0facc;
    ram_cell[   11946] = 32'hfa8065b5;
    ram_cell[   11947] = 32'h7f33da10;
    ram_cell[   11948] = 32'hdf5b5bc3;
    ram_cell[   11949] = 32'h2595a561;
    ram_cell[   11950] = 32'h1f9491e6;
    ram_cell[   11951] = 32'h7f76819c;
    ram_cell[   11952] = 32'h2f593fe7;
    ram_cell[   11953] = 32'h9dcc052a;
    ram_cell[   11954] = 32'h94e4b512;
    ram_cell[   11955] = 32'h1b57519e;
    ram_cell[   11956] = 32'h75737cd5;
    ram_cell[   11957] = 32'h7246c9fc;
    ram_cell[   11958] = 32'h254c82c5;
    ram_cell[   11959] = 32'hc2e56564;
    ram_cell[   11960] = 32'h97d2b7b7;
    ram_cell[   11961] = 32'h26e4fa97;
    ram_cell[   11962] = 32'h0d492703;
    ram_cell[   11963] = 32'hfc0027f5;
    ram_cell[   11964] = 32'h4ebb3010;
    ram_cell[   11965] = 32'h85718915;
    ram_cell[   11966] = 32'h9a5da4e2;
    ram_cell[   11967] = 32'h456ed79e;
    ram_cell[   11968] = 32'ha20b575c;
    ram_cell[   11969] = 32'h5afbfc0e;
    ram_cell[   11970] = 32'ha8407bfa;
    ram_cell[   11971] = 32'hb2639e48;
    ram_cell[   11972] = 32'ha4d26070;
    ram_cell[   11973] = 32'hd99350fb;
    ram_cell[   11974] = 32'hbf37212a;
    ram_cell[   11975] = 32'h3f501fc1;
    ram_cell[   11976] = 32'h91e149bf;
    ram_cell[   11977] = 32'h14b6df37;
    ram_cell[   11978] = 32'h24c271ec;
    ram_cell[   11979] = 32'he3902054;
    ram_cell[   11980] = 32'h093bbed7;
    ram_cell[   11981] = 32'h11bb4eb9;
    ram_cell[   11982] = 32'ha5cece1d;
    ram_cell[   11983] = 32'h6d23b8e8;
    ram_cell[   11984] = 32'h864ee6ef;
    ram_cell[   11985] = 32'h8901970f;
    ram_cell[   11986] = 32'hce9709cd;
    ram_cell[   11987] = 32'h81473fb3;
    ram_cell[   11988] = 32'h9862139e;
    ram_cell[   11989] = 32'he353b581;
    ram_cell[   11990] = 32'hcf0e7f77;
    ram_cell[   11991] = 32'h98f1dacc;
    ram_cell[   11992] = 32'h174dcd0a;
    ram_cell[   11993] = 32'h4639eb99;
    ram_cell[   11994] = 32'hb98f64e9;
    ram_cell[   11995] = 32'h0f6225fc;
    ram_cell[   11996] = 32'hfd5207ce;
    ram_cell[   11997] = 32'h2b106613;
    ram_cell[   11998] = 32'h74490fab;
    ram_cell[   11999] = 32'ha4393f66;
    ram_cell[   12000] = 32'h39b61a4c;
    ram_cell[   12001] = 32'hd7848c7d;
    ram_cell[   12002] = 32'h53aad312;
    ram_cell[   12003] = 32'ha10850f6;
    ram_cell[   12004] = 32'h1b320fc3;
    ram_cell[   12005] = 32'hca4057e0;
    ram_cell[   12006] = 32'hc655978b;
    ram_cell[   12007] = 32'hb610b4dc;
    ram_cell[   12008] = 32'h2a1bc519;
    ram_cell[   12009] = 32'h05f1375a;
    ram_cell[   12010] = 32'hdf7bb056;
    ram_cell[   12011] = 32'h70d998fc;
    ram_cell[   12012] = 32'hbf2e2066;
    ram_cell[   12013] = 32'ha6daf508;
    ram_cell[   12014] = 32'h04ab0978;
    ram_cell[   12015] = 32'he2f35bf7;
    ram_cell[   12016] = 32'hd3c7fe3d;
    ram_cell[   12017] = 32'h23d4ebd2;
    ram_cell[   12018] = 32'h63b0f911;
    ram_cell[   12019] = 32'h0b1bb34b;
    ram_cell[   12020] = 32'h66bd9e1b;
    ram_cell[   12021] = 32'h182deec8;
    ram_cell[   12022] = 32'h53fe820e;
    ram_cell[   12023] = 32'ha22c34f1;
    ram_cell[   12024] = 32'hcb4380e6;
    ram_cell[   12025] = 32'ha43b8dd8;
    ram_cell[   12026] = 32'hefb3df76;
    ram_cell[   12027] = 32'ha58a6186;
    ram_cell[   12028] = 32'h79e273e0;
    ram_cell[   12029] = 32'hf1a8c632;
    ram_cell[   12030] = 32'h9e2f6149;
    ram_cell[   12031] = 32'h3beee95b;
    ram_cell[   12032] = 32'hce503d4b;
    ram_cell[   12033] = 32'h9dd6cb89;
    ram_cell[   12034] = 32'hc777e8cc;
    ram_cell[   12035] = 32'hf6b561b5;
    ram_cell[   12036] = 32'hf7310e73;
    ram_cell[   12037] = 32'hed0b5227;
    ram_cell[   12038] = 32'h5ec1783d;
    ram_cell[   12039] = 32'h96f5c96c;
    ram_cell[   12040] = 32'h730827d8;
    ram_cell[   12041] = 32'h90e5cd04;
    ram_cell[   12042] = 32'he422c14f;
    ram_cell[   12043] = 32'hcfb8b6d6;
    ram_cell[   12044] = 32'h8f564f69;
    ram_cell[   12045] = 32'h9abc4333;
    ram_cell[   12046] = 32'h44e9bafd;
    ram_cell[   12047] = 32'h84857224;
    ram_cell[   12048] = 32'ha25fa616;
    ram_cell[   12049] = 32'ha555d13c;
    ram_cell[   12050] = 32'h043670d0;
    ram_cell[   12051] = 32'h808124af;
    ram_cell[   12052] = 32'h62ef2d0b;
    ram_cell[   12053] = 32'hbb9ee59a;
    ram_cell[   12054] = 32'hfee56054;
    ram_cell[   12055] = 32'h1773854c;
    ram_cell[   12056] = 32'h57a02331;
    ram_cell[   12057] = 32'h0446cd5f;
    ram_cell[   12058] = 32'h757d31c1;
    ram_cell[   12059] = 32'h2e5359c7;
    ram_cell[   12060] = 32'h6ccdce8d;
    ram_cell[   12061] = 32'h3c942e49;
    ram_cell[   12062] = 32'h6a590329;
    ram_cell[   12063] = 32'h36175936;
    ram_cell[   12064] = 32'h6a237595;
    ram_cell[   12065] = 32'h9e5cadd2;
    ram_cell[   12066] = 32'h2e81f505;
    ram_cell[   12067] = 32'hc695fd9f;
    ram_cell[   12068] = 32'h62a2dd0c;
    ram_cell[   12069] = 32'h48af5691;
    ram_cell[   12070] = 32'h2439c8fa;
    ram_cell[   12071] = 32'hfa470e99;
    ram_cell[   12072] = 32'h3e1cdb83;
    ram_cell[   12073] = 32'h986f807b;
    ram_cell[   12074] = 32'hac6b638c;
    ram_cell[   12075] = 32'h0b77dfb4;
    ram_cell[   12076] = 32'hfddb3538;
    ram_cell[   12077] = 32'hf4d4b978;
    ram_cell[   12078] = 32'h4ac80dd4;
    ram_cell[   12079] = 32'hfd36b783;
    ram_cell[   12080] = 32'he16c6edd;
    ram_cell[   12081] = 32'hba2398ce;
    ram_cell[   12082] = 32'h53756fff;
    ram_cell[   12083] = 32'h439b69d0;
    ram_cell[   12084] = 32'h78a1042a;
    ram_cell[   12085] = 32'hd2f2cee7;
    ram_cell[   12086] = 32'h2a89a688;
    ram_cell[   12087] = 32'h116821e4;
    ram_cell[   12088] = 32'h1c52aa51;
    ram_cell[   12089] = 32'h73cbdeb6;
    ram_cell[   12090] = 32'he25cd06c;
    ram_cell[   12091] = 32'had42768c;
    ram_cell[   12092] = 32'h822526f7;
    ram_cell[   12093] = 32'h140d9197;
    ram_cell[   12094] = 32'h031db9a7;
    ram_cell[   12095] = 32'h9e772f88;
    ram_cell[   12096] = 32'h7b69efb1;
    ram_cell[   12097] = 32'h14ccdc2b;
    ram_cell[   12098] = 32'h9f465792;
    ram_cell[   12099] = 32'hcb68dbad;
    ram_cell[   12100] = 32'h86c47b64;
    ram_cell[   12101] = 32'h3816451f;
    ram_cell[   12102] = 32'hbcbb5f90;
    ram_cell[   12103] = 32'hd97ef8e2;
    ram_cell[   12104] = 32'hfd3e6cee;
    ram_cell[   12105] = 32'h72ed1be0;
    ram_cell[   12106] = 32'h64b05fc8;
    ram_cell[   12107] = 32'hef0c50ad;
    ram_cell[   12108] = 32'hce8c103d;
    ram_cell[   12109] = 32'h11262a73;
    ram_cell[   12110] = 32'h43b8471b;
    ram_cell[   12111] = 32'h38f89505;
    ram_cell[   12112] = 32'h364e1fce;
    ram_cell[   12113] = 32'h429e1229;
    ram_cell[   12114] = 32'hfb638f6f;
    ram_cell[   12115] = 32'h167341d8;
    ram_cell[   12116] = 32'hb0096d50;
    ram_cell[   12117] = 32'h1b483d75;
    ram_cell[   12118] = 32'h089df873;
    ram_cell[   12119] = 32'hcc94b8e6;
    ram_cell[   12120] = 32'hca4551a2;
    ram_cell[   12121] = 32'h26160730;
    ram_cell[   12122] = 32'h34bb3a9b;
    ram_cell[   12123] = 32'h96bea44a;
    ram_cell[   12124] = 32'hece04e1a;
    ram_cell[   12125] = 32'h81020404;
    ram_cell[   12126] = 32'hb1c0034d;
    ram_cell[   12127] = 32'h1b0007ce;
    ram_cell[   12128] = 32'h7889154c;
    ram_cell[   12129] = 32'hc09ee817;
    ram_cell[   12130] = 32'h703c11b1;
    ram_cell[   12131] = 32'h0740103c;
    ram_cell[   12132] = 32'he508dd6c;
    ram_cell[   12133] = 32'h210c9b75;
    ram_cell[   12134] = 32'h86efc43b;
    ram_cell[   12135] = 32'h6ea859ba;
    ram_cell[   12136] = 32'hedb0d0a9;
    ram_cell[   12137] = 32'h054d48ed;
    ram_cell[   12138] = 32'hc938a9a1;
    ram_cell[   12139] = 32'hb64bdf71;
    ram_cell[   12140] = 32'h41b73cb3;
    ram_cell[   12141] = 32'h50cf0d0f;
    ram_cell[   12142] = 32'h057388c7;
    ram_cell[   12143] = 32'h009ba632;
    ram_cell[   12144] = 32'h71f81bde;
    ram_cell[   12145] = 32'h15f1a6d3;
    ram_cell[   12146] = 32'h54672c9c;
    ram_cell[   12147] = 32'h34e3142e;
    ram_cell[   12148] = 32'h5e4b60b9;
    ram_cell[   12149] = 32'h85163d44;
    ram_cell[   12150] = 32'h282623ac;
    ram_cell[   12151] = 32'hd5c7f33b;
    ram_cell[   12152] = 32'hd3f962e1;
    ram_cell[   12153] = 32'ha974ce54;
    ram_cell[   12154] = 32'hd491b368;
    ram_cell[   12155] = 32'hf85cded5;
    ram_cell[   12156] = 32'h30ce534f;
    ram_cell[   12157] = 32'h42e3080c;
    ram_cell[   12158] = 32'h508c051c;
    ram_cell[   12159] = 32'hf1773115;
    ram_cell[   12160] = 32'hb89d7a81;
    ram_cell[   12161] = 32'h9234ef36;
    ram_cell[   12162] = 32'h291e8799;
    ram_cell[   12163] = 32'h434c87bd;
    ram_cell[   12164] = 32'h7e3214c8;
    ram_cell[   12165] = 32'h87cd528a;
    ram_cell[   12166] = 32'h7ad0673a;
    ram_cell[   12167] = 32'h037b7272;
    ram_cell[   12168] = 32'h53aa9ab3;
    ram_cell[   12169] = 32'hb984a792;
    ram_cell[   12170] = 32'h6ffc6baf;
    ram_cell[   12171] = 32'hb2e440ce;
    ram_cell[   12172] = 32'h6a7724b3;
    ram_cell[   12173] = 32'h2079e97c;
    ram_cell[   12174] = 32'h04e8fd97;
    ram_cell[   12175] = 32'h990b598b;
    ram_cell[   12176] = 32'hb8546cbb;
    ram_cell[   12177] = 32'h030b8fc6;
    ram_cell[   12178] = 32'hc9149436;
    ram_cell[   12179] = 32'hf8f9dff1;
    ram_cell[   12180] = 32'hb7b61c2c;
    ram_cell[   12181] = 32'h9079013c;
    ram_cell[   12182] = 32'hb2694309;
    ram_cell[   12183] = 32'hd277a199;
    ram_cell[   12184] = 32'h694fc890;
    ram_cell[   12185] = 32'hfaf10b97;
    ram_cell[   12186] = 32'h8b019a6d;
    ram_cell[   12187] = 32'h3f6994d1;
    ram_cell[   12188] = 32'hda2824c9;
    ram_cell[   12189] = 32'hda9b9299;
    ram_cell[   12190] = 32'hf4a0a78c;
    ram_cell[   12191] = 32'h344d35fb;
    ram_cell[   12192] = 32'h45db9333;
    ram_cell[   12193] = 32'haa7591ba;
    ram_cell[   12194] = 32'h078c87f8;
    ram_cell[   12195] = 32'h37f72f35;
    ram_cell[   12196] = 32'h97a9a7c4;
    ram_cell[   12197] = 32'h2f28c8ee;
    ram_cell[   12198] = 32'h1f32ee51;
    ram_cell[   12199] = 32'haa8b7e2e;
    ram_cell[   12200] = 32'ha7382cf3;
    ram_cell[   12201] = 32'h9cda7c2f;
    ram_cell[   12202] = 32'ha07c064b;
    ram_cell[   12203] = 32'h5a751bbc;
    ram_cell[   12204] = 32'h6ec8ab6b;
    ram_cell[   12205] = 32'h9a4fae99;
    ram_cell[   12206] = 32'h83825314;
    ram_cell[   12207] = 32'h7ba9c94c;
    ram_cell[   12208] = 32'hd3e6f1e1;
    ram_cell[   12209] = 32'h89af4b22;
    ram_cell[   12210] = 32'h2019b7f8;
    ram_cell[   12211] = 32'hf2c5b547;
    ram_cell[   12212] = 32'h628344ad;
    ram_cell[   12213] = 32'ha812ed36;
    ram_cell[   12214] = 32'h4864c03c;
    ram_cell[   12215] = 32'h6c612496;
    ram_cell[   12216] = 32'hd44517f1;
    ram_cell[   12217] = 32'h9bc7effc;
    ram_cell[   12218] = 32'hbe2cb38c;
    ram_cell[   12219] = 32'h059159fa;
    ram_cell[   12220] = 32'h82a06fbd;
    ram_cell[   12221] = 32'h8bbbc4d4;
    ram_cell[   12222] = 32'h0af1e2c0;
    ram_cell[   12223] = 32'h357700c5;
    ram_cell[   12224] = 32'h94fe29fa;
    ram_cell[   12225] = 32'he6487528;
    ram_cell[   12226] = 32'h32d76961;
    ram_cell[   12227] = 32'h7b9a10d2;
    ram_cell[   12228] = 32'h201af49d;
    ram_cell[   12229] = 32'hbe385573;
    ram_cell[   12230] = 32'h403685eb;
    ram_cell[   12231] = 32'h9f2f7916;
    ram_cell[   12232] = 32'h347b7b28;
    ram_cell[   12233] = 32'h5fa8523a;
    ram_cell[   12234] = 32'h03407989;
    ram_cell[   12235] = 32'h8ae5b64e;
    ram_cell[   12236] = 32'h7ab4cb6e;
    ram_cell[   12237] = 32'h550230df;
    ram_cell[   12238] = 32'hd58dd897;
    ram_cell[   12239] = 32'hd70b3f6d;
    ram_cell[   12240] = 32'h1d0a5738;
    ram_cell[   12241] = 32'h5abdbdcb;
    ram_cell[   12242] = 32'hc89d3978;
    ram_cell[   12243] = 32'h76ab8edc;
    ram_cell[   12244] = 32'h8f067590;
    ram_cell[   12245] = 32'he4dfe51c;
    ram_cell[   12246] = 32'h80e104f1;
    ram_cell[   12247] = 32'h7af887dd;
    ram_cell[   12248] = 32'hfd599914;
    ram_cell[   12249] = 32'hd163872e;
    ram_cell[   12250] = 32'habe84d12;
    ram_cell[   12251] = 32'h4f94489f;
    ram_cell[   12252] = 32'h9c447854;
    ram_cell[   12253] = 32'hc33a8ecf;
    ram_cell[   12254] = 32'he3394b27;
    ram_cell[   12255] = 32'h3446c482;
    ram_cell[   12256] = 32'haae41f65;
    ram_cell[   12257] = 32'hf80f603e;
    ram_cell[   12258] = 32'h40dc3727;
    ram_cell[   12259] = 32'hf4f5ba33;
    ram_cell[   12260] = 32'he06db2d0;
    ram_cell[   12261] = 32'h332e3c31;
    ram_cell[   12262] = 32'he88c4152;
    ram_cell[   12263] = 32'h4546ff8b;
    ram_cell[   12264] = 32'haab42a88;
    ram_cell[   12265] = 32'h8b1be1de;
    ram_cell[   12266] = 32'h42ef7997;
    ram_cell[   12267] = 32'hf5ac362e;
    ram_cell[   12268] = 32'h5b3cc95b;
    ram_cell[   12269] = 32'h07cee79e;
    ram_cell[   12270] = 32'h8678ac32;
    ram_cell[   12271] = 32'hefd34f18;
    ram_cell[   12272] = 32'ha98b9b72;
    ram_cell[   12273] = 32'h97f6d92c;
    ram_cell[   12274] = 32'he60bcbcf;
    ram_cell[   12275] = 32'h6f545889;
    ram_cell[   12276] = 32'h8cffa5f2;
    ram_cell[   12277] = 32'h9b13035b;
    ram_cell[   12278] = 32'hf2940e6d;
    ram_cell[   12279] = 32'hcb810daa;
    ram_cell[   12280] = 32'hed91cf5b;
    ram_cell[   12281] = 32'hb7c0735b;
    ram_cell[   12282] = 32'h014c7124;
    ram_cell[   12283] = 32'h4347b776;
    ram_cell[   12284] = 32'h5e57e2f0;
    ram_cell[   12285] = 32'h8ee43bd9;
    ram_cell[   12286] = 32'h76864859;
    ram_cell[   12287] = 32'h99196678;
end

endmodule

