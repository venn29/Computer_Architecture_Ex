
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hc8742729;
    ram_cell[       1] = 32'h0;  // 32'hb44b5467;
    ram_cell[       2] = 32'h0;  // 32'hcb714f65;
    ram_cell[       3] = 32'h0;  // 32'h3d172c8e;
    ram_cell[       4] = 32'h0;  // 32'h43ea6a7f;
    ram_cell[       5] = 32'h0;  // 32'h42a5a64a;
    ram_cell[       6] = 32'h0;  // 32'h8fc97f0b;
    ram_cell[       7] = 32'h0;  // 32'hb4eaf273;
    ram_cell[       8] = 32'h0;  // 32'h11dbef86;
    ram_cell[       9] = 32'h0;  // 32'h03fa4828;
    ram_cell[      10] = 32'h0;  // 32'h867d31bf;
    ram_cell[      11] = 32'h0;  // 32'h839fc462;
    ram_cell[      12] = 32'h0;  // 32'hfa1cec32;
    ram_cell[      13] = 32'h0;  // 32'h751bf489;
    ram_cell[      14] = 32'h0;  // 32'hb6de3a9e;
    ram_cell[      15] = 32'h0;  // 32'h2044f4e8;
    ram_cell[      16] = 32'h0;  // 32'hcc2b2738;
    ram_cell[      17] = 32'h0;  // 32'h1dc26fd8;
    ram_cell[      18] = 32'h0;  // 32'h6d14a405;
    ram_cell[      19] = 32'h0;  // 32'h0b7ca264;
    ram_cell[      20] = 32'h0;  // 32'h3f3158b1;
    ram_cell[      21] = 32'h0;  // 32'h156e0988;
    ram_cell[      22] = 32'h0;  // 32'h5cb7a295;
    ram_cell[      23] = 32'h0;  // 32'h54b92301;
    ram_cell[      24] = 32'h0;  // 32'h202c2596;
    ram_cell[      25] = 32'h0;  // 32'h00c510e6;
    ram_cell[      26] = 32'h0;  // 32'hfe5ef80a;
    ram_cell[      27] = 32'h0;  // 32'hd82d41cd;
    ram_cell[      28] = 32'h0;  // 32'h0e5958e1;
    ram_cell[      29] = 32'h0;  // 32'h16ca0c10;
    ram_cell[      30] = 32'h0;  // 32'hde8aec8f;
    ram_cell[      31] = 32'h0;  // 32'h35da2bac;
    ram_cell[      32] = 32'h0;  // 32'h369ee5b6;
    ram_cell[      33] = 32'h0;  // 32'h7b602b99;
    ram_cell[      34] = 32'h0;  // 32'hbd6571e2;
    ram_cell[      35] = 32'h0;  // 32'h5d66f17a;
    ram_cell[      36] = 32'h0;  // 32'hf427e8ec;
    ram_cell[      37] = 32'h0;  // 32'hb9c8fb57;
    ram_cell[      38] = 32'h0;  // 32'h240f3858;
    ram_cell[      39] = 32'h0;  // 32'h5e9657e8;
    ram_cell[      40] = 32'h0;  // 32'h3e63353e;
    ram_cell[      41] = 32'h0;  // 32'h5ad43e0c;
    ram_cell[      42] = 32'h0;  // 32'h547d37ec;
    ram_cell[      43] = 32'h0;  // 32'h772feac3;
    ram_cell[      44] = 32'h0;  // 32'h0a6ee2c0;
    ram_cell[      45] = 32'h0;  // 32'hce286adc;
    ram_cell[      46] = 32'h0;  // 32'h63d5c8ac;
    ram_cell[      47] = 32'h0;  // 32'h4d962a71;
    ram_cell[      48] = 32'h0;  // 32'hf8e5357a;
    ram_cell[      49] = 32'h0;  // 32'h5debbf4b;
    ram_cell[      50] = 32'h0;  // 32'h79695841;
    ram_cell[      51] = 32'h0;  // 32'ha12c8725;
    ram_cell[      52] = 32'h0;  // 32'h3870fca7;
    ram_cell[      53] = 32'h0;  // 32'h29bc1947;
    ram_cell[      54] = 32'h0;  // 32'h192542a4;
    ram_cell[      55] = 32'h0;  // 32'h2e47514a;
    ram_cell[      56] = 32'h0;  // 32'heb6a0c03;
    ram_cell[      57] = 32'h0;  // 32'h9847170d;
    ram_cell[      58] = 32'h0;  // 32'h107288aa;
    ram_cell[      59] = 32'h0;  // 32'h5a1a4171;
    ram_cell[      60] = 32'h0;  // 32'h49074f4e;
    ram_cell[      61] = 32'h0;  // 32'h728bdad4;
    ram_cell[      62] = 32'h0;  // 32'h6f16d0f9;
    ram_cell[      63] = 32'h0;  // 32'h77365d07;
    ram_cell[      64] = 32'h0;  // 32'hf1ebab94;
    ram_cell[      65] = 32'h0;  // 32'h09926be7;
    ram_cell[      66] = 32'h0;  // 32'h1ac005ac;
    ram_cell[      67] = 32'h0;  // 32'h6aa6bccc;
    ram_cell[      68] = 32'h0;  // 32'hda4ceba4;
    ram_cell[      69] = 32'h0;  // 32'h44d4b289;
    ram_cell[      70] = 32'h0;  // 32'hd0a6eb93;
    ram_cell[      71] = 32'h0;  // 32'hdde4939d;
    ram_cell[      72] = 32'h0;  // 32'hb84f9747;
    ram_cell[      73] = 32'h0;  // 32'h2a57151d;
    ram_cell[      74] = 32'h0;  // 32'h353b9f00;
    ram_cell[      75] = 32'h0;  // 32'h922f2778;
    ram_cell[      76] = 32'h0;  // 32'h3f6f42b6;
    ram_cell[      77] = 32'h0;  // 32'hff80c873;
    ram_cell[      78] = 32'h0;  // 32'h5cb85244;
    ram_cell[      79] = 32'h0;  // 32'h42017f8a;
    ram_cell[      80] = 32'h0;  // 32'h313fda42;
    ram_cell[      81] = 32'h0;  // 32'h04582cb6;
    ram_cell[      82] = 32'h0;  // 32'hddaa013b;
    ram_cell[      83] = 32'h0;  // 32'hc927adb9;
    ram_cell[      84] = 32'h0;  // 32'hfecb4d20;
    ram_cell[      85] = 32'h0;  // 32'he8133dd4;
    ram_cell[      86] = 32'h0;  // 32'h83e60aa5;
    ram_cell[      87] = 32'h0;  // 32'h95f8d6a5;
    ram_cell[      88] = 32'h0;  // 32'hb8bf69d4;
    ram_cell[      89] = 32'h0;  // 32'hb4114e08;
    ram_cell[      90] = 32'h0;  // 32'ha0205d7f;
    ram_cell[      91] = 32'h0;  // 32'h471444cc;
    ram_cell[      92] = 32'h0;  // 32'hc9de6b79;
    ram_cell[      93] = 32'h0;  // 32'h35d446d9;
    ram_cell[      94] = 32'h0;  // 32'h74b5673c;
    ram_cell[      95] = 32'h0;  // 32'hfca9ad97;
    ram_cell[      96] = 32'h0;  // 32'h1989f9af;
    ram_cell[      97] = 32'h0;  // 32'hd987e186;
    ram_cell[      98] = 32'h0;  // 32'h615611c5;
    ram_cell[      99] = 32'h0;  // 32'h4068c5da;
    ram_cell[     100] = 32'h0;  // 32'h3a45372d;
    ram_cell[     101] = 32'h0;  // 32'hfffc1b5c;
    ram_cell[     102] = 32'h0;  // 32'h8da4b6fc;
    ram_cell[     103] = 32'h0;  // 32'h4fbd32a4;
    ram_cell[     104] = 32'h0;  // 32'h67281444;
    ram_cell[     105] = 32'h0;  // 32'hcbf02c00;
    ram_cell[     106] = 32'h0;  // 32'hf2066377;
    ram_cell[     107] = 32'h0;  // 32'h6b3c5d41;
    ram_cell[     108] = 32'h0;  // 32'hb9b7b0da;
    ram_cell[     109] = 32'h0;  // 32'h642a42df;
    ram_cell[     110] = 32'h0;  // 32'h5b94a7cd;
    ram_cell[     111] = 32'h0;  // 32'h732cbe09;
    ram_cell[     112] = 32'h0;  // 32'h811be51e;
    ram_cell[     113] = 32'h0;  // 32'h10bb4be6;
    ram_cell[     114] = 32'h0;  // 32'h1548d2f3;
    ram_cell[     115] = 32'h0;  // 32'h072826db;
    ram_cell[     116] = 32'h0;  // 32'h5e93fe75;
    ram_cell[     117] = 32'h0;  // 32'hf8341929;
    ram_cell[     118] = 32'h0;  // 32'hd4380251;
    ram_cell[     119] = 32'h0;  // 32'h7b605f39;
    ram_cell[     120] = 32'h0;  // 32'h48b903f4;
    ram_cell[     121] = 32'h0;  // 32'hf7e99d5b;
    ram_cell[     122] = 32'h0;  // 32'hfe5c29cc;
    ram_cell[     123] = 32'h0;  // 32'h0aa5de3d;
    ram_cell[     124] = 32'h0;  // 32'h360c0702;
    ram_cell[     125] = 32'h0;  // 32'hc5238cf6;
    ram_cell[     126] = 32'h0;  // 32'hc9ebbb66;
    ram_cell[     127] = 32'h0;  // 32'h2b845981;
    ram_cell[     128] = 32'h0;  // 32'he263312f;
    ram_cell[     129] = 32'h0;  // 32'h84ccc853;
    ram_cell[     130] = 32'h0;  // 32'hf45d18f4;
    ram_cell[     131] = 32'h0;  // 32'h3700ca7c;
    ram_cell[     132] = 32'h0;  // 32'h1d97be76;
    ram_cell[     133] = 32'h0;  // 32'hae0ceb54;
    ram_cell[     134] = 32'h0;  // 32'hc866f9e0;
    ram_cell[     135] = 32'h0;  // 32'hbb76b464;
    ram_cell[     136] = 32'h0;  // 32'hbc1cc7aa;
    ram_cell[     137] = 32'h0;  // 32'h13deffa0;
    ram_cell[     138] = 32'h0;  // 32'hfb6466e4;
    ram_cell[     139] = 32'h0;  // 32'h7eb4f59c;
    ram_cell[     140] = 32'h0;  // 32'hada82af2;
    ram_cell[     141] = 32'h0;  // 32'hafef981d;
    ram_cell[     142] = 32'h0;  // 32'haa5910d9;
    ram_cell[     143] = 32'h0;  // 32'h889f437e;
    ram_cell[     144] = 32'h0;  // 32'h9407a5cf;
    ram_cell[     145] = 32'h0;  // 32'hfdd1884b;
    ram_cell[     146] = 32'h0;  // 32'h5bedec40;
    ram_cell[     147] = 32'h0;  // 32'h828d234d;
    ram_cell[     148] = 32'h0;  // 32'h17f0352a;
    ram_cell[     149] = 32'h0;  // 32'haa22bf04;
    ram_cell[     150] = 32'h0;  // 32'h10c9d301;
    ram_cell[     151] = 32'h0;  // 32'hf025bfb2;
    ram_cell[     152] = 32'h0;  // 32'hfca1ff43;
    ram_cell[     153] = 32'h0;  // 32'h2c8722ec;
    ram_cell[     154] = 32'h0;  // 32'hd073943d;
    ram_cell[     155] = 32'h0;  // 32'hb9f5dc7f;
    ram_cell[     156] = 32'h0;  // 32'hf04d273b;
    ram_cell[     157] = 32'h0;  // 32'h595b2a5e;
    ram_cell[     158] = 32'h0;  // 32'h07ca363d;
    ram_cell[     159] = 32'h0;  // 32'h2db03d64;
    ram_cell[     160] = 32'h0;  // 32'h4a67038b;
    ram_cell[     161] = 32'h0;  // 32'h11ddea7e;
    ram_cell[     162] = 32'h0;  // 32'h8740f68d;
    ram_cell[     163] = 32'h0;  // 32'h9b334255;
    ram_cell[     164] = 32'h0;  // 32'h09e8fa82;
    ram_cell[     165] = 32'h0;  // 32'h89a4487d;
    ram_cell[     166] = 32'h0;  // 32'hce94c8c3;
    ram_cell[     167] = 32'h0;  // 32'ha90019e0;
    ram_cell[     168] = 32'h0;  // 32'h009343a5;
    ram_cell[     169] = 32'h0;  // 32'h5474bc40;
    ram_cell[     170] = 32'h0;  // 32'h49972940;
    ram_cell[     171] = 32'h0;  // 32'h83a7e133;
    ram_cell[     172] = 32'h0;  // 32'h513e978b;
    ram_cell[     173] = 32'h0;  // 32'h96fcb0fa;
    ram_cell[     174] = 32'h0;  // 32'haddbe85a;
    ram_cell[     175] = 32'h0;  // 32'hf51920af;
    ram_cell[     176] = 32'h0;  // 32'h1edb2fc9;
    ram_cell[     177] = 32'h0;  // 32'h3b43c89e;
    ram_cell[     178] = 32'h0;  // 32'haff63188;
    ram_cell[     179] = 32'h0;  // 32'hc0555f64;
    ram_cell[     180] = 32'h0;  // 32'h97cbae36;
    ram_cell[     181] = 32'h0;  // 32'h5ad36e20;
    ram_cell[     182] = 32'h0;  // 32'he3db5042;
    ram_cell[     183] = 32'h0;  // 32'h9fd20c66;
    ram_cell[     184] = 32'h0;  // 32'ha78cf01f;
    ram_cell[     185] = 32'h0;  // 32'h59632d7b;
    ram_cell[     186] = 32'h0;  // 32'h5f689636;
    ram_cell[     187] = 32'h0;  // 32'h6ddb1aef;
    ram_cell[     188] = 32'h0;  // 32'hfbb2d210;
    ram_cell[     189] = 32'h0;  // 32'hc20ee16d;
    ram_cell[     190] = 32'h0;  // 32'h7a0d7b78;
    ram_cell[     191] = 32'h0;  // 32'h187b97aa;
    ram_cell[     192] = 32'h0;  // 32'ha2e9e213;
    ram_cell[     193] = 32'h0;  // 32'h61f4dc14;
    ram_cell[     194] = 32'h0;  // 32'hdf566017;
    ram_cell[     195] = 32'h0;  // 32'hed19403c;
    ram_cell[     196] = 32'h0;  // 32'h02f08141;
    ram_cell[     197] = 32'h0;  // 32'h9be3fa27;
    ram_cell[     198] = 32'h0;  // 32'h66ceda34;
    ram_cell[     199] = 32'h0;  // 32'h86c5b39a;
    ram_cell[     200] = 32'h0;  // 32'hc81cb35f;
    ram_cell[     201] = 32'h0;  // 32'heb66ae46;
    ram_cell[     202] = 32'h0;  // 32'hf317836f;
    ram_cell[     203] = 32'h0;  // 32'h66c9983d;
    ram_cell[     204] = 32'h0;  // 32'h997f14b7;
    ram_cell[     205] = 32'h0;  // 32'h0bcfce7e;
    ram_cell[     206] = 32'h0;  // 32'h57fad9c1;
    ram_cell[     207] = 32'h0;  // 32'hf693df4e;
    ram_cell[     208] = 32'h0;  // 32'h72c6e2ac;
    ram_cell[     209] = 32'h0;  // 32'h45fe2d43;
    ram_cell[     210] = 32'h0;  // 32'h52886c76;
    ram_cell[     211] = 32'h0;  // 32'h66f05f67;
    ram_cell[     212] = 32'h0;  // 32'haf194783;
    ram_cell[     213] = 32'h0;  // 32'h565d6368;
    ram_cell[     214] = 32'h0;  // 32'haa7ddc22;
    ram_cell[     215] = 32'h0;  // 32'h34cd0631;
    ram_cell[     216] = 32'h0;  // 32'h7c033607;
    ram_cell[     217] = 32'h0;  // 32'hb99f9ddd;
    ram_cell[     218] = 32'h0;  // 32'h01734a88;
    ram_cell[     219] = 32'h0;  // 32'he820b0a8;
    ram_cell[     220] = 32'h0;  // 32'hab2d68b9;
    ram_cell[     221] = 32'h0;  // 32'h4906ae01;
    ram_cell[     222] = 32'h0;  // 32'had914160;
    ram_cell[     223] = 32'h0;  // 32'hec5f0e92;
    ram_cell[     224] = 32'h0;  // 32'hfdedaf10;
    ram_cell[     225] = 32'h0;  // 32'ha8c864b8;
    ram_cell[     226] = 32'h0;  // 32'h570933de;
    ram_cell[     227] = 32'h0;  // 32'h3cb9cc1d;
    ram_cell[     228] = 32'h0;  // 32'h9a611dce;
    ram_cell[     229] = 32'h0;  // 32'h6c90a0d4;
    ram_cell[     230] = 32'h0;  // 32'hbc668a4a;
    ram_cell[     231] = 32'h0;  // 32'h5a515151;
    ram_cell[     232] = 32'h0;  // 32'hbacd34e9;
    ram_cell[     233] = 32'h0;  // 32'hf37cd221;
    ram_cell[     234] = 32'h0;  // 32'h0df7dc60;
    ram_cell[     235] = 32'h0;  // 32'ha5fa8d7b;
    ram_cell[     236] = 32'h0;  // 32'h1956032a;
    ram_cell[     237] = 32'h0;  // 32'hd82336b1;
    ram_cell[     238] = 32'h0;  // 32'h3ac4bf16;
    ram_cell[     239] = 32'h0;  // 32'he4e35693;
    ram_cell[     240] = 32'h0;  // 32'h96755e74;
    ram_cell[     241] = 32'h0;  // 32'ha1215197;
    ram_cell[     242] = 32'h0;  // 32'h6d231197;
    ram_cell[     243] = 32'h0;  // 32'h2b374abd;
    ram_cell[     244] = 32'h0;  // 32'he23f3763;
    ram_cell[     245] = 32'h0;  // 32'h82819494;
    ram_cell[     246] = 32'h0;  // 32'hea563a96;
    ram_cell[     247] = 32'h0;  // 32'h30683771;
    ram_cell[     248] = 32'h0;  // 32'h1070613a;
    ram_cell[     249] = 32'h0;  // 32'hc69880b6;
    ram_cell[     250] = 32'h0;  // 32'hdc3c673f;
    ram_cell[     251] = 32'h0;  // 32'hed39cc99;
    ram_cell[     252] = 32'h0;  // 32'hd87c19cb;
    ram_cell[     253] = 32'h0;  // 32'heabccef4;
    ram_cell[     254] = 32'h0;  // 32'h265ae689;
    ram_cell[     255] = 32'h0;  // 32'h1c50f057;
    ram_cell[     256] = 32'h0;  // 32'ha2a842bc;
    ram_cell[     257] = 32'h0;  // 32'hf3aec7e9;
    ram_cell[     258] = 32'h0;  // 32'h82f4ad11;
    ram_cell[     259] = 32'h0;  // 32'hbf134ca9;
    ram_cell[     260] = 32'h0;  // 32'h24d668b8;
    ram_cell[     261] = 32'h0;  // 32'h9b7b247a;
    ram_cell[     262] = 32'h0;  // 32'hc80292be;
    ram_cell[     263] = 32'h0;  // 32'h7619b1c5;
    ram_cell[     264] = 32'h0;  // 32'h7a3cdd0d;
    ram_cell[     265] = 32'h0;  // 32'h9b07a5b8;
    ram_cell[     266] = 32'h0;  // 32'h87b3dc19;
    ram_cell[     267] = 32'h0;  // 32'h5838d3f9;
    ram_cell[     268] = 32'h0;  // 32'hbf898bab;
    ram_cell[     269] = 32'h0;  // 32'h1eccf2df;
    ram_cell[     270] = 32'h0;  // 32'h4ec417d4;
    ram_cell[     271] = 32'h0;  // 32'h4704c997;
    ram_cell[     272] = 32'h0;  // 32'h83c4d87a;
    ram_cell[     273] = 32'h0;  // 32'hca41a82c;
    ram_cell[     274] = 32'h0;  // 32'h269371d0;
    ram_cell[     275] = 32'h0;  // 32'hb3f3afc2;
    ram_cell[     276] = 32'h0;  // 32'h969b9fe9;
    ram_cell[     277] = 32'h0;  // 32'h491ad5bd;
    ram_cell[     278] = 32'h0;  // 32'h5d9ec639;
    ram_cell[     279] = 32'h0;  // 32'hb207b691;
    ram_cell[     280] = 32'h0;  // 32'h0afbb90a;
    ram_cell[     281] = 32'h0;  // 32'hb3a39971;
    ram_cell[     282] = 32'h0;  // 32'h43b29612;
    ram_cell[     283] = 32'h0;  // 32'hd3de650a;
    ram_cell[     284] = 32'h0;  // 32'h341ebf37;
    ram_cell[     285] = 32'h0;  // 32'h734a1ec9;
    ram_cell[     286] = 32'h0;  // 32'h5398d894;
    ram_cell[     287] = 32'h0;  // 32'hd9803715;
    ram_cell[     288] = 32'h0;  // 32'hb8f68c45;
    ram_cell[     289] = 32'h0;  // 32'h4b0ce352;
    ram_cell[     290] = 32'h0;  // 32'h973bc33c;
    ram_cell[     291] = 32'h0;  // 32'hf8aa92cb;
    ram_cell[     292] = 32'h0;  // 32'h61b6442c;
    ram_cell[     293] = 32'h0;  // 32'h010e4c3a;
    ram_cell[     294] = 32'h0;  // 32'h5d78e307;
    ram_cell[     295] = 32'h0;  // 32'hd7dcad64;
    ram_cell[     296] = 32'h0;  // 32'h398279b8;
    ram_cell[     297] = 32'h0;  // 32'h58dee8ad;
    ram_cell[     298] = 32'h0;  // 32'ha262aee2;
    ram_cell[     299] = 32'h0;  // 32'ha7dfa6b3;
    ram_cell[     300] = 32'h0;  // 32'ha2da6889;
    ram_cell[     301] = 32'h0;  // 32'h8c3cebaf;
    ram_cell[     302] = 32'h0;  // 32'h1261423b;
    ram_cell[     303] = 32'h0;  // 32'h2c33534e;
    ram_cell[     304] = 32'h0;  // 32'h23e50d20;
    ram_cell[     305] = 32'h0;  // 32'h401a63b4;
    ram_cell[     306] = 32'h0;  // 32'h94f3ea29;
    ram_cell[     307] = 32'h0;  // 32'hcf0b402f;
    ram_cell[     308] = 32'h0;  // 32'hf8bfe1ff;
    ram_cell[     309] = 32'h0;  // 32'h36db66ce;
    ram_cell[     310] = 32'h0;  // 32'hac5e3dc9;
    ram_cell[     311] = 32'h0;  // 32'h0432c1f9;
    ram_cell[     312] = 32'h0;  // 32'hb8971a14;
    ram_cell[     313] = 32'h0;  // 32'h66bf2331;
    ram_cell[     314] = 32'h0;  // 32'hb3f7e76c;
    ram_cell[     315] = 32'h0;  // 32'hd148bb22;
    ram_cell[     316] = 32'h0;  // 32'h46bf9469;
    ram_cell[     317] = 32'h0;  // 32'ha112c306;
    ram_cell[     318] = 32'h0;  // 32'hdbc8192b;
    ram_cell[     319] = 32'h0;  // 32'hb3012728;
    ram_cell[     320] = 32'h0;  // 32'h9cf244f7;
    ram_cell[     321] = 32'h0;  // 32'hb46e023e;
    ram_cell[     322] = 32'h0;  // 32'he518594f;
    ram_cell[     323] = 32'h0;  // 32'h92d6ad14;
    ram_cell[     324] = 32'h0;  // 32'h27c84d5e;
    ram_cell[     325] = 32'h0;  // 32'ha4fe0a1a;
    ram_cell[     326] = 32'h0;  // 32'h83616910;
    ram_cell[     327] = 32'h0;  // 32'h2d352ad7;
    ram_cell[     328] = 32'h0;  // 32'h75336073;
    ram_cell[     329] = 32'h0;  // 32'h6b2f8632;
    ram_cell[     330] = 32'h0;  // 32'h535040a3;
    ram_cell[     331] = 32'h0;  // 32'hb1e1800a;
    ram_cell[     332] = 32'h0;  // 32'h13332cff;
    ram_cell[     333] = 32'h0;  // 32'hf303ad7b;
    ram_cell[     334] = 32'h0;  // 32'h77bb0aec;
    ram_cell[     335] = 32'h0;  // 32'hc9bfde75;
    ram_cell[     336] = 32'h0;  // 32'h9bb66857;
    ram_cell[     337] = 32'h0;  // 32'h3b3eea06;
    ram_cell[     338] = 32'h0;  // 32'hbe38addd;
    ram_cell[     339] = 32'h0;  // 32'hce06b9ac;
    ram_cell[     340] = 32'h0;  // 32'he6f959aa;
    ram_cell[     341] = 32'h0;  // 32'haa979495;
    ram_cell[     342] = 32'h0;  // 32'hec82d329;
    ram_cell[     343] = 32'h0;  // 32'he49b876d;
    ram_cell[     344] = 32'h0;  // 32'h320d8bfa;
    ram_cell[     345] = 32'h0;  // 32'h43a88bd8;
    ram_cell[     346] = 32'h0;  // 32'h6722000a;
    ram_cell[     347] = 32'h0;  // 32'h72ab7dfb;
    ram_cell[     348] = 32'h0;  // 32'h156c75ce;
    ram_cell[     349] = 32'h0;  // 32'hd90ca22c;
    ram_cell[     350] = 32'h0;  // 32'h55210e6a;
    ram_cell[     351] = 32'h0;  // 32'h9d227dec;
    ram_cell[     352] = 32'h0;  // 32'h322818ab;
    ram_cell[     353] = 32'h0;  // 32'h861e5331;
    ram_cell[     354] = 32'h0;  // 32'hf19f077c;
    ram_cell[     355] = 32'h0;  // 32'hd2a1c6e0;
    ram_cell[     356] = 32'h0;  // 32'h00af9c90;
    ram_cell[     357] = 32'h0;  // 32'h142aa3e8;
    ram_cell[     358] = 32'h0;  // 32'hc75efbc4;
    ram_cell[     359] = 32'h0;  // 32'hc88c55d2;
    ram_cell[     360] = 32'h0;  // 32'h41d8e22d;
    ram_cell[     361] = 32'h0;  // 32'hfd28d534;
    ram_cell[     362] = 32'h0;  // 32'h235ab62c;
    ram_cell[     363] = 32'h0;  // 32'h9341076a;
    ram_cell[     364] = 32'h0;  // 32'h9bc5de92;
    ram_cell[     365] = 32'h0;  // 32'h46b50aa4;
    ram_cell[     366] = 32'h0;  // 32'h7b60be23;
    ram_cell[     367] = 32'h0;  // 32'hb77bcace;
    ram_cell[     368] = 32'h0;  // 32'h65dcbf0e;
    ram_cell[     369] = 32'h0;  // 32'h22507340;
    ram_cell[     370] = 32'h0;  // 32'hc73f161a;
    ram_cell[     371] = 32'h0;  // 32'h66803daf;
    ram_cell[     372] = 32'h0;  // 32'h2437b2b9;
    ram_cell[     373] = 32'h0;  // 32'h361cdc29;
    ram_cell[     374] = 32'h0;  // 32'hfc732ea9;
    ram_cell[     375] = 32'h0;  // 32'h1a64d8d4;
    ram_cell[     376] = 32'h0;  // 32'h78251f4a;
    ram_cell[     377] = 32'h0;  // 32'h200f48b7;
    ram_cell[     378] = 32'h0;  // 32'h46b552ab;
    ram_cell[     379] = 32'h0;  // 32'hc0c8cccb;
    ram_cell[     380] = 32'h0;  // 32'h0c9f8eb9;
    ram_cell[     381] = 32'h0;  // 32'h3eead140;
    ram_cell[     382] = 32'h0;  // 32'h8e319a20;
    ram_cell[     383] = 32'h0;  // 32'h9f7f498e;
    ram_cell[     384] = 32'h0;  // 32'h7eb1ffcc;
    ram_cell[     385] = 32'h0;  // 32'h30e23778;
    ram_cell[     386] = 32'h0;  // 32'hd4d07f33;
    ram_cell[     387] = 32'h0;  // 32'h74d8e136;
    ram_cell[     388] = 32'h0;  // 32'hc699a8b4;
    ram_cell[     389] = 32'h0;  // 32'h1f42ff62;
    ram_cell[     390] = 32'h0;  // 32'ha368f7e0;
    ram_cell[     391] = 32'h0;  // 32'h48be6a4d;
    ram_cell[     392] = 32'h0;  // 32'h3ab54520;
    ram_cell[     393] = 32'h0;  // 32'h64b913f7;
    ram_cell[     394] = 32'h0;  // 32'hf65e103d;
    ram_cell[     395] = 32'h0;  // 32'hbca5bb24;
    ram_cell[     396] = 32'h0;  // 32'h0880e351;
    ram_cell[     397] = 32'h0;  // 32'h85086df6;
    ram_cell[     398] = 32'h0;  // 32'hc955e3c5;
    ram_cell[     399] = 32'h0;  // 32'h3da187ce;
    ram_cell[     400] = 32'h0;  // 32'hc0f81522;
    ram_cell[     401] = 32'h0;  // 32'hf354ce18;
    ram_cell[     402] = 32'h0;  // 32'h22efdd53;
    ram_cell[     403] = 32'h0;  // 32'h52f07f9d;
    ram_cell[     404] = 32'h0;  // 32'h3bb2ef25;
    ram_cell[     405] = 32'h0;  // 32'he8b2ebb4;
    ram_cell[     406] = 32'h0;  // 32'haa653b0d;
    ram_cell[     407] = 32'h0;  // 32'h127c89fa;
    ram_cell[     408] = 32'h0;  // 32'h947365c2;
    ram_cell[     409] = 32'h0;  // 32'he38e8010;
    ram_cell[     410] = 32'h0;  // 32'hf75f5591;
    ram_cell[     411] = 32'h0;  // 32'hd4836af5;
    ram_cell[     412] = 32'h0;  // 32'hbdbc2158;
    ram_cell[     413] = 32'h0;  // 32'h61df1b9e;
    ram_cell[     414] = 32'h0;  // 32'h411d575a;
    ram_cell[     415] = 32'h0;  // 32'hb31cdff8;
    ram_cell[     416] = 32'h0;  // 32'h29d051eb;
    ram_cell[     417] = 32'h0;  // 32'hf1ec0979;
    ram_cell[     418] = 32'h0;  // 32'he2b2eaec;
    ram_cell[     419] = 32'h0;  // 32'h7af90f66;
    ram_cell[     420] = 32'h0;  // 32'h2f4f7bab;
    ram_cell[     421] = 32'h0;  // 32'h0f7763b7;
    ram_cell[     422] = 32'h0;  // 32'he3a0fd26;
    ram_cell[     423] = 32'h0;  // 32'h31642b28;
    ram_cell[     424] = 32'h0;  // 32'h50b7f1c6;
    ram_cell[     425] = 32'h0;  // 32'h5a8f9249;
    ram_cell[     426] = 32'h0;  // 32'h853054d4;
    ram_cell[     427] = 32'h0;  // 32'h060939e4;
    ram_cell[     428] = 32'h0;  // 32'hbe404ce0;
    ram_cell[     429] = 32'h0;  // 32'h3ec9dec6;
    ram_cell[     430] = 32'h0;  // 32'hd167c9d0;
    ram_cell[     431] = 32'h0;  // 32'h6ffb205f;
    ram_cell[     432] = 32'h0;  // 32'h13d965e1;
    ram_cell[     433] = 32'h0;  // 32'h57e63319;
    ram_cell[     434] = 32'h0;  // 32'hd7c17d7a;
    ram_cell[     435] = 32'h0;  // 32'hda76b538;
    ram_cell[     436] = 32'h0;  // 32'h2fb25c25;
    ram_cell[     437] = 32'h0;  // 32'ha7f29793;
    ram_cell[     438] = 32'h0;  // 32'h8661946d;
    ram_cell[     439] = 32'h0;  // 32'he504e500;
    ram_cell[     440] = 32'h0;  // 32'h3225a3a6;
    ram_cell[     441] = 32'h0;  // 32'h0bb756f9;
    ram_cell[     442] = 32'h0;  // 32'hc149c357;
    ram_cell[     443] = 32'h0;  // 32'h2bdb0691;
    ram_cell[     444] = 32'h0;  // 32'h9b7f62d1;
    ram_cell[     445] = 32'h0;  // 32'ha3ad12e6;
    ram_cell[     446] = 32'h0;  // 32'h58999438;
    ram_cell[     447] = 32'h0;  // 32'hd1f14760;
    ram_cell[     448] = 32'h0;  // 32'hca2ff92c;
    ram_cell[     449] = 32'h0;  // 32'h1df1815a;
    ram_cell[     450] = 32'h0;  // 32'hb4e36454;
    ram_cell[     451] = 32'h0;  // 32'hd5bdcd18;
    ram_cell[     452] = 32'h0;  // 32'h608aea87;
    ram_cell[     453] = 32'h0;  // 32'hc10b0ace;
    ram_cell[     454] = 32'h0;  // 32'h0d1b011e;
    ram_cell[     455] = 32'h0;  // 32'h5148b5c8;
    ram_cell[     456] = 32'h0;  // 32'hf92d9943;
    ram_cell[     457] = 32'h0;  // 32'h1b43966c;
    ram_cell[     458] = 32'h0;  // 32'h178b3ab0;
    ram_cell[     459] = 32'h0;  // 32'hd361f9c2;
    ram_cell[     460] = 32'h0;  // 32'hcf5fe749;
    ram_cell[     461] = 32'h0;  // 32'h7e96bf09;
    ram_cell[     462] = 32'h0;  // 32'h2a713d90;
    ram_cell[     463] = 32'h0;  // 32'ha60b953f;
    ram_cell[     464] = 32'h0;  // 32'hc476c4b1;
    ram_cell[     465] = 32'h0;  // 32'hab38e034;
    ram_cell[     466] = 32'h0;  // 32'h5d04a28a;
    ram_cell[     467] = 32'h0;  // 32'h6a170f6c;
    ram_cell[     468] = 32'h0;  // 32'h1bba1dbb;
    ram_cell[     469] = 32'h0;  // 32'hccdd41cb;
    ram_cell[     470] = 32'h0;  // 32'h2b6d4b8b;
    ram_cell[     471] = 32'h0;  // 32'h45468d5c;
    ram_cell[     472] = 32'h0;  // 32'hc070b0ec;
    ram_cell[     473] = 32'h0;  // 32'hc2aad5bc;
    ram_cell[     474] = 32'h0;  // 32'h345f8b02;
    ram_cell[     475] = 32'h0;  // 32'h53eb2731;
    ram_cell[     476] = 32'h0;  // 32'he832457e;
    ram_cell[     477] = 32'h0;  // 32'heda8a70a;
    ram_cell[     478] = 32'h0;  // 32'hd8c5d79d;
    ram_cell[     479] = 32'h0;  // 32'h0bbb7a37;
    ram_cell[     480] = 32'h0;  // 32'h22627e6e;
    ram_cell[     481] = 32'h0;  // 32'hbf89fcf5;
    ram_cell[     482] = 32'h0;  // 32'h808218f6;
    ram_cell[     483] = 32'h0;  // 32'hbbe62b40;
    ram_cell[     484] = 32'h0;  // 32'h70f04137;
    ram_cell[     485] = 32'h0;  // 32'h0ce6859e;
    ram_cell[     486] = 32'h0;  // 32'h2b3cc402;
    ram_cell[     487] = 32'h0;  // 32'ha31c22c1;
    ram_cell[     488] = 32'h0;  // 32'hf345d1b3;
    ram_cell[     489] = 32'h0;  // 32'he4e468f7;
    ram_cell[     490] = 32'h0;  // 32'hbdd2783d;
    ram_cell[     491] = 32'h0;  // 32'h4b63888e;
    ram_cell[     492] = 32'h0;  // 32'h0b212119;
    ram_cell[     493] = 32'h0;  // 32'h15913767;
    ram_cell[     494] = 32'h0;  // 32'h6469e49d;
    ram_cell[     495] = 32'h0;  // 32'h796f51df;
    ram_cell[     496] = 32'h0;  // 32'h341d9611;
    ram_cell[     497] = 32'h0;  // 32'h8520dcae;
    ram_cell[     498] = 32'h0;  // 32'h8c05a5d3;
    ram_cell[     499] = 32'h0;  // 32'h658c9e9e;
    ram_cell[     500] = 32'h0;  // 32'h61c5176c;
    ram_cell[     501] = 32'h0;  // 32'hde10c832;
    ram_cell[     502] = 32'h0;  // 32'hdd677bfc;
    ram_cell[     503] = 32'h0;  // 32'h8ce4195d;
    ram_cell[     504] = 32'h0;  // 32'hfc62ebbb;
    ram_cell[     505] = 32'h0;  // 32'h2b910ad3;
    ram_cell[     506] = 32'h0;  // 32'h9b28ae40;
    ram_cell[     507] = 32'h0;  // 32'hfa765132;
    ram_cell[     508] = 32'h0;  // 32'hf187839b;
    ram_cell[     509] = 32'h0;  // 32'h52c034c9;
    ram_cell[     510] = 32'h0;  // 32'h4fa288a3;
    ram_cell[     511] = 32'h0;  // 32'hfee41faf;
    ram_cell[     512] = 32'h0;  // 32'h322a8d81;
    ram_cell[     513] = 32'h0;  // 32'h3adf5408;
    ram_cell[     514] = 32'h0;  // 32'hdd067931;
    ram_cell[     515] = 32'h0;  // 32'ha2211a63;
    ram_cell[     516] = 32'h0;  // 32'h9854d9c6;
    ram_cell[     517] = 32'h0;  // 32'hdc47aefa;
    ram_cell[     518] = 32'h0;  // 32'h47b4059c;
    ram_cell[     519] = 32'h0;  // 32'hb27368bc;
    ram_cell[     520] = 32'h0;  // 32'h41c880b4;
    ram_cell[     521] = 32'h0;  // 32'h4a6889c7;
    ram_cell[     522] = 32'h0;  // 32'h61e21f2c;
    ram_cell[     523] = 32'h0;  // 32'h0c00ead3;
    ram_cell[     524] = 32'h0;  // 32'h724bb0b8;
    ram_cell[     525] = 32'h0;  // 32'h83cd27f3;
    ram_cell[     526] = 32'h0;  // 32'h7821debd;
    ram_cell[     527] = 32'h0;  // 32'hb0080d0d;
    ram_cell[     528] = 32'h0;  // 32'h4bdc43fc;
    ram_cell[     529] = 32'h0;  // 32'hc0d78969;
    ram_cell[     530] = 32'h0;  // 32'h565dbb6b;
    ram_cell[     531] = 32'h0;  // 32'hc9d2099c;
    ram_cell[     532] = 32'h0;  // 32'hc823132b;
    ram_cell[     533] = 32'h0;  // 32'h5770c335;
    ram_cell[     534] = 32'h0;  // 32'hdf95f3ba;
    ram_cell[     535] = 32'h0;  // 32'h1b5b564e;
    ram_cell[     536] = 32'h0;  // 32'h3b887fc1;
    ram_cell[     537] = 32'h0;  // 32'h1e0e63d3;
    ram_cell[     538] = 32'h0;  // 32'hc0a40535;
    ram_cell[     539] = 32'h0;  // 32'hc7bcd47c;
    ram_cell[     540] = 32'h0;  // 32'h61572cfe;
    ram_cell[     541] = 32'h0;  // 32'h011d3cd9;
    ram_cell[     542] = 32'h0;  // 32'h6f0e3947;
    ram_cell[     543] = 32'h0;  // 32'h73687783;
    ram_cell[     544] = 32'h0;  // 32'h1a55e098;
    ram_cell[     545] = 32'h0;  // 32'h56c97067;
    ram_cell[     546] = 32'h0;  // 32'h1d302aaa;
    ram_cell[     547] = 32'h0;  // 32'h3f8b78a7;
    ram_cell[     548] = 32'h0;  // 32'h802ce10d;
    ram_cell[     549] = 32'h0;  // 32'h0281a811;
    ram_cell[     550] = 32'h0;  // 32'h9c816533;
    ram_cell[     551] = 32'h0;  // 32'hb62747be;
    ram_cell[     552] = 32'h0;  // 32'h396d50e0;
    ram_cell[     553] = 32'h0;  // 32'hfb5aa37d;
    ram_cell[     554] = 32'h0;  // 32'hd59d7303;
    ram_cell[     555] = 32'h0;  // 32'h3d3bd25d;
    ram_cell[     556] = 32'h0;  // 32'hb9959362;
    ram_cell[     557] = 32'h0;  // 32'hb848261e;
    ram_cell[     558] = 32'h0;  // 32'hbb94bdca;
    ram_cell[     559] = 32'h0;  // 32'h9904b076;
    ram_cell[     560] = 32'h0;  // 32'h16dca012;
    ram_cell[     561] = 32'h0;  // 32'h7ffc2dcb;
    ram_cell[     562] = 32'h0;  // 32'h93b4efd0;
    ram_cell[     563] = 32'h0;  // 32'h47395ba8;
    ram_cell[     564] = 32'h0;  // 32'h38fa0705;
    ram_cell[     565] = 32'h0;  // 32'hc92e4b7c;
    ram_cell[     566] = 32'h0;  // 32'h7f5483eb;
    ram_cell[     567] = 32'h0;  // 32'hd57bfed5;
    ram_cell[     568] = 32'h0;  // 32'ha08f2087;
    ram_cell[     569] = 32'h0;  // 32'hccee7f0b;
    ram_cell[     570] = 32'h0;  // 32'h812d494b;
    ram_cell[     571] = 32'h0;  // 32'h34d7a531;
    ram_cell[     572] = 32'h0;  // 32'hc99c0b33;
    ram_cell[     573] = 32'h0;  // 32'h79736fb0;
    ram_cell[     574] = 32'h0;  // 32'h6298128b;
    ram_cell[     575] = 32'h0;  // 32'h71069af6;
    ram_cell[     576] = 32'h0;  // 32'hcb31c723;
    ram_cell[     577] = 32'h0;  // 32'h5c1a2dfd;
    ram_cell[     578] = 32'h0;  // 32'ha5364ef2;
    ram_cell[     579] = 32'h0;  // 32'hd7ec423a;
    ram_cell[     580] = 32'h0;  // 32'h63b7658a;
    ram_cell[     581] = 32'h0;  // 32'h8beaba5b;
    ram_cell[     582] = 32'h0;  // 32'h68b2c2d6;
    ram_cell[     583] = 32'h0;  // 32'hc777d860;
    ram_cell[     584] = 32'h0;  // 32'h33272d2e;
    ram_cell[     585] = 32'h0;  // 32'h87a36ae8;
    ram_cell[     586] = 32'h0;  // 32'h52e47124;
    ram_cell[     587] = 32'h0;  // 32'h7151343b;
    ram_cell[     588] = 32'h0;  // 32'h5b6cb8ce;
    ram_cell[     589] = 32'h0;  // 32'hfc3f916e;
    ram_cell[     590] = 32'h0;  // 32'hcfef2848;
    ram_cell[     591] = 32'h0;  // 32'hdb7e545e;
    ram_cell[     592] = 32'h0;  // 32'h40acd1f5;
    ram_cell[     593] = 32'h0;  // 32'hda752383;
    ram_cell[     594] = 32'h0;  // 32'hfeb53f1e;
    ram_cell[     595] = 32'h0;  // 32'h0ecf40bd;
    ram_cell[     596] = 32'h0;  // 32'h7cf28026;
    ram_cell[     597] = 32'h0;  // 32'ha844683b;
    ram_cell[     598] = 32'h0;  // 32'ha8509cae;
    ram_cell[     599] = 32'h0;  // 32'h9a8838e8;
    ram_cell[     600] = 32'h0;  // 32'hc0479b38;
    ram_cell[     601] = 32'h0;  // 32'hbc2d2609;
    ram_cell[     602] = 32'h0;  // 32'h290dde29;
    ram_cell[     603] = 32'h0;  // 32'hbd95b02d;
    ram_cell[     604] = 32'h0;  // 32'hfbdeb470;
    ram_cell[     605] = 32'h0;  // 32'h9eb7ca18;
    ram_cell[     606] = 32'h0;  // 32'hc05c71b6;
    ram_cell[     607] = 32'h0;  // 32'hb81b06b9;
    ram_cell[     608] = 32'h0;  // 32'h0c7c8d88;
    ram_cell[     609] = 32'h0;  // 32'he6339369;
    ram_cell[     610] = 32'h0;  // 32'hc1650153;
    ram_cell[     611] = 32'h0;  // 32'hb948a366;
    ram_cell[     612] = 32'h0;  // 32'h60d94f0b;
    ram_cell[     613] = 32'h0;  // 32'h6f649b91;
    ram_cell[     614] = 32'h0;  // 32'h60c9b93e;
    ram_cell[     615] = 32'h0;  // 32'hb8c64ef9;
    ram_cell[     616] = 32'h0;  // 32'h3da0b577;
    ram_cell[     617] = 32'h0;  // 32'hcad55da7;
    ram_cell[     618] = 32'h0;  // 32'h21bcbf1d;
    ram_cell[     619] = 32'h0;  // 32'hb91d51a6;
    ram_cell[     620] = 32'h0;  // 32'h82793f81;
    ram_cell[     621] = 32'h0;  // 32'ha77636af;
    ram_cell[     622] = 32'h0;  // 32'h5fef737d;
    ram_cell[     623] = 32'h0;  // 32'h178a5d27;
    ram_cell[     624] = 32'h0;  // 32'h2bb862c6;
    ram_cell[     625] = 32'h0;  // 32'h29818f1c;
    ram_cell[     626] = 32'h0;  // 32'h3c497c2c;
    ram_cell[     627] = 32'h0;  // 32'h964ffa79;
    ram_cell[     628] = 32'h0;  // 32'h894b100a;
    ram_cell[     629] = 32'h0;  // 32'h605a24df;
    ram_cell[     630] = 32'h0;  // 32'hd0f2aacf;
    ram_cell[     631] = 32'h0;  // 32'hd075e2cf;
    ram_cell[     632] = 32'h0;  // 32'he27a628c;
    ram_cell[     633] = 32'h0;  // 32'habdf66a3;
    ram_cell[     634] = 32'h0;  // 32'hc4a1a4a4;
    ram_cell[     635] = 32'h0;  // 32'hf54e5c5c;
    ram_cell[     636] = 32'h0;  // 32'hd35d8647;
    ram_cell[     637] = 32'h0;  // 32'hd8613611;
    ram_cell[     638] = 32'h0;  // 32'h2cb27735;
    ram_cell[     639] = 32'h0;  // 32'hb7927a82;
    ram_cell[     640] = 32'h0;  // 32'h0f7416e5;
    ram_cell[     641] = 32'h0;  // 32'h5f2ecd57;
    ram_cell[     642] = 32'h0;  // 32'h67344f07;
    ram_cell[     643] = 32'h0;  // 32'hd9e57882;
    ram_cell[     644] = 32'h0;  // 32'ha31b2387;
    ram_cell[     645] = 32'h0;  // 32'hd89bbf6a;
    ram_cell[     646] = 32'h0;  // 32'h0a7c27ec;
    ram_cell[     647] = 32'h0;  // 32'haf8cf2db;
    ram_cell[     648] = 32'h0;  // 32'hcc31a9de;
    ram_cell[     649] = 32'h0;  // 32'h8d1acc9f;
    ram_cell[     650] = 32'h0;  // 32'h60dae9cb;
    ram_cell[     651] = 32'h0;  // 32'h512ea73c;
    ram_cell[     652] = 32'h0;  // 32'h6dc26fa0;
    ram_cell[     653] = 32'h0;  // 32'h82b418d1;
    ram_cell[     654] = 32'h0;  // 32'hf322adea;
    ram_cell[     655] = 32'h0;  // 32'hd73818c5;
    ram_cell[     656] = 32'h0;  // 32'h04dc95ee;
    ram_cell[     657] = 32'h0;  // 32'h60555c83;
    ram_cell[     658] = 32'h0;  // 32'h3caa00aa;
    ram_cell[     659] = 32'h0;  // 32'hb74d2292;
    ram_cell[     660] = 32'h0;  // 32'hf481e249;
    ram_cell[     661] = 32'h0;  // 32'h9df12e6f;
    ram_cell[     662] = 32'h0;  // 32'h2bd2c0ba;
    ram_cell[     663] = 32'h0;  // 32'h0bec0fe9;
    ram_cell[     664] = 32'h0;  // 32'h0cf8534f;
    ram_cell[     665] = 32'h0;  // 32'he5086f08;
    ram_cell[     666] = 32'h0;  // 32'h63cd6876;
    ram_cell[     667] = 32'h0;  // 32'h5461f06b;
    ram_cell[     668] = 32'h0;  // 32'h1784aab9;
    ram_cell[     669] = 32'h0;  // 32'hd28fb0ec;
    ram_cell[     670] = 32'h0;  // 32'h7097aacb;
    ram_cell[     671] = 32'h0;  // 32'h17aedf0d;
    ram_cell[     672] = 32'h0;  // 32'h7914a21f;
    ram_cell[     673] = 32'h0;  // 32'ha47c1b2b;
    ram_cell[     674] = 32'h0;  // 32'h0384282c;
    ram_cell[     675] = 32'h0;  // 32'h7825c10e;
    ram_cell[     676] = 32'h0;  // 32'h016d6d18;
    ram_cell[     677] = 32'h0;  // 32'hf1519dc8;
    ram_cell[     678] = 32'h0;  // 32'hdf879a03;
    ram_cell[     679] = 32'h0;  // 32'hbadd9dba;
    ram_cell[     680] = 32'h0;  // 32'haf3fac06;
    ram_cell[     681] = 32'h0;  // 32'h700408b5;
    ram_cell[     682] = 32'h0;  // 32'h918d2059;
    ram_cell[     683] = 32'h0;  // 32'h8038c7d6;
    ram_cell[     684] = 32'h0;  // 32'hcd80e773;
    ram_cell[     685] = 32'h0;  // 32'h2235a612;
    ram_cell[     686] = 32'h0;  // 32'h5073242d;
    ram_cell[     687] = 32'h0;  // 32'hfd4100ed;
    ram_cell[     688] = 32'h0;  // 32'h9c868c22;
    ram_cell[     689] = 32'h0;  // 32'h24ff74d0;
    ram_cell[     690] = 32'h0;  // 32'ha25269f9;
    ram_cell[     691] = 32'h0;  // 32'hfd7340b2;
    ram_cell[     692] = 32'h0;  // 32'hcd6cb41f;
    ram_cell[     693] = 32'h0;  // 32'hcca8ff65;
    ram_cell[     694] = 32'h0;  // 32'h9f490e62;
    ram_cell[     695] = 32'h0;  // 32'h7634162e;
    ram_cell[     696] = 32'h0;  // 32'h940aec63;
    ram_cell[     697] = 32'h0;  // 32'h1631659a;
    ram_cell[     698] = 32'h0;  // 32'h989bbe19;
    ram_cell[     699] = 32'h0;  // 32'hf420c56e;
    ram_cell[     700] = 32'h0;  // 32'h0623be52;
    ram_cell[     701] = 32'h0;  // 32'h7ac86292;
    ram_cell[     702] = 32'h0;  // 32'h879bdb11;
    ram_cell[     703] = 32'h0;  // 32'hc521fe1f;
    ram_cell[     704] = 32'h0;  // 32'h77d0f688;
    ram_cell[     705] = 32'h0;  // 32'he4101a2d;
    ram_cell[     706] = 32'h0;  // 32'hceda482b;
    ram_cell[     707] = 32'h0;  // 32'hdee5c44f;
    ram_cell[     708] = 32'h0;  // 32'hfdd7abd7;
    ram_cell[     709] = 32'h0;  // 32'h302aa140;
    ram_cell[     710] = 32'h0;  // 32'haaf56088;
    ram_cell[     711] = 32'h0;  // 32'h98c95b99;
    ram_cell[     712] = 32'h0;  // 32'h9f88f25a;
    ram_cell[     713] = 32'h0;  // 32'hb69f2e9d;
    ram_cell[     714] = 32'h0;  // 32'hac8a9052;
    ram_cell[     715] = 32'h0;  // 32'hddf1aed9;
    ram_cell[     716] = 32'h0;  // 32'h4d505023;
    ram_cell[     717] = 32'h0;  // 32'hd1bd3741;
    ram_cell[     718] = 32'h0;  // 32'hb802d361;
    ram_cell[     719] = 32'h0;  // 32'h4646c149;
    ram_cell[     720] = 32'h0;  // 32'hbe699f05;
    ram_cell[     721] = 32'h0;  // 32'h6a3b95dc;
    ram_cell[     722] = 32'h0;  // 32'hb0a775fd;
    ram_cell[     723] = 32'h0;  // 32'h2bdce8ae;
    ram_cell[     724] = 32'h0;  // 32'h2f15cfc5;
    ram_cell[     725] = 32'h0;  // 32'habbef784;
    ram_cell[     726] = 32'h0;  // 32'hc92e35f4;
    ram_cell[     727] = 32'h0;  // 32'h93ed7948;
    ram_cell[     728] = 32'h0;  // 32'he8dda7a6;
    ram_cell[     729] = 32'h0;  // 32'h67350e28;
    ram_cell[     730] = 32'h0;  // 32'h932731fc;
    ram_cell[     731] = 32'h0;  // 32'h0ed08b0a;
    ram_cell[     732] = 32'h0;  // 32'h3c12841b;
    ram_cell[     733] = 32'h0;  // 32'hc9839c4d;
    ram_cell[     734] = 32'h0;  // 32'h7a84ed11;
    ram_cell[     735] = 32'h0;  // 32'hcaa095a2;
    ram_cell[     736] = 32'h0;  // 32'h39b9daba;
    ram_cell[     737] = 32'h0;  // 32'ha652f98d;
    ram_cell[     738] = 32'h0;  // 32'h6ff23987;
    ram_cell[     739] = 32'h0;  // 32'h6be49152;
    ram_cell[     740] = 32'h0;  // 32'h5881fb14;
    ram_cell[     741] = 32'h0;  // 32'h2fc4b19f;
    ram_cell[     742] = 32'h0;  // 32'h2cccc2f8;
    ram_cell[     743] = 32'h0;  // 32'h7e4b78fc;
    ram_cell[     744] = 32'h0;  // 32'hfdf7d024;
    ram_cell[     745] = 32'h0;  // 32'h14b95c7e;
    ram_cell[     746] = 32'h0;  // 32'h04fc4853;
    ram_cell[     747] = 32'h0;  // 32'h6cdd56dd;
    ram_cell[     748] = 32'h0;  // 32'h19b75b62;
    ram_cell[     749] = 32'h0;  // 32'h3f92e5fe;
    ram_cell[     750] = 32'h0;  // 32'h2a91ccc2;
    ram_cell[     751] = 32'h0;  // 32'h52b8dccb;
    ram_cell[     752] = 32'h0;  // 32'h519b4df8;
    ram_cell[     753] = 32'h0;  // 32'he1fdb040;
    ram_cell[     754] = 32'h0;  // 32'hf0bd3ec7;
    ram_cell[     755] = 32'h0;  // 32'h230af1e9;
    ram_cell[     756] = 32'h0;  // 32'h7efcaf37;
    ram_cell[     757] = 32'h0;  // 32'hc745eccf;
    ram_cell[     758] = 32'h0;  // 32'h445ed664;
    ram_cell[     759] = 32'h0;  // 32'h4a28e566;
    ram_cell[     760] = 32'h0;  // 32'hfc68511d;
    ram_cell[     761] = 32'h0;  // 32'h0855b1f7;
    ram_cell[     762] = 32'h0;  // 32'h9547e4cc;
    ram_cell[     763] = 32'h0;  // 32'h7dad1aef;
    ram_cell[     764] = 32'h0;  // 32'h6b34325a;
    ram_cell[     765] = 32'h0;  // 32'h8fd420f1;
    ram_cell[     766] = 32'h0;  // 32'h20d72b9a;
    ram_cell[     767] = 32'h0;  // 32'hbee080bf;
    ram_cell[     768] = 32'h0;  // 32'h8d5bfc44;
    ram_cell[     769] = 32'h0;  // 32'h4b952457;
    ram_cell[     770] = 32'h0;  // 32'h47aceb2a;
    ram_cell[     771] = 32'h0;  // 32'h51884867;
    ram_cell[     772] = 32'h0;  // 32'h576fd8cd;
    ram_cell[     773] = 32'h0;  // 32'h48871ef5;
    ram_cell[     774] = 32'h0;  // 32'ha8fbb4b6;
    ram_cell[     775] = 32'h0;  // 32'hb0c71e51;
    ram_cell[     776] = 32'h0;  // 32'h1db08cfe;
    ram_cell[     777] = 32'h0;  // 32'h5e722926;
    ram_cell[     778] = 32'h0;  // 32'ha7888746;
    ram_cell[     779] = 32'h0;  // 32'h528f196c;
    ram_cell[     780] = 32'h0;  // 32'h675d0c07;
    ram_cell[     781] = 32'h0;  // 32'h89d07fa7;
    ram_cell[     782] = 32'h0;  // 32'h3ac68f63;
    ram_cell[     783] = 32'h0;  // 32'he6472ed1;
    ram_cell[     784] = 32'h0;  // 32'h1188b9f6;
    ram_cell[     785] = 32'h0;  // 32'h6952d7f1;
    ram_cell[     786] = 32'h0;  // 32'h39c621de;
    ram_cell[     787] = 32'h0;  // 32'h3796631e;
    ram_cell[     788] = 32'h0;  // 32'hbe977755;
    ram_cell[     789] = 32'h0;  // 32'hcd01777d;
    ram_cell[     790] = 32'h0;  // 32'h14bbf48a;
    ram_cell[     791] = 32'h0;  // 32'h3963cb24;
    ram_cell[     792] = 32'h0;  // 32'h38be4930;
    ram_cell[     793] = 32'h0;  // 32'hf49016db;
    ram_cell[     794] = 32'h0;  // 32'h891148f2;
    ram_cell[     795] = 32'h0;  // 32'hfe212186;
    ram_cell[     796] = 32'h0;  // 32'h497669e2;
    ram_cell[     797] = 32'h0;  // 32'h26a24561;
    ram_cell[     798] = 32'h0;  // 32'h024680a0;
    ram_cell[     799] = 32'h0;  // 32'h79b5524f;
    ram_cell[     800] = 32'h0;  // 32'h2ca40899;
    ram_cell[     801] = 32'h0;  // 32'h24d9d5d8;
    ram_cell[     802] = 32'h0;  // 32'h840de786;
    ram_cell[     803] = 32'h0;  // 32'hc1f3ec1f;
    ram_cell[     804] = 32'h0;  // 32'h00961800;
    ram_cell[     805] = 32'h0;  // 32'h88dc18cf;
    ram_cell[     806] = 32'h0;  // 32'hdff9d8d5;
    ram_cell[     807] = 32'h0;  // 32'h8b23a69a;
    ram_cell[     808] = 32'h0;  // 32'hd8d540ca;
    ram_cell[     809] = 32'h0;  // 32'h746a3ebd;
    ram_cell[     810] = 32'h0;  // 32'ha392bc66;
    ram_cell[     811] = 32'h0;  // 32'h15823ae0;
    ram_cell[     812] = 32'h0;  // 32'h0a2b095f;
    ram_cell[     813] = 32'h0;  // 32'hdfd7a342;
    ram_cell[     814] = 32'h0;  // 32'ha84bd366;
    ram_cell[     815] = 32'h0;  // 32'h03bfb23f;
    ram_cell[     816] = 32'h0;  // 32'h43cd8ae9;
    ram_cell[     817] = 32'h0;  // 32'hac382c70;
    ram_cell[     818] = 32'h0;  // 32'hd20acd76;
    ram_cell[     819] = 32'h0;  // 32'he5b5a30f;
    ram_cell[     820] = 32'h0;  // 32'h56913f8b;
    ram_cell[     821] = 32'h0;  // 32'hd557dbd1;
    ram_cell[     822] = 32'h0;  // 32'h47dae410;
    ram_cell[     823] = 32'h0;  // 32'h3f36a20d;
    ram_cell[     824] = 32'h0;  // 32'h293f5f09;
    ram_cell[     825] = 32'h0;  // 32'h9fd5bcbf;
    ram_cell[     826] = 32'h0;  // 32'hd7f663eb;
    ram_cell[     827] = 32'h0;  // 32'h48f2c2e9;
    ram_cell[     828] = 32'h0;  // 32'hfa1ff78b;
    ram_cell[     829] = 32'h0;  // 32'hf21b9e77;
    ram_cell[     830] = 32'h0;  // 32'hf22ee630;
    ram_cell[     831] = 32'h0;  // 32'h86279220;
    ram_cell[     832] = 32'h0;  // 32'h16fe37ce;
    ram_cell[     833] = 32'h0;  // 32'h636f775d;
    ram_cell[     834] = 32'h0;  // 32'h457b35fe;
    ram_cell[     835] = 32'h0;  // 32'h942bbdc7;
    ram_cell[     836] = 32'h0;  // 32'h045d6eef;
    ram_cell[     837] = 32'h0;  // 32'hd496fb95;
    ram_cell[     838] = 32'h0;  // 32'hc2052a5a;
    ram_cell[     839] = 32'h0;  // 32'h5df2b992;
    ram_cell[     840] = 32'h0;  // 32'h728ab97f;
    ram_cell[     841] = 32'h0;  // 32'hb0fc9cfb;
    ram_cell[     842] = 32'h0;  // 32'h380399a1;
    ram_cell[     843] = 32'h0;  // 32'h23956cbe;
    ram_cell[     844] = 32'h0;  // 32'h4f45b299;
    ram_cell[     845] = 32'h0;  // 32'h478a4b24;
    ram_cell[     846] = 32'h0;  // 32'h36f78ff9;
    ram_cell[     847] = 32'h0;  // 32'h79a61787;
    ram_cell[     848] = 32'h0;  // 32'hd21e0df5;
    ram_cell[     849] = 32'h0;  // 32'h40e74c52;
    ram_cell[     850] = 32'h0;  // 32'hbebbadd5;
    ram_cell[     851] = 32'h0;  // 32'h55d1d23a;
    ram_cell[     852] = 32'h0;  // 32'h52de5474;
    ram_cell[     853] = 32'h0;  // 32'ha163f297;
    ram_cell[     854] = 32'h0;  // 32'ha6371148;
    ram_cell[     855] = 32'h0;  // 32'hd7c991a9;
    ram_cell[     856] = 32'h0;  // 32'hd4d44b63;
    ram_cell[     857] = 32'h0;  // 32'hf251c255;
    ram_cell[     858] = 32'h0;  // 32'h4c75fc95;
    ram_cell[     859] = 32'h0;  // 32'h1800963d;
    ram_cell[     860] = 32'h0;  // 32'hbc537d2a;
    ram_cell[     861] = 32'h0;  // 32'h9b64f4ec;
    ram_cell[     862] = 32'h0;  // 32'h2c4087f3;
    ram_cell[     863] = 32'h0;  // 32'h0bff682c;
    ram_cell[     864] = 32'h0;  // 32'ha78dd43f;
    ram_cell[     865] = 32'h0;  // 32'h4e148216;
    ram_cell[     866] = 32'h0;  // 32'h26be9bae;
    ram_cell[     867] = 32'h0;  // 32'hfd38e854;
    ram_cell[     868] = 32'h0;  // 32'h66fd7153;
    ram_cell[     869] = 32'h0;  // 32'h97eecd11;
    ram_cell[     870] = 32'h0;  // 32'he5e6dfae;
    ram_cell[     871] = 32'h0;  // 32'h6b4c9a7b;
    ram_cell[     872] = 32'h0;  // 32'hc738e5f8;
    ram_cell[     873] = 32'h0;  // 32'h03628a20;
    ram_cell[     874] = 32'h0;  // 32'hef577610;
    ram_cell[     875] = 32'h0;  // 32'hb8e95924;
    ram_cell[     876] = 32'h0;  // 32'hc340081f;
    ram_cell[     877] = 32'h0;  // 32'hffb54c7f;
    ram_cell[     878] = 32'h0;  // 32'hcd009f76;
    ram_cell[     879] = 32'h0;  // 32'h92f7869d;
    ram_cell[     880] = 32'h0;  // 32'hd4f12493;
    ram_cell[     881] = 32'h0;  // 32'h7e095ecc;
    ram_cell[     882] = 32'h0;  // 32'h75afa250;
    ram_cell[     883] = 32'h0;  // 32'hf11dad6c;
    ram_cell[     884] = 32'h0;  // 32'h77a94b62;
    ram_cell[     885] = 32'h0;  // 32'h198238a2;
    ram_cell[     886] = 32'h0;  // 32'h1beb2a0f;
    ram_cell[     887] = 32'h0;  // 32'h36b96bf0;
    ram_cell[     888] = 32'h0;  // 32'hfcbfe2b2;
    ram_cell[     889] = 32'h0;  // 32'hdece9572;
    ram_cell[     890] = 32'h0;  // 32'h2964b836;
    ram_cell[     891] = 32'h0;  // 32'hbc2c5126;
    ram_cell[     892] = 32'h0;  // 32'hfd0339cb;
    ram_cell[     893] = 32'h0;  // 32'h3b133cba;
    ram_cell[     894] = 32'h0;  // 32'h1a572804;
    ram_cell[     895] = 32'h0;  // 32'h5b3cb3b5;
    ram_cell[     896] = 32'h0;  // 32'heaa5e74f;
    ram_cell[     897] = 32'h0;  // 32'h0f0cfea3;
    ram_cell[     898] = 32'h0;  // 32'hf824b350;
    ram_cell[     899] = 32'h0;  // 32'h544341c7;
    ram_cell[     900] = 32'h0;  // 32'h8602a060;
    ram_cell[     901] = 32'h0;  // 32'h05972016;
    ram_cell[     902] = 32'h0;  // 32'h2f8ade90;
    ram_cell[     903] = 32'h0;  // 32'h5ca48608;
    ram_cell[     904] = 32'h0;  // 32'h6e494e2d;
    ram_cell[     905] = 32'h0;  // 32'hd491af5d;
    ram_cell[     906] = 32'h0;  // 32'he2816b04;
    ram_cell[     907] = 32'h0;  // 32'hf52b6cc7;
    ram_cell[     908] = 32'h0;  // 32'hc4b7b105;
    ram_cell[     909] = 32'h0;  // 32'hb3bd812d;
    ram_cell[     910] = 32'h0;  // 32'haa5a297a;
    ram_cell[     911] = 32'h0;  // 32'h25dd7407;
    ram_cell[     912] = 32'h0;  // 32'h0c659498;
    ram_cell[     913] = 32'h0;  // 32'h5fa662da;
    ram_cell[     914] = 32'h0;  // 32'he19d7746;
    ram_cell[     915] = 32'h0;  // 32'h9eb08b25;
    ram_cell[     916] = 32'h0;  // 32'hdc8cabad;
    ram_cell[     917] = 32'h0;  // 32'ha143ab78;
    ram_cell[     918] = 32'h0;  // 32'h29091894;
    ram_cell[     919] = 32'h0;  // 32'hdf7e80d2;
    ram_cell[     920] = 32'h0;  // 32'hb5ef037e;
    ram_cell[     921] = 32'h0;  // 32'had0d3843;
    ram_cell[     922] = 32'h0;  // 32'h0608aca2;
    ram_cell[     923] = 32'h0;  // 32'h45b602cc;
    ram_cell[     924] = 32'h0;  // 32'h07801431;
    ram_cell[     925] = 32'h0;  // 32'hf57061dc;
    ram_cell[     926] = 32'h0;  // 32'ha4063473;
    ram_cell[     927] = 32'h0;  // 32'hf1351790;
    ram_cell[     928] = 32'h0;  // 32'hb1f08715;
    ram_cell[     929] = 32'h0;  // 32'hc2c022cf;
    ram_cell[     930] = 32'h0;  // 32'h5008d76d;
    ram_cell[     931] = 32'h0;  // 32'h563ce8bc;
    ram_cell[     932] = 32'h0;  // 32'h47e89ede;
    ram_cell[     933] = 32'h0;  // 32'hd9f817d1;
    ram_cell[     934] = 32'h0;  // 32'h392ae8f6;
    ram_cell[     935] = 32'h0;  // 32'h2b7d4775;
    ram_cell[     936] = 32'h0;  // 32'he0de1536;
    ram_cell[     937] = 32'h0;  // 32'h8085b689;
    ram_cell[     938] = 32'h0;  // 32'ha22f093c;
    ram_cell[     939] = 32'h0;  // 32'h635aa697;
    ram_cell[     940] = 32'h0;  // 32'h9966585d;
    ram_cell[     941] = 32'h0;  // 32'hc20ff688;
    ram_cell[     942] = 32'h0;  // 32'hdec25cc7;
    ram_cell[     943] = 32'h0;  // 32'hd8fab380;
    ram_cell[     944] = 32'h0;  // 32'h4a44e575;
    ram_cell[     945] = 32'h0;  // 32'h632951ea;
    ram_cell[     946] = 32'h0;  // 32'h6fdac324;
    ram_cell[     947] = 32'h0;  // 32'h66c9e6b9;
    ram_cell[     948] = 32'h0;  // 32'h2d4cc44f;
    ram_cell[     949] = 32'h0;  // 32'h3dbf5e59;
    ram_cell[     950] = 32'h0;  // 32'h68b57e19;
    ram_cell[     951] = 32'h0;  // 32'hb1fb583b;
    ram_cell[     952] = 32'h0;  // 32'h9208a503;
    ram_cell[     953] = 32'h0;  // 32'h7df8ae3d;
    ram_cell[     954] = 32'h0;  // 32'h4245bae3;
    ram_cell[     955] = 32'h0;  // 32'hf7b00dce;
    ram_cell[     956] = 32'h0;  // 32'h15266d3a;
    ram_cell[     957] = 32'h0;  // 32'he4997d18;
    ram_cell[     958] = 32'h0;  // 32'hd7a6bd88;
    ram_cell[     959] = 32'h0;  // 32'ha1e0c4a1;
    ram_cell[     960] = 32'h0;  // 32'ha273bd5c;
    ram_cell[     961] = 32'h0;  // 32'ha68b5434;
    ram_cell[     962] = 32'h0;  // 32'h22c45b90;
    ram_cell[     963] = 32'h0;  // 32'heeff0144;
    ram_cell[     964] = 32'h0;  // 32'hca999012;
    ram_cell[     965] = 32'h0;  // 32'h79fb4e8c;
    ram_cell[     966] = 32'h0;  // 32'ha52d47cb;
    ram_cell[     967] = 32'h0;  // 32'hf7682970;
    ram_cell[     968] = 32'h0;  // 32'hb4fddc43;
    ram_cell[     969] = 32'h0;  // 32'hca021880;
    ram_cell[     970] = 32'h0;  // 32'h21917fec;
    ram_cell[     971] = 32'h0;  // 32'h275ed211;
    ram_cell[     972] = 32'h0;  // 32'hf7503187;
    ram_cell[     973] = 32'h0;  // 32'hd721bca4;
    ram_cell[     974] = 32'h0;  // 32'h5b63a38f;
    ram_cell[     975] = 32'h0;  // 32'h014d8d3e;
    ram_cell[     976] = 32'h0;  // 32'h03267ec4;
    ram_cell[     977] = 32'h0;  // 32'h6a12e388;
    ram_cell[     978] = 32'h0;  // 32'hf3aad3a1;
    ram_cell[     979] = 32'h0;  // 32'heeee9550;
    ram_cell[     980] = 32'h0;  // 32'hb905b2d8;
    ram_cell[     981] = 32'h0;  // 32'he2a6c883;
    ram_cell[     982] = 32'h0;  // 32'h7be6f282;
    ram_cell[     983] = 32'h0;  // 32'ha67ef9af;
    ram_cell[     984] = 32'h0;  // 32'hbf3b4559;
    ram_cell[     985] = 32'h0;  // 32'h20e38558;
    ram_cell[     986] = 32'h0;  // 32'h058083bb;
    ram_cell[     987] = 32'h0;  // 32'h04104e9d;
    ram_cell[     988] = 32'h0;  // 32'he2ca2d16;
    ram_cell[     989] = 32'h0;  // 32'h65b92ad0;
    ram_cell[     990] = 32'h0;  // 32'h9b26e134;
    ram_cell[     991] = 32'h0;  // 32'h3590f10e;
    ram_cell[     992] = 32'h0;  // 32'hda659e61;
    ram_cell[     993] = 32'h0;  // 32'haa035ad5;
    ram_cell[     994] = 32'h0;  // 32'hd40887ff;
    ram_cell[     995] = 32'h0;  // 32'habaa4569;
    ram_cell[     996] = 32'h0;  // 32'hae44535d;
    ram_cell[     997] = 32'h0;  // 32'hf8d328b1;
    ram_cell[     998] = 32'h0;  // 32'h44ba8314;
    ram_cell[     999] = 32'h0;  // 32'he6a06149;
    ram_cell[    1000] = 32'h0;  // 32'h4402fbc7;
    ram_cell[    1001] = 32'h0;  // 32'hb59deb4a;
    ram_cell[    1002] = 32'h0;  // 32'h6299d18f;
    ram_cell[    1003] = 32'h0;  // 32'h295ff631;
    ram_cell[    1004] = 32'h0;  // 32'h1851c92c;
    ram_cell[    1005] = 32'h0;  // 32'h930ab40f;
    ram_cell[    1006] = 32'h0;  // 32'h3f13755c;
    ram_cell[    1007] = 32'h0;  // 32'h173035a8;
    ram_cell[    1008] = 32'h0;  // 32'hcf22a3fe;
    ram_cell[    1009] = 32'h0;  // 32'h38e2a511;
    ram_cell[    1010] = 32'h0;  // 32'h0c24a6d7;
    ram_cell[    1011] = 32'h0;  // 32'hc96b8d3e;
    ram_cell[    1012] = 32'h0;  // 32'hca4b307d;
    ram_cell[    1013] = 32'h0;  // 32'hb1c603ac;
    ram_cell[    1014] = 32'h0;  // 32'hb8d326e5;
    ram_cell[    1015] = 32'h0;  // 32'hd245c92e;
    ram_cell[    1016] = 32'h0;  // 32'h959f0982;
    ram_cell[    1017] = 32'h0;  // 32'hb3ea7823;
    ram_cell[    1018] = 32'h0;  // 32'hae693fd1;
    ram_cell[    1019] = 32'h0;  // 32'hdaeb58de;
    ram_cell[    1020] = 32'h0;  // 32'h64308c9c;
    ram_cell[    1021] = 32'h0;  // 32'hc0e0362b;
    ram_cell[    1022] = 32'h0;  // 32'hfe436ffe;
    ram_cell[    1023] = 32'h0;  // 32'h61315105;
    // src matrix A
    ram_cell[    1024] = 32'h45dbb061;
    ram_cell[    1025] = 32'h8d8c4ecd;
    ram_cell[    1026] = 32'h35da3b54;
    ram_cell[    1027] = 32'h61a1ae0b;
    ram_cell[    1028] = 32'h3c23f7c5;
    ram_cell[    1029] = 32'h2bb4ab76;
    ram_cell[    1030] = 32'h79383ff7;
    ram_cell[    1031] = 32'hbd35d287;
    ram_cell[    1032] = 32'h02be0ae7;
    ram_cell[    1033] = 32'hb00bf1a4;
    ram_cell[    1034] = 32'h45f1f2fa;
    ram_cell[    1035] = 32'h860c4922;
    ram_cell[    1036] = 32'ha1a6cc5e;
    ram_cell[    1037] = 32'h05c64068;
    ram_cell[    1038] = 32'h8902228b;
    ram_cell[    1039] = 32'h3f654f03;
    ram_cell[    1040] = 32'h399aa357;
    ram_cell[    1041] = 32'h91c99682;
    ram_cell[    1042] = 32'h3e71cb37;
    ram_cell[    1043] = 32'h21ca37f0;
    ram_cell[    1044] = 32'h33a33a98;
    ram_cell[    1045] = 32'h04a0f8f1;
    ram_cell[    1046] = 32'ha48a3958;
    ram_cell[    1047] = 32'hced85758;
    ram_cell[    1048] = 32'he9c20a5b;
    ram_cell[    1049] = 32'hb01ada82;
    ram_cell[    1050] = 32'h2ae93c56;
    ram_cell[    1051] = 32'h16a0183b;
    ram_cell[    1052] = 32'h72cfcf46;
    ram_cell[    1053] = 32'h20066fba;
    ram_cell[    1054] = 32'h3171487e;
    ram_cell[    1055] = 32'he680e70f;
    ram_cell[    1056] = 32'hd28767ee;
    ram_cell[    1057] = 32'h006aa410;
    ram_cell[    1058] = 32'hc20388ee;
    ram_cell[    1059] = 32'h292cb5b5;
    ram_cell[    1060] = 32'h2e1dc238;
    ram_cell[    1061] = 32'h1daf6948;
    ram_cell[    1062] = 32'hd6d3718a;
    ram_cell[    1063] = 32'ha1aa41df;
    ram_cell[    1064] = 32'h69678946;
    ram_cell[    1065] = 32'h6aaa20c5;
    ram_cell[    1066] = 32'hafef316c;
    ram_cell[    1067] = 32'hc044b2ba;
    ram_cell[    1068] = 32'hc34104d4;
    ram_cell[    1069] = 32'hf2becd91;
    ram_cell[    1070] = 32'ha4dfaa7c;
    ram_cell[    1071] = 32'h75513f19;
    ram_cell[    1072] = 32'hd279c7c6;
    ram_cell[    1073] = 32'hd98fb35e;
    ram_cell[    1074] = 32'h3ef99787;
    ram_cell[    1075] = 32'h45dead1f;
    ram_cell[    1076] = 32'h62643a8a;
    ram_cell[    1077] = 32'h139b2a3c;
    ram_cell[    1078] = 32'hcaf3a6a6;
    ram_cell[    1079] = 32'h317ae471;
    ram_cell[    1080] = 32'hcd8b2ea0;
    ram_cell[    1081] = 32'h799be92f;
    ram_cell[    1082] = 32'h763f8b5d;
    ram_cell[    1083] = 32'haf430cbd;
    ram_cell[    1084] = 32'h7a78a73e;
    ram_cell[    1085] = 32'h4d95a40b;
    ram_cell[    1086] = 32'h0c5973bf;
    ram_cell[    1087] = 32'h4a26357b;
    ram_cell[    1088] = 32'h38cd7780;
    ram_cell[    1089] = 32'hcec09caf;
    ram_cell[    1090] = 32'h7f418f69;
    ram_cell[    1091] = 32'he5cddfa0;
    ram_cell[    1092] = 32'hb0efb94d;
    ram_cell[    1093] = 32'h782bb7e8;
    ram_cell[    1094] = 32'h3639dadb;
    ram_cell[    1095] = 32'hc23b0f57;
    ram_cell[    1096] = 32'h597ede8f;
    ram_cell[    1097] = 32'h099885f6;
    ram_cell[    1098] = 32'h30b786bd;
    ram_cell[    1099] = 32'hd401e588;
    ram_cell[    1100] = 32'h55694827;
    ram_cell[    1101] = 32'hdc522b5d;
    ram_cell[    1102] = 32'h03550e4f;
    ram_cell[    1103] = 32'hd65eb27d;
    ram_cell[    1104] = 32'h9088a851;
    ram_cell[    1105] = 32'h308acfe4;
    ram_cell[    1106] = 32'h46bb665e;
    ram_cell[    1107] = 32'h39c6663a;
    ram_cell[    1108] = 32'h34b23d65;
    ram_cell[    1109] = 32'h4422eb9a;
    ram_cell[    1110] = 32'hae768724;
    ram_cell[    1111] = 32'hd19ba169;
    ram_cell[    1112] = 32'h9bb0c223;
    ram_cell[    1113] = 32'h6a2b52c5;
    ram_cell[    1114] = 32'h929ad86f;
    ram_cell[    1115] = 32'hd4ae05fa;
    ram_cell[    1116] = 32'hdcd665c7;
    ram_cell[    1117] = 32'hcd25da4a;
    ram_cell[    1118] = 32'h1f0e4022;
    ram_cell[    1119] = 32'hf5f0c8f2;
    ram_cell[    1120] = 32'h2c87f685;
    ram_cell[    1121] = 32'hff5ee25a;
    ram_cell[    1122] = 32'hc8f6beed;
    ram_cell[    1123] = 32'h32154e08;
    ram_cell[    1124] = 32'h44980aab;
    ram_cell[    1125] = 32'h05c39779;
    ram_cell[    1126] = 32'h1d4c706e;
    ram_cell[    1127] = 32'h5bb69cce;
    ram_cell[    1128] = 32'h98e40607;
    ram_cell[    1129] = 32'h674fc79a;
    ram_cell[    1130] = 32'h672c2489;
    ram_cell[    1131] = 32'h19f3fde0;
    ram_cell[    1132] = 32'hd11a614d;
    ram_cell[    1133] = 32'h90527a0a;
    ram_cell[    1134] = 32'h392ec918;
    ram_cell[    1135] = 32'h5e229107;
    ram_cell[    1136] = 32'hea973ade;
    ram_cell[    1137] = 32'hd15a1192;
    ram_cell[    1138] = 32'h45807e0a;
    ram_cell[    1139] = 32'h3b4fbcaf;
    ram_cell[    1140] = 32'hce35e0dc;
    ram_cell[    1141] = 32'hd8d414a3;
    ram_cell[    1142] = 32'hbb19bf5f;
    ram_cell[    1143] = 32'hf78574ef;
    ram_cell[    1144] = 32'h448ea46f;
    ram_cell[    1145] = 32'h11220f75;
    ram_cell[    1146] = 32'hc87c9113;
    ram_cell[    1147] = 32'h9b8a9dfa;
    ram_cell[    1148] = 32'hf3d524c2;
    ram_cell[    1149] = 32'hbda002d0;
    ram_cell[    1150] = 32'h1adb8b34;
    ram_cell[    1151] = 32'h8e37dd9d;
    ram_cell[    1152] = 32'h54713206;
    ram_cell[    1153] = 32'ha58a5e35;
    ram_cell[    1154] = 32'h386d6e9c;
    ram_cell[    1155] = 32'h998d0b1a;
    ram_cell[    1156] = 32'h297b326d;
    ram_cell[    1157] = 32'h5f129318;
    ram_cell[    1158] = 32'hbb3248e0;
    ram_cell[    1159] = 32'h2bbb0466;
    ram_cell[    1160] = 32'h4cfda1b1;
    ram_cell[    1161] = 32'h4a18a06d;
    ram_cell[    1162] = 32'h66804fcd;
    ram_cell[    1163] = 32'h49ed166e;
    ram_cell[    1164] = 32'h1e708e68;
    ram_cell[    1165] = 32'ha95c9886;
    ram_cell[    1166] = 32'h4f21f863;
    ram_cell[    1167] = 32'h20b5ba94;
    ram_cell[    1168] = 32'h95a677ef;
    ram_cell[    1169] = 32'h70438798;
    ram_cell[    1170] = 32'h7551e0d9;
    ram_cell[    1171] = 32'hafc56591;
    ram_cell[    1172] = 32'h068d0477;
    ram_cell[    1173] = 32'h885907f0;
    ram_cell[    1174] = 32'h9c0e86cd;
    ram_cell[    1175] = 32'hc8530ce0;
    ram_cell[    1176] = 32'h61c5d035;
    ram_cell[    1177] = 32'h9589a6c2;
    ram_cell[    1178] = 32'h7a4e325b;
    ram_cell[    1179] = 32'hc06ec99f;
    ram_cell[    1180] = 32'hb3ea074d;
    ram_cell[    1181] = 32'hd9400ffc;
    ram_cell[    1182] = 32'h34ec28f9;
    ram_cell[    1183] = 32'hda03928f;
    ram_cell[    1184] = 32'he4eb37ce;
    ram_cell[    1185] = 32'he38abf0c;
    ram_cell[    1186] = 32'h80801508;
    ram_cell[    1187] = 32'h6819644f;
    ram_cell[    1188] = 32'h1bc55a90;
    ram_cell[    1189] = 32'h4fd3d731;
    ram_cell[    1190] = 32'hbc066a8a;
    ram_cell[    1191] = 32'h272a262e;
    ram_cell[    1192] = 32'h920d5acc;
    ram_cell[    1193] = 32'hd328fc08;
    ram_cell[    1194] = 32'hf66dd972;
    ram_cell[    1195] = 32'h4c3c9a22;
    ram_cell[    1196] = 32'h3dae427d;
    ram_cell[    1197] = 32'h8c20c8a0;
    ram_cell[    1198] = 32'h1af70ff0;
    ram_cell[    1199] = 32'h2ed30d26;
    ram_cell[    1200] = 32'ha8c3351c;
    ram_cell[    1201] = 32'h2aa19e19;
    ram_cell[    1202] = 32'hf93e9260;
    ram_cell[    1203] = 32'hfb93cc24;
    ram_cell[    1204] = 32'h48e114ea;
    ram_cell[    1205] = 32'ha5b91b50;
    ram_cell[    1206] = 32'h96fb0206;
    ram_cell[    1207] = 32'hfa385cbe;
    ram_cell[    1208] = 32'h3d28bd22;
    ram_cell[    1209] = 32'hdd3b1bae;
    ram_cell[    1210] = 32'hc598ba91;
    ram_cell[    1211] = 32'h74926c18;
    ram_cell[    1212] = 32'hb04efa82;
    ram_cell[    1213] = 32'h411e8dcc;
    ram_cell[    1214] = 32'hadf1a616;
    ram_cell[    1215] = 32'h716f007e;
    ram_cell[    1216] = 32'h5ddc39b4;
    ram_cell[    1217] = 32'h8bbdb02a;
    ram_cell[    1218] = 32'h81f82da2;
    ram_cell[    1219] = 32'hfb179eda;
    ram_cell[    1220] = 32'h8b52c7f4;
    ram_cell[    1221] = 32'h4f356ed2;
    ram_cell[    1222] = 32'h6a32beea;
    ram_cell[    1223] = 32'h4d4c0f4e;
    ram_cell[    1224] = 32'h30aa0e6d;
    ram_cell[    1225] = 32'h390ead73;
    ram_cell[    1226] = 32'h9854414b;
    ram_cell[    1227] = 32'h291ab948;
    ram_cell[    1228] = 32'haa0e66d6;
    ram_cell[    1229] = 32'h9598ef42;
    ram_cell[    1230] = 32'h2ba199b7;
    ram_cell[    1231] = 32'hd45c8404;
    ram_cell[    1232] = 32'h29d07fbd;
    ram_cell[    1233] = 32'hdd1473b1;
    ram_cell[    1234] = 32'h2122cb81;
    ram_cell[    1235] = 32'hc34c8aeb;
    ram_cell[    1236] = 32'hbe807def;
    ram_cell[    1237] = 32'h8a910d76;
    ram_cell[    1238] = 32'hebcf0270;
    ram_cell[    1239] = 32'hdf512015;
    ram_cell[    1240] = 32'h36bf8e04;
    ram_cell[    1241] = 32'h5005cd77;
    ram_cell[    1242] = 32'h7661b6fb;
    ram_cell[    1243] = 32'he72ee719;
    ram_cell[    1244] = 32'h713a913e;
    ram_cell[    1245] = 32'hed81df69;
    ram_cell[    1246] = 32'he9deec0f;
    ram_cell[    1247] = 32'haa9eb7c2;
    ram_cell[    1248] = 32'h1ba3e4d6;
    ram_cell[    1249] = 32'h33913abd;
    ram_cell[    1250] = 32'h73b3ea12;
    ram_cell[    1251] = 32'h5348ffc4;
    ram_cell[    1252] = 32'hbaf38a6e;
    ram_cell[    1253] = 32'h1cd4b1d0;
    ram_cell[    1254] = 32'h06c09e1a;
    ram_cell[    1255] = 32'hfad07458;
    ram_cell[    1256] = 32'hcdd87c97;
    ram_cell[    1257] = 32'ha51f51aa;
    ram_cell[    1258] = 32'ha9589a99;
    ram_cell[    1259] = 32'hb783e34a;
    ram_cell[    1260] = 32'h7af40103;
    ram_cell[    1261] = 32'h8daea9ef;
    ram_cell[    1262] = 32'hefb02d64;
    ram_cell[    1263] = 32'ha139ecb9;
    ram_cell[    1264] = 32'h58018bba;
    ram_cell[    1265] = 32'hf1745141;
    ram_cell[    1266] = 32'h7885717a;
    ram_cell[    1267] = 32'h5e7b2ded;
    ram_cell[    1268] = 32'h4afa2c72;
    ram_cell[    1269] = 32'h144b3efd;
    ram_cell[    1270] = 32'hb2a58bf3;
    ram_cell[    1271] = 32'h47542f46;
    ram_cell[    1272] = 32'he5bcdb88;
    ram_cell[    1273] = 32'h7e86cf25;
    ram_cell[    1274] = 32'h49f0e085;
    ram_cell[    1275] = 32'h802d5da9;
    ram_cell[    1276] = 32'hcb0a7027;
    ram_cell[    1277] = 32'hcbd7b5e9;
    ram_cell[    1278] = 32'h6c8129f4;
    ram_cell[    1279] = 32'he5cffe9c;
    ram_cell[    1280] = 32'h7db7d6a8;
    ram_cell[    1281] = 32'h89727616;
    ram_cell[    1282] = 32'h5a431c52;
    ram_cell[    1283] = 32'he4330730;
    ram_cell[    1284] = 32'h8d096771;
    ram_cell[    1285] = 32'h84e167a5;
    ram_cell[    1286] = 32'hd76e0981;
    ram_cell[    1287] = 32'h2d86c9af;
    ram_cell[    1288] = 32'h6fd7d30d;
    ram_cell[    1289] = 32'h586892aa;
    ram_cell[    1290] = 32'h001e3fe9;
    ram_cell[    1291] = 32'h103d5b83;
    ram_cell[    1292] = 32'h0d2eb89b;
    ram_cell[    1293] = 32'hb851be8f;
    ram_cell[    1294] = 32'hb1587105;
    ram_cell[    1295] = 32'h9aef93a3;
    ram_cell[    1296] = 32'h0ae5a4a6;
    ram_cell[    1297] = 32'h04fcc63c;
    ram_cell[    1298] = 32'hd5328871;
    ram_cell[    1299] = 32'h5ecf8e74;
    ram_cell[    1300] = 32'h819fcb32;
    ram_cell[    1301] = 32'hdaf81396;
    ram_cell[    1302] = 32'h5678ed98;
    ram_cell[    1303] = 32'hc237088c;
    ram_cell[    1304] = 32'h31eb5b7c;
    ram_cell[    1305] = 32'h7d4b0cba;
    ram_cell[    1306] = 32'hda3d0727;
    ram_cell[    1307] = 32'hb5fed57d;
    ram_cell[    1308] = 32'h5e9ee458;
    ram_cell[    1309] = 32'hea19f4fc;
    ram_cell[    1310] = 32'h24ceb3ff;
    ram_cell[    1311] = 32'h57df473e;
    ram_cell[    1312] = 32'h08aa0420;
    ram_cell[    1313] = 32'h7da079ef;
    ram_cell[    1314] = 32'h54fbb0a4;
    ram_cell[    1315] = 32'ha4e0446f;
    ram_cell[    1316] = 32'h62176cc5;
    ram_cell[    1317] = 32'h2a559fd8;
    ram_cell[    1318] = 32'h9d8700af;
    ram_cell[    1319] = 32'h9d73fa58;
    ram_cell[    1320] = 32'h42745cd8;
    ram_cell[    1321] = 32'ha8fe7a0c;
    ram_cell[    1322] = 32'hb45c097c;
    ram_cell[    1323] = 32'h55fe1ec1;
    ram_cell[    1324] = 32'h90b7cc57;
    ram_cell[    1325] = 32'hce64b355;
    ram_cell[    1326] = 32'he4c011dc;
    ram_cell[    1327] = 32'h6728a3e0;
    ram_cell[    1328] = 32'h087409e2;
    ram_cell[    1329] = 32'h331c5d7a;
    ram_cell[    1330] = 32'h759152d5;
    ram_cell[    1331] = 32'h57751fbd;
    ram_cell[    1332] = 32'ha272ad01;
    ram_cell[    1333] = 32'hb325d38f;
    ram_cell[    1334] = 32'hc34e1d4f;
    ram_cell[    1335] = 32'hb7af786b;
    ram_cell[    1336] = 32'h963bf337;
    ram_cell[    1337] = 32'hd2f021e1;
    ram_cell[    1338] = 32'he366823c;
    ram_cell[    1339] = 32'ha188e39b;
    ram_cell[    1340] = 32'hd896759b;
    ram_cell[    1341] = 32'h86841acf;
    ram_cell[    1342] = 32'h7cba5233;
    ram_cell[    1343] = 32'h17e38fa9;
    ram_cell[    1344] = 32'hc7c6c70f;
    ram_cell[    1345] = 32'h802136d0;
    ram_cell[    1346] = 32'h4a230335;
    ram_cell[    1347] = 32'hf23e79ae;
    ram_cell[    1348] = 32'h5ac21b5a;
    ram_cell[    1349] = 32'h22f2dae7;
    ram_cell[    1350] = 32'h47463075;
    ram_cell[    1351] = 32'h5c38f18e;
    ram_cell[    1352] = 32'h35bd3145;
    ram_cell[    1353] = 32'h62f2face;
    ram_cell[    1354] = 32'hff9147e9;
    ram_cell[    1355] = 32'h1be0727a;
    ram_cell[    1356] = 32'h6721074b;
    ram_cell[    1357] = 32'h2ecfa4d0;
    ram_cell[    1358] = 32'hcc4b04c8;
    ram_cell[    1359] = 32'h69fb50ab;
    ram_cell[    1360] = 32'h85d9b55a;
    ram_cell[    1361] = 32'hf47ffaa2;
    ram_cell[    1362] = 32'ha01826ab;
    ram_cell[    1363] = 32'hef6824ea;
    ram_cell[    1364] = 32'h8fa7cfba;
    ram_cell[    1365] = 32'h3fab151f;
    ram_cell[    1366] = 32'h54cf1417;
    ram_cell[    1367] = 32'ha5de9ac2;
    ram_cell[    1368] = 32'hbae65114;
    ram_cell[    1369] = 32'h896d4f5c;
    ram_cell[    1370] = 32'h0b4af590;
    ram_cell[    1371] = 32'h3c431fd6;
    ram_cell[    1372] = 32'hf45e0ea8;
    ram_cell[    1373] = 32'h73d05fe3;
    ram_cell[    1374] = 32'ha50f9242;
    ram_cell[    1375] = 32'he52b73e4;
    ram_cell[    1376] = 32'hf9411fd2;
    ram_cell[    1377] = 32'hb7f9eab8;
    ram_cell[    1378] = 32'h8141557a;
    ram_cell[    1379] = 32'h4d819168;
    ram_cell[    1380] = 32'hc996ab9f;
    ram_cell[    1381] = 32'h2e350507;
    ram_cell[    1382] = 32'h30f6c5df;
    ram_cell[    1383] = 32'h884201c8;
    ram_cell[    1384] = 32'h46aecd90;
    ram_cell[    1385] = 32'h815856ed;
    ram_cell[    1386] = 32'ha6e4205b;
    ram_cell[    1387] = 32'hec0a6dbc;
    ram_cell[    1388] = 32'ha0f8bb5b;
    ram_cell[    1389] = 32'hd6d74cdc;
    ram_cell[    1390] = 32'he80a8935;
    ram_cell[    1391] = 32'h9003b81f;
    ram_cell[    1392] = 32'h2cac604f;
    ram_cell[    1393] = 32'h8732798b;
    ram_cell[    1394] = 32'h08546106;
    ram_cell[    1395] = 32'h9380995d;
    ram_cell[    1396] = 32'h616b8843;
    ram_cell[    1397] = 32'hc4634fd0;
    ram_cell[    1398] = 32'h1420f514;
    ram_cell[    1399] = 32'h355b6afe;
    ram_cell[    1400] = 32'h19df768e;
    ram_cell[    1401] = 32'h7f2cf91b;
    ram_cell[    1402] = 32'hf7cb5a5d;
    ram_cell[    1403] = 32'h05146f7b;
    ram_cell[    1404] = 32'heca5be29;
    ram_cell[    1405] = 32'h8af6a094;
    ram_cell[    1406] = 32'h626f2b1d;
    ram_cell[    1407] = 32'h471e64de;
    ram_cell[    1408] = 32'h21346d75;
    ram_cell[    1409] = 32'hf7d0778b;
    ram_cell[    1410] = 32'h0b1e1fc9;
    ram_cell[    1411] = 32'h9eacd5e5;
    ram_cell[    1412] = 32'ha779a557;
    ram_cell[    1413] = 32'hc977cd17;
    ram_cell[    1414] = 32'he2bd4ebf;
    ram_cell[    1415] = 32'h1742ceaf;
    ram_cell[    1416] = 32'hfee82de5;
    ram_cell[    1417] = 32'h80c4f2d3;
    ram_cell[    1418] = 32'hb5f26c6b;
    ram_cell[    1419] = 32'h2369076b;
    ram_cell[    1420] = 32'hdd74fea5;
    ram_cell[    1421] = 32'h180b66a4;
    ram_cell[    1422] = 32'h8e61532d;
    ram_cell[    1423] = 32'h515f3eeb;
    ram_cell[    1424] = 32'h1c1355f6;
    ram_cell[    1425] = 32'h972fbec1;
    ram_cell[    1426] = 32'h81ada239;
    ram_cell[    1427] = 32'hbae7e8fd;
    ram_cell[    1428] = 32'h31025c5e;
    ram_cell[    1429] = 32'h85d091a0;
    ram_cell[    1430] = 32'h87fd03c3;
    ram_cell[    1431] = 32'h6299d39e;
    ram_cell[    1432] = 32'hdf5fbe59;
    ram_cell[    1433] = 32'hedce7cab;
    ram_cell[    1434] = 32'h874d79ab;
    ram_cell[    1435] = 32'h0320c0c8;
    ram_cell[    1436] = 32'h0e8bbab6;
    ram_cell[    1437] = 32'ha8ac1ab5;
    ram_cell[    1438] = 32'hb5f0f89f;
    ram_cell[    1439] = 32'h5951c891;
    ram_cell[    1440] = 32'hf7ad6bca;
    ram_cell[    1441] = 32'hfe66bf17;
    ram_cell[    1442] = 32'hce6e79dc;
    ram_cell[    1443] = 32'hb1cf20ea;
    ram_cell[    1444] = 32'hdb566391;
    ram_cell[    1445] = 32'h76b1d711;
    ram_cell[    1446] = 32'h6cdf5993;
    ram_cell[    1447] = 32'had321f24;
    ram_cell[    1448] = 32'hc17fce0d;
    ram_cell[    1449] = 32'h03cd6467;
    ram_cell[    1450] = 32'h887737f2;
    ram_cell[    1451] = 32'hc73f6c11;
    ram_cell[    1452] = 32'h72c8f0bb;
    ram_cell[    1453] = 32'h82120dac;
    ram_cell[    1454] = 32'hd0cc986a;
    ram_cell[    1455] = 32'h45381e7b;
    ram_cell[    1456] = 32'h28e1b388;
    ram_cell[    1457] = 32'h7e2e701d;
    ram_cell[    1458] = 32'h4ec0ec0e;
    ram_cell[    1459] = 32'hdfcc60bb;
    ram_cell[    1460] = 32'h83ff08c7;
    ram_cell[    1461] = 32'h35c8d464;
    ram_cell[    1462] = 32'h32602620;
    ram_cell[    1463] = 32'h5e9fa210;
    ram_cell[    1464] = 32'hbd884b3b;
    ram_cell[    1465] = 32'h05125d34;
    ram_cell[    1466] = 32'h8b0ed87e;
    ram_cell[    1467] = 32'he2fa3ee0;
    ram_cell[    1468] = 32'h46e2a457;
    ram_cell[    1469] = 32'hbfe1479e;
    ram_cell[    1470] = 32'h2d734493;
    ram_cell[    1471] = 32'h147aa2f8;
    ram_cell[    1472] = 32'he445e6ea;
    ram_cell[    1473] = 32'hf8b1cbe4;
    ram_cell[    1474] = 32'hc30924d6;
    ram_cell[    1475] = 32'haf906281;
    ram_cell[    1476] = 32'hed4b23f8;
    ram_cell[    1477] = 32'he527be66;
    ram_cell[    1478] = 32'h0f015da3;
    ram_cell[    1479] = 32'heec2197d;
    ram_cell[    1480] = 32'hc68fb55e;
    ram_cell[    1481] = 32'h315476f2;
    ram_cell[    1482] = 32'h6272d600;
    ram_cell[    1483] = 32'h5737b8a2;
    ram_cell[    1484] = 32'hcd640a45;
    ram_cell[    1485] = 32'h3c23c4ea;
    ram_cell[    1486] = 32'h27fca22d;
    ram_cell[    1487] = 32'hd42b0343;
    ram_cell[    1488] = 32'hb1b5cb74;
    ram_cell[    1489] = 32'h9fb9a569;
    ram_cell[    1490] = 32'hd30f77dd;
    ram_cell[    1491] = 32'h71f6aba4;
    ram_cell[    1492] = 32'h0ddfa752;
    ram_cell[    1493] = 32'h7b90df8b;
    ram_cell[    1494] = 32'hc1adfcb1;
    ram_cell[    1495] = 32'hb135c789;
    ram_cell[    1496] = 32'h77f1484f;
    ram_cell[    1497] = 32'h4ed9b5f6;
    ram_cell[    1498] = 32'h084949cf;
    ram_cell[    1499] = 32'hf97e3db9;
    ram_cell[    1500] = 32'h7aff7795;
    ram_cell[    1501] = 32'h358d368e;
    ram_cell[    1502] = 32'hf5a8a451;
    ram_cell[    1503] = 32'h3b1dcea6;
    ram_cell[    1504] = 32'hb09eeff5;
    ram_cell[    1505] = 32'hfc44771d;
    ram_cell[    1506] = 32'h5251869b;
    ram_cell[    1507] = 32'ha0f90d7b;
    ram_cell[    1508] = 32'h3e7bf593;
    ram_cell[    1509] = 32'hf4d896bb;
    ram_cell[    1510] = 32'hbd437f9f;
    ram_cell[    1511] = 32'head9537a;
    ram_cell[    1512] = 32'h232d3d7e;
    ram_cell[    1513] = 32'h6ac1299c;
    ram_cell[    1514] = 32'h8dc8309f;
    ram_cell[    1515] = 32'h40df2a39;
    ram_cell[    1516] = 32'h3cf2c319;
    ram_cell[    1517] = 32'hf875ee91;
    ram_cell[    1518] = 32'h116d70e4;
    ram_cell[    1519] = 32'hd77840b8;
    ram_cell[    1520] = 32'h59067d1c;
    ram_cell[    1521] = 32'h1bba4d7c;
    ram_cell[    1522] = 32'hd2b99cc3;
    ram_cell[    1523] = 32'hb2985250;
    ram_cell[    1524] = 32'hacb66513;
    ram_cell[    1525] = 32'h4156bfee;
    ram_cell[    1526] = 32'hbf8270a4;
    ram_cell[    1527] = 32'h16fbc117;
    ram_cell[    1528] = 32'hf51100ac;
    ram_cell[    1529] = 32'h0d73c362;
    ram_cell[    1530] = 32'hffe13e30;
    ram_cell[    1531] = 32'h1ae5bd19;
    ram_cell[    1532] = 32'h429206d1;
    ram_cell[    1533] = 32'ha62d3d7c;
    ram_cell[    1534] = 32'h37906c51;
    ram_cell[    1535] = 32'hb49e6392;
    ram_cell[    1536] = 32'heb2007b0;
    ram_cell[    1537] = 32'hefa66680;
    ram_cell[    1538] = 32'h2d05b6e4;
    ram_cell[    1539] = 32'ha7e55672;
    ram_cell[    1540] = 32'h28b414f0;
    ram_cell[    1541] = 32'hed2a97b3;
    ram_cell[    1542] = 32'h324b3ab2;
    ram_cell[    1543] = 32'h70537fec;
    ram_cell[    1544] = 32'h7e400a85;
    ram_cell[    1545] = 32'h29a5b397;
    ram_cell[    1546] = 32'h0292dda0;
    ram_cell[    1547] = 32'h3ad55b5b;
    ram_cell[    1548] = 32'h2a9d3833;
    ram_cell[    1549] = 32'ha857a9d5;
    ram_cell[    1550] = 32'h40034a15;
    ram_cell[    1551] = 32'h575bca51;
    ram_cell[    1552] = 32'h0c8cfbd2;
    ram_cell[    1553] = 32'hd4a00971;
    ram_cell[    1554] = 32'hba84b588;
    ram_cell[    1555] = 32'ha0b33915;
    ram_cell[    1556] = 32'hbe0ca09d;
    ram_cell[    1557] = 32'h51c89b25;
    ram_cell[    1558] = 32'hbdb83a1c;
    ram_cell[    1559] = 32'hf6a7964c;
    ram_cell[    1560] = 32'h4f58fd56;
    ram_cell[    1561] = 32'h57c47d60;
    ram_cell[    1562] = 32'h7e258a72;
    ram_cell[    1563] = 32'hcaf73a9e;
    ram_cell[    1564] = 32'hac3deb30;
    ram_cell[    1565] = 32'h27d5c70a;
    ram_cell[    1566] = 32'hc55ba477;
    ram_cell[    1567] = 32'hf5ed2f8b;
    ram_cell[    1568] = 32'h83a42160;
    ram_cell[    1569] = 32'h9d3045be;
    ram_cell[    1570] = 32'hf6f6f41f;
    ram_cell[    1571] = 32'hf0916341;
    ram_cell[    1572] = 32'hf146aa1b;
    ram_cell[    1573] = 32'hd22c43d4;
    ram_cell[    1574] = 32'h51538fd8;
    ram_cell[    1575] = 32'hc354c44f;
    ram_cell[    1576] = 32'h86e087fc;
    ram_cell[    1577] = 32'hf7677a6d;
    ram_cell[    1578] = 32'h6afb8138;
    ram_cell[    1579] = 32'hba57ef6c;
    ram_cell[    1580] = 32'h595c1818;
    ram_cell[    1581] = 32'h171d32b3;
    ram_cell[    1582] = 32'hae9e8bac;
    ram_cell[    1583] = 32'ha03c0396;
    ram_cell[    1584] = 32'h4892e017;
    ram_cell[    1585] = 32'h98e17f1b;
    ram_cell[    1586] = 32'h303167dc;
    ram_cell[    1587] = 32'hc83ea84b;
    ram_cell[    1588] = 32'h988ae72b;
    ram_cell[    1589] = 32'h223a054c;
    ram_cell[    1590] = 32'h35ee835b;
    ram_cell[    1591] = 32'he670d384;
    ram_cell[    1592] = 32'h9e0483d0;
    ram_cell[    1593] = 32'hbb03d0a6;
    ram_cell[    1594] = 32'hd1d3e148;
    ram_cell[    1595] = 32'h2c127e1c;
    ram_cell[    1596] = 32'h52e069be;
    ram_cell[    1597] = 32'h0fe3d011;
    ram_cell[    1598] = 32'h32ddd366;
    ram_cell[    1599] = 32'hbc5a040d;
    ram_cell[    1600] = 32'hda5a3d30;
    ram_cell[    1601] = 32'hf958e174;
    ram_cell[    1602] = 32'ha80c4cea;
    ram_cell[    1603] = 32'hf39040e3;
    ram_cell[    1604] = 32'h5a0031f7;
    ram_cell[    1605] = 32'h5e56454b;
    ram_cell[    1606] = 32'h5dccb001;
    ram_cell[    1607] = 32'hd698fec6;
    ram_cell[    1608] = 32'h640d5f99;
    ram_cell[    1609] = 32'hec3f98ad;
    ram_cell[    1610] = 32'he1ecf270;
    ram_cell[    1611] = 32'hb007b788;
    ram_cell[    1612] = 32'hc624ea71;
    ram_cell[    1613] = 32'h0cd7d805;
    ram_cell[    1614] = 32'hc9b9c153;
    ram_cell[    1615] = 32'h20d2cf79;
    ram_cell[    1616] = 32'h86c12269;
    ram_cell[    1617] = 32'hbd721713;
    ram_cell[    1618] = 32'ha25a83b4;
    ram_cell[    1619] = 32'hc67e3545;
    ram_cell[    1620] = 32'h27076fe3;
    ram_cell[    1621] = 32'h089aca67;
    ram_cell[    1622] = 32'hf8605b3b;
    ram_cell[    1623] = 32'h699181e4;
    ram_cell[    1624] = 32'h61d4f86c;
    ram_cell[    1625] = 32'h209232f4;
    ram_cell[    1626] = 32'hfed95dd6;
    ram_cell[    1627] = 32'hba3502c7;
    ram_cell[    1628] = 32'h0429cb98;
    ram_cell[    1629] = 32'hc3fd8078;
    ram_cell[    1630] = 32'h6e4d1b9a;
    ram_cell[    1631] = 32'h0b114e05;
    ram_cell[    1632] = 32'h5f03d508;
    ram_cell[    1633] = 32'h5693dde3;
    ram_cell[    1634] = 32'h7b9585c5;
    ram_cell[    1635] = 32'h4d84c375;
    ram_cell[    1636] = 32'h9dd38377;
    ram_cell[    1637] = 32'h274a3d04;
    ram_cell[    1638] = 32'hdd61d114;
    ram_cell[    1639] = 32'h48c10102;
    ram_cell[    1640] = 32'hf35f9ff0;
    ram_cell[    1641] = 32'hd182963a;
    ram_cell[    1642] = 32'h57a03abf;
    ram_cell[    1643] = 32'h0f280204;
    ram_cell[    1644] = 32'he411c731;
    ram_cell[    1645] = 32'hb65c8858;
    ram_cell[    1646] = 32'h5ab4458f;
    ram_cell[    1647] = 32'h273cb010;
    ram_cell[    1648] = 32'h5202e534;
    ram_cell[    1649] = 32'h09404015;
    ram_cell[    1650] = 32'h8b1241ff;
    ram_cell[    1651] = 32'h85fb4f42;
    ram_cell[    1652] = 32'h47ae93e6;
    ram_cell[    1653] = 32'ha0c59854;
    ram_cell[    1654] = 32'h3970ffac;
    ram_cell[    1655] = 32'h2350262d;
    ram_cell[    1656] = 32'h24c235cf;
    ram_cell[    1657] = 32'h4d920f2c;
    ram_cell[    1658] = 32'h4e673bb2;
    ram_cell[    1659] = 32'h686d0625;
    ram_cell[    1660] = 32'h6803612d;
    ram_cell[    1661] = 32'h7be1bf0b;
    ram_cell[    1662] = 32'hfe9891a1;
    ram_cell[    1663] = 32'h653cc649;
    ram_cell[    1664] = 32'h2411e314;
    ram_cell[    1665] = 32'h79217ba3;
    ram_cell[    1666] = 32'hc5443af9;
    ram_cell[    1667] = 32'hb02ba9e2;
    ram_cell[    1668] = 32'h26c81b15;
    ram_cell[    1669] = 32'hbdc54282;
    ram_cell[    1670] = 32'h2e286980;
    ram_cell[    1671] = 32'h9e222f96;
    ram_cell[    1672] = 32'h304d5913;
    ram_cell[    1673] = 32'h7bc8c0dd;
    ram_cell[    1674] = 32'h182c674e;
    ram_cell[    1675] = 32'hfb42a513;
    ram_cell[    1676] = 32'h6752a7c8;
    ram_cell[    1677] = 32'h157fcf62;
    ram_cell[    1678] = 32'h933fa826;
    ram_cell[    1679] = 32'h5f38b782;
    ram_cell[    1680] = 32'hde92b402;
    ram_cell[    1681] = 32'h9f2f9f30;
    ram_cell[    1682] = 32'h4a7a2424;
    ram_cell[    1683] = 32'h2777a40e;
    ram_cell[    1684] = 32'h8fd3ebdb;
    ram_cell[    1685] = 32'h1eac84e7;
    ram_cell[    1686] = 32'hcbd65658;
    ram_cell[    1687] = 32'h338ab387;
    ram_cell[    1688] = 32'hdee3a052;
    ram_cell[    1689] = 32'h13c0dbe9;
    ram_cell[    1690] = 32'hc28b4e51;
    ram_cell[    1691] = 32'haf53edb6;
    ram_cell[    1692] = 32'h7ffaa07d;
    ram_cell[    1693] = 32'h62b0112a;
    ram_cell[    1694] = 32'h48a6232d;
    ram_cell[    1695] = 32'h9710871e;
    ram_cell[    1696] = 32'h4a5fd64b;
    ram_cell[    1697] = 32'hf1038f35;
    ram_cell[    1698] = 32'h87ff1ae7;
    ram_cell[    1699] = 32'h5f0ce737;
    ram_cell[    1700] = 32'h61d4cdc0;
    ram_cell[    1701] = 32'he50269f5;
    ram_cell[    1702] = 32'h6f67e4e4;
    ram_cell[    1703] = 32'h92e02653;
    ram_cell[    1704] = 32'h08456e31;
    ram_cell[    1705] = 32'h38c7cb1e;
    ram_cell[    1706] = 32'h423839bb;
    ram_cell[    1707] = 32'hed46f7ac;
    ram_cell[    1708] = 32'h3dd1cd00;
    ram_cell[    1709] = 32'he8b1fe22;
    ram_cell[    1710] = 32'h399c053c;
    ram_cell[    1711] = 32'ha08ed44a;
    ram_cell[    1712] = 32'h47856d39;
    ram_cell[    1713] = 32'h7993c4f3;
    ram_cell[    1714] = 32'hd60d3a4c;
    ram_cell[    1715] = 32'h13a81192;
    ram_cell[    1716] = 32'h4f17a018;
    ram_cell[    1717] = 32'ha9f394c1;
    ram_cell[    1718] = 32'h1c91e164;
    ram_cell[    1719] = 32'haf722679;
    ram_cell[    1720] = 32'hb5d87279;
    ram_cell[    1721] = 32'hc0877ad9;
    ram_cell[    1722] = 32'h6bb9636b;
    ram_cell[    1723] = 32'h19e31c8c;
    ram_cell[    1724] = 32'hdbed596f;
    ram_cell[    1725] = 32'he2e9a360;
    ram_cell[    1726] = 32'h0e657666;
    ram_cell[    1727] = 32'h87c0b6e1;
    ram_cell[    1728] = 32'h2096fbe1;
    ram_cell[    1729] = 32'hacbb49ea;
    ram_cell[    1730] = 32'h4317b41d;
    ram_cell[    1731] = 32'h257306e4;
    ram_cell[    1732] = 32'h5fa59ec5;
    ram_cell[    1733] = 32'hc9e0ee71;
    ram_cell[    1734] = 32'h17ccab3a;
    ram_cell[    1735] = 32'h9c874ad5;
    ram_cell[    1736] = 32'hb0d80437;
    ram_cell[    1737] = 32'he7777723;
    ram_cell[    1738] = 32'hde5bf1a3;
    ram_cell[    1739] = 32'h072149d1;
    ram_cell[    1740] = 32'h1bf99604;
    ram_cell[    1741] = 32'h72080746;
    ram_cell[    1742] = 32'h0d514fad;
    ram_cell[    1743] = 32'hd5eebad6;
    ram_cell[    1744] = 32'hea755f62;
    ram_cell[    1745] = 32'h32fee869;
    ram_cell[    1746] = 32'h9eb3de79;
    ram_cell[    1747] = 32'h4828c291;
    ram_cell[    1748] = 32'h5ad10097;
    ram_cell[    1749] = 32'h7d15b5fe;
    ram_cell[    1750] = 32'h5943bee6;
    ram_cell[    1751] = 32'hbf752342;
    ram_cell[    1752] = 32'h6e8c7c1a;
    ram_cell[    1753] = 32'h5f24e4c7;
    ram_cell[    1754] = 32'hcffb8c93;
    ram_cell[    1755] = 32'hdf3168ca;
    ram_cell[    1756] = 32'hb8f8f9d2;
    ram_cell[    1757] = 32'h2c55a2f8;
    ram_cell[    1758] = 32'hb6469d44;
    ram_cell[    1759] = 32'hcf8bbaf4;
    ram_cell[    1760] = 32'h74b6116e;
    ram_cell[    1761] = 32'h6caa791d;
    ram_cell[    1762] = 32'h64d79efc;
    ram_cell[    1763] = 32'h96437971;
    ram_cell[    1764] = 32'he8f4f84a;
    ram_cell[    1765] = 32'h0f6c35ad;
    ram_cell[    1766] = 32'ha8c099a8;
    ram_cell[    1767] = 32'h100ec2e3;
    ram_cell[    1768] = 32'hebe79289;
    ram_cell[    1769] = 32'h28bcf4c9;
    ram_cell[    1770] = 32'h6f08866c;
    ram_cell[    1771] = 32'he39d710d;
    ram_cell[    1772] = 32'hddd812c4;
    ram_cell[    1773] = 32'h2325e22f;
    ram_cell[    1774] = 32'hdfd03177;
    ram_cell[    1775] = 32'hc3452abb;
    ram_cell[    1776] = 32'h41864438;
    ram_cell[    1777] = 32'h1cbc265e;
    ram_cell[    1778] = 32'h5853c70d;
    ram_cell[    1779] = 32'h39f5eb24;
    ram_cell[    1780] = 32'h5cc94957;
    ram_cell[    1781] = 32'hf2116324;
    ram_cell[    1782] = 32'h1a248867;
    ram_cell[    1783] = 32'h56a1f79e;
    ram_cell[    1784] = 32'hb5384019;
    ram_cell[    1785] = 32'h17dcd635;
    ram_cell[    1786] = 32'hfcbcbb5a;
    ram_cell[    1787] = 32'hcdbdd447;
    ram_cell[    1788] = 32'h6340b953;
    ram_cell[    1789] = 32'h3b35e6db;
    ram_cell[    1790] = 32'h7ec1abb3;
    ram_cell[    1791] = 32'h1daea24d;
    ram_cell[    1792] = 32'hed068de0;
    ram_cell[    1793] = 32'hfd78e124;
    ram_cell[    1794] = 32'h05b096b6;
    ram_cell[    1795] = 32'hb06499eb;
    ram_cell[    1796] = 32'hcbd4bf1b;
    ram_cell[    1797] = 32'h232c77fd;
    ram_cell[    1798] = 32'hde330d9c;
    ram_cell[    1799] = 32'h44f42af6;
    ram_cell[    1800] = 32'h7876b0aa;
    ram_cell[    1801] = 32'hfa5ecfc8;
    ram_cell[    1802] = 32'he7a3f1bd;
    ram_cell[    1803] = 32'h4fb506d3;
    ram_cell[    1804] = 32'hf6adcb69;
    ram_cell[    1805] = 32'h41cf7395;
    ram_cell[    1806] = 32'h0b93e4af;
    ram_cell[    1807] = 32'h416e58cf;
    ram_cell[    1808] = 32'hc4d82d24;
    ram_cell[    1809] = 32'h8a50a344;
    ram_cell[    1810] = 32'h2760b257;
    ram_cell[    1811] = 32'h46771bee;
    ram_cell[    1812] = 32'h079cd30b;
    ram_cell[    1813] = 32'h0d615149;
    ram_cell[    1814] = 32'h4a11a04a;
    ram_cell[    1815] = 32'hbf0283ce;
    ram_cell[    1816] = 32'h822416de;
    ram_cell[    1817] = 32'hc4295d2c;
    ram_cell[    1818] = 32'he8891fb3;
    ram_cell[    1819] = 32'h581243c5;
    ram_cell[    1820] = 32'h9f23b894;
    ram_cell[    1821] = 32'hf4d81906;
    ram_cell[    1822] = 32'h99d9ddd9;
    ram_cell[    1823] = 32'h28ccc630;
    ram_cell[    1824] = 32'h5d8c89b4;
    ram_cell[    1825] = 32'h5247252e;
    ram_cell[    1826] = 32'h791e99ed;
    ram_cell[    1827] = 32'hee5bd111;
    ram_cell[    1828] = 32'h3d0a276a;
    ram_cell[    1829] = 32'hff5c0521;
    ram_cell[    1830] = 32'hab52dd68;
    ram_cell[    1831] = 32'he6ca8f07;
    ram_cell[    1832] = 32'h1dcc613b;
    ram_cell[    1833] = 32'hd4cb003c;
    ram_cell[    1834] = 32'he2192d6a;
    ram_cell[    1835] = 32'h02f1856d;
    ram_cell[    1836] = 32'h9de8ce80;
    ram_cell[    1837] = 32'h6569210e;
    ram_cell[    1838] = 32'h0db909b0;
    ram_cell[    1839] = 32'hce81c27b;
    ram_cell[    1840] = 32'hed7bae92;
    ram_cell[    1841] = 32'h5cc6cb05;
    ram_cell[    1842] = 32'h8049f1ec;
    ram_cell[    1843] = 32'ha8f1e04f;
    ram_cell[    1844] = 32'h0dfd6953;
    ram_cell[    1845] = 32'h868a8600;
    ram_cell[    1846] = 32'h1f553bf9;
    ram_cell[    1847] = 32'h461748c6;
    ram_cell[    1848] = 32'h93b6d9f3;
    ram_cell[    1849] = 32'ha1bb312f;
    ram_cell[    1850] = 32'h6dca561b;
    ram_cell[    1851] = 32'hb8593005;
    ram_cell[    1852] = 32'ha5f48876;
    ram_cell[    1853] = 32'h9df533f4;
    ram_cell[    1854] = 32'h7e9ef7cd;
    ram_cell[    1855] = 32'h7bb9d930;
    ram_cell[    1856] = 32'h002eec49;
    ram_cell[    1857] = 32'hbddc0d92;
    ram_cell[    1858] = 32'h46427b0d;
    ram_cell[    1859] = 32'hd7a11923;
    ram_cell[    1860] = 32'h7bc2fc5a;
    ram_cell[    1861] = 32'hafa22a2e;
    ram_cell[    1862] = 32'hcf8d7169;
    ram_cell[    1863] = 32'hf9f2cb49;
    ram_cell[    1864] = 32'he287543f;
    ram_cell[    1865] = 32'hd1eada3a;
    ram_cell[    1866] = 32'hb1f47e4d;
    ram_cell[    1867] = 32'h818a5a7b;
    ram_cell[    1868] = 32'h6473b2d9;
    ram_cell[    1869] = 32'h97f5e97c;
    ram_cell[    1870] = 32'h3e2b6a2e;
    ram_cell[    1871] = 32'h668e4ba1;
    ram_cell[    1872] = 32'h789191ec;
    ram_cell[    1873] = 32'h543b6a21;
    ram_cell[    1874] = 32'hb5caf38f;
    ram_cell[    1875] = 32'h29429e27;
    ram_cell[    1876] = 32'h9d92ae3d;
    ram_cell[    1877] = 32'he4270aea;
    ram_cell[    1878] = 32'hdd9f3e59;
    ram_cell[    1879] = 32'h47998fc7;
    ram_cell[    1880] = 32'h492dd85c;
    ram_cell[    1881] = 32'h7e13ed53;
    ram_cell[    1882] = 32'h22aa30c9;
    ram_cell[    1883] = 32'h48c90e7b;
    ram_cell[    1884] = 32'ha9cf6909;
    ram_cell[    1885] = 32'hbefba4b6;
    ram_cell[    1886] = 32'h0f241895;
    ram_cell[    1887] = 32'hbbc23f77;
    ram_cell[    1888] = 32'hfad67dcc;
    ram_cell[    1889] = 32'hd53b4352;
    ram_cell[    1890] = 32'h421323a7;
    ram_cell[    1891] = 32'h776f3094;
    ram_cell[    1892] = 32'hde710dec;
    ram_cell[    1893] = 32'hfb415c1f;
    ram_cell[    1894] = 32'h4d7f2d94;
    ram_cell[    1895] = 32'hf0771cb2;
    ram_cell[    1896] = 32'hd668c9d6;
    ram_cell[    1897] = 32'h1454f07d;
    ram_cell[    1898] = 32'h0d9f2dc7;
    ram_cell[    1899] = 32'h6235bca0;
    ram_cell[    1900] = 32'h8feb6d99;
    ram_cell[    1901] = 32'h98ca5220;
    ram_cell[    1902] = 32'h219fcca3;
    ram_cell[    1903] = 32'h5ad358b3;
    ram_cell[    1904] = 32'heef290f0;
    ram_cell[    1905] = 32'hf0c4fdd1;
    ram_cell[    1906] = 32'h1d1b7009;
    ram_cell[    1907] = 32'hcdeaedda;
    ram_cell[    1908] = 32'hf18d430a;
    ram_cell[    1909] = 32'h46e83269;
    ram_cell[    1910] = 32'h73929c2a;
    ram_cell[    1911] = 32'h37f29d8a;
    ram_cell[    1912] = 32'hd6f8e9ed;
    ram_cell[    1913] = 32'hc63e7884;
    ram_cell[    1914] = 32'h903d958f;
    ram_cell[    1915] = 32'h7f341b82;
    ram_cell[    1916] = 32'h1938eee0;
    ram_cell[    1917] = 32'hd4d99179;
    ram_cell[    1918] = 32'h38e652e5;
    ram_cell[    1919] = 32'h3aa6edb7;
    ram_cell[    1920] = 32'h9bf3b3a3;
    ram_cell[    1921] = 32'h257d8963;
    ram_cell[    1922] = 32'h22f545ae;
    ram_cell[    1923] = 32'hc9d23283;
    ram_cell[    1924] = 32'hdbc52341;
    ram_cell[    1925] = 32'hc45d7e97;
    ram_cell[    1926] = 32'hc0efec22;
    ram_cell[    1927] = 32'h92e7deca;
    ram_cell[    1928] = 32'h55e8d905;
    ram_cell[    1929] = 32'ha30a7b27;
    ram_cell[    1930] = 32'h679a7256;
    ram_cell[    1931] = 32'h7822d1f4;
    ram_cell[    1932] = 32'h2d3cfbe7;
    ram_cell[    1933] = 32'he5f0fcdc;
    ram_cell[    1934] = 32'ha2992b9e;
    ram_cell[    1935] = 32'h072a9baf;
    ram_cell[    1936] = 32'h0e494000;
    ram_cell[    1937] = 32'h96b8a8fb;
    ram_cell[    1938] = 32'h2b27e61e;
    ram_cell[    1939] = 32'h2c3cc87c;
    ram_cell[    1940] = 32'h2d8116c9;
    ram_cell[    1941] = 32'hf8502b75;
    ram_cell[    1942] = 32'h8dd54896;
    ram_cell[    1943] = 32'h02c5e181;
    ram_cell[    1944] = 32'hb834d055;
    ram_cell[    1945] = 32'hc8323017;
    ram_cell[    1946] = 32'hd29c0a78;
    ram_cell[    1947] = 32'h6010f28f;
    ram_cell[    1948] = 32'h674adbaf;
    ram_cell[    1949] = 32'h27dfda5a;
    ram_cell[    1950] = 32'hc61b86a5;
    ram_cell[    1951] = 32'h30711653;
    ram_cell[    1952] = 32'hbceeb823;
    ram_cell[    1953] = 32'h4f6d14db;
    ram_cell[    1954] = 32'h3fdd73e7;
    ram_cell[    1955] = 32'haa818247;
    ram_cell[    1956] = 32'hd4da43ef;
    ram_cell[    1957] = 32'hd03d0fae;
    ram_cell[    1958] = 32'h7c0966fd;
    ram_cell[    1959] = 32'h406a9cb3;
    ram_cell[    1960] = 32'h1f35be19;
    ram_cell[    1961] = 32'h03493253;
    ram_cell[    1962] = 32'h73503101;
    ram_cell[    1963] = 32'h4013f876;
    ram_cell[    1964] = 32'hddcdf84e;
    ram_cell[    1965] = 32'hebf6e485;
    ram_cell[    1966] = 32'ha1c6f552;
    ram_cell[    1967] = 32'h71bf8cac;
    ram_cell[    1968] = 32'h35b0e48f;
    ram_cell[    1969] = 32'ha29ddfc9;
    ram_cell[    1970] = 32'h4981392c;
    ram_cell[    1971] = 32'hc887719f;
    ram_cell[    1972] = 32'hc81df036;
    ram_cell[    1973] = 32'h2b94dee7;
    ram_cell[    1974] = 32'had205cc4;
    ram_cell[    1975] = 32'h5bdab47b;
    ram_cell[    1976] = 32'h3c86194b;
    ram_cell[    1977] = 32'h0e67cfe9;
    ram_cell[    1978] = 32'h7d80bf85;
    ram_cell[    1979] = 32'hf00eb1dc;
    ram_cell[    1980] = 32'h6c68b8de;
    ram_cell[    1981] = 32'h5f4c6f64;
    ram_cell[    1982] = 32'he5655fe6;
    ram_cell[    1983] = 32'h3129ee4e;
    ram_cell[    1984] = 32'hd3881ad4;
    ram_cell[    1985] = 32'hd5e62d87;
    ram_cell[    1986] = 32'h95bdb0be;
    ram_cell[    1987] = 32'h491648a0;
    ram_cell[    1988] = 32'h5a253a8e;
    ram_cell[    1989] = 32'h2888f41f;
    ram_cell[    1990] = 32'h7d3e32a1;
    ram_cell[    1991] = 32'h0f2b014e;
    ram_cell[    1992] = 32'hf61c83cf;
    ram_cell[    1993] = 32'hb4ca85f2;
    ram_cell[    1994] = 32'h9c988495;
    ram_cell[    1995] = 32'hf1ec9bc7;
    ram_cell[    1996] = 32'h12f9df84;
    ram_cell[    1997] = 32'hc4e4c9f5;
    ram_cell[    1998] = 32'h3ab1405e;
    ram_cell[    1999] = 32'h91464fb9;
    ram_cell[    2000] = 32'h42bc9142;
    ram_cell[    2001] = 32'hc3e2a158;
    ram_cell[    2002] = 32'h04b0df81;
    ram_cell[    2003] = 32'h7d8f905f;
    ram_cell[    2004] = 32'h5decc6a8;
    ram_cell[    2005] = 32'hc248cd6e;
    ram_cell[    2006] = 32'he9ee9ab0;
    ram_cell[    2007] = 32'h24ac5f82;
    ram_cell[    2008] = 32'hd96f74be;
    ram_cell[    2009] = 32'h0270336b;
    ram_cell[    2010] = 32'h9f96294f;
    ram_cell[    2011] = 32'h8ee4970b;
    ram_cell[    2012] = 32'he073aefe;
    ram_cell[    2013] = 32'h9d6bae2c;
    ram_cell[    2014] = 32'hb28ee152;
    ram_cell[    2015] = 32'h9eaa475a;
    ram_cell[    2016] = 32'h6f8240fd;
    ram_cell[    2017] = 32'hd1be4e55;
    ram_cell[    2018] = 32'hf29b0e2c;
    ram_cell[    2019] = 32'h073dc576;
    ram_cell[    2020] = 32'h409d97a1;
    ram_cell[    2021] = 32'h1d1623af;
    ram_cell[    2022] = 32'h29d1fc9b;
    ram_cell[    2023] = 32'haeac58ea;
    ram_cell[    2024] = 32'h94f5b25e;
    ram_cell[    2025] = 32'h7e523bdf;
    ram_cell[    2026] = 32'h405612e8;
    ram_cell[    2027] = 32'he07e10e9;
    ram_cell[    2028] = 32'ha5f1c815;
    ram_cell[    2029] = 32'h5b2683c7;
    ram_cell[    2030] = 32'h4e838337;
    ram_cell[    2031] = 32'h3e6c95db;
    ram_cell[    2032] = 32'h6ad0eb70;
    ram_cell[    2033] = 32'h9cce40cb;
    ram_cell[    2034] = 32'h6de7b74d;
    ram_cell[    2035] = 32'h15726079;
    ram_cell[    2036] = 32'hf0dbb225;
    ram_cell[    2037] = 32'h6200ff73;
    ram_cell[    2038] = 32'h30c22182;
    ram_cell[    2039] = 32'he116706c;
    ram_cell[    2040] = 32'hed461acf;
    ram_cell[    2041] = 32'h496b3e05;
    ram_cell[    2042] = 32'h44f7ed64;
    ram_cell[    2043] = 32'hb5df74d1;
    ram_cell[    2044] = 32'h89257420;
    ram_cell[    2045] = 32'hbeb65faa;
    ram_cell[    2046] = 32'hec913939;
    ram_cell[    2047] = 32'h31961820;
    // src matrix B
    ram_cell[    2048] = 32'h7ccdd257;
    ram_cell[    2049] = 32'hfa6255a0;
    ram_cell[    2050] = 32'h38014a49;
    ram_cell[    2051] = 32'hd7e39371;
    ram_cell[    2052] = 32'hcc62a62d;
    ram_cell[    2053] = 32'h18ac2e3d;
    ram_cell[    2054] = 32'h68d2664e;
    ram_cell[    2055] = 32'h9ff93968;
    ram_cell[    2056] = 32'h5f50811b;
    ram_cell[    2057] = 32'h0cddbbb9;
    ram_cell[    2058] = 32'h6883d2a4;
    ram_cell[    2059] = 32'h21bc4da3;
    ram_cell[    2060] = 32'h7de474be;
    ram_cell[    2061] = 32'haea8deb9;
    ram_cell[    2062] = 32'hea38f067;
    ram_cell[    2063] = 32'ha6270087;
    ram_cell[    2064] = 32'h8bf9c800;
    ram_cell[    2065] = 32'h756ebdb9;
    ram_cell[    2066] = 32'h05146c4b;
    ram_cell[    2067] = 32'h5df7a3e5;
    ram_cell[    2068] = 32'hdac7b3ca;
    ram_cell[    2069] = 32'heba94291;
    ram_cell[    2070] = 32'h304306df;
    ram_cell[    2071] = 32'he849a2e2;
    ram_cell[    2072] = 32'h8e89bdce;
    ram_cell[    2073] = 32'hfc8ea3ec;
    ram_cell[    2074] = 32'hbe5a18d0;
    ram_cell[    2075] = 32'h772fb8d4;
    ram_cell[    2076] = 32'ha8a3e408;
    ram_cell[    2077] = 32'h95b59de0;
    ram_cell[    2078] = 32'h76cc6d3e;
    ram_cell[    2079] = 32'h6ffbe7ed;
    ram_cell[    2080] = 32'hd8d65252;
    ram_cell[    2081] = 32'hcfc190aa;
    ram_cell[    2082] = 32'h9acbb625;
    ram_cell[    2083] = 32'ha73c77d3;
    ram_cell[    2084] = 32'h35ee4b35;
    ram_cell[    2085] = 32'ha7692248;
    ram_cell[    2086] = 32'ha618ce76;
    ram_cell[    2087] = 32'h0793ae28;
    ram_cell[    2088] = 32'h4e8a72af;
    ram_cell[    2089] = 32'hcb171718;
    ram_cell[    2090] = 32'h2c7ea5d4;
    ram_cell[    2091] = 32'h5fff70de;
    ram_cell[    2092] = 32'h377e6f39;
    ram_cell[    2093] = 32'h3f20b1c6;
    ram_cell[    2094] = 32'h8e6bb7fe;
    ram_cell[    2095] = 32'ha4a39ec6;
    ram_cell[    2096] = 32'h77eaf198;
    ram_cell[    2097] = 32'h90598e24;
    ram_cell[    2098] = 32'h93f9b132;
    ram_cell[    2099] = 32'h4aa10ff4;
    ram_cell[    2100] = 32'hd85f0530;
    ram_cell[    2101] = 32'h5e951740;
    ram_cell[    2102] = 32'hfbdf2f47;
    ram_cell[    2103] = 32'ha0b0fcd7;
    ram_cell[    2104] = 32'h38f02605;
    ram_cell[    2105] = 32'h70018715;
    ram_cell[    2106] = 32'ha92f8aaa;
    ram_cell[    2107] = 32'h2145c5d2;
    ram_cell[    2108] = 32'h068cceae;
    ram_cell[    2109] = 32'hef1ff7a8;
    ram_cell[    2110] = 32'hcae16607;
    ram_cell[    2111] = 32'hd3be0a65;
    ram_cell[    2112] = 32'h3659a6d4;
    ram_cell[    2113] = 32'h6eabc882;
    ram_cell[    2114] = 32'hf240a1fa;
    ram_cell[    2115] = 32'hd443997b;
    ram_cell[    2116] = 32'h6c64df76;
    ram_cell[    2117] = 32'h16b1e34f;
    ram_cell[    2118] = 32'hb8be07ca;
    ram_cell[    2119] = 32'hd7fbd6ac;
    ram_cell[    2120] = 32'h3ac2d722;
    ram_cell[    2121] = 32'hfa1c643b;
    ram_cell[    2122] = 32'h5dd58ba1;
    ram_cell[    2123] = 32'h63d20d5b;
    ram_cell[    2124] = 32'hade5fdd2;
    ram_cell[    2125] = 32'ha71c088d;
    ram_cell[    2126] = 32'h08c41083;
    ram_cell[    2127] = 32'h4ac2c367;
    ram_cell[    2128] = 32'hf66ebf21;
    ram_cell[    2129] = 32'h1d2736a3;
    ram_cell[    2130] = 32'h680e5fe6;
    ram_cell[    2131] = 32'hbb4d4494;
    ram_cell[    2132] = 32'hd94f86cd;
    ram_cell[    2133] = 32'h9209bb2e;
    ram_cell[    2134] = 32'h61c98e78;
    ram_cell[    2135] = 32'hf800606d;
    ram_cell[    2136] = 32'h52eab98f;
    ram_cell[    2137] = 32'he24c7f82;
    ram_cell[    2138] = 32'hb3915851;
    ram_cell[    2139] = 32'hd433e02f;
    ram_cell[    2140] = 32'hda3cb04e;
    ram_cell[    2141] = 32'h4aa046ef;
    ram_cell[    2142] = 32'h05b166ad;
    ram_cell[    2143] = 32'hcaf55bbe;
    ram_cell[    2144] = 32'h6dee176e;
    ram_cell[    2145] = 32'hc164d9d5;
    ram_cell[    2146] = 32'h8622f721;
    ram_cell[    2147] = 32'hd17f9f3d;
    ram_cell[    2148] = 32'hea7c7ce0;
    ram_cell[    2149] = 32'h38d1ebd2;
    ram_cell[    2150] = 32'hcbcb4f39;
    ram_cell[    2151] = 32'hbdddfb5b;
    ram_cell[    2152] = 32'hc9a1694e;
    ram_cell[    2153] = 32'h29882713;
    ram_cell[    2154] = 32'h7c724ffa;
    ram_cell[    2155] = 32'hf773641d;
    ram_cell[    2156] = 32'h1909b379;
    ram_cell[    2157] = 32'h8b55ce97;
    ram_cell[    2158] = 32'h55ed68ec;
    ram_cell[    2159] = 32'h5933ee03;
    ram_cell[    2160] = 32'h064b4ab1;
    ram_cell[    2161] = 32'h8ce77745;
    ram_cell[    2162] = 32'h20cbcb7f;
    ram_cell[    2163] = 32'hf33a7f15;
    ram_cell[    2164] = 32'ha87c29c1;
    ram_cell[    2165] = 32'h99e649bb;
    ram_cell[    2166] = 32'hfb843f6b;
    ram_cell[    2167] = 32'h47fd5576;
    ram_cell[    2168] = 32'he3ecbeef;
    ram_cell[    2169] = 32'h32edef16;
    ram_cell[    2170] = 32'h4c2e2336;
    ram_cell[    2171] = 32'h1d696c31;
    ram_cell[    2172] = 32'h67a22c46;
    ram_cell[    2173] = 32'h73b693b7;
    ram_cell[    2174] = 32'h6fa9cf40;
    ram_cell[    2175] = 32'hd87b099e;
    ram_cell[    2176] = 32'hfdef2bad;
    ram_cell[    2177] = 32'hfa55ba0d;
    ram_cell[    2178] = 32'h3b646780;
    ram_cell[    2179] = 32'ha253118b;
    ram_cell[    2180] = 32'h7bb2bfef;
    ram_cell[    2181] = 32'h32d041e8;
    ram_cell[    2182] = 32'hd478ab50;
    ram_cell[    2183] = 32'hf9f93dd2;
    ram_cell[    2184] = 32'h6d5465fa;
    ram_cell[    2185] = 32'h0555436e;
    ram_cell[    2186] = 32'h800f0d95;
    ram_cell[    2187] = 32'hd88344d2;
    ram_cell[    2188] = 32'h28e55e80;
    ram_cell[    2189] = 32'hf4ef89ca;
    ram_cell[    2190] = 32'h29d9ff47;
    ram_cell[    2191] = 32'heff48a76;
    ram_cell[    2192] = 32'h5ce44f98;
    ram_cell[    2193] = 32'h41a21e70;
    ram_cell[    2194] = 32'hf5beaf05;
    ram_cell[    2195] = 32'h03fe2081;
    ram_cell[    2196] = 32'hacf6c562;
    ram_cell[    2197] = 32'h8f49634b;
    ram_cell[    2198] = 32'he2059f58;
    ram_cell[    2199] = 32'h09e72adf;
    ram_cell[    2200] = 32'h19f7727d;
    ram_cell[    2201] = 32'h8cf1f27e;
    ram_cell[    2202] = 32'hffa582a3;
    ram_cell[    2203] = 32'h8a2b17ae;
    ram_cell[    2204] = 32'h11784555;
    ram_cell[    2205] = 32'he2b74a77;
    ram_cell[    2206] = 32'h9fa04dd5;
    ram_cell[    2207] = 32'hdc755a1b;
    ram_cell[    2208] = 32'h47cec220;
    ram_cell[    2209] = 32'h52d0bde0;
    ram_cell[    2210] = 32'h753ad620;
    ram_cell[    2211] = 32'h3cc16585;
    ram_cell[    2212] = 32'hc31db591;
    ram_cell[    2213] = 32'haaec9861;
    ram_cell[    2214] = 32'h59b375b8;
    ram_cell[    2215] = 32'h69bb5e3d;
    ram_cell[    2216] = 32'h2877acd2;
    ram_cell[    2217] = 32'h0d870f28;
    ram_cell[    2218] = 32'h6db6b11e;
    ram_cell[    2219] = 32'h3af18dc0;
    ram_cell[    2220] = 32'ha0d8cbe8;
    ram_cell[    2221] = 32'h107357d3;
    ram_cell[    2222] = 32'h3911d285;
    ram_cell[    2223] = 32'hc7cafb9d;
    ram_cell[    2224] = 32'hed1821cc;
    ram_cell[    2225] = 32'h82dfcb67;
    ram_cell[    2226] = 32'h4081afe9;
    ram_cell[    2227] = 32'h0197eaa8;
    ram_cell[    2228] = 32'h306237c9;
    ram_cell[    2229] = 32'hf49b89c1;
    ram_cell[    2230] = 32'h65d501df;
    ram_cell[    2231] = 32'hab7fe113;
    ram_cell[    2232] = 32'h03636827;
    ram_cell[    2233] = 32'h7dd4fc50;
    ram_cell[    2234] = 32'hcbe1728a;
    ram_cell[    2235] = 32'h2f73164c;
    ram_cell[    2236] = 32'h4dd3522e;
    ram_cell[    2237] = 32'ha27f2605;
    ram_cell[    2238] = 32'ha5692aaa;
    ram_cell[    2239] = 32'h7f08bb08;
    ram_cell[    2240] = 32'h8dd74c9a;
    ram_cell[    2241] = 32'h7b1c4201;
    ram_cell[    2242] = 32'h45fdad85;
    ram_cell[    2243] = 32'h42f3ad8a;
    ram_cell[    2244] = 32'h85aabd48;
    ram_cell[    2245] = 32'h31cd2e8e;
    ram_cell[    2246] = 32'h2d0771e4;
    ram_cell[    2247] = 32'h32fba61c;
    ram_cell[    2248] = 32'h083ca987;
    ram_cell[    2249] = 32'h6c7bc597;
    ram_cell[    2250] = 32'h80c5f1bc;
    ram_cell[    2251] = 32'h861c8baf;
    ram_cell[    2252] = 32'h852798cb;
    ram_cell[    2253] = 32'haa3a3681;
    ram_cell[    2254] = 32'h30b15e3a;
    ram_cell[    2255] = 32'hf1c1e912;
    ram_cell[    2256] = 32'habff960f;
    ram_cell[    2257] = 32'h92d1d89d;
    ram_cell[    2258] = 32'hfb167776;
    ram_cell[    2259] = 32'h6659bb24;
    ram_cell[    2260] = 32'hacb150db;
    ram_cell[    2261] = 32'hb599a5f4;
    ram_cell[    2262] = 32'hd902aed0;
    ram_cell[    2263] = 32'h3d7f0a1a;
    ram_cell[    2264] = 32'h2b944682;
    ram_cell[    2265] = 32'h7f4406ee;
    ram_cell[    2266] = 32'h2c78827f;
    ram_cell[    2267] = 32'h501170ab;
    ram_cell[    2268] = 32'h6deeb58f;
    ram_cell[    2269] = 32'h33ee52b9;
    ram_cell[    2270] = 32'h06048c7d;
    ram_cell[    2271] = 32'h0c9296a8;
    ram_cell[    2272] = 32'haf6214d4;
    ram_cell[    2273] = 32'h85cb1114;
    ram_cell[    2274] = 32'ha852ef68;
    ram_cell[    2275] = 32'hfe5dae1e;
    ram_cell[    2276] = 32'hf4cb6931;
    ram_cell[    2277] = 32'h9d06f615;
    ram_cell[    2278] = 32'h66c45df5;
    ram_cell[    2279] = 32'h4ea06242;
    ram_cell[    2280] = 32'h79ae3e45;
    ram_cell[    2281] = 32'h8691c498;
    ram_cell[    2282] = 32'h03224870;
    ram_cell[    2283] = 32'h357b9db4;
    ram_cell[    2284] = 32'heb0a8d79;
    ram_cell[    2285] = 32'h4862d07f;
    ram_cell[    2286] = 32'habcda148;
    ram_cell[    2287] = 32'h956375d3;
    ram_cell[    2288] = 32'h05c79667;
    ram_cell[    2289] = 32'h6dbcdee4;
    ram_cell[    2290] = 32'h19e3610b;
    ram_cell[    2291] = 32'hbc5ae265;
    ram_cell[    2292] = 32'h0a4c2d04;
    ram_cell[    2293] = 32'hfb09f578;
    ram_cell[    2294] = 32'haa1ec871;
    ram_cell[    2295] = 32'hf57a9ad9;
    ram_cell[    2296] = 32'h4cb43b69;
    ram_cell[    2297] = 32'h9343bd94;
    ram_cell[    2298] = 32'h71cc01ab;
    ram_cell[    2299] = 32'h397c7b16;
    ram_cell[    2300] = 32'h69ad3605;
    ram_cell[    2301] = 32'hdae336c2;
    ram_cell[    2302] = 32'h38ddc069;
    ram_cell[    2303] = 32'h81046abf;
    ram_cell[    2304] = 32'h414e9a8f;
    ram_cell[    2305] = 32'h6945b1a4;
    ram_cell[    2306] = 32'h15c0dc95;
    ram_cell[    2307] = 32'hcd3e0a6f;
    ram_cell[    2308] = 32'h03f40824;
    ram_cell[    2309] = 32'h8f51e6de;
    ram_cell[    2310] = 32'h4a135375;
    ram_cell[    2311] = 32'hd544ab36;
    ram_cell[    2312] = 32'h50b9ecc0;
    ram_cell[    2313] = 32'hd86a9d4c;
    ram_cell[    2314] = 32'hcbc62cf0;
    ram_cell[    2315] = 32'hedf10229;
    ram_cell[    2316] = 32'h57501ab3;
    ram_cell[    2317] = 32'h0d020f38;
    ram_cell[    2318] = 32'h8d09abbf;
    ram_cell[    2319] = 32'h5dc5e221;
    ram_cell[    2320] = 32'h2406cca8;
    ram_cell[    2321] = 32'h26bd99c6;
    ram_cell[    2322] = 32'he7d479e1;
    ram_cell[    2323] = 32'hfee14536;
    ram_cell[    2324] = 32'h6c72aa31;
    ram_cell[    2325] = 32'h7ec70902;
    ram_cell[    2326] = 32'h88809995;
    ram_cell[    2327] = 32'he7a86f62;
    ram_cell[    2328] = 32'ha8882897;
    ram_cell[    2329] = 32'he45b8bf0;
    ram_cell[    2330] = 32'hfc1f2198;
    ram_cell[    2331] = 32'h816c502b;
    ram_cell[    2332] = 32'hde5896f3;
    ram_cell[    2333] = 32'h99edbf83;
    ram_cell[    2334] = 32'h7209cf66;
    ram_cell[    2335] = 32'hab1e38b5;
    ram_cell[    2336] = 32'h5805a181;
    ram_cell[    2337] = 32'h48c3eab1;
    ram_cell[    2338] = 32'h9004d0fc;
    ram_cell[    2339] = 32'h6a9766ed;
    ram_cell[    2340] = 32'hfb84daaf;
    ram_cell[    2341] = 32'h5de9a6f6;
    ram_cell[    2342] = 32'hce46c89c;
    ram_cell[    2343] = 32'h9df9b9cb;
    ram_cell[    2344] = 32'hb8bfbee8;
    ram_cell[    2345] = 32'he28ba66b;
    ram_cell[    2346] = 32'hece3f2a0;
    ram_cell[    2347] = 32'h42b42c39;
    ram_cell[    2348] = 32'hf0b90362;
    ram_cell[    2349] = 32'h2419e818;
    ram_cell[    2350] = 32'h870a74fc;
    ram_cell[    2351] = 32'hd526f602;
    ram_cell[    2352] = 32'h845fcabf;
    ram_cell[    2353] = 32'ha4e51e23;
    ram_cell[    2354] = 32'hd92bfc5a;
    ram_cell[    2355] = 32'h2468f061;
    ram_cell[    2356] = 32'hee53be14;
    ram_cell[    2357] = 32'h68c6495c;
    ram_cell[    2358] = 32'h3c074b1d;
    ram_cell[    2359] = 32'h4d94e622;
    ram_cell[    2360] = 32'hd89cc464;
    ram_cell[    2361] = 32'hb51f4646;
    ram_cell[    2362] = 32'h091633cb;
    ram_cell[    2363] = 32'h9eda8820;
    ram_cell[    2364] = 32'hc5222de4;
    ram_cell[    2365] = 32'h5e9a4506;
    ram_cell[    2366] = 32'hf5512561;
    ram_cell[    2367] = 32'h268b5a1b;
    ram_cell[    2368] = 32'h250151a7;
    ram_cell[    2369] = 32'h31d94771;
    ram_cell[    2370] = 32'hb7293f25;
    ram_cell[    2371] = 32'had663d14;
    ram_cell[    2372] = 32'hb7fe7814;
    ram_cell[    2373] = 32'hf74ca643;
    ram_cell[    2374] = 32'hc56e6ead;
    ram_cell[    2375] = 32'hb59c8a0a;
    ram_cell[    2376] = 32'h347a0520;
    ram_cell[    2377] = 32'hb557c3dc;
    ram_cell[    2378] = 32'h0236847a;
    ram_cell[    2379] = 32'h95765182;
    ram_cell[    2380] = 32'h392b1e12;
    ram_cell[    2381] = 32'h1e6ceebc;
    ram_cell[    2382] = 32'hc185a02d;
    ram_cell[    2383] = 32'h6544cdff;
    ram_cell[    2384] = 32'hcfe2e68c;
    ram_cell[    2385] = 32'h918674d3;
    ram_cell[    2386] = 32'h3559dd93;
    ram_cell[    2387] = 32'h63c3239b;
    ram_cell[    2388] = 32'h8d0abbfb;
    ram_cell[    2389] = 32'h6340f6cf;
    ram_cell[    2390] = 32'h0c4dd192;
    ram_cell[    2391] = 32'h9e766c51;
    ram_cell[    2392] = 32'h71c295b8;
    ram_cell[    2393] = 32'h375db63c;
    ram_cell[    2394] = 32'hdf6c372c;
    ram_cell[    2395] = 32'hbef98f96;
    ram_cell[    2396] = 32'hb9b243d3;
    ram_cell[    2397] = 32'h0818ee76;
    ram_cell[    2398] = 32'h7e1824c3;
    ram_cell[    2399] = 32'hcdd6ab76;
    ram_cell[    2400] = 32'h0ef8cf73;
    ram_cell[    2401] = 32'hfab56b07;
    ram_cell[    2402] = 32'h3b2806b6;
    ram_cell[    2403] = 32'h7eb0796d;
    ram_cell[    2404] = 32'h9624ce2c;
    ram_cell[    2405] = 32'h10a283b2;
    ram_cell[    2406] = 32'h2c424ae5;
    ram_cell[    2407] = 32'ha22e4a63;
    ram_cell[    2408] = 32'h8b2a6629;
    ram_cell[    2409] = 32'h11462084;
    ram_cell[    2410] = 32'h57924135;
    ram_cell[    2411] = 32'h52173c43;
    ram_cell[    2412] = 32'hb253e227;
    ram_cell[    2413] = 32'h51ff2a81;
    ram_cell[    2414] = 32'hdc48499b;
    ram_cell[    2415] = 32'h0bb45ab3;
    ram_cell[    2416] = 32'h726f1308;
    ram_cell[    2417] = 32'h81a40913;
    ram_cell[    2418] = 32'h0249c0af;
    ram_cell[    2419] = 32'ha666f6b8;
    ram_cell[    2420] = 32'h9fb5a615;
    ram_cell[    2421] = 32'he45299d5;
    ram_cell[    2422] = 32'h074e8995;
    ram_cell[    2423] = 32'h213b6b8f;
    ram_cell[    2424] = 32'h115fb7d4;
    ram_cell[    2425] = 32'hebc08cc5;
    ram_cell[    2426] = 32'hffc8e689;
    ram_cell[    2427] = 32'h7cc63789;
    ram_cell[    2428] = 32'h8003ba9e;
    ram_cell[    2429] = 32'h06fc01e3;
    ram_cell[    2430] = 32'hb62167d6;
    ram_cell[    2431] = 32'h8e5b8492;
    ram_cell[    2432] = 32'h86d904a7;
    ram_cell[    2433] = 32'h99c88491;
    ram_cell[    2434] = 32'hf2e2a324;
    ram_cell[    2435] = 32'hda8c2dfb;
    ram_cell[    2436] = 32'h4d045541;
    ram_cell[    2437] = 32'hef89e8b4;
    ram_cell[    2438] = 32'hfa54cd5a;
    ram_cell[    2439] = 32'h834e09a0;
    ram_cell[    2440] = 32'h7e4975a5;
    ram_cell[    2441] = 32'h457e1e8b;
    ram_cell[    2442] = 32'h5b827c23;
    ram_cell[    2443] = 32'h8b431d14;
    ram_cell[    2444] = 32'hbb2f810b;
    ram_cell[    2445] = 32'he8c83db0;
    ram_cell[    2446] = 32'hd818cf43;
    ram_cell[    2447] = 32'hf31daf58;
    ram_cell[    2448] = 32'h87319dc7;
    ram_cell[    2449] = 32'h1e84e006;
    ram_cell[    2450] = 32'hce8b6ee0;
    ram_cell[    2451] = 32'h0a648b2b;
    ram_cell[    2452] = 32'hde3a43bb;
    ram_cell[    2453] = 32'h351e978b;
    ram_cell[    2454] = 32'h909f8ab3;
    ram_cell[    2455] = 32'heb775639;
    ram_cell[    2456] = 32'hb765cf32;
    ram_cell[    2457] = 32'hd1da4248;
    ram_cell[    2458] = 32'h47d8f9f5;
    ram_cell[    2459] = 32'hc99e23d1;
    ram_cell[    2460] = 32'hd9676e04;
    ram_cell[    2461] = 32'h513a28ae;
    ram_cell[    2462] = 32'h33279878;
    ram_cell[    2463] = 32'h7826a03e;
    ram_cell[    2464] = 32'h71832c19;
    ram_cell[    2465] = 32'h3c78e265;
    ram_cell[    2466] = 32'hc7c553b0;
    ram_cell[    2467] = 32'hd2e9977b;
    ram_cell[    2468] = 32'he4211167;
    ram_cell[    2469] = 32'hd60ac0d9;
    ram_cell[    2470] = 32'h1f225bdc;
    ram_cell[    2471] = 32'h39fba48d;
    ram_cell[    2472] = 32'h2d88c8f1;
    ram_cell[    2473] = 32'h3d654d3a;
    ram_cell[    2474] = 32'h47eb1c1a;
    ram_cell[    2475] = 32'haac6113e;
    ram_cell[    2476] = 32'hd332ecf8;
    ram_cell[    2477] = 32'h0f56ab59;
    ram_cell[    2478] = 32'h6b8aa049;
    ram_cell[    2479] = 32'h8bd5e008;
    ram_cell[    2480] = 32'h2324cb79;
    ram_cell[    2481] = 32'he16ef9b1;
    ram_cell[    2482] = 32'h22c94acf;
    ram_cell[    2483] = 32'h917879f6;
    ram_cell[    2484] = 32'hd193312b;
    ram_cell[    2485] = 32'hcfa564d5;
    ram_cell[    2486] = 32'h1580a88b;
    ram_cell[    2487] = 32'hc0246681;
    ram_cell[    2488] = 32'h1c68c141;
    ram_cell[    2489] = 32'h06d8ccad;
    ram_cell[    2490] = 32'h23db6dec;
    ram_cell[    2491] = 32'hb307e84f;
    ram_cell[    2492] = 32'h8deee2b7;
    ram_cell[    2493] = 32'h842d15fe;
    ram_cell[    2494] = 32'hf3f1171b;
    ram_cell[    2495] = 32'h01436c1b;
    ram_cell[    2496] = 32'h89b57d46;
    ram_cell[    2497] = 32'h50527819;
    ram_cell[    2498] = 32'hf15e24b1;
    ram_cell[    2499] = 32'h661b7cfb;
    ram_cell[    2500] = 32'he728668e;
    ram_cell[    2501] = 32'h9ae7f287;
    ram_cell[    2502] = 32'hc18273cf;
    ram_cell[    2503] = 32'h1fdcc377;
    ram_cell[    2504] = 32'h6a9c5dae;
    ram_cell[    2505] = 32'h838e89d9;
    ram_cell[    2506] = 32'h45d56f96;
    ram_cell[    2507] = 32'ha429cd0f;
    ram_cell[    2508] = 32'he8b817c3;
    ram_cell[    2509] = 32'hb82298ff;
    ram_cell[    2510] = 32'h98fa31ca;
    ram_cell[    2511] = 32'h546fda20;
    ram_cell[    2512] = 32'had47aebb;
    ram_cell[    2513] = 32'h41fae862;
    ram_cell[    2514] = 32'he93cd3f3;
    ram_cell[    2515] = 32'h3bbf3e2d;
    ram_cell[    2516] = 32'h2bf9d068;
    ram_cell[    2517] = 32'h63b8ed61;
    ram_cell[    2518] = 32'h7579328d;
    ram_cell[    2519] = 32'hbd986077;
    ram_cell[    2520] = 32'h9c39bfcf;
    ram_cell[    2521] = 32'h7cabf587;
    ram_cell[    2522] = 32'ha0be5326;
    ram_cell[    2523] = 32'hbbec1594;
    ram_cell[    2524] = 32'h49dc853a;
    ram_cell[    2525] = 32'h081ffe6d;
    ram_cell[    2526] = 32'he9151203;
    ram_cell[    2527] = 32'hdd877954;
    ram_cell[    2528] = 32'h01d9e0d7;
    ram_cell[    2529] = 32'h8d07438c;
    ram_cell[    2530] = 32'h785c2160;
    ram_cell[    2531] = 32'h85873711;
    ram_cell[    2532] = 32'ha91bae94;
    ram_cell[    2533] = 32'h7463dd3a;
    ram_cell[    2534] = 32'ha73aaba1;
    ram_cell[    2535] = 32'hc4873246;
    ram_cell[    2536] = 32'hf6437857;
    ram_cell[    2537] = 32'hb91ff865;
    ram_cell[    2538] = 32'hc8a1dbc2;
    ram_cell[    2539] = 32'hf6816595;
    ram_cell[    2540] = 32'h642cdb38;
    ram_cell[    2541] = 32'h9af10106;
    ram_cell[    2542] = 32'hf3894670;
    ram_cell[    2543] = 32'hb65981e0;
    ram_cell[    2544] = 32'ha28bc92e;
    ram_cell[    2545] = 32'h1aa67671;
    ram_cell[    2546] = 32'h3ad86ec5;
    ram_cell[    2547] = 32'h3b0a571c;
    ram_cell[    2548] = 32'h02985b5e;
    ram_cell[    2549] = 32'he2796233;
    ram_cell[    2550] = 32'h15e5c538;
    ram_cell[    2551] = 32'h04cb1c46;
    ram_cell[    2552] = 32'h25913a39;
    ram_cell[    2553] = 32'h3b1338fa;
    ram_cell[    2554] = 32'ha6f87b3c;
    ram_cell[    2555] = 32'hf72af81c;
    ram_cell[    2556] = 32'h44ee1578;
    ram_cell[    2557] = 32'h557eae3c;
    ram_cell[    2558] = 32'h9b5191d9;
    ram_cell[    2559] = 32'hed525d51;
    ram_cell[    2560] = 32'hdd5fcdcd;
    ram_cell[    2561] = 32'h936ce66b;
    ram_cell[    2562] = 32'hc877a73b;
    ram_cell[    2563] = 32'h9ac3eb3e;
    ram_cell[    2564] = 32'hf75ced6c;
    ram_cell[    2565] = 32'hf15747e7;
    ram_cell[    2566] = 32'hbb2e8d93;
    ram_cell[    2567] = 32'h12be51e0;
    ram_cell[    2568] = 32'h237d8800;
    ram_cell[    2569] = 32'hd277a470;
    ram_cell[    2570] = 32'h706c7447;
    ram_cell[    2571] = 32'h478ee480;
    ram_cell[    2572] = 32'hc91bac38;
    ram_cell[    2573] = 32'h890b41b0;
    ram_cell[    2574] = 32'h86bd25c4;
    ram_cell[    2575] = 32'h94a339bc;
    ram_cell[    2576] = 32'h459c7897;
    ram_cell[    2577] = 32'h26aa303b;
    ram_cell[    2578] = 32'hc0206db9;
    ram_cell[    2579] = 32'hd2915a2e;
    ram_cell[    2580] = 32'h43aed1d9;
    ram_cell[    2581] = 32'h66ff7d49;
    ram_cell[    2582] = 32'hef6ca195;
    ram_cell[    2583] = 32'heee5eebd;
    ram_cell[    2584] = 32'h2bdccde4;
    ram_cell[    2585] = 32'hef1d445e;
    ram_cell[    2586] = 32'h6f1eb2ce;
    ram_cell[    2587] = 32'h711c2d78;
    ram_cell[    2588] = 32'h722377cf;
    ram_cell[    2589] = 32'hba5cf5c8;
    ram_cell[    2590] = 32'hd70b24ec;
    ram_cell[    2591] = 32'hdebfb50c;
    ram_cell[    2592] = 32'h44049084;
    ram_cell[    2593] = 32'h3451f480;
    ram_cell[    2594] = 32'hbc061e46;
    ram_cell[    2595] = 32'h17e054ee;
    ram_cell[    2596] = 32'hec641a67;
    ram_cell[    2597] = 32'h85f6128e;
    ram_cell[    2598] = 32'h0f0f977d;
    ram_cell[    2599] = 32'h4042beb7;
    ram_cell[    2600] = 32'hcef22cd2;
    ram_cell[    2601] = 32'h6f590916;
    ram_cell[    2602] = 32'h28de9fbe;
    ram_cell[    2603] = 32'h1431bf5b;
    ram_cell[    2604] = 32'haeb786d9;
    ram_cell[    2605] = 32'hcdad40cb;
    ram_cell[    2606] = 32'h0fd6aaf7;
    ram_cell[    2607] = 32'h2518f762;
    ram_cell[    2608] = 32'hd5d7580f;
    ram_cell[    2609] = 32'hbc0b8671;
    ram_cell[    2610] = 32'h2913dd59;
    ram_cell[    2611] = 32'he330df77;
    ram_cell[    2612] = 32'h73d8585f;
    ram_cell[    2613] = 32'h9d25f376;
    ram_cell[    2614] = 32'h7326af6a;
    ram_cell[    2615] = 32'h72ee9a19;
    ram_cell[    2616] = 32'h7e41efa8;
    ram_cell[    2617] = 32'h67509661;
    ram_cell[    2618] = 32'h790b572e;
    ram_cell[    2619] = 32'h5c330ffa;
    ram_cell[    2620] = 32'h0325467c;
    ram_cell[    2621] = 32'h22d0fc9d;
    ram_cell[    2622] = 32'haea41885;
    ram_cell[    2623] = 32'h7509d488;
    ram_cell[    2624] = 32'hcdfc2960;
    ram_cell[    2625] = 32'hd898f253;
    ram_cell[    2626] = 32'hf82c67b3;
    ram_cell[    2627] = 32'h19617e98;
    ram_cell[    2628] = 32'h0cdf50cb;
    ram_cell[    2629] = 32'h675fbefb;
    ram_cell[    2630] = 32'hbf54a7c4;
    ram_cell[    2631] = 32'hb532c609;
    ram_cell[    2632] = 32'h850af88e;
    ram_cell[    2633] = 32'haec4d345;
    ram_cell[    2634] = 32'h1e311e5f;
    ram_cell[    2635] = 32'h6a1b3689;
    ram_cell[    2636] = 32'heffd3693;
    ram_cell[    2637] = 32'ha47c2402;
    ram_cell[    2638] = 32'h13966642;
    ram_cell[    2639] = 32'h97390a97;
    ram_cell[    2640] = 32'hadeb7acf;
    ram_cell[    2641] = 32'h873b3597;
    ram_cell[    2642] = 32'hcd0748c0;
    ram_cell[    2643] = 32'h5a7c12eb;
    ram_cell[    2644] = 32'h6fbf0c0a;
    ram_cell[    2645] = 32'h22c37c98;
    ram_cell[    2646] = 32'h342c840b;
    ram_cell[    2647] = 32'h35a86d9f;
    ram_cell[    2648] = 32'h6695254e;
    ram_cell[    2649] = 32'h72e47cfd;
    ram_cell[    2650] = 32'h307e9b21;
    ram_cell[    2651] = 32'hd3f452c6;
    ram_cell[    2652] = 32'hc0182680;
    ram_cell[    2653] = 32'h127b8818;
    ram_cell[    2654] = 32'h41e47f5d;
    ram_cell[    2655] = 32'h6e37d648;
    ram_cell[    2656] = 32'h3f80c1b4;
    ram_cell[    2657] = 32'h4ada63a2;
    ram_cell[    2658] = 32'h8ec0209c;
    ram_cell[    2659] = 32'ha4014f8e;
    ram_cell[    2660] = 32'h72809eb4;
    ram_cell[    2661] = 32'h4f6b0b1d;
    ram_cell[    2662] = 32'hd6240934;
    ram_cell[    2663] = 32'hf08c4a3f;
    ram_cell[    2664] = 32'hcd45de8d;
    ram_cell[    2665] = 32'h5a30708c;
    ram_cell[    2666] = 32'hd60f8287;
    ram_cell[    2667] = 32'hf4b84e43;
    ram_cell[    2668] = 32'h35d2b5f8;
    ram_cell[    2669] = 32'ha0ff932c;
    ram_cell[    2670] = 32'h7f87bbb7;
    ram_cell[    2671] = 32'h04305fc4;
    ram_cell[    2672] = 32'haf649016;
    ram_cell[    2673] = 32'h82a44b43;
    ram_cell[    2674] = 32'h53425468;
    ram_cell[    2675] = 32'h7d79b318;
    ram_cell[    2676] = 32'h39ab516f;
    ram_cell[    2677] = 32'he080efcf;
    ram_cell[    2678] = 32'h51f7d8a9;
    ram_cell[    2679] = 32'h3170cd34;
    ram_cell[    2680] = 32'ha942f4b7;
    ram_cell[    2681] = 32'h1e0b10d1;
    ram_cell[    2682] = 32'had57d724;
    ram_cell[    2683] = 32'hcec54ab7;
    ram_cell[    2684] = 32'h6345d836;
    ram_cell[    2685] = 32'h675ca1d5;
    ram_cell[    2686] = 32'he66f13c3;
    ram_cell[    2687] = 32'h50d88efb;
    ram_cell[    2688] = 32'haa0b735b;
    ram_cell[    2689] = 32'hd4dbca44;
    ram_cell[    2690] = 32'ha1b1dd78;
    ram_cell[    2691] = 32'h4896848f;
    ram_cell[    2692] = 32'hdf12fad4;
    ram_cell[    2693] = 32'hefd4a6bc;
    ram_cell[    2694] = 32'h14315829;
    ram_cell[    2695] = 32'h20e2dbeb;
    ram_cell[    2696] = 32'h7bce467d;
    ram_cell[    2697] = 32'he8ecea63;
    ram_cell[    2698] = 32'hb40e8cba;
    ram_cell[    2699] = 32'h0070f29d;
    ram_cell[    2700] = 32'hec78df7a;
    ram_cell[    2701] = 32'habab234e;
    ram_cell[    2702] = 32'h64d3fae4;
    ram_cell[    2703] = 32'h7f98d20a;
    ram_cell[    2704] = 32'hecad073f;
    ram_cell[    2705] = 32'h4e32a7c0;
    ram_cell[    2706] = 32'h7dcd164d;
    ram_cell[    2707] = 32'h78810afa;
    ram_cell[    2708] = 32'h0e516f8c;
    ram_cell[    2709] = 32'h28a335a5;
    ram_cell[    2710] = 32'hebabc19d;
    ram_cell[    2711] = 32'hcd21caee;
    ram_cell[    2712] = 32'h176f1490;
    ram_cell[    2713] = 32'hc34cfee8;
    ram_cell[    2714] = 32'hec00ce1c;
    ram_cell[    2715] = 32'hffcb0ecd;
    ram_cell[    2716] = 32'hb2ea9ce0;
    ram_cell[    2717] = 32'h3a1c1e01;
    ram_cell[    2718] = 32'h86b3f08a;
    ram_cell[    2719] = 32'h8b92ad01;
    ram_cell[    2720] = 32'hf6e6089c;
    ram_cell[    2721] = 32'hc049a584;
    ram_cell[    2722] = 32'h09353634;
    ram_cell[    2723] = 32'hd68f3645;
    ram_cell[    2724] = 32'hc396c9ac;
    ram_cell[    2725] = 32'h35e5377e;
    ram_cell[    2726] = 32'heeae7560;
    ram_cell[    2727] = 32'h3d03de6a;
    ram_cell[    2728] = 32'ha89dad4a;
    ram_cell[    2729] = 32'h838cb38b;
    ram_cell[    2730] = 32'h2617184d;
    ram_cell[    2731] = 32'h2f93bf4f;
    ram_cell[    2732] = 32'h73617946;
    ram_cell[    2733] = 32'hfcc3ce1b;
    ram_cell[    2734] = 32'h6c94327c;
    ram_cell[    2735] = 32'h113a8de9;
    ram_cell[    2736] = 32'h2e09c340;
    ram_cell[    2737] = 32'h2fbbfe1d;
    ram_cell[    2738] = 32'h22368b42;
    ram_cell[    2739] = 32'hdc75199c;
    ram_cell[    2740] = 32'h3c5564e7;
    ram_cell[    2741] = 32'hc244f122;
    ram_cell[    2742] = 32'h9ccb403b;
    ram_cell[    2743] = 32'h9ecb212a;
    ram_cell[    2744] = 32'h450374e3;
    ram_cell[    2745] = 32'he756aa9e;
    ram_cell[    2746] = 32'h6236aa88;
    ram_cell[    2747] = 32'h9a3e414a;
    ram_cell[    2748] = 32'hce66458c;
    ram_cell[    2749] = 32'h9cd7dcda;
    ram_cell[    2750] = 32'hab7faefa;
    ram_cell[    2751] = 32'h63ea0283;
    ram_cell[    2752] = 32'hef84e5e0;
    ram_cell[    2753] = 32'h3f749475;
    ram_cell[    2754] = 32'h1d3cc146;
    ram_cell[    2755] = 32'h8e7a9d39;
    ram_cell[    2756] = 32'h4348a2c0;
    ram_cell[    2757] = 32'he7e63026;
    ram_cell[    2758] = 32'h29e99c0a;
    ram_cell[    2759] = 32'hd8951717;
    ram_cell[    2760] = 32'he5287fd5;
    ram_cell[    2761] = 32'h7472443e;
    ram_cell[    2762] = 32'h6facf595;
    ram_cell[    2763] = 32'hc3eb88fb;
    ram_cell[    2764] = 32'h60b1afa5;
    ram_cell[    2765] = 32'h96e77a9a;
    ram_cell[    2766] = 32'h87eaba0b;
    ram_cell[    2767] = 32'h6224b651;
    ram_cell[    2768] = 32'h0cfae662;
    ram_cell[    2769] = 32'hce47f976;
    ram_cell[    2770] = 32'h9573fc31;
    ram_cell[    2771] = 32'h7541b26e;
    ram_cell[    2772] = 32'hef0eaf69;
    ram_cell[    2773] = 32'hd8e66634;
    ram_cell[    2774] = 32'he88627d5;
    ram_cell[    2775] = 32'hcd4c265a;
    ram_cell[    2776] = 32'h7174f337;
    ram_cell[    2777] = 32'haec6b622;
    ram_cell[    2778] = 32'h0f88aa5a;
    ram_cell[    2779] = 32'h762fb806;
    ram_cell[    2780] = 32'hfd0e9a76;
    ram_cell[    2781] = 32'hb956b480;
    ram_cell[    2782] = 32'hd8fe18c4;
    ram_cell[    2783] = 32'h3a63b3c9;
    ram_cell[    2784] = 32'h74cff772;
    ram_cell[    2785] = 32'h7cac39d8;
    ram_cell[    2786] = 32'hf3d1de82;
    ram_cell[    2787] = 32'h81b6d621;
    ram_cell[    2788] = 32'h66ca12d7;
    ram_cell[    2789] = 32'ha75059b9;
    ram_cell[    2790] = 32'he0e316ff;
    ram_cell[    2791] = 32'h519ecf90;
    ram_cell[    2792] = 32'hf7fe7fdf;
    ram_cell[    2793] = 32'h73745485;
    ram_cell[    2794] = 32'ha659c039;
    ram_cell[    2795] = 32'hd9ff883f;
    ram_cell[    2796] = 32'h433b0642;
    ram_cell[    2797] = 32'h57915072;
    ram_cell[    2798] = 32'h8a433116;
    ram_cell[    2799] = 32'h7dfa2469;
    ram_cell[    2800] = 32'hc2031e1f;
    ram_cell[    2801] = 32'ha6fdf316;
    ram_cell[    2802] = 32'h83755814;
    ram_cell[    2803] = 32'hdcef52a7;
    ram_cell[    2804] = 32'h2e6f0502;
    ram_cell[    2805] = 32'hbebfec45;
    ram_cell[    2806] = 32'hf06f8c47;
    ram_cell[    2807] = 32'h6983aa70;
    ram_cell[    2808] = 32'hea355fef;
    ram_cell[    2809] = 32'h8b30a314;
    ram_cell[    2810] = 32'h6c49c285;
    ram_cell[    2811] = 32'h1d9b1ead;
    ram_cell[    2812] = 32'hd6b740ed;
    ram_cell[    2813] = 32'h72cb81d5;
    ram_cell[    2814] = 32'h0ad863f6;
    ram_cell[    2815] = 32'h75295d76;
    ram_cell[    2816] = 32'hcb75fdd3;
    ram_cell[    2817] = 32'h5734bef9;
    ram_cell[    2818] = 32'ha3d0f9a6;
    ram_cell[    2819] = 32'hfe0317d6;
    ram_cell[    2820] = 32'h1ab4eb7c;
    ram_cell[    2821] = 32'h9a03c2cd;
    ram_cell[    2822] = 32'h57f08050;
    ram_cell[    2823] = 32'h20ce67d5;
    ram_cell[    2824] = 32'h504b03f2;
    ram_cell[    2825] = 32'h920ee571;
    ram_cell[    2826] = 32'hd8eb2f05;
    ram_cell[    2827] = 32'he4f1ade0;
    ram_cell[    2828] = 32'h3bed4a46;
    ram_cell[    2829] = 32'h62edf8e2;
    ram_cell[    2830] = 32'h425a7313;
    ram_cell[    2831] = 32'hf3222c8f;
    ram_cell[    2832] = 32'hfcb28d3a;
    ram_cell[    2833] = 32'h90f3450e;
    ram_cell[    2834] = 32'he49b6e4c;
    ram_cell[    2835] = 32'he614fd63;
    ram_cell[    2836] = 32'h71dff7b3;
    ram_cell[    2837] = 32'h199ae819;
    ram_cell[    2838] = 32'h6768f73e;
    ram_cell[    2839] = 32'h4cdb4968;
    ram_cell[    2840] = 32'h8c21bebc;
    ram_cell[    2841] = 32'h98fecd62;
    ram_cell[    2842] = 32'h9ff4b023;
    ram_cell[    2843] = 32'he0973dec;
    ram_cell[    2844] = 32'hb84d4ccb;
    ram_cell[    2845] = 32'h13769a14;
    ram_cell[    2846] = 32'he6abac12;
    ram_cell[    2847] = 32'h1dd9f603;
    ram_cell[    2848] = 32'h18cd7143;
    ram_cell[    2849] = 32'h9f3d9d93;
    ram_cell[    2850] = 32'h393e8f60;
    ram_cell[    2851] = 32'h221779e8;
    ram_cell[    2852] = 32'h7bd9da0f;
    ram_cell[    2853] = 32'h6b19ba16;
    ram_cell[    2854] = 32'h427d9afa;
    ram_cell[    2855] = 32'h6ee324ba;
    ram_cell[    2856] = 32'ha562da4b;
    ram_cell[    2857] = 32'h262c8f21;
    ram_cell[    2858] = 32'hafac13fc;
    ram_cell[    2859] = 32'h85366726;
    ram_cell[    2860] = 32'h4bb22591;
    ram_cell[    2861] = 32'h3d4e89f7;
    ram_cell[    2862] = 32'hc4abb86f;
    ram_cell[    2863] = 32'h09c3252e;
    ram_cell[    2864] = 32'h534ea556;
    ram_cell[    2865] = 32'h9e5d1ece;
    ram_cell[    2866] = 32'hfc7e1f14;
    ram_cell[    2867] = 32'h9feec6df;
    ram_cell[    2868] = 32'hd00f67ec;
    ram_cell[    2869] = 32'hbeb6ff9d;
    ram_cell[    2870] = 32'hd722d2c5;
    ram_cell[    2871] = 32'h969d63d2;
    ram_cell[    2872] = 32'h8aa6f01c;
    ram_cell[    2873] = 32'h40834941;
    ram_cell[    2874] = 32'h114d4163;
    ram_cell[    2875] = 32'h35e04a0a;
    ram_cell[    2876] = 32'h2c877dfb;
    ram_cell[    2877] = 32'h46fcf2da;
    ram_cell[    2878] = 32'hb1acb393;
    ram_cell[    2879] = 32'h3fd0b92b;
    ram_cell[    2880] = 32'h115987c2;
    ram_cell[    2881] = 32'hf75bfa00;
    ram_cell[    2882] = 32'h33c1277e;
    ram_cell[    2883] = 32'h5a1d2c66;
    ram_cell[    2884] = 32'h0b09b92f;
    ram_cell[    2885] = 32'ha6994bc8;
    ram_cell[    2886] = 32'h01c2ebc1;
    ram_cell[    2887] = 32'hfab00615;
    ram_cell[    2888] = 32'h6d889d18;
    ram_cell[    2889] = 32'h6d3b0fec;
    ram_cell[    2890] = 32'he74d39a1;
    ram_cell[    2891] = 32'h49fde469;
    ram_cell[    2892] = 32'h0797026e;
    ram_cell[    2893] = 32'hb1bf7085;
    ram_cell[    2894] = 32'h1ab287eb;
    ram_cell[    2895] = 32'ha0b38ed1;
    ram_cell[    2896] = 32'h5d40a6f8;
    ram_cell[    2897] = 32'ha187aa55;
    ram_cell[    2898] = 32'hd461c9c7;
    ram_cell[    2899] = 32'h21692ed5;
    ram_cell[    2900] = 32'hbfe98d9e;
    ram_cell[    2901] = 32'h3d075c85;
    ram_cell[    2902] = 32'ha0e90401;
    ram_cell[    2903] = 32'h15eb26f3;
    ram_cell[    2904] = 32'h50043395;
    ram_cell[    2905] = 32'h84d4846a;
    ram_cell[    2906] = 32'hfb9e7d3f;
    ram_cell[    2907] = 32'he2fcc8b5;
    ram_cell[    2908] = 32'ha855429c;
    ram_cell[    2909] = 32'h08a94c48;
    ram_cell[    2910] = 32'hfeb87fe5;
    ram_cell[    2911] = 32'h2d73ee8c;
    ram_cell[    2912] = 32'h92e94db4;
    ram_cell[    2913] = 32'h58e099e6;
    ram_cell[    2914] = 32'h730e72a3;
    ram_cell[    2915] = 32'h57441960;
    ram_cell[    2916] = 32'hd3fdafc0;
    ram_cell[    2917] = 32'h4f39c011;
    ram_cell[    2918] = 32'h918aef26;
    ram_cell[    2919] = 32'h348507f4;
    ram_cell[    2920] = 32'hde350834;
    ram_cell[    2921] = 32'h428c897a;
    ram_cell[    2922] = 32'he5664676;
    ram_cell[    2923] = 32'he2f1ed8a;
    ram_cell[    2924] = 32'h25b46899;
    ram_cell[    2925] = 32'habc93d36;
    ram_cell[    2926] = 32'h91b67f41;
    ram_cell[    2927] = 32'hcaa6b13a;
    ram_cell[    2928] = 32'h072aa9c7;
    ram_cell[    2929] = 32'h9f978783;
    ram_cell[    2930] = 32'he2fecf4a;
    ram_cell[    2931] = 32'he3b367b6;
    ram_cell[    2932] = 32'h089fb0a7;
    ram_cell[    2933] = 32'h5af01733;
    ram_cell[    2934] = 32'hbfa1038f;
    ram_cell[    2935] = 32'hced5ecd2;
    ram_cell[    2936] = 32'hf95191e6;
    ram_cell[    2937] = 32'h1dc4cdc6;
    ram_cell[    2938] = 32'h9d5665fe;
    ram_cell[    2939] = 32'hfa85692d;
    ram_cell[    2940] = 32'h36198d37;
    ram_cell[    2941] = 32'ha69c87e7;
    ram_cell[    2942] = 32'h718cca03;
    ram_cell[    2943] = 32'h794c06e0;
    ram_cell[    2944] = 32'h6c4d9588;
    ram_cell[    2945] = 32'hade32976;
    ram_cell[    2946] = 32'h3e6bb722;
    ram_cell[    2947] = 32'ha53d8842;
    ram_cell[    2948] = 32'hda2b0338;
    ram_cell[    2949] = 32'h835bd647;
    ram_cell[    2950] = 32'h9c8752b0;
    ram_cell[    2951] = 32'h9c6d73bc;
    ram_cell[    2952] = 32'hfe81c612;
    ram_cell[    2953] = 32'ha08fb5e0;
    ram_cell[    2954] = 32'h8daf5999;
    ram_cell[    2955] = 32'h83292bc8;
    ram_cell[    2956] = 32'h4c24538b;
    ram_cell[    2957] = 32'h3cd222a2;
    ram_cell[    2958] = 32'h6274d277;
    ram_cell[    2959] = 32'hc6c41b25;
    ram_cell[    2960] = 32'hcf529a17;
    ram_cell[    2961] = 32'hfcd8cdf5;
    ram_cell[    2962] = 32'he1e46d97;
    ram_cell[    2963] = 32'h0d149d90;
    ram_cell[    2964] = 32'hcb128f70;
    ram_cell[    2965] = 32'h9f647d0c;
    ram_cell[    2966] = 32'h50aff31e;
    ram_cell[    2967] = 32'hf6242d05;
    ram_cell[    2968] = 32'he073f956;
    ram_cell[    2969] = 32'h33ba6fa4;
    ram_cell[    2970] = 32'h98203912;
    ram_cell[    2971] = 32'h267c1be4;
    ram_cell[    2972] = 32'h5ad4d3df;
    ram_cell[    2973] = 32'hccc5be02;
    ram_cell[    2974] = 32'h8937897b;
    ram_cell[    2975] = 32'h791c0728;
    ram_cell[    2976] = 32'hbff59146;
    ram_cell[    2977] = 32'h45b7405b;
    ram_cell[    2978] = 32'h816312c6;
    ram_cell[    2979] = 32'h870061ee;
    ram_cell[    2980] = 32'h8b98fe7a;
    ram_cell[    2981] = 32'h8129b54f;
    ram_cell[    2982] = 32'h084105bb;
    ram_cell[    2983] = 32'h13dc8b80;
    ram_cell[    2984] = 32'hf6ec9dfc;
    ram_cell[    2985] = 32'hfeec56a9;
    ram_cell[    2986] = 32'ha76272d8;
    ram_cell[    2987] = 32'h46a0ba3e;
    ram_cell[    2988] = 32'hf4b589c2;
    ram_cell[    2989] = 32'heec8fe08;
    ram_cell[    2990] = 32'habaf5d29;
    ram_cell[    2991] = 32'h56b5646b;
    ram_cell[    2992] = 32'h0302d201;
    ram_cell[    2993] = 32'hc79ff968;
    ram_cell[    2994] = 32'h32cda979;
    ram_cell[    2995] = 32'hfa09908a;
    ram_cell[    2996] = 32'h956668fa;
    ram_cell[    2997] = 32'hdc494680;
    ram_cell[    2998] = 32'hef0c12fa;
    ram_cell[    2999] = 32'h47543a1e;
    ram_cell[    3000] = 32'h771a4e68;
    ram_cell[    3001] = 32'hd34ed513;
    ram_cell[    3002] = 32'hea3d64de;
    ram_cell[    3003] = 32'h665d7405;
    ram_cell[    3004] = 32'hc250a4f7;
    ram_cell[    3005] = 32'h282bd0da;
    ram_cell[    3006] = 32'h6c1b3d3f;
    ram_cell[    3007] = 32'h1e4c10d7;
    ram_cell[    3008] = 32'hc680a297;
    ram_cell[    3009] = 32'hdd1dba9d;
    ram_cell[    3010] = 32'h6ea27c33;
    ram_cell[    3011] = 32'h53c52751;
    ram_cell[    3012] = 32'hd76456f3;
    ram_cell[    3013] = 32'h432c7729;
    ram_cell[    3014] = 32'h8fdfb8fb;
    ram_cell[    3015] = 32'h55126073;
    ram_cell[    3016] = 32'hcd278a69;
    ram_cell[    3017] = 32'hf8e50c4d;
    ram_cell[    3018] = 32'hc0d5902e;
    ram_cell[    3019] = 32'hef1c13ca;
    ram_cell[    3020] = 32'h421ccad1;
    ram_cell[    3021] = 32'h0a716b02;
    ram_cell[    3022] = 32'hb4eaff9b;
    ram_cell[    3023] = 32'h620db296;
    ram_cell[    3024] = 32'hb299a977;
    ram_cell[    3025] = 32'h86927ae3;
    ram_cell[    3026] = 32'h0e003938;
    ram_cell[    3027] = 32'h95c8c15f;
    ram_cell[    3028] = 32'hb0035931;
    ram_cell[    3029] = 32'h80c8c9c1;
    ram_cell[    3030] = 32'h2b04b013;
    ram_cell[    3031] = 32'hf563e93f;
    ram_cell[    3032] = 32'h98cbc98c;
    ram_cell[    3033] = 32'h7b7879d1;
    ram_cell[    3034] = 32'he88ae51f;
    ram_cell[    3035] = 32'h873a1539;
    ram_cell[    3036] = 32'hcc02036e;
    ram_cell[    3037] = 32'h01eb6776;
    ram_cell[    3038] = 32'h8fe5f1de;
    ram_cell[    3039] = 32'h9615a1b2;
    ram_cell[    3040] = 32'h95c11d05;
    ram_cell[    3041] = 32'h50ab9d0e;
    ram_cell[    3042] = 32'hd6096fa8;
    ram_cell[    3043] = 32'h618e9140;
    ram_cell[    3044] = 32'ha6a54788;
    ram_cell[    3045] = 32'ha494fee1;
    ram_cell[    3046] = 32'h1a21b33f;
    ram_cell[    3047] = 32'h4025915b;
    ram_cell[    3048] = 32'h24d777b1;
    ram_cell[    3049] = 32'hcb7d1a86;
    ram_cell[    3050] = 32'h1a67a190;
    ram_cell[    3051] = 32'h192f5a08;
    ram_cell[    3052] = 32'h35d3fcb0;
    ram_cell[    3053] = 32'hac59478b;
    ram_cell[    3054] = 32'h1559d145;
    ram_cell[    3055] = 32'h50699f09;
    ram_cell[    3056] = 32'hfa8930fb;
    ram_cell[    3057] = 32'h401fc9b4;
    ram_cell[    3058] = 32'ha7735fdf;
    ram_cell[    3059] = 32'h3e5d591f;
    ram_cell[    3060] = 32'h7f7f9b8e;
    ram_cell[    3061] = 32'h5bcce02e;
    ram_cell[    3062] = 32'h82bd1d85;
    ram_cell[    3063] = 32'he7a7af85;
    ram_cell[    3064] = 32'h189d8168;
    ram_cell[    3065] = 32'ha7f66bc1;
    ram_cell[    3066] = 32'hcc266875;
    ram_cell[    3067] = 32'hb2ce006f;
    ram_cell[    3068] = 32'h1fa640f6;
    ram_cell[    3069] = 32'hfdadcc24;
    ram_cell[    3070] = 32'hcd6fff35;
    ram_cell[    3071] = 32'hfcf26c46;
end

endmodule

