`timescale 1ns/100ps
//correct read result:
// 00000042 0000161a 0000142c 00000c3c 00000c86 000004fb 00001064 00000f20 000001a3 000004ef 000019eb 0000086f 00001f14 00001b9b 00000e73 00000e13 00000c17 00001570 0000011e 00000512 00000b8a 000008b8 00000858 000004d1 00001082 0000156c 00000665 00000979 000019d3 00000967 0000127b 00001f06 00001f25 00001766 00000c2a 000010f4 0000078a 00000ae5 000016db 0000131c 000010db 0000127e 000017d8 000011c7 00001219 00000ede 00001842 00001c84 0000107a 00001474 0000197f 00000f15 00000cf0 00001e4e 00001b60 00000107 00001449 00001147 00000997 00000008 000012de 00001e74 00000f07 000005a1 0000069f 00000d73 00001cab 00001002 0000140c 00001e3d 000011eb 00001126 00001d92 000019bc 00001a2e 00000b99 00001a60 000018eb 0000179d 00001969 00000ce7 000000a3 00001724 00000453 00001d70 00000315 00000cd9 00001516 000006ae 000007c2 00000618 00000ac7 0000062f 00000600 000016d9 00001881 00000a68 0000187f 00000902 0000143d 00001590 00000746 00000616 00001220 00001783 000018e4 000017e0 0000050f 000007bc 00000f69 00000ae3 0000023d 000009ec 00000e08 00000cdb 00001dd3 00001eac 00001aa8 00001088 00001aca 000001d1 000011f3 000004eb 0000180b 00000dd4 00000760 00001f2e 000007d7 00000176 000004a1 0000185e 00000326 00000e3b 00000551 00000de0 000017cd 000009b8 00000f51 00000bc1 00001632 00000579 00001b0f 0000134c 00001d37 00000243 00001631 000019e8 000018cc 00000bc1 00001352 00000c51 00000e23 0000118f 0000009c 00000070 00000d92 00001629 000002bc 00001777 00001098 00001da0 00001326 00000de2 0000066a 00001648 00000405 00000325 00000fb7 00000ac4 0000107f 00000261 00000e39 000001f8 00001884 00000261 00000aa4 00000e4a 00000ef3 00000902 00000885 00000fde 00001f2c 00001035 000004d5 0000140c 00000dc8 000015e4 00001350 000009c0 000011a4 00000d91 00001ab1 000007a0 0000188e 000008f9 00000aff 0000019b 00000c12 00001aa0 00000fd7 00000327 00001cf3 000017f8 00001e03 000012e7 000009d0 00000654 000000fe 000010d0 00001e0f 00001c18 00000000 00001b42 00001b70 0000016d 000013d4 00000462 00000872 00001d6f 00000c0a 00000cb6 000019a4 00001aa0 00000f7b 00000ca4 00000eaa 000010aa 000007c1 00001c15 000012fb 00000212 00000238 00000c98 00001a43 000009ef 0000023d 000008d8 00001216 00001924 0000137d 00001b29 00000279 00000462 00001b38 00000041 00001247 00000e78 00001689 00000578 000019aa 00000488 00000f56 000002c5 00001902 0000013a 00000fe8 00001ccb 00001c2a 000017d3 0000170f 000004ab 00000c48 000003b3 000019ce 00001ebf 00000f8d 00001f0d 000014f8 00001bfe 000015cb 00001abd 0000145f 00001502 00000a55 00001095 0000058f 00000096 00000eb3 000015ff 00001be4 0000136d 000015e8 0000014e 00000656 00000e71 0000159e 00000f1c 00001be4 0000172a 00001d12 00000de2 0000055d 00001285 0000075e 00000e25 000010a4 00000541 00000635 00001b11 00000dad 00001d05 00000cff 00000dfc 0000063c 00000f02 00000416 0000193a 00001b6b 00001ce1 000013b0 00000bc3 00001aa7 00001847 00001dbb 00000769 00001c24 000017d3 000008f6 00000662 0000039b 0000042a 000007f6 000004dd 00001173 00000020 00001b15 000000e4 00001a7a 00000d53 0000144a 000017c3 0000173c 000008bc 00000c2e 00001377 00001169 00001092 00000a68 00000510 00001838 000013f7 00001bd2 00001b43 0000124f 0000016f 0000104e 000002c0 00000db7 00001e3e 00001a77 00000e41 00001581 00000246 00001053 00000b0f 00000cc4 00000ad5 00001783 000009c9 00000ab0 00000964 00000c53 000017a9 00000ee6 0000103a 000016c6 00001979 00001e01 000011f5 00000d8f 000010ff 00000f53 0000146e 00000ee4 00000009 0000149c 00000682 000007c9 00000115 00000609 00001b14 000005d3 00000692 000002e6 000005e8 0000194a 000010e3 0000039b 00001cc8 00001c8b 00000591 00000765 00000dda 000002cf 00001227 00000b94 00001861 00000cce 0000057b 0000110e 000008c8 00001278 00000d4b 000007c8 000000d2 000001ec 00001d2a 00001957 00001510 000009f6 000019c8 0000125e 000004a8 00000eba 000015dc 00000c42 0000111d 00000e2b 0000153d 00000b0d 00001c73 000012cf 000007ac 00001d43 00001595 00000d29 00001979 000013fe 00001119 00001ad3 00000472 000016fe 00001783 00001bd3 000004df 00001507 00000266 000002dd 00000afc 00000dfc 00000e5c 000018e0 00001609 00001c28 00000afd 0000154e 00001146 00001d89 00001dbd 00001177 00000b7c 000011e9 0000190e 00001cd2 0000022c 00000dfe 000010ad 00000509 00001bf3 0000146e 00001e69 00001cf5 00001d52 000002ad 000001a2 000001a7 0000132d 00001dd4 00000ea4 00001188 00001820 0000101a 000007ef 00001646 00001aa1 0000158b 0000185e 000006c5 000013d7 00001a48 00000d39 000000b1 000006a9 00000ac5 00000877 00000532 00001d5d 000012a9 00001020 00000d22 00000934 00000171 000003fc 00001c31 00001154 00001c9a 000003a5 00001dbd 00001065 00001f27 000003bf 0000072b 0000062c 00000f80 0000156b 00001d2d 000001c4 00000785 00000133 0000095d 000000f3 00001327 00000d56 00000cad 000015f5 00000256 000004cc 00000e5b 000019be 00000320 000011ae 000003cf 000017cd 00000ef4 0000035c 00000902 00000b92 000010f9 00001693 0000134c 00000355 00000748 000008b9 00000fd7 000013fa 00000eb8 00000051 00001b75 000003cd 0000038a 00001731 00001b85 00001bac 00000e2b 00000491 000009b9 00000249 00001d9a 000005c2 00000226 00001cbf 00001e8d 00001b33 000015ac 000016cc 00001a47 00001463 0000046b 00000013 00001a9e 000009e7 00001483 00001bbc 000014e2 00000a59 000014fe 00001df3 0000150d 000004c0 00001e72 0000056e 0000164f 000016ca 000019f9 00000e89 00000fa4 00000165 00001558 000011e1 00001800 000016ac 00000418 00001d61 00000ce2 00000d21 0000070a 00001b3d 00000fa5 00000f0f 00001ef0 00001c11 000003af 00000279 000015d0 00001851 00001c3b 000002ee 00001c14 00000217 000014d9 00001c64 00000379 000019b5 000014e4 00000f0a 00000dc9 00001ba0 00000e3d 000018d2 00001872 00001d77 00001171 00001bd2 0000076f 0000057b 00000fc0 00000293 00000fef 0000030e 00001bf8 00001506 0000119b 00001866 000001be 00000d7e 00000444 00001aa5 00001970 00001030 00000a68 00000cf2 00001284 0000045b 0000148f 00000b4d 000008c6 00000e4f 00001e50 00001ca3 000006d0 000001d6 00000aee 00001c95 000009b1 00001526 0000113f 000011b3 0000125d 00000497 000009b5 000014d8 0000173c 0000143d 00000ff9 0000197c 00001cda 0000077a 000015ad 0000013e 0000163a 00001183 00001340 0000166f 000001f9 000003e1 00000ba2 00000bc9 00001758 00001619 00000b7f 000013af 00000cac 00001755 00000022 00001c8a 0000090f 00000aa7 00000a1d 00000755 000012d0 00000090 00001675 000014cc 00000ddc 0000110c 00000513 00000b76 000003f7 00000a02 00001eb6 00001640 00001ccd 00001c8f 000001b3 000010a7 00001d4a 00001932 000007f7 000009b1 0000028f 000019e8 00000f66 0000141e 00000a9d 0000140c 0000177b 00001e5c 00000dd6 00000a29 00000ceb 00000805 00001c3d 00001ae8 000001b2 0000064f 000014a7 000015d6 00000d88 00001946 000000ff 000003f1 00001441 00001047 00000631 0000076c 00001464 00000b45 0000141d 00000e66 0000012b 000008dc 00001403 00000b59 00001ae9 0000147e 000012e3 00001dde 00000092 000012d3 00001e38 0000127e 00000dde 0000011d 00000f01 00000887 0000014b 00001df2 000017b5 00001ba1 00001393 000009b0 00000c2c 00000846 00001b78 00001dcd 00000bc6 00001b24 00000a8f 00000da3 0000145d 0000142c 000018ad 00001828 0000163f 00000a6a 000007dc 00001d45 00000634 00001913 00000fa9 000014fa 00001cec 0000016a 0000044c 000001d0 000012fe 00000663 000004b4 00000af9 00001e05 000015dc 00001a24 00001a2f 00001b06 00001c5b 00001217 00001813 000011b4 00001eb3 00000d1d 00000c83 00001bcc 00000c61 000008c3 0000173e 0000132b 0000015d 0000196b 000007af 00000817 00001307 000007fc 0000137b 0000071b 00000dab 000013ea 000016e8 00000077 00000aad 00001dc1 00001577 00000e9b 00001d92 00000405 0000122c 00000eca 000011cd 0000088c 00000c31 00001e6f 000002ee 00000173 00000b14 0000078f 00001c37 000012c9 00001c5f 00000abb 00001acc 00000e58 00001da1 00000075 00001de4 00000d52 00000dd8 00000197 00001b3c 000010fb 00000baf 000014f2 0000084d 00000ae8 00000206 0000181a 0000126a 000019fa 00000b7f 00001b4d 000002ec 00000d2b 00000851 000015bd 00000750 00000c25 00001abe 00001c5a 00001445 00001ecf 000012ef 000000e6 00001426 00000186 00000dd6 00000a6c 0000020b 00000e79 00000f1b 00001e5a 00000fb2 00000786 00000f07 0000074f 00001dcb 0000137d 00000979 00000182 00001a11 00000b0a 00000291 0000021a 000003a9 000017f6 0000044a 00000b43 00000200 000008ec 00001017 00001ed1 00000175 00001a9a 00001592 00000ffd 00000356 00000b73 00000c62 00001245 000009b6 00001ae3 0000075f 00000385 000011f4 0000029a 000012c4 0000170c 00000f95 00001e76 000012b5 000016ce 00001322 000014b2 00000b64 0000004f 000007fa 00001974 00001267 00001271 000005e6 00000c47 00001677 000002a1 00001700 000015e8 00001864 00000ac6 000007ea 00001359 000001a4 00000536 000010a6 00001294 00000173 00000ed7 00000e42 00000a7a 00000e8a 0000057e 000005ec 00001391 000013d1 0000128a 00000bda 0000048e 0000138e 0000047a 00001bea 0000040d 00001437 0000018b 00000f8e 000011af 000001d5 0000109b 00001a90 000009b6 00001f1c 0000082a 000011b9 000009dd 000006df 000001b5 0000113e 00000d0f 00000c40 000002e3 000003e3 00000f7b 00000c9c 0000017f 00000345 00001c59 00001460 00001725 0000037a 000010a5 00000edb 00000923 00001254 00000748 000019dc 00001cae 00000dec 0000072d 00000491 00000fa1 00001358 0000156f 00000ea5 000007ab 00001893 00000bc1 00000b08 0000011b 00000187 000016ea 00000b93 0000132a 00001d99 0000157f 0000104b 000017de 0000196a 000000c9 00000f42 00000298 00000f91 00001604 00001ad7 00000984 00000a99 00001af7 00001f3a 000006a5 0000105c 000019e5 00000c31 00001f03 00000fd5 000017f0 00001df1 00001a75 00000bfc 00000f4f 00000df4 000004a1 00000f40 000009f3 00001e2f 00000183 000010f8 00001a5a 00000537 00001bfc 00000779 00001df6 000013aa 00000075 0000098c 00001c38 000018ee 0000166e 0000126f 00000620 00000839 000014f1 0000128c 00000af6 000011f3 00001d31 000018de 00000ff7 0000064b 0000036f 00000556 00001ce6 0000041c 00000668 00000616 0000130c 00001304 000019f9 00001559 00000675 00000956 00001d67 000001fa 00001139 00001edd 0000006a 00001d69 00001ac6 00001783 00001b0e 00000b66 00001991 000001e7 0000186b 00000a79 00001ccd 00001b59 0000128b 00001380 0000157e 0000036e 000007cc 0000121b 000015c9 000004b3 00001852 0000003c 00000077 000000dd 00000bd2 00000440 0000098d 000015fb 000008d2 00000984 00000a00 00000fdf 00001b52 000001df 00000834 00001457 00000159 00001a85 00001c6a 00000e61 000004ee 00001635 00000c96 0000156d 00000078 00000a39 00000fc6 000013d3 00001b1f 000014f0 00000db6 0000151f 0000095b 000000a2 00000116 00001ad4 00001e77 00001935 000005ac 00001d78 00001269 0000131e 000009b3 00000dbc 00000926 0000081c 00001c84 00000e52 00000a95 000009f1 00000a25 00000979 00001b9a 00000ccf 0000110b 00000862 00000561 0000184a 00000303 00001c07 00001e87 000013a8 00001d3b 0000184e 00001068 000013ed 00000061 00001033 000010e1 000019c6 0000048b 00000acc 00001eef 000016de 000009c0 00001d9f 00000be6 00000589 00001b92 000005c8 0000084a 00000fd2 00000c72 00000ce3 00000bdb 00001b1c 0000166f 00000905 0000171d 0000068b 00000171 00000449 00000a7b 0000192e 000017db 00000b20 00001ee5 000001de 00000d05 000004a5 00001345 00000864 0000059a 00001537 00001dd3 00001143 00000639 000004e4 0000156e 000002f6 00001e20 00001f0d 00000ceb 00000853 00000466 00000abf 00001834 00001e5c 0000059e 000014e0 00001d7c 0000162d 0000132b 0000159b 000009d0 000000bc 00000cff 00000581 00000732 000010c2 000006c0 0000188f 0000115f 0000016b 00000f82 000003ea 00001df2 00001e10 00001cd1 00000a79 00000cc5 000001b1 000019a5 00001c32 00000389 00001b61 000019a2 0000169d 00000a2c 00000fc8 0000021a 00000108 00000dfc 00001748 00000b94 000011e2 00000613 00001838 000014e3 0000166f 000010ed 0000044e 000007fe 000012c5 0000071c 0000144e 000000eb 000010db 0000066d 00001edc 00001ca8 00001b39 00001bd1 00001579 0000070d 00000f47 000000b7 00000655 00000320 000013d6 000017cf 000012d4 00001549 00000204 0000152f 000004c7 00000d45 00000b9b 0000174d 00000400 000012e2 00001c23 0000133f 00001ddd 0000001f 000002a7 000008e3 00000484 00000c4a 00000e51 00000012 00000e6c 000009dc 00001864 000017f9 00001b32 00000260 00001784 00001c7f 00001698 00001905 000012b0 000014c5 00001def 00001588 00000b84 000000af 00000192 00001d89 00000a01 000002c4 00001a01 00001f1e 00001c91 00000d53 0000158f 00000536 00001985 00001db0 0000089d 00001215 000009b5 00000310 0000111e 00001474 00001323 00000954 00001036 00001b34 00001d88 00001bcb 000010bb 000004ad 0000047f 000014d6 00000983 000016bc 00000a3e 00001004 00001d2c 00001015 00000eee 000002f1 0000132b 00001083 000009fa 00000a1f 00001ca7 000009e0 00001355 0000133f 000003ed 0000053d 00000fca 00000bf6 00001605 000006ea 000007a8 00001b39 00000d7a 00001732 00000b6f 0000038d 000013e5 0000192d 00000015 000007ea 00000efa 00001ec1 00000fad 00000a30 00001548 00001102 000005bf 00001b72 00000b55 00000247 000004bf 00001631 00001815 000004fb 00001841 00000ae8 000005c7 0000008a 000018e5 00001e70 000000dc 00001c81 00000de4 000001be 00000054 00001349 000008d5 0000175e 00001890 0000139c 00001437 00000008 0000109d 0000097e 00000411 00001cad 000009e4 000013c6 0000188e 00001068 0000178d 00001e06 0000061a 00001d2e 000010ac 000005ae 00000dbc 00000339 000002ee 00001db6 00000755 000000d5 00000acb 000007e0 00001a47 00001404 00001878 0000005a 0000080b 0000084b 00001e30 00001450 00000533 00001760 00001f3b 000014f4 00000926 00000180 00000e8b 00001a1e 00001442 00000691 00000cee 00000dbf 000017ed 00001826 000002e3 00001515 0000101a 00001ac0 0000162a 00000f1f 00001898 00000f19 000018e8 00001d8f 00000ae2 00001eaf 00001c94 00001918 00000847 00000bd6 0000111b 0000009e 00001aa3 0000117a 000015aa 0000012b 00001d1e 00001a5b 00001d57 0000039f 000005be 00001dc8 00000754 000013e8 000000a0 00001859 0000095f 00001a1d 000011cd 00000cda 00001d93 00000cf1 000004e0 00000a23 00000cee 0000004f 00001270 00000ac8 00000b79 00000cfe 000000ab 000012ea 000004e4 00001559 0000042c 0000052f 000019b0 00000ac7 00000f62 000018e2 000000b2 0000172d 000011d1 00000c16 00000d38 00000f15 00001da8 00001d3a 000010f7 00001dbf 00001871 00000a68 0000139d 00001e89 000011e3 00001cc5 000004a6 00000baf 000008a7 000000f7 000001ed 00000abe 00001314 0000118d 00000250 0000062d 000009f8 000012c5 0000116a 00001713 000011b0 000003d5 000015c5 00000a69 000012e3 0000137b 00001952 000001b3 000015f8 0000046e 000007eb 0000061b 00001bdc 00000ab6 0000012a 00000196 00000234 00001b94 00000557 00001d81 0000048c 00001d36 00001a6d 0000108d 00000446 0000075f 00000873 00000797 00001763 00001b45 00001879 000014c7 00000ec7 00000845 00000028 0000142a 00000df9 000009b1 00000ece 00000bdb 0000181b 00001d33 00001bda 000000df 000000a9 00000501 00001a99 00001b27 00001e00 00000578 000000ec 00001e8d 0000091f 00001468 0000078a 0000062c 00000052 00000a95 00000824 000012bb 000013d3 00000ba7 0000141e 00001d2d 000014eb 0000093a 00000d14 0000087d 00000a30 000006ac 00001ee8 0000140e 00000d99 00000b6d 0000076d 00001bbd 00001dcf 0000013d 00000926 000010dc 00000f0b 00001d26 00000871 00001200 00001349 00001406 00000114 00000095 00001436 000019ba 00001801 00000cba 0000137c 00001abe 00000254 0000085f 00000452 00001cae 0000068f 0000090c 0000057b 000013a8 00000319 00001d95 000019cb 00000e4b 00000694 0000174e 00001ee5 000000fe 00000271 00000d2e 00000ca3 00000be7 00000622 000001df 00000db8 00001c5d 00001f0c 00001188 00001908 000010b9 00000ba9 000016c3 000004ad 00000681 00001e90 00001069 000015b2 00000456 0000096e 000010e8 0000123e 000018f3 00001094 0000006c 00000a4a 00000e5f 00001878 000001cd 000015b6 00001b72 00000150 00001a84 00001f16 00001044 00000b64 000012c5 000006fc 000007e2 00000fe7 00000da6 00000b48 0000011d 00001776 00000a54 000013cd 00001457 0000176a 00001054 000000c6 00000d4c 00000f6b 00001909 00001d32 00001705 000008e4 00001084 00001dcd 00000d8f 0000047b 00000987 00000f8e 000002cd 000001e9 00001933 00001d2c 00000778 00001aab 00001a41 00000651 00000d4b 00001223 000011e9 000018a5 00000456 00001c0e 0000123c 00001e3b 00000209 0000013f 000009f8 00000889 000014b8 0000157c 000017d3 00001103 00000abb 000012a5 000013fd 00001c84 000016f7 00000257 00001f05 000001e7 00001a0c 0000020f 00000777 00000394 00000254 00000e43 00001015 00001ec3 00000c57 00001bba 000008b2 00001076 00000a28 000003bd 00000027 0000151c 000016fa 0000052f 0000199f 0000015e 0000154d 00001199 00000843 00000cab 00001350 000011d7 00001ec3 00000eab 00001c92 00001671 0000096a 000005ed 000008ad 00001dd5 00001dc1 000010d6 00001cea 00000848 00001d5e 00000e3e 00000ada 000006f3 000011ca 000002a7 00001c6f 00000eb5 0000169c 000009fb 00000c83 00001c8b 00001928 0000159c 00000c15 00000b12 0000190d 00000ac4 000006c1 000012bc 00001338 00000dc7 0000093f 000006db 000018fe 00001576 00000efb 00000cb6 000004e4 00001a19 00000168 00000bee 00000068 00000cc0 0000155d 000001cc 00000053 00000f17 0000191a 0000095d 00000da1 00001192 00001b7d 00000024 000001f5 000010d2 00000b87 00000670 00001e60 000008e4 00001ec8 000015e8 00000429 00000bd2 000017c3 00001d44 00001994 00000bae 00000a69 00000916 00000b5f 00001516 00000c4b 000009e0 00000eb9 00001f39 000017d8 00000e04 00001664 00000951 00000cdb 000009e7 0000049f 000011c0 00001ac7 00001734 00001064 00000a85 00000d18 000000f7 00001040 00000433 00000406 00001da2 0000153f 00001380 000001b3 00001a32 00000a46 00001c2b 000017ab 00000f0b 0000130c 00000052 00001944 000014da 000011eb 00000b8f 000011e2 00000932 0000191a 00001d2e 00000529 00000e9f 00000e43 0000178f 000011a1 000006af 000012a2 00001690 00000b53 00000620 00001794 00001900 0000072c 000016c6 0000060b 00000fa7 000009d6 00001712 0000169c 00001afb 00001e75 0000083d 00001f11 00001c11 0000069b 000013bd 00000625 00001172 00000790 00001574 00000e4e 000005bc 0000124a 00000654 00000b7c 00001a72 00000a72 000013fa 0000084f 0000037d 000011ac 000014c2 000000e5 00000083 00000975 00001934 0000135b 00001728 0000012c 000000d4 000004ae 00000d2d 00001b54 00000dd8 000000d2 00000f22 00000b01 000001ec 00001a53 00000b40 000007b5 00001d2e 00000169 00001d27 00000eea 00000254 00000665 0000177f 00000411 00001c70 00000123 00001de9 00001bd6 00001c18 00001a9d 00000f45 000000eb 0000151e 000016a6 000011cd 00001285 0000117c 00001805 00000131 00000746 00001b1e 0000050c 000013ee 00000ca0 00001a04 00001ad0 0000171c 000002e1 00000e3a 00001d58 00001770 00000a2a 00000e7d 00001339 00001488 00001793 0000108e 00001661 00000665 000003c2 00000785 00001c91 0000157a 00001bf4 00001c2c 00001110 00000e67 000015d0 00001a0e 0000056a 0000008d 00001b6d 00001629 00000523 00000b99 0000067b 00000496 00000160 00001810 00001148 0000045f 0000017d 0000054e 00001427

module cache_tb();

`define DATA_COUNT (2000)
`define RDWR_COUNT (6*`DATA_COUNT)

reg wr_cycle           [`RDWR_COUNT];
reg rd_cycle           [`RDWR_COUNT];
reg [31:0] addr_rom    [`RDWR_COUNT];
reg [31:0] wr_data_rom [`RDWR_COUNT];
reg [31:0] validation_data [`DATA_COUNT];

initial begin
    // 2000 sequence write cycles
    rd_cycle[    0] = 1'b0;  wr_cycle[    0] = 1'b1;  addr_rom[    0]='h00000000;  wr_data_rom[    0]='h00000042;
    rd_cycle[    1] = 1'b0;  wr_cycle[    1] = 1'b1;  addr_rom[    1]='h00000004;  wr_data_rom[    1]='h000004f8;
    rd_cycle[    2] = 1'b0;  wr_cycle[    2] = 1'b1;  addr_rom[    2]='h00000008;  wr_data_rom[    2]='h000011e6;
    rd_cycle[    3] = 1'b0;  wr_cycle[    3] = 1'b1;  addr_rom[    3]='h0000000c;  wr_data_rom[    3]='h00000c3c;
    rd_cycle[    4] = 1'b0;  wr_cycle[    4] = 1'b1;  addr_rom[    4]='h00000010;  wr_data_rom[    4]='h00000666;
    rd_cycle[    5] = 1'b0;  wr_cycle[    5] = 1'b1;  addr_rom[    5]='h00000014;  wr_data_rom[    5]='h0000077e;
    rd_cycle[    6] = 1'b0;  wr_cycle[    6] = 1'b1;  addr_rom[    6]='h00000018;  wr_data_rom[    6]='h00001064;
    rd_cycle[    7] = 1'b0;  wr_cycle[    7] = 1'b1;  addr_rom[    7]='h0000001c;  wr_data_rom[    7]='h00000fb1;
    rd_cycle[    8] = 1'b0;  wr_cycle[    8] = 1'b1;  addr_rom[    8]='h00000020;  wr_data_rom[    8]='h000001a3;
    rd_cycle[    9] = 1'b0;  wr_cycle[    9] = 1'b1;  addr_rom[    9]='h00000024;  wr_data_rom[    9]='h000004ef;
    rd_cycle[   10] = 1'b0;  wr_cycle[   10] = 1'b1;  addr_rom[   10]='h00000028;  wr_data_rom[   10]='h000019eb;
    rd_cycle[   11] = 1'b0;  wr_cycle[   11] = 1'b1;  addr_rom[   11]='h0000002c;  wr_data_rom[   11]='h000007c6;
    rd_cycle[   12] = 1'b0;  wr_cycle[   12] = 1'b1;  addr_rom[   12]='h00000030;  wr_data_rom[   12]='h00000b9b;
    rd_cycle[   13] = 1'b0;  wr_cycle[   13] = 1'b1;  addr_rom[   13]='h00000034;  wr_data_rom[   13]='h00001807;
    rd_cycle[   14] = 1'b0;  wr_cycle[   14] = 1'b1;  addr_rom[   14]='h00000038;  wr_data_rom[   14]='h00001e4b;
    rd_cycle[   15] = 1'b0;  wr_cycle[   15] = 1'b1;  addr_rom[   15]='h0000003c;  wr_data_rom[   15]='h000002f0;
    rd_cycle[   16] = 1'b0;  wr_cycle[   16] = 1'b1;  addr_rom[   16]='h00000040;  wr_data_rom[   16]='h00000e7f;
    rd_cycle[   17] = 1'b0;  wr_cycle[   17] = 1'b1;  addr_rom[   17]='h00000044;  wr_data_rom[   17]='h000008e4;
    rd_cycle[   18] = 1'b0;  wr_cycle[   18] = 1'b1;  addr_rom[   18]='h00000048;  wr_data_rom[   18]='h0000152a;
    rd_cycle[   19] = 1'b0;  wr_cycle[   19] = 1'b1;  addr_rom[   19]='h0000004c;  wr_data_rom[   19]='h00000512;
    rd_cycle[   20] = 1'b0;  wr_cycle[   20] = 1'b1;  addr_rom[   20]='h00000050;  wr_data_rom[   20]='h000000e7;
    rd_cycle[   21] = 1'b0;  wr_cycle[   21] = 1'b1;  addr_rom[   21]='h00000054;  wr_data_rom[   21]='h00001366;
    rd_cycle[   22] = 1'b0;  wr_cycle[   22] = 1'b1;  addr_rom[   22]='h00000058;  wr_data_rom[   22]='h000019d5;
    rd_cycle[   23] = 1'b0;  wr_cycle[   23] = 1'b1;  addr_rom[   23]='h0000005c;  wr_data_rom[   23]='h000012d4;
    rd_cycle[   24] = 1'b0;  wr_cycle[   24] = 1'b1;  addr_rom[   24]='h00000060;  wr_data_rom[   24]='h00001082;
    rd_cycle[   25] = 1'b0;  wr_cycle[   25] = 1'b1;  addr_rom[   25]='h00000064;  wr_data_rom[   25]='h00001407;
    rd_cycle[   26] = 1'b0;  wr_cycle[   26] = 1'b1;  addr_rom[   26]='h00000068;  wr_data_rom[   26]='h00001e13;
    rd_cycle[   27] = 1'b0;  wr_cycle[   27] = 1'b1;  addr_rom[   27]='h0000006c;  wr_data_rom[   27]='h00000979;
    rd_cycle[   28] = 1'b0;  wr_cycle[   28] = 1'b1;  addr_rom[   28]='h00000070;  wr_data_rom[   28]='h00000a69;
    rd_cycle[   29] = 1'b0;  wr_cycle[   29] = 1'b1;  addr_rom[   29]='h00000074;  wr_data_rom[   29]='h0000038c;
    rd_cycle[   30] = 1'b0;  wr_cycle[   30] = 1'b1;  addr_rom[   30]='h00000078;  wr_data_rom[   30]='h0000010c;
    rd_cycle[   31] = 1'b0;  wr_cycle[   31] = 1'b1;  addr_rom[   31]='h0000007c;  wr_data_rom[   31]='h00000545;
    rd_cycle[   32] = 1'b0;  wr_cycle[   32] = 1'b1;  addr_rom[   32]='h00000080;  wr_data_rom[   32]='h00001f25;
    rd_cycle[   33] = 1'b0;  wr_cycle[   33] = 1'b1;  addr_rom[   33]='h00000084;  wr_data_rom[   33]='h00001826;
    rd_cycle[   34] = 1'b0;  wr_cycle[   34] = 1'b1;  addr_rom[   34]='h00000088;  wr_data_rom[   34]='h0000003b;
    rd_cycle[   35] = 1'b0;  wr_cycle[   35] = 1'b1;  addr_rom[   35]='h0000008c;  wr_data_rom[   35]='h00001e63;
    rd_cycle[   36] = 1'b0;  wr_cycle[   36] = 1'b1;  addr_rom[   36]='h00000090;  wr_data_rom[   36]='h00001039;
    rd_cycle[   37] = 1'b0;  wr_cycle[   37] = 1'b1;  addr_rom[   37]='h00000094;  wr_data_rom[   37]='h00001156;
    rd_cycle[   38] = 1'b0;  wr_cycle[   38] = 1'b1;  addr_rom[   38]='h00000098;  wr_data_rom[   38]='h00001daa;
    rd_cycle[   39] = 1'b0;  wr_cycle[   39] = 1'b1;  addr_rom[   39]='h0000009c;  wr_data_rom[   39]='h00000bed;
    rd_cycle[   40] = 1'b0;  wr_cycle[   40] = 1'b1;  addr_rom[   40]='h000000a0;  wr_data_rom[   40]='h000010db;
    rd_cycle[   41] = 1'b0;  wr_cycle[   41] = 1'b1;  addr_rom[   41]='h000000a4;  wr_data_rom[   41]='h0000127e;
    rd_cycle[   42] = 1'b0;  wr_cycle[   42] = 1'b1;  addr_rom[   42]='h000000a8;  wr_data_rom[   42]='h000017d8;
    rd_cycle[   43] = 1'b0;  wr_cycle[   43] = 1'b1;  addr_rom[   43]='h000000ac;  wr_data_rom[   43]='h00001c64;
    rd_cycle[   44] = 1'b0;  wr_cycle[   44] = 1'b1;  addr_rom[   44]='h000000b0;  wr_data_rom[   44]='h000018aa;
    rd_cycle[   45] = 1'b0;  wr_cycle[   45] = 1'b1;  addr_rom[   45]='h000000b4;  wr_data_rom[   45]='h00000b5d;
    rd_cycle[   46] = 1'b0;  wr_cycle[   46] = 1'b1;  addr_rom[   46]='h000000b8;  wr_data_rom[   46]='h00001842;
    rd_cycle[   47] = 1'b0;  wr_cycle[   47] = 1'b1;  addr_rom[   47]='h000000bc;  wr_data_rom[   47]='h00001c84;
    rd_cycle[   48] = 1'b0;  wr_cycle[   48] = 1'b1;  addr_rom[   48]='h000000c0;  wr_data_rom[   48]='h00000731;
    rd_cycle[   49] = 1'b0;  wr_cycle[   49] = 1'b1;  addr_rom[   49]='h000000c4;  wr_data_rom[   49]='h00001474;
    rd_cycle[   50] = 1'b0;  wr_cycle[   50] = 1'b1;  addr_rom[   50]='h000000c8;  wr_data_rom[   50]='h0000122d;
    rd_cycle[   51] = 1'b0;  wr_cycle[   51] = 1'b1;  addr_rom[   51]='h000000cc;  wr_data_rom[   51]='h0000172e;
    rd_cycle[   52] = 1'b0;  wr_cycle[   52] = 1'b1;  addr_rom[   52]='h000000d0;  wr_data_rom[   52]='h0000029a;
    rd_cycle[   53] = 1'b0;  wr_cycle[   53] = 1'b1;  addr_rom[   53]='h000000d4;  wr_data_rom[   53]='h00001b2e;
    rd_cycle[   54] = 1'b0;  wr_cycle[   54] = 1'b1;  addr_rom[   54]='h000000d8;  wr_data_rom[   54]='h00001b60;
    rd_cycle[   55] = 1'b0;  wr_cycle[   55] = 1'b1;  addr_rom[   55]='h000000dc;  wr_data_rom[   55]='h0000099a;
    rd_cycle[   56] = 1'b0;  wr_cycle[   56] = 1'b1;  addr_rom[   56]='h000000e0;  wr_data_rom[   56]='h00001802;
    rd_cycle[   57] = 1'b0;  wr_cycle[   57] = 1'b1;  addr_rom[   57]='h000000e4;  wr_data_rom[   57]='h00001157;
    rd_cycle[   58] = 1'b0;  wr_cycle[   58] = 1'b1;  addr_rom[   58]='h000000e8;  wr_data_rom[   58]='h00001e11;
    rd_cycle[   59] = 1'b0;  wr_cycle[   59] = 1'b1;  addr_rom[   59]='h000000ec;  wr_data_rom[   59]='h00001b7f;
    rd_cycle[   60] = 1'b0;  wr_cycle[   60] = 1'b1;  addr_rom[   60]='h000000f0;  wr_data_rom[   60]='h00001340;
    rd_cycle[   61] = 1'b0;  wr_cycle[   61] = 1'b1;  addr_rom[   61]='h000000f4;  wr_data_rom[   61]='h00000042;
    rd_cycle[   62] = 1'b0;  wr_cycle[   62] = 1'b1;  addr_rom[   62]='h000000f8;  wr_data_rom[   62]='h00000cdb;
    rd_cycle[   63] = 1'b0;  wr_cycle[   63] = 1'b1;  addr_rom[   63]='h000000fc;  wr_data_rom[   63]='h000016fb;
    rd_cycle[   64] = 1'b0;  wr_cycle[   64] = 1'b1;  addr_rom[   64]='h00000100;  wr_data_rom[   64]='h0000069f;
    rd_cycle[   65] = 1'b0;  wr_cycle[   65] = 1'b1;  addr_rom[   65]='h00000104;  wr_data_rom[   65]='h00001c6e;
    rd_cycle[   66] = 1'b0;  wr_cycle[   66] = 1'b1;  addr_rom[   66]='h00000108;  wr_data_rom[   66]='h00001cab;
    rd_cycle[   67] = 1'b0;  wr_cycle[   67] = 1'b1;  addr_rom[   67]='h0000010c;  wr_data_rom[   67]='h0000008c;
    rd_cycle[   68] = 1'b0;  wr_cycle[   68] = 1'b1;  addr_rom[   68]='h00000110;  wr_data_rom[   68]='h0000166d;
    rd_cycle[   69] = 1'b0;  wr_cycle[   69] = 1'b1;  addr_rom[   69]='h00000114;  wr_data_rom[   69]='h00001e3d;
    rd_cycle[   70] = 1'b0;  wr_cycle[   70] = 1'b1;  addr_rom[   70]='h00000118;  wr_data_rom[   70]='h000011eb;
    rd_cycle[   71] = 1'b0;  wr_cycle[   71] = 1'b1;  addr_rom[   71]='h0000011c;  wr_data_rom[   71]='h0000151a;
    rd_cycle[   72] = 1'b0;  wr_cycle[   72] = 1'b1;  addr_rom[   72]='h00000120;  wr_data_rom[   72]='h00001d92;
    rd_cycle[   73] = 1'b0;  wr_cycle[   73] = 1'b1;  addr_rom[   73]='h00000124;  wr_data_rom[   73]='h000015a1;
    rd_cycle[   74] = 1'b0;  wr_cycle[   74] = 1'b1;  addr_rom[   74]='h00000128;  wr_data_rom[   74]='h000002e7;
    rd_cycle[   75] = 1'b0;  wr_cycle[   75] = 1'b1;  addr_rom[   75]='h0000012c;  wr_data_rom[   75]='h00000588;
    rd_cycle[   76] = 1'b0;  wr_cycle[   76] = 1'b1;  addr_rom[   76]='h00000130;  wr_data_rom[   76]='h000012ed;
    rd_cycle[   77] = 1'b0;  wr_cycle[   77] = 1'b1;  addr_rom[   77]='h00000134;  wr_data_rom[   77]='h000011ea;
    rd_cycle[   78] = 1'b0;  wr_cycle[   78] = 1'b1;  addr_rom[   78]='h00000138;  wr_data_rom[   78]='h0000179d;
    rd_cycle[   79] = 1'b0;  wr_cycle[   79] = 1'b1;  addr_rom[   79]='h0000013c;  wr_data_rom[   79]='h00001969;
    rd_cycle[   80] = 1'b0;  wr_cycle[   80] = 1'b1;  addr_rom[   80]='h00000140;  wr_data_rom[   80]='h00000ce7;
    rd_cycle[   81] = 1'b0;  wr_cycle[   81] = 1'b1;  addr_rom[   81]='h00000144;  wr_data_rom[   81]='h000000a3;
    rd_cycle[   82] = 1'b0;  wr_cycle[   82] = 1'b1;  addr_rom[   82]='h00000148;  wr_data_rom[   82]='h0000160e;
    rd_cycle[   83] = 1'b0;  wr_cycle[   83] = 1'b1;  addr_rom[   83]='h0000014c;  wr_data_rom[   83]='h00000453;
    rd_cycle[   84] = 1'b0;  wr_cycle[   84] = 1'b1;  addr_rom[   84]='h00000150;  wr_data_rom[   84]='h00001d70;
    rd_cycle[   85] = 1'b0;  wr_cycle[   85] = 1'b1;  addr_rom[   85]='h00000154;  wr_data_rom[   85]='h00000315;
    rd_cycle[   86] = 1'b0;  wr_cycle[   86] = 1'b1;  addr_rom[   86]='h00000158;  wr_data_rom[   86]='h00000af6;
    rd_cycle[   87] = 1'b0;  wr_cycle[   87] = 1'b1;  addr_rom[   87]='h0000015c;  wr_data_rom[   87]='h000005a8;
    rd_cycle[   88] = 1'b0;  wr_cycle[   88] = 1'b1;  addr_rom[   88]='h00000160;  wr_data_rom[   88]='h00000066;
    rd_cycle[   89] = 1'b0;  wr_cycle[   89] = 1'b1;  addr_rom[   89]='h00000164;  wr_data_rom[   89]='h0000097c;
    rd_cycle[   90] = 1'b0;  wr_cycle[   90] = 1'b1;  addr_rom[   90]='h00000168;  wr_data_rom[   90]='h00001e4c;
    rd_cycle[   91] = 1'b0;  wr_cycle[   91] = 1'b1;  addr_rom[   91]='h0000016c;  wr_data_rom[   91]='h00000ac7;
    rd_cycle[   92] = 1'b0;  wr_cycle[   92] = 1'b1;  addr_rom[   92]='h00000170;  wr_data_rom[   92]='h00001128;
    rd_cycle[   93] = 1'b0;  wr_cycle[   93] = 1'b1;  addr_rom[   93]='h00000174;  wr_data_rom[   93]='h00000d54;
    rd_cycle[   94] = 1'b0;  wr_cycle[   94] = 1'b1;  addr_rom[   94]='h00000178;  wr_data_rom[   94]='h00000ed1;
    rd_cycle[   95] = 1'b0;  wr_cycle[   95] = 1'b1;  addr_rom[   95]='h0000017c;  wr_data_rom[   95]='h000016dd;
    rd_cycle[   96] = 1'b0;  wr_cycle[   96] = 1'b1;  addr_rom[   96]='h00000180;  wr_data_rom[   96]='h00001dd4;
    rd_cycle[   97] = 1'b0;  wr_cycle[   97] = 1'b1;  addr_rom[   97]='h00000184;  wr_data_rom[   97]='h000004d5;
    rd_cycle[   98] = 1'b0;  wr_cycle[   98] = 1'b1;  addr_rom[   98]='h00000188;  wr_data_rom[   98]='h00000946;
    rd_cycle[   99] = 1'b0;  wr_cycle[   99] = 1'b1;  addr_rom[   99]='h0000018c;  wr_data_rom[   99]='h00000461;
    rd_cycle[  100] = 1'b0;  wr_cycle[  100] = 1'b1;  addr_rom[  100]='h00000190;  wr_data_rom[  100]='h00001d74;
    rd_cycle[  101] = 1'b0;  wr_cycle[  101] = 1'b1;  addr_rom[  101]='h00000194;  wr_data_rom[  101]='h00000746;
    rd_cycle[  102] = 1'b0;  wr_cycle[  102] = 1'b1;  addr_rom[  102]='h00000198;  wr_data_rom[  102]='h00001907;
    rd_cycle[  103] = 1'b0;  wr_cycle[  103] = 1'b1;  addr_rom[  103]='h0000019c;  wr_data_rom[  103]='h000007ed;
    rd_cycle[  104] = 1'b0;  wr_cycle[  104] = 1'b1;  addr_rom[  104]='h000001a0;  wr_data_rom[  104]='h00001783;
    rd_cycle[  105] = 1'b0;  wr_cycle[  105] = 1'b1;  addr_rom[  105]='h000001a4;  wr_data_rom[  105]='h000009b6;
    rd_cycle[  106] = 1'b0;  wr_cycle[  106] = 1'b1;  addr_rom[  106]='h000001a8;  wr_data_rom[  106]='h0000042b;
    rd_cycle[  107] = 1'b0;  wr_cycle[  107] = 1'b1;  addr_rom[  107]='h000001ac;  wr_data_rom[  107]='h000002c7;
    rd_cycle[  108] = 1'b0;  wr_cycle[  108] = 1'b1;  addr_rom[  108]='h000001b0;  wr_data_rom[  108]='h000007bc;
    rd_cycle[  109] = 1'b0;  wr_cycle[  109] = 1'b1;  addr_rom[  109]='h000001b4;  wr_data_rom[  109]='h00000c91;
    rd_cycle[  110] = 1'b0;  wr_cycle[  110] = 1'b1;  addr_rom[  110]='h000001b8;  wr_data_rom[  110]='h00001a53;
    rd_cycle[  111] = 1'b0;  wr_cycle[  111] = 1'b1;  addr_rom[  111]='h000001bc;  wr_data_rom[  111]='h00001d92;
    rd_cycle[  112] = 1'b0;  wr_cycle[  112] = 1'b1;  addr_rom[  112]='h000001c0;  wr_data_rom[  112]='h00000e32;
    rd_cycle[  113] = 1'b0;  wr_cycle[  113] = 1'b1;  addr_rom[  113]='h000001c4;  wr_data_rom[  113]='h00000e08;
    rd_cycle[  114] = 1'b0;  wr_cycle[  114] = 1'b1;  addr_rom[  114]='h000001c8;  wr_data_rom[  114]='h00000cdb;
    rd_cycle[  115] = 1'b0;  wr_cycle[  115] = 1'b1;  addr_rom[  115]='h000001cc;  wr_data_rom[  115]='h00001cbd;
    rd_cycle[  116] = 1'b0;  wr_cycle[  116] = 1'b1;  addr_rom[  116]='h000001d0;  wr_data_rom[  116]='h00001c03;
    rd_cycle[  117] = 1'b0;  wr_cycle[  117] = 1'b1;  addr_rom[  117]='h000001d4;  wr_data_rom[  117]='h00001aa8;
    rd_cycle[  118] = 1'b0;  wr_cycle[  118] = 1'b1;  addr_rom[  118]='h000001d8;  wr_data_rom[  118]='h00001088;
    rd_cycle[  119] = 1'b0;  wr_cycle[  119] = 1'b1;  addr_rom[  119]='h000001dc;  wr_data_rom[  119]='h00001196;
    rd_cycle[  120] = 1'b0;  wr_cycle[  120] = 1'b1;  addr_rom[  120]='h000001e0;  wr_data_rom[  120]='h00000a78;
    rd_cycle[  121] = 1'b0;  wr_cycle[  121] = 1'b1;  addr_rom[  121]='h000001e4;  wr_data_rom[  121]='h000002de;
    rd_cycle[  122] = 1'b0;  wr_cycle[  122] = 1'b1;  addr_rom[  122]='h000001e8;  wr_data_rom[  122]='h000015d1;
    rd_cycle[  123] = 1'b0;  wr_cycle[  123] = 1'b1;  addr_rom[  123]='h000001ec;  wr_data_rom[  123]='h000000c0;
    rd_cycle[  124] = 1'b0;  wr_cycle[  124] = 1'b1;  addr_rom[  124]='h000001f0;  wr_data_rom[  124]='h000009e4;
    rd_cycle[  125] = 1'b0;  wr_cycle[  125] = 1'b1;  addr_rom[  125]='h000001f4;  wr_data_rom[  125]='h00000760;
    rd_cycle[  126] = 1'b0;  wr_cycle[  126] = 1'b1;  addr_rom[  126]='h000001f8;  wr_data_rom[  126]='h00000b12;
    rd_cycle[  127] = 1'b0;  wr_cycle[  127] = 1'b1;  addr_rom[  127]='h000001fc;  wr_data_rom[  127]='h0000165b;
    rd_cycle[  128] = 1'b0;  wr_cycle[  128] = 1'b1;  addr_rom[  128]='h00000200;  wr_data_rom[  128]='h00000677;
    rd_cycle[  129] = 1'b0;  wr_cycle[  129] = 1'b1;  addr_rom[  129]='h00000204;  wr_data_rom[  129]='h00000de4;
    rd_cycle[  130] = 1'b0;  wr_cycle[  130] = 1'b1;  addr_rom[  130]='h00000208;  wr_data_rom[  130]='h000019d1;
    rd_cycle[  131] = 1'b0;  wr_cycle[  131] = 1'b1;  addr_rom[  131]='h0000020c;  wr_data_rom[  131]='h00001b0a;
    rd_cycle[  132] = 1'b0;  wr_cycle[  132] = 1'b1;  addr_rom[  132]='h00000210;  wr_data_rom[  132]='h000005a1;
    rd_cycle[  133] = 1'b0;  wr_cycle[  133] = 1'b1;  addr_rom[  133]='h00000214;  wr_data_rom[  133]='h000013d3;
    rd_cycle[  134] = 1'b0;  wr_cycle[  134] = 1'b1;  addr_rom[  134]='h00000218;  wr_data_rom[  134]='h00001f0a;
    rd_cycle[  135] = 1'b0;  wr_cycle[  135] = 1'b1;  addr_rom[  135]='h0000021c;  wr_data_rom[  135]='h00001ba2;
    rd_cycle[  136] = 1'b0;  wr_cycle[  136] = 1'b1;  addr_rom[  136]='h00000220;  wr_data_rom[  136]='h00000903;
    rd_cycle[  137] = 1'b0;  wr_cycle[  137] = 1'b1;  addr_rom[  137]='h00000224;  wr_data_rom[  137]='h00001458;
    rd_cycle[  138] = 1'b0;  wr_cycle[  138] = 1'b1;  addr_rom[  138]='h00000228;  wr_data_rom[  138]='h000016a5;
    rd_cycle[  139] = 1'b0;  wr_cycle[  139] = 1'b1;  addr_rom[  139]='h0000022c;  wr_data_rom[  139]='h00000a69;
    rd_cycle[  140] = 1'b0;  wr_cycle[  140] = 1'b1;  addr_rom[  140]='h00000230;  wr_data_rom[  140]='h0000127f;
    rd_cycle[  141] = 1'b0;  wr_cycle[  141] = 1'b1;  addr_rom[  141]='h00000234;  wr_data_rom[  141]='h0000052d;
    rd_cycle[  142] = 1'b0;  wr_cycle[  142] = 1'b1;  addr_rom[  142]='h00000238;  wr_data_rom[  142]='h00000fb3;
    rd_cycle[  143] = 1'b0;  wr_cycle[  143] = 1'b1;  addr_rom[  143]='h0000023c;  wr_data_rom[  143]='h000012a6;
    rd_cycle[  144] = 1'b0;  wr_cycle[  144] = 1'b1;  addr_rom[  144]='h00000240;  wr_data_rom[  144]='h00001a10;
    rd_cycle[  145] = 1'b0;  wr_cycle[  145] = 1'b1;  addr_rom[  145]='h00000244;  wr_data_rom[  145]='h00001631;
    rd_cycle[  146] = 1'b0;  wr_cycle[  146] = 1'b1;  addr_rom[  146]='h00000248;  wr_data_rom[  146]='h00001b8d;
    rd_cycle[  147] = 1'b0;  wr_cycle[  147] = 1'b1;  addr_rom[  147]='h0000024c;  wr_data_rom[  147]='h000002e2;
    rd_cycle[  148] = 1'b0;  wr_cycle[  148] = 1'b1;  addr_rom[  148]='h00000250;  wr_data_rom[  148]='h0000132c;
    rd_cycle[  149] = 1'b0;  wr_cycle[  149] = 1'b1;  addr_rom[  149]='h00000254;  wr_data_rom[  149]='h0000035d;
    rd_cycle[  150] = 1'b0;  wr_cycle[  150] = 1'b1;  addr_rom[  150]='h00000258;  wr_data_rom[  150]='h00001e21;
    rd_cycle[  151] = 1'b0;  wr_cycle[  151] = 1'b1;  addr_rom[  151]='h0000025c;  wr_data_rom[  151]='h00000e23;
    rd_cycle[  152] = 1'b0;  wr_cycle[  152] = 1'b1;  addr_rom[  152]='h00000260;  wr_data_rom[  152]='h000013d7;
    rd_cycle[  153] = 1'b0;  wr_cycle[  153] = 1'b1;  addr_rom[  153]='h00000264;  wr_data_rom[  153]='h00001d4a;
    rd_cycle[  154] = 1'b0;  wr_cycle[  154] = 1'b1;  addr_rom[  154]='h00000268;  wr_data_rom[  154]='h00000720;
    rd_cycle[  155] = 1'b0;  wr_cycle[  155] = 1'b1;  addr_rom[  155]='h0000026c;  wr_data_rom[  155]='h00000de1;
    rd_cycle[  156] = 1'b0;  wr_cycle[  156] = 1'b1;  addr_rom[  156]='h00000270;  wr_data_rom[  156]='h00000aa6;
    rd_cycle[  157] = 1'b0;  wr_cycle[  157] = 1'b1;  addr_rom[  157]='h00000274;  wr_data_rom[  157]='h0000040e;
    rd_cycle[  158] = 1'b0;  wr_cycle[  158] = 1'b1;  addr_rom[  158]='h00000278;  wr_data_rom[  158]='h00001dea;
    rd_cycle[  159] = 1'b0;  wr_cycle[  159] = 1'b1;  addr_rom[  159]='h0000027c;  wr_data_rom[  159]='h00001b78;
    rd_cycle[  160] = 1'b0;  wr_cycle[  160] = 1'b1;  addr_rom[  160]='h00000280;  wr_data_rom[  160]='h0000110c;
    rd_cycle[  161] = 1'b0;  wr_cycle[  161] = 1'b1;  addr_rom[  161]='h00000284;  wr_data_rom[  161]='h00000bf7;
    rd_cycle[  162] = 1'b0;  wr_cycle[  162] = 1'b1;  addr_rom[  162]='h00000288;  wr_data_rom[  162]='h0000140d;
    rd_cycle[  163] = 1'b0;  wr_cycle[  163] = 1'b1;  addr_rom[  163]='h0000028c;  wr_data_rom[  163]='h00001f2c;
    rd_cycle[  164] = 1'b0;  wr_cycle[  164] = 1'b1;  addr_rom[  164]='h00000290;  wr_data_rom[  164]='h00001648;
    rd_cycle[  165] = 1'b0;  wr_cycle[  165] = 1'b1;  addr_rom[  165]='h00000294;  wr_data_rom[  165]='h000010ea;
    rd_cycle[  166] = 1'b0;  wr_cycle[  166] = 1'b1;  addr_rom[  166]='h00000298;  wr_data_rom[  166]='h00000f4d;
    rd_cycle[  167] = 1'b0;  wr_cycle[  167] = 1'b1;  addr_rom[  167]='h0000029c;  wr_data_rom[  167]='h000011fc;
    rd_cycle[  168] = 1'b0;  wr_cycle[  168] = 1'b1;  addr_rom[  168]='h000002a0;  wr_data_rom[  168]='h00000ecd;
    rd_cycle[  169] = 1'b0;  wr_cycle[  169] = 1'b1;  addr_rom[  169]='h000002a4;  wr_data_rom[  169]='h000019f7;
    rd_cycle[  170] = 1'b0;  wr_cycle[  170] = 1'b1;  addr_rom[  170]='h000002a8;  wr_data_rom[  170]='h000013f9;
    rd_cycle[  171] = 1'b0;  wr_cycle[  171] = 1'b1;  addr_rom[  171]='h000002ac;  wr_data_rom[  171]='h000000b3;
    rd_cycle[  172] = 1'b0;  wr_cycle[  172] = 1'b1;  addr_rom[  172]='h000002b0;  wr_data_rom[  172]='h000001f8;
    rd_cycle[  173] = 1'b0;  wr_cycle[  173] = 1'b1;  addr_rom[  173]='h000002b4;  wr_data_rom[  173]='h00000263;
    rd_cycle[  174] = 1'b0;  wr_cycle[  174] = 1'b1;  addr_rom[  174]='h000002b8;  wr_data_rom[  174]='h00000a26;
    rd_cycle[  175] = 1'b0;  wr_cycle[  175] = 1'b1;  addr_rom[  175]='h000002bc;  wr_data_rom[  175]='h000014a1;
    rd_cycle[  176] = 1'b0;  wr_cycle[  176] = 1'b1;  addr_rom[  176]='h000002c0;  wr_data_rom[  176]='h00000fc8;
    rd_cycle[  177] = 1'b0;  wr_cycle[  177] = 1'b1;  addr_rom[  177]='h000002c4;  wr_data_rom[  177]='h0000010b;
    rd_cycle[  178] = 1'b0;  wr_cycle[  178] = 1'b1;  addr_rom[  178]='h000002c8;  wr_data_rom[  178]='h00000549;
    rd_cycle[  179] = 1'b0;  wr_cycle[  179] = 1'b1;  addr_rom[  179]='h000002cc;  wr_data_rom[  179]='h00000425;
    rd_cycle[  180] = 1'b0;  wr_cycle[  180] = 1'b1;  addr_rom[  180]='h000002d0;  wr_data_rom[  180]='h000014e3;
    rd_cycle[  181] = 1'b0;  wr_cycle[  181] = 1'b1;  addr_rom[  181]='h000002d4;  wr_data_rom[  181]='h00001f2c;
    rd_cycle[  182] = 1'b0;  wr_cycle[  182] = 1'b1;  addr_rom[  182]='h000002d8;  wr_data_rom[  182]='h0000051c;
    rd_cycle[  183] = 1'b0;  wr_cycle[  183] = 1'b1;  addr_rom[  183]='h000002dc;  wr_data_rom[  183]='h00000cb5;
    rd_cycle[  184] = 1'b0;  wr_cycle[  184] = 1'b1;  addr_rom[  184]='h000002e0;  wr_data_rom[  184]='h00000637;
    rd_cycle[  185] = 1'b0;  wr_cycle[  185] = 1'b1;  addr_rom[  185]='h000002e4;  wr_data_rom[  185]='h00000dc8;
    rd_cycle[  186] = 1'b0;  wr_cycle[  186] = 1'b1;  addr_rom[  186]='h000002e8;  wr_data_rom[  186]='h000015e4;
    rd_cycle[  187] = 1'b0;  wr_cycle[  187] = 1'b1;  addr_rom[  187]='h000002ec;  wr_data_rom[  187]='h00000681;
    rd_cycle[  188] = 1'b0;  wr_cycle[  188] = 1'b1;  addr_rom[  188]='h000002f0;  wr_data_rom[  188]='h0000015f;
    rd_cycle[  189] = 1'b0;  wr_cycle[  189] = 1'b1;  addr_rom[  189]='h000002f4;  wr_data_rom[  189]='h000011a4;
    rd_cycle[  190] = 1'b0;  wr_cycle[  190] = 1'b1;  addr_rom[  190]='h000002f8;  wr_data_rom[  190]='h000005c6;
    rd_cycle[  191] = 1'b0;  wr_cycle[  191] = 1'b1;  addr_rom[  191]='h000002fc;  wr_data_rom[  191]='h0000135c;
    rd_cycle[  192] = 1'b0;  wr_cycle[  192] = 1'b1;  addr_rom[  192]='h00000300;  wr_data_rom[  192]='h00000f0c;
    rd_cycle[  193] = 1'b0;  wr_cycle[  193] = 1'b1;  addr_rom[  193]='h00000304;  wr_data_rom[  193]='h00000174;
    rd_cycle[  194] = 1'b0;  wr_cycle[  194] = 1'b1;  addr_rom[  194]='h00000308;  wr_data_rom[  194]='h00001c34;
    rd_cycle[  195] = 1'b0;  wr_cycle[  195] = 1'b1;  addr_rom[  195]='h0000030c;  wr_data_rom[  195]='h00001c12;
    rd_cycle[  196] = 1'b0;  wr_cycle[  196] = 1'b1;  addr_rom[  196]='h00000310;  wr_data_rom[  196]='h000001e3;
    rd_cycle[  197] = 1'b0;  wr_cycle[  197] = 1'b1;  addr_rom[  197]='h00000314;  wr_data_rom[  197]='h00000255;
    rd_cycle[  198] = 1'b0;  wr_cycle[  198] = 1'b1;  addr_rom[  198]='h00000318;  wr_data_rom[  198]='h000001e7;
    rd_cycle[  199] = 1'b0;  wr_cycle[  199] = 1'b1;  addr_rom[  199]='h0000031c;  wr_data_rom[  199]='h00001433;
    rd_cycle[  200] = 1'b0;  wr_cycle[  200] = 1'b1;  addr_rom[  200]='h00000320;  wr_data_rom[  200]='h000017e4;
    rd_cycle[  201] = 1'b0;  wr_cycle[  201] = 1'b1;  addr_rom[  201]='h00000324;  wr_data_rom[  201]='h00000f1f;
    rd_cycle[  202] = 1'b0;  wr_cycle[  202] = 1'b1;  addr_rom[  202]='h00000328;  wr_data_rom[  202]='h00000367;
    rd_cycle[  203] = 1'b0;  wr_cycle[  203] = 1'b1;  addr_rom[  203]='h0000032c;  wr_data_rom[  203]='h0000155d;
    rd_cycle[  204] = 1'b0;  wr_cycle[  204] = 1'b1;  addr_rom[  204]='h00000330;  wr_data_rom[  204]='h000012e7;
    rd_cycle[  205] = 1'b0;  wr_cycle[  205] = 1'b1;  addr_rom[  205]='h00000334;  wr_data_rom[  205]='h000015f4;
    rd_cycle[  206] = 1'b0;  wr_cycle[  206] = 1'b1;  addr_rom[  206]='h00000338;  wr_data_rom[  206]='h00000a62;
    rd_cycle[  207] = 1'b0;  wr_cycle[  207] = 1'b1;  addr_rom[  207]='h0000033c;  wr_data_rom[  207]='h00000b4c;
    rd_cycle[  208] = 1'b0;  wr_cycle[  208] = 1'b1;  addr_rom[  208]='h00000340;  wr_data_rom[  208]='h000000ce;
    rd_cycle[  209] = 1'b0;  wr_cycle[  209] = 1'b1;  addr_rom[  209]='h00000344;  wr_data_rom[  209]='h000008c1;
    rd_cycle[  210] = 1'b0;  wr_cycle[  210] = 1'b1;  addr_rom[  210]='h00000348;  wr_data_rom[  210]='h00001c18;
    rd_cycle[  211] = 1'b0;  wr_cycle[  211] = 1'b1;  addr_rom[  211]='h0000034c;  wr_data_rom[  211]='h0000002b;
    rd_cycle[  212] = 1'b0;  wr_cycle[  212] = 1'b1;  addr_rom[  212]='h00000350;  wr_data_rom[  212]='h00000c4d;
    rd_cycle[  213] = 1'b0;  wr_cycle[  213] = 1'b1;  addr_rom[  213]='h00000354;  wr_data_rom[  213]='h00001b70;
    rd_cycle[  214] = 1'b0;  wr_cycle[  214] = 1'b1;  addr_rom[  214]='h00000358;  wr_data_rom[  214]='h0000016d;
    rd_cycle[  215] = 1'b0;  wr_cycle[  215] = 1'b1;  addr_rom[  215]='h0000035c;  wr_data_rom[  215]='h00001092;
    rd_cycle[  216] = 1'b0;  wr_cycle[  216] = 1'b1;  addr_rom[  216]='h00000360;  wr_data_rom[  216]='h000006d6;
    rd_cycle[  217] = 1'b0;  wr_cycle[  217] = 1'b1;  addr_rom[  217]='h00000364;  wr_data_rom[  217]='h00000872;
    rd_cycle[  218] = 1'b0;  wr_cycle[  218] = 1'b1;  addr_rom[  218]='h00000368;  wr_data_rom[  218]='h0000064a;
    rd_cycle[  219] = 1'b0;  wr_cycle[  219] = 1'b1;  addr_rom[  219]='h0000036c;  wr_data_rom[  219]='h00000bc3;
    rd_cycle[  220] = 1'b0;  wr_cycle[  220] = 1'b1;  addr_rom[  220]='h00000370;  wr_data_rom[  220]='h000013f4;
    rd_cycle[  221] = 1'b0;  wr_cycle[  221] = 1'b1;  addr_rom[  221]='h00000374;  wr_data_rom[  221]='h00000393;
    rd_cycle[  222] = 1'b0;  wr_cycle[  222] = 1'b1;  addr_rom[  222]='h00000378;  wr_data_rom[  222]='h00001c5e;
    rd_cycle[  223] = 1'b0;  wr_cycle[  223] = 1'b1;  addr_rom[  223]='h0000037c;  wr_data_rom[  223]='h00000362;
    rd_cycle[  224] = 1'b0;  wr_cycle[  224] = 1'b1;  addr_rom[  224]='h00000380;  wr_data_rom[  224]='h00001221;
    rd_cycle[  225] = 1'b0;  wr_cycle[  225] = 1'b1;  addr_rom[  225]='h00000384;  wr_data_rom[  225]='h00000eaa;
    rd_cycle[  226] = 1'b0;  wr_cycle[  226] = 1'b1;  addr_rom[  226]='h00000388;  wr_data_rom[  226]='h00001452;
    rd_cycle[  227] = 1'b0;  wr_cycle[  227] = 1'b1;  addr_rom[  227]='h0000038c;  wr_data_rom[  227]='h00001dbc;
    rd_cycle[  228] = 1'b0;  wr_cycle[  228] = 1'b1;  addr_rom[  228]='h00000390;  wr_data_rom[  228]='h00001c15;
    rd_cycle[  229] = 1'b0;  wr_cycle[  229] = 1'b1;  addr_rom[  229]='h00000394;  wr_data_rom[  229]='h00001262;
    rd_cycle[  230] = 1'b0;  wr_cycle[  230] = 1'b1;  addr_rom[  230]='h00000398;  wr_data_rom[  230]='h00001f38;
    rd_cycle[  231] = 1'b0;  wr_cycle[  231] = 1'b1;  addr_rom[  231]='h0000039c;  wr_data_rom[  231]='h00001082;
    rd_cycle[  232] = 1'b0;  wr_cycle[  232] = 1'b1;  addr_rom[  232]='h000003a0;  wr_data_rom[  232]='h00000c98;
    rd_cycle[  233] = 1'b0;  wr_cycle[  233] = 1'b1;  addr_rom[  233]='h000003a4;  wr_data_rom[  233]='h000008ca;
    rd_cycle[  234] = 1'b0;  wr_cycle[  234] = 1'b1;  addr_rom[  234]='h000003a8;  wr_data_rom[  234]='h00000407;
    rd_cycle[  235] = 1'b0;  wr_cycle[  235] = 1'b1;  addr_rom[  235]='h000003ac;  wr_data_rom[  235]='h000011fc;
    rd_cycle[  236] = 1'b0;  wr_cycle[  236] = 1'b1;  addr_rom[  236]='h000003b0;  wr_data_rom[  236]='h000017b6;
    rd_cycle[  237] = 1'b0;  wr_cycle[  237] = 1'b1;  addr_rom[  237]='h000003b4;  wr_data_rom[  237]='h000001a4;
    rd_cycle[  238] = 1'b0;  wr_cycle[  238] = 1'b1;  addr_rom[  238]='h000003b8;  wr_data_rom[  238]='h00001034;
    rd_cycle[  239] = 1'b0;  wr_cycle[  239] = 1'b1;  addr_rom[  239]='h000003bc;  wr_data_rom[  239]='h00001ee7;
    rd_cycle[  240] = 1'b0;  wr_cycle[  240] = 1'b1;  addr_rom[  240]='h000003c0;  wr_data_rom[  240]='h00000533;
    rd_cycle[  241] = 1'b0;  wr_cycle[  241] = 1'b1;  addr_rom[  241]='h000003c4;  wr_data_rom[  241]='h00001d56;
    rd_cycle[  242] = 1'b0;  wr_cycle[  242] = 1'b1;  addr_rom[  242]='h000003c8;  wr_data_rom[  242]='h000014f7;
    rd_cycle[  243] = 1'b0;  wr_cycle[  243] = 1'b1;  addr_rom[  243]='h000003cc;  wr_data_rom[  243]='h0000180c;
    rd_cycle[  244] = 1'b0;  wr_cycle[  244] = 1'b1;  addr_rom[  244]='h000003d0;  wr_data_rom[  244]='h00000f78;
    rd_cycle[  245] = 1'b0;  wr_cycle[  245] = 1'b1;  addr_rom[  245]='h000003d4;  wr_data_rom[  245]='h00000f83;
    rd_cycle[  246] = 1'b0;  wr_cycle[  246] = 1'b1;  addr_rom[  246]='h000003d8;  wr_data_rom[  246]='h00000735;
    rd_cycle[  247] = 1'b0;  wr_cycle[  247] = 1'b1;  addr_rom[  247]='h000003dc;  wr_data_rom[  247]='h0000094e;
    rd_cycle[  248] = 1'b0;  wr_cycle[  248] = 1'b1;  addr_rom[  248]='h000003e0;  wr_data_rom[  248]='h00000bce;
    rd_cycle[  249] = 1'b0;  wr_cycle[  249] = 1'b1;  addr_rom[  249]='h000003e4;  wr_data_rom[  249]='h000019aa;
    rd_cycle[  250] = 1'b0;  wr_cycle[  250] = 1'b1;  addr_rom[  250]='h000003e8;  wr_data_rom[  250]='h00001846;
    rd_cycle[  251] = 1'b0;  wr_cycle[  251] = 1'b1;  addr_rom[  251]='h000003ec;  wr_data_rom[  251]='h00001178;
    rd_cycle[  252] = 1'b0;  wr_cycle[  252] = 1'b1;  addr_rom[  252]='h000003f0;  wr_data_rom[  252]='h000010fd;
    rd_cycle[  253] = 1'b0;  wr_cycle[  253] = 1'b1;  addr_rom[  253]='h000003f4;  wr_data_rom[  253]='h00001954;
    rd_cycle[  254] = 1'b0;  wr_cycle[  254] = 1'b1;  addr_rom[  254]='h000003f8;  wr_data_rom[  254]='h0000070a;
    rd_cycle[  255] = 1'b0;  wr_cycle[  255] = 1'b1;  addr_rom[  255]='h000003fc;  wr_data_rom[  255]='h00000fe8;
    rd_cycle[  256] = 1'b0;  wr_cycle[  256] = 1'b1;  addr_rom[  256]='h00000400;  wr_data_rom[  256]='h00000e1c;
    rd_cycle[  257] = 1'b0;  wr_cycle[  257] = 1'b1;  addr_rom[  257]='h00000404;  wr_data_rom[  257]='h00001e65;
    rd_cycle[  258] = 1'b0;  wr_cycle[  258] = 1'b1;  addr_rom[  258]='h00000408;  wr_data_rom[  258]='h00001bd0;
    rd_cycle[  259] = 1'b0;  wr_cycle[  259] = 1'b1;  addr_rom[  259]='h0000040c;  wr_data_rom[  259]='h00001bcd;
    rd_cycle[  260] = 1'b0;  wr_cycle[  260] = 1'b1;  addr_rom[  260]='h00000410;  wr_data_rom[  260]='h00000a51;
    rd_cycle[  261] = 1'b0;  wr_cycle[  261] = 1'b1;  addr_rom[  261]='h00000414;  wr_data_rom[  261]='h00000e9a;
    rd_cycle[  262] = 1'b0;  wr_cycle[  262] = 1'b1;  addr_rom[  262]='h00000418;  wr_data_rom[  262]='h000003b3;
    rd_cycle[  263] = 1'b0;  wr_cycle[  263] = 1'b1;  addr_rom[  263]='h0000041c;  wr_data_rom[  263]='h00000c8c;
    rd_cycle[  264] = 1'b0;  wr_cycle[  264] = 1'b1;  addr_rom[  264]='h00000420;  wr_data_rom[  264]='h000018b7;
    rd_cycle[  265] = 1'b0;  wr_cycle[  265] = 1'b1;  addr_rom[  265]='h00000424;  wr_data_rom[  265]='h00000f8d;
    rd_cycle[  266] = 1'b0;  wr_cycle[  266] = 1'b1;  addr_rom[  266]='h00000428;  wr_data_rom[  266]='h00001f0d;
    rd_cycle[  267] = 1'b0;  wr_cycle[  267] = 1'b1;  addr_rom[  267]='h0000042c;  wr_data_rom[  267]='h0000115e;
    rd_cycle[  268] = 1'b0;  wr_cycle[  268] = 1'b1;  addr_rom[  268]='h00000430;  wr_data_rom[  268]='h00001bfe;
    rd_cycle[  269] = 1'b0;  wr_cycle[  269] = 1'b1;  addr_rom[  269]='h00000434;  wr_data_rom[  269]='h00000db1;
    rd_cycle[  270] = 1'b0;  wr_cycle[  270] = 1'b1;  addr_rom[  270]='h00000438;  wr_data_rom[  270]='h00000e07;
    rd_cycle[  271] = 1'b0;  wr_cycle[  271] = 1'b1;  addr_rom[  271]='h0000043c;  wr_data_rom[  271]='h00000109;
    rd_cycle[  272] = 1'b0;  wr_cycle[  272] = 1'b1;  addr_rom[  272]='h00000440;  wr_data_rom[  272]='h0000193f;
    rd_cycle[  273] = 1'b0;  wr_cycle[  273] = 1'b1;  addr_rom[  273]='h00000444;  wr_data_rom[  273]='h00000a55;
    rd_cycle[  274] = 1'b0;  wr_cycle[  274] = 1'b1;  addr_rom[  274]='h00000448;  wr_data_rom[  274]='h00000fbd;
    rd_cycle[  275] = 1'b0;  wr_cycle[  275] = 1'b1;  addr_rom[  275]='h0000044c;  wr_data_rom[  275]='h0000114d;
    rd_cycle[  276] = 1'b0;  wr_cycle[  276] = 1'b1;  addr_rom[  276]='h00000450;  wr_data_rom[  276]='h00000b69;
    rd_cycle[  277] = 1'b0;  wr_cycle[  277] = 1'b1;  addr_rom[  277]='h00000454;  wr_data_rom[  277]='h00001a47;
    rd_cycle[  278] = 1'b0;  wr_cycle[  278] = 1'b1;  addr_rom[  278]='h00000458;  wr_data_rom[  278]='h00001d41;
    rd_cycle[  279] = 1'b0;  wr_cycle[  279] = 1'b1;  addr_rom[  279]='h0000045c;  wr_data_rom[  279]='h000017cf;
    rd_cycle[  280] = 1'b0;  wr_cycle[  280] = 1'b1;  addr_rom[  280]='h00000460;  wr_data_rom[  280]='h000006ad;
    rd_cycle[  281] = 1'b0;  wr_cycle[  281] = 1'b1;  addr_rom[  281]='h00000464;  wr_data_rom[  281]='h0000066d;
    rd_cycle[  282] = 1'b0;  wr_cycle[  282] = 1'b1;  addr_rom[  282]='h00000468;  wr_data_rom[  282]='h0000014e;
    rd_cycle[  283] = 1'b0;  wr_cycle[  283] = 1'b1;  addr_rom[  283]='h0000046c;  wr_data_rom[  283]='h00000656;
    rd_cycle[  284] = 1'b0;  wr_cycle[  284] = 1'b1;  addr_rom[  284]='h00000470;  wr_data_rom[  284]='h00000e71;
    rd_cycle[  285] = 1'b0;  wr_cycle[  285] = 1'b1;  addr_rom[  285]='h00000474;  wr_data_rom[  285]='h0000089f;
    rd_cycle[  286] = 1'b0;  wr_cycle[  286] = 1'b1;  addr_rom[  286]='h00000478;  wr_data_rom[  286]='h00001f1e;
    rd_cycle[  287] = 1'b0;  wr_cycle[  287] = 1'b1;  addr_rom[  287]='h0000047c;  wr_data_rom[  287]='h000014c8;
    rd_cycle[  288] = 1'b0;  wr_cycle[  288] = 1'b1;  addr_rom[  288]='h00000480;  wr_data_rom[  288]='h00001a63;
    rd_cycle[  289] = 1'b0;  wr_cycle[  289] = 1'b1;  addr_rom[  289]='h00000484;  wr_data_rom[  289]='h00001d12;
    rd_cycle[  290] = 1'b0;  wr_cycle[  290] = 1'b1;  addr_rom[  290]='h00000488;  wr_data_rom[  290]='h00001eb2;
    rd_cycle[  291] = 1'b0;  wr_cycle[  291] = 1'b1;  addr_rom[  291]='h0000048c;  wr_data_rom[  291]='h0000183c;
    rd_cycle[  292] = 1'b0;  wr_cycle[  292] = 1'b1;  addr_rom[  292]='h00000490;  wr_data_rom[  292]='h00001d85;
    rd_cycle[  293] = 1'b0;  wr_cycle[  293] = 1'b1;  addr_rom[  293]='h00000494;  wr_data_rom[  293]='h000010ce;
    rd_cycle[  294] = 1'b0;  wr_cycle[  294] = 1'b1;  addr_rom[  294]='h00000498;  wr_data_rom[  294]='h0000022f;
    rd_cycle[  295] = 1'b0;  wr_cycle[  295] = 1'b1;  addr_rom[  295]='h0000049c;  wr_data_rom[  295]='h0000041d;
    rd_cycle[  296] = 1'b0;  wr_cycle[  296] = 1'b1;  addr_rom[  296]='h000004a0;  wr_data_rom[  296]='h00000541;
    rd_cycle[  297] = 1'b0;  wr_cycle[  297] = 1'b1;  addr_rom[  297]='h000004a4;  wr_data_rom[  297]='h0000099b;
    rd_cycle[  298] = 1'b0;  wr_cycle[  298] = 1'b1;  addr_rom[  298]='h000004a8;  wr_data_rom[  298]='h00000dde;
    rd_cycle[  299] = 1'b0;  wr_cycle[  299] = 1'b1;  addr_rom[  299]='h000004ac;  wr_data_rom[  299]='h00000dad;
    rd_cycle[  300] = 1'b0;  wr_cycle[  300] = 1'b1;  addr_rom[  300]='h000004b0;  wr_data_rom[  300]='h0000027e;
    rd_cycle[  301] = 1'b0;  wr_cycle[  301] = 1'b1;  addr_rom[  301]='h000004b4;  wr_data_rom[  301]='h00000f7f;
    rd_cycle[  302] = 1'b0;  wr_cycle[  302] = 1'b1;  addr_rom[  302]='h000004b8;  wr_data_rom[  302]='h00000384;
    rd_cycle[  303] = 1'b0;  wr_cycle[  303] = 1'b1;  addr_rom[  303]='h000004bc;  wr_data_rom[  303]='h00001185;
    rd_cycle[  304] = 1'b0;  wr_cycle[  304] = 1'b1;  addr_rom[  304]='h000004c0;  wr_data_rom[  304]='h0000051c;
    rd_cycle[  305] = 1'b0;  wr_cycle[  305] = 1'b1;  addr_rom[  305]='h000004c4;  wr_data_rom[  305]='h00000cf4;
    rd_cycle[  306] = 1'b0;  wr_cycle[  306] = 1'b1;  addr_rom[  306]='h000004c8;  wr_data_rom[  306]='h00000bfd;
    rd_cycle[  307] = 1'b0;  wr_cycle[  307] = 1'b1;  addr_rom[  307]='h000004cc;  wr_data_rom[  307]='h00001b6b;
    rd_cycle[  308] = 1'b0;  wr_cycle[  308] = 1'b1;  addr_rom[  308]='h000004d0;  wr_data_rom[  308]='h00001a69;
    rd_cycle[  309] = 1'b0;  wr_cycle[  309] = 1'b1;  addr_rom[  309]='h000004d4;  wr_data_rom[  309]='h000013b0;
    rd_cycle[  310] = 1'b0;  wr_cycle[  310] = 1'b1;  addr_rom[  310]='h000004d8;  wr_data_rom[  310]='h000007ee;
    rd_cycle[  311] = 1'b0;  wr_cycle[  311] = 1'b1;  addr_rom[  311]='h000004dc;  wr_data_rom[  311]='h00000488;
    rd_cycle[  312] = 1'b0;  wr_cycle[  312] = 1'b1;  addr_rom[  312]='h000004e0;  wr_data_rom[  312]='h0000167b;
    rd_cycle[  313] = 1'b0;  wr_cycle[  313] = 1'b1;  addr_rom[  313]='h000004e4;  wr_data_rom[  313]='h00001dbb;
    rd_cycle[  314] = 1'b0;  wr_cycle[  314] = 1'b1;  addr_rom[  314]='h000004e8;  wr_data_rom[  314]='h00000396;
    rd_cycle[  315] = 1'b0;  wr_cycle[  315] = 1'b1;  addr_rom[  315]='h000004ec;  wr_data_rom[  315]='h0000033c;
    rd_cycle[  316] = 1'b0;  wr_cycle[  316] = 1'b1;  addr_rom[  316]='h000004f0;  wr_data_rom[  316]='h000001d9;
    rd_cycle[  317] = 1'b0;  wr_cycle[  317] = 1'b1;  addr_rom[  317]='h000004f4;  wr_data_rom[  317]='h000013b9;
    rd_cycle[  318] = 1'b0;  wr_cycle[  318] = 1'b1;  addr_rom[  318]='h000004f8;  wr_data_rom[  318]='h000012ef;
    rd_cycle[  319] = 1'b0;  wr_cycle[  319] = 1'b1;  addr_rom[  319]='h000004fc;  wr_data_rom[  319]='h00000fac;
    rd_cycle[  320] = 1'b0;  wr_cycle[  320] = 1'b1;  addr_rom[  320]='h00000500;  wr_data_rom[  320]='h0000002a;
    rd_cycle[  321] = 1'b0;  wr_cycle[  321] = 1'b1;  addr_rom[  321]='h00000504;  wr_data_rom[  321]='h00000c9e;
    rd_cycle[  322] = 1'b0;  wr_cycle[  322] = 1'b1;  addr_rom[  322]='h00000508;  wr_data_rom[  322]='h00000d7a;
    rd_cycle[  323] = 1'b0;  wr_cycle[  323] = 1'b1;  addr_rom[  323]='h0000050c;  wr_data_rom[  323]='h00000832;
    rd_cycle[  324] = 1'b0;  wr_cycle[  324] = 1'b1;  addr_rom[  324]='h00000510;  wr_data_rom[  324]='h00000977;
    rd_cycle[  325] = 1'b0;  wr_cycle[  325] = 1'b1;  addr_rom[  325]='h00000514;  wr_data_rom[  325]='h00001b15;
    rd_cycle[  326] = 1'b0;  wr_cycle[  326] = 1'b1;  addr_rom[  326]='h00000518;  wr_data_rom[  326]='h00000f72;
    rd_cycle[  327] = 1'b0;  wr_cycle[  327] = 1'b1;  addr_rom[  327]='h0000051c;  wr_data_rom[  327]='h0000184f;
    rd_cycle[  328] = 1'b0;  wr_cycle[  328] = 1'b1;  addr_rom[  328]='h00000520;  wr_data_rom[  328]='h000008f6;
    rd_cycle[  329] = 1'b0;  wr_cycle[  329] = 1'b1;  addr_rom[  329]='h00000524;  wr_data_rom[  329]='h0000070f;
    rd_cycle[  330] = 1'b0;  wr_cycle[  330] = 1'b1;  addr_rom[  330]='h00000528;  wr_data_rom[  330]='h00000ef8;
    rd_cycle[  331] = 1'b0;  wr_cycle[  331] = 1'b1;  addr_rom[  331]='h0000052c;  wr_data_rom[  331]='h00001756;
    rd_cycle[  332] = 1'b0;  wr_cycle[  332] = 1'b1;  addr_rom[  332]='h00000530;  wr_data_rom[  332]='h000008bc;
    rd_cycle[  333] = 1'b0;  wr_cycle[  333] = 1'b1;  addr_rom[  333]='h00000534;  wr_data_rom[  333]='h00000c2e;
    rd_cycle[  334] = 1'b0;  wr_cycle[  334] = 1'b1;  addr_rom[  334]='h00000538;  wr_data_rom[  334]='h00001377;
    rd_cycle[  335] = 1'b0;  wr_cycle[  335] = 1'b1;  addr_rom[  335]='h0000053c;  wr_data_rom[  335]='h0000135c;
    rd_cycle[  336] = 1'b0;  wr_cycle[  336] = 1'b1;  addr_rom[  336]='h00000540;  wr_data_rom[  336]='h00001cc4;
    rd_cycle[  337] = 1'b0;  wr_cycle[  337] = 1'b1;  addr_rom[  337]='h00000544;  wr_data_rom[  337]='h00001943;
    rd_cycle[  338] = 1'b0;  wr_cycle[  338] = 1'b1;  addr_rom[  338]='h00000548;  wr_data_rom[  338]='h00000510;
    rd_cycle[  339] = 1'b0;  wr_cycle[  339] = 1'b1;  addr_rom[  339]='h0000054c;  wr_data_rom[  339]='h00000957;
    rd_cycle[  340] = 1'b0;  wr_cycle[  340] = 1'b1;  addr_rom[  340]='h00000550;  wr_data_rom[  340]='h0000147e;
    rd_cycle[  341] = 1'b0;  wr_cycle[  341] = 1'b1;  addr_rom[  341]='h00000554;  wr_data_rom[  341]='h000016e6;
    rd_cycle[  342] = 1'b0;  wr_cycle[  342] = 1'b1;  addr_rom[  342]='h00000558;  wr_data_rom[  342]='h00001b43;
    rd_cycle[  343] = 1'b0;  wr_cycle[  343] = 1'b1;  addr_rom[  343]='h0000055c;  wr_data_rom[  343]='h0000124f;
    rd_cycle[  344] = 1'b0;  wr_cycle[  344] = 1'b1;  addr_rom[  344]='h00000560;  wr_data_rom[  344]='h0000016f;
    rd_cycle[  345] = 1'b0;  wr_cycle[  345] = 1'b1;  addr_rom[  345]='h00000564;  wr_data_rom[  345]='h0000104e;
    rd_cycle[  346] = 1'b0;  wr_cycle[  346] = 1'b1;  addr_rom[  346]='h00000568;  wr_data_rom[  346]='h000002c0;
    rd_cycle[  347] = 1'b0;  wr_cycle[  347] = 1'b1;  addr_rom[  347]='h0000056c;  wr_data_rom[  347]='h0000099c;
    rd_cycle[  348] = 1'b0;  wr_cycle[  348] = 1'b1;  addr_rom[  348]='h00000570;  wr_data_rom[  348]='h00001e3e;
    rd_cycle[  349] = 1'b0;  wr_cycle[  349] = 1'b1;  addr_rom[  349]='h00000574;  wr_data_rom[  349]='h00001a77;
    rd_cycle[  350] = 1'b0;  wr_cycle[  350] = 1'b1;  addr_rom[  350]='h00000578;  wr_data_rom[  350]='h000002e2;
    rd_cycle[  351] = 1'b0;  wr_cycle[  351] = 1'b1;  addr_rom[  351]='h0000057c;  wr_data_rom[  351]='h000017bd;
    rd_cycle[  352] = 1'b0;  wr_cycle[  352] = 1'b1;  addr_rom[  352]='h00000580;  wr_data_rom[  352]='h00000572;
    rd_cycle[  353] = 1'b0;  wr_cycle[  353] = 1'b1;  addr_rom[  353]='h00000584;  wr_data_rom[  353]='h000003f5;
    rd_cycle[  354] = 1'b0;  wr_cycle[  354] = 1'b1;  addr_rom[  354]='h00000588;  wr_data_rom[  354]='h00000a34;
    rd_cycle[  355] = 1'b0;  wr_cycle[  355] = 1'b1;  addr_rom[  355]='h0000058c;  wr_data_rom[  355]='h000015f6;
    rd_cycle[  356] = 1'b0;  wr_cycle[  356] = 1'b1;  addr_rom[  356]='h00000590;  wr_data_rom[  356]='h00000ad5;
    rd_cycle[  357] = 1'b0;  wr_cycle[  357] = 1'b1;  addr_rom[  357]='h00000594;  wr_data_rom[  357]='h000006fd;
    rd_cycle[  358] = 1'b0;  wr_cycle[  358] = 1'b1;  addr_rom[  358]='h00000598;  wr_data_rom[  358]='h00001049;
    rd_cycle[  359] = 1'b0;  wr_cycle[  359] = 1'b1;  addr_rom[  359]='h0000059c;  wr_data_rom[  359]='h000019e8;
    rd_cycle[  360] = 1'b0;  wr_cycle[  360] = 1'b1;  addr_rom[  360]='h000005a0;  wr_data_rom[  360]='h00000964;
    rd_cycle[  361] = 1'b0;  wr_cycle[  361] = 1'b1;  addr_rom[  361]='h000005a4;  wr_data_rom[  361]='h000006a5;
    rd_cycle[  362] = 1'b0;  wr_cycle[  362] = 1'b1;  addr_rom[  362]='h000005a8;  wr_data_rom[  362]='h000017a9;
    rd_cycle[  363] = 1'b0;  wr_cycle[  363] = 1'b1;  addr_rom[  363]='h000005ac;  wr_data_rom[  363]='h0000075a;
    rd_cycle[  364] = 1'b0;  wr_cycle[  364] = 1'b1;  addr_rom[  364]='h000005b0;  wr_data_rom[  364]='h00001048;
    rd_cycle[  365] = 1'b0;  wr_cycle[  365] = 1'b1;  addr_rom[  365]='h000005b4;  wr_data_rom[  365]='h00000e5d;
    rd_cycle[  366] = 1'b0;  wr_cycle[  366] = 1'b1;  addr_rom[  366]='h000005b8;  wr_data_rom[  366]='h0000116b;
    rd_cycle[  367] = 1'b0;  wr_cycle[  367] = 1'b1;  addr_rom[  367]='h000005bc;  wr_data_rom[  367]='h00001e01;
    rd_cycle[  368] = 1'b0;  wr_cycle[  368] = 1'b1;  addr_rom[  368]='h000005c0;  wr_data_rom[  368]='h00001e46;
    rd_cycle[  369] = 1'b0;  wr_cycle[  369] = 1'b1;  addr_rom[  369]='h000005c4;  wr_data_rom[  369]='h000002bf;
    rd_cycle[  370] = 1'b0;  wr_cycle[  370] = 1'b1;  addr_rom[  370]='h000005c8;  wr_data_rom[  370]='h00000a15;
    rd_cycle[  371] = 1'b0;  wr_cycle[  371] = 1'b1;  addr_rom[  371]='h000005cc;  wr_data_rom[  371]='h00000cfd;
    rd_cycle[  372] = 1'b0;  wr_cycle[  372] = 1'b1;  addr_rom[  372]='h000005d0;  wr_data_rom[  372]='h000018b9;
    rd_cycle[  373] = 1'b0;  wr_cycle[  373] = 1'b1;  addr_rom[  373]='h000005d4;  wr_data_rom[  373]='h00000ee4;
    rd_cycle[  374] = 1'b0;  wr_cycle[  374] = 1'b1;  addr_rom[  374]='h000005d8;  wr_data_rom[  374]='h000019bd;
    rd_cycle[  375] = 1'b0;  wr_cycle[  375] = 1'b1;  addr_rom[  375]='h000005dc;  wr_data_rom[  375]='h0000149c;
    rd_cycle[  376] = 1'b0;  wr_cycle[  376] = 1'b1;  addr_rom[  376]='h000005e0;  wr_data_rom[  376]='h000005d5;
    rd_cycle[  377] = 1'b0;  wr_cycle[  377] = 1'b1;  addr_rom[  377]='h000005e4;  wr_data_rom[  377]='h0000100b;
    rd_cycle[  378] = 1'b0;  wr_cycle[  378] = 1'b1;  addr_rom[  378]='h000005e8;  wr_data_rom[  378]='h00001d8a;
    rd_cycle[  379] = 1'b0;  wr_cycle[  379] = 1'b1;  addr_rom[  379]='h000005ec;  wr_data_rom[  379]='h00001ea8;
    rd_cycle[  380] = 1'b0;  wr_cycle[  380] = 1'b1;  addr_rom[  380]='h000005f0;  wr_data_rom[  380]='h00001c34;
    rd_cycle[  381] = 1'b0;  wr_cycle[  381] = 1'b1;  addr_rom[  381]='h000005f4;  wr_data_rom[  381]='h00000119;
    rd_cycle[  382] = 1'b0;  wr_cycle[  382] = 1'b1;  addr_rom[  382]='h000005f8;  wr_data_rom[  382]='h00001696;
    rd_cycle[  383] = 1'b0;  wr_cycle[  383] = 1'b1;  addr_rom[  383]='h000005fc;  wr_data_rom[  383]='h0000016d;
    rd_cycle[  384] = 1'b0;  wr_cycle[  384] = 1'b1;  addr_rom[  384]='h00000600;  wr_data_rom[  384]='h000011e9;
    rd_cycle[  385] = 1'b0;  wr_cycle[  385] = 1'b1;  addr_rom[  385]='h00000604;  wr_data_rom[  385]='h00000d08;
    rd_cycle[  386] = 1'b0;  wr_cycle[  386] = 1'b1;  addr_rom[  386]='h00000608;  wr_data_rom[  386]='h0000166f;
    rd_cycle[  387] = 1'b0;  wr_cycle[  387] = 1'b1;  addr_rom[  387]='h0000060c;  wr_data_rom[  387]='h00001e0b;
    rd_cycle[  388] = 1'b0;  wr_cycle[  388] = 1'b1;  addr_rom[  388]='h00000610;  wr_data_rom[  388]='h00001cc8;
    rd_cycle[  389] = 1'b0;  wr_cycle[  389] = 1'b1;  addr_rom[  389]='h00000614;  wr_data_rom[  389]='h00000dda;
    rd_cycle[  390] = 1'b0;  wr_cycle[  390] = 1'b1;  addr_rom[  390]='h00000618;  wr_data_rom[  390]='h00001ce0;
    rd_cycle[  391] = 1'b0;  wr_cycle[  391] = 1'b1;  addr_rom[  391]='h0000061c;  wr_data_rom[  391]='h00001915;
    rd_cycle[  392] = 1'b0;  wr_cycle[  392] = 1'b1;  addr_rom[  392]='h00000620;  wr_data_rom[  392]='h00001c42;
    rd_cycle[  393] = 1'b0;  wr_cycle[  393] = 1'b1;  addr_rom[  393]='h00000624;  wr_data_rom[  393]='h000002ee;
    rd_cycle[  394] = 1'b0;  wr_cycle[  394] = 1'b1;  addr_rom[  394]='h00000628;  wr_data_rom[  394]='h00000c7e;
    rd_cycle[  395] = 1'b0;  wr_cycle[  395] = 1'b1;  addr_rom[  395]='h0000062c;  wr_data_rom[  395]='h00000b94;
    rd_cycle[  396] = 1'b0;  wr_cycle[  396] = 1'b1;  addr_rom[  396]='h00000630;  wr_data_rom[  396]='h00001936;
    rd_cycle[  397] = 1'b0;  wr_cycle[  397] = 1'b1;  addr_rom[  397]='h00000634;  wr_data_rom[  397]='h00001e78;
    rd_cycle[  398] = 1'b0;  wr_cycle[  398] = 1'b1;  addr_rom[  398]='h00000638;  wr_data_rom[  398]='h00001b76;
    rd_cycle[  399] = 1'b0;  wr_cycle[  399] = 1'b1;  addr_rom[  399]='h0000063c;  wr_data_rom[  399]='h00001875;
    rd_cycle[  400] = 1'b0;  wr_cycle[  400] = 1'b1;  addr_rom[  400]='h00000640;  wr_data_rom[  400]='h00000544;
    rd_cycle[  401] = 1'b0;  wr_cycle[  401] = 1'b1;  addr_rom[  401]='h00000644;  wr_data_rom[  401]='h00000331;
    rd_cycle[  402] = 1'b0;  wr_cycle[  402] = 1'b1;  addr_rom[  402]='h00000648;  wr_data_rom[  402]='h000011c5;
    rd_cycle[  403] = 1'b0;  wr_cycle[  403] = 1'b1;  addr_rom[  403]='h0000064c;  wr_data_rom[  403]='h0000009a;
    rd_cycle[  404] = 1'b0;  wr_cycle[  404] = 1'b1;  addr_rom[  404]='h00000650;  wr_data_rom[  404]='h00000c53;
    rd_cycle[  405] = 1'b0;  wr_cycle[  405] = 1'b1;  addr_rom[  405]='h00000654;  wr_data_rom[  405]='h000009ba;
    rd_cycle[  406] = 1'b0;  wr_cycle[  406] = 1'b1;  addr_rom[  406]='h00000658;  wr_data_rom[  406]='h0000141f;
    rd_cycle[  407] = 1'b0;  wr_cycle[  407] = 1'b1;  addr_rom[  407]='h0000065c;  wr_data_rom[  407]='h00000f22;
    rd_cycle[  408] = 1'b0;  wr_cycle[  408] = 1'b1;  addr_rom[  408]='h00000660;  wr_data_rom[  408]='h00001510;
    rd_cycle[  409] = 1'b0;  wr_cycle[  409] = 1'b1;  addr_rom[  409]='h00000664;  wr_data_rom[  409]='h00000e17;
    rd_cycle[  410] = 1'b0;  wr_cycle[  410] = 1'b1;  addr_rom[  410]='h00000668;  wr_data_rom[  410]='h000019c8;
    rd_cycle[  411] = 1'b0;  wr_cycle[  411] = 1'b1;  addr_rom[  411]='h0000066c;  wr_data_rom[  411]='h000004a4;
    rd_cycle[  412] = 1'b0;  wr_cycle[  412] = 1'b1;  addr_rom[  412]='h00000670;  wr_data_rom[  412]='h000019b5;
    rd_cycle[  413] = 1'b0;  wr_cycle[  413] = 1'b1;  addr_rom[  413]='h00000674;  wr_data_rom[  413]='h00001b6f;
    rd_cycle[  414] = 1'b0;  wr_cycle[  414] = 1'b1;  addr_rom[  414]='h00000678;  wr_data_rom[  414]='h000015dc;
    rd_cycle[  415] = 1'b0;  wr_cycle[  415] = 1'b1;  addr_rom[  415]='h0000067c;  wr_data_rom[  415]='h00000c42;
    rd_cycle[  416] = 1'b0;  wr_cycle[  416] = 1'b1;  addr_rom[  416]='h00000680;  wr_data_rom[  416]='h00000480;
    rd_cycle[  417] = 1'b0;  wr_cycle[  417] = 1'b1;  addr_rom[  417]='h00000684;  wr_data_rom[  417]='h00000e2b;
    rd_cycle[  418] = 1'b0;  wr_cycle[  418] = 1'b1;  addr_rom[  418]='h00000688;  wr_data_rom[  418]='h000010af;
    rd_cycle[  419] = 1'b0;  wr_cycle[  419] = 1'b1;  addr_rom[  419]='h0000068c;  wr_data_rom[  419]='h0000029a;
    rd_cycle[  420] = 1'b0;  wr_cycle[  420] = 1'b1;  addr_rom[  420]='h00000690;  wr_data_rom[  420]='h00000b92;
    rd_cycle[  421] = 1'b0;  wr_cycle[  421] = 1'b1;  addr_rom[  421]='h00000694;  wr_data_rom[  421]='h00001dff;
    rd_cycle[  422] = 1'b0;  wr_cycle[  422] = 1'b1;  addr_rom[  422]='h00000698;  wr_data_rom[  422]='h000013ef;
    rd_cycle[  423] = 1'b0;  wr_cycle[  423] = 1'b1;  addr_rom[  423]='h0000069c;  wr_data_rom[  423]='h000006b3;
    rd_cycle[  424] = 1'b0;  wr_cycle[  424] = 1'b1;  addr_rom[  424]='h000006a0;  wr_data_rom[  424]='h000009e8;
    rd_cycle[  425] = 1'b0;  wr_cycle[  425] = 1'b1;  addr_rom[  425]='h000006a4;  wr_data_rom[  425]='h00001bcc;
    rd_cycle[  426] = 1'b0;  wr_cycle[  426] = 1'b1;  addr_rom[  426]='h000006a8;  wr_data_rom[  426]='h00001cdf;
    rd_cycle[  427] = 1'b0;  wr_cycle[  427] = 1'b1;  addr_rom[  427]='h000006ac;  wr_data_rom[  427]='h00001e04;
    rd_cycle[  428] = 1'b0;  wr_cycle[  428] = 1'b1;  addr_rom[  428]='h000006b0;  wr_data_rom[  428]='h000015ff;
    rd_cycle[  429] = 1'b0;  wr_cycle[  429] = 1'b1;  addr_rom[  429]='h000006b4;  wr_data_rom[  429]='h00001ad3;
    rd_cycle[  430] = 1'b0;  wr_cycle[  430] = 1'b1;  addr_rom[  430]='h000006b8;  wr_data_rom[  430]='h00000472;
    rd_cycle[  431] = 1'b0;  wr_cycle[  431] = 1'b1;  addr_rom[  431]='h000006bc;  wr_data_rom[  431]='h000008a8;
    rd_cycle[  432] = 1'b0;  wr_cycle[  432] = 1'b1;  addr_rom[  432]='h000006c0;  wr_data_rom[  432]='h0000154c;
    rd_cycle[  433] = 1'b0;  wr_cycle[  433] = 1'b1;  addr_rom[  433]='h000006c4;  wr_data_rom[  433]='h000001bc;
    rd_cycle[  434] = 1'b0;  wr_cycle[  434] = 1'b1;  addr_rom[  434]='h000006c8;  wr_data_rom[  434]='h000004ac;
    rd_cycle[  435] = 1'b0;  wr_cycle[  435] = 1'b1;  addr_rom[  435]='h000006cc;  wr_data_rom[  435]='h00000a04;
    rd_cycle[  436] = 1'b0;  wr_cycle[  436] = 1'b1;  addr_rom[  436]='h000006d0;  wr_data_rom[  436]='h00000266;
    rd_cycle[  437] = 1'b0;  wr_cycle[  437] = 1'b1;  addr_rom[  437]='h000006d4;  wr_data_rom[  437]='h000009a9;
    rd_cycle[  438] = 1'b0;  wr_cycle[  438] = 1'b1;  addr_rom[  438]='h000006d8;  wr_data_rom[  438]='h00000eb3;
    rd_cycle[  439] = 1'b0;  wr_cycle[  439] = 1'b1;  addr_rom[  439]='h000006dc;  wr_data_rom[  439]='h000010fd;
    rd_cycle[  440] = 1'b0;  wr_cycle[  440] = 1'b1;  addr_rom[  440]='h000006e0;  wr_data_rom[  440]='h0000075d;
    rd_cycle[  441] = 1'b0;  wr_cycle[  441] = 1'b1;  addr_rom[  441]='h000006e4;  wr_data_rom[  441]='h00001971;
    rd_cycle[  442] = 1'b0;  wr_cycle[  442] = 1'b1;  addr_rom[  442]='h000006e8;  wr_data_rom[  442]='h00001609;
    rd_cycle[  443] = 1'b0;  wr_cycle[  443] = 1'b1;  addr_rom[  443]='h000006ec;  wr_data_rom[  443]='h00001232;
    rd_cycle[  444] = 1'b0;  wr_cycle[  444] = 1'b1;  addr_rom[  444]='h000006f0;  wr_data_rom[  444]='h000005a5;
    rd_cycle[  445] = 1'b0;  wr_cycle[  445] = 1'b1;  addr_rom[  445]='h000006f4;  wr_data_rom[  445]='h00000987;
    rd_cycle[  446] = 1'b0;  wr_cycle[  446] = 1'b1;  addr_rom[  446]='h000006f8;  wr_data_rom[  446]='h00001879;
    rd_cycle[  447] = 1'b0;  wr_cycle[  447] = 1'b1;  addr_rom[  447]='h000006fc;  wr_data_rom[  447]='h00001d89;
    rd_cycle[  448] = 1'b0;  wr_cycle[  448] = 1'b1;  addr_rom[  448]='h00000700;  wr_data_rom[  448]='h000001fc;
    rd_cycle[  449] = 1'b0;  wr_cycle[  449] = 1'b1;  addr_rom[  449]='h00000704;  wr_data_rom[  449]='h00001177;
    rd_cycle[  450] = 1'b0;  wr_cycle[  450] = 1'b1;  addr_rom[  450]='h00000708;  wr_data_rom[  450]='h0000124b;
    rd_cycle[  451] = 1'b0;  wr_cycle[  451] = 1'b1;  addr_rom[  451]='h0000070c;  wr_data_rom[  451]='h00000dc0;
    rd_cycle[  452] = 1'b0;  wr_cycle[  452] = 1'b1;  addr_rom[  452]='h00000710;  wr_data_rom[  452]='h00001bdc;
    rd_cycle[  453] = 1'b0;  wr_cycle[  453] = 1'b1;  addr_rom[  453]='h00000714;  wr_data_rom[  453]='h00001cd2;
    rd_cycle[  454] = 1'b0;  wr_cycle[  454] = 1'b1;  addr_rom[  454]='h00000718;  wr_data_rom[  454]='h000012ac;
    rd_cycle[  455] = 1'b0;  wr_cycle[  455] = 1'b1;  addr_rom[  455]='h0000071c;  wr_data_rom[  455]='h00001491;
    rd_cycle[  456] = 1'b0;  wr_cycle[  456] = 1'b1;  addr_rom[  456]='h00000720;  wr_data_rom[  456]='h000010ad;
    rd_cycle[  457] = 1'b0;  wr_cycle[  457] = 1'b1;  addr_rom[  457]='h00000724;  wr_data_rom[  457]='h00001617;
    rd_cycle[  458] = 1'b0;  wr_cycle[  458] = 1'b1;  addr_rom[  458]='h00000728;  wr_data_rom[  458]='h00000028;
    rd_cycle[  459] = 1'b0;  wr_cycle[  459] = 1'b1;  addr_rom[  459]='h0000072c;  wr_data_rom[  459]='h00001d00;
    rd_cycle[  460] = 1'b0;  wr_cycle[  460] = 1'b1;  addr_rom[  460]='h00000730;  wr_data_rom[  460]='h0000057f;
    rd_cycle[  461] = 1'b0;  wr_cycle[  461] = 1'b1;  addr_rom[  461]='h00000734;  wr_data_rom[  461]='h0000115f;
    rd_cycle[  462] = 1'b0;  wr_cycle[  462] = 1'b1;  addr_rom[  462]='h00000738;  wr_data_rom[  462]='h00001d52;
    rd_cycle[  463] = 1'b0;  wr_cycle[  463] = 1'b1;  addr_rom[  463]='h0000073c;  wr_data_rom[  463]='h00000662;
    rd_cycle[  464] = 1'b0;  wr_cycle[  464] = 1'b1;  addr_rom[  464]='h00000740;  wr_data_rom[  464]='h000007ff;
    rd_cycle[  465] = 1'b0;  wr_cycle[  465] = 1'b1;  addr_rom[  465]='h00000744;  wr_data_rom[  465]='h00001ba7;
    rd_cycle[  466] = 1'b0;  wr_cycle[  466] = 1'b1;  addr_rom[  466]='h00000748;  wr_data_rom[  466]='h00000348;
    rd_cycle[  467] = 1'b0;  wr_cycle[  467] = 1'b1;  addr_rom[  467]='h0000074c;  wr_data_rom[  467]='h00000a59;
    rd_cycle[  468] = 1'b0;  wr_cycle[  468] = 1'b1;  addr_rom[  468]='h00000750;  wr_data_rom[  468]='h000009db;
    rd_cycle[  469] = 1'b0;  wr_cycle[  469] = 1'b1;  addr_rom[  469]='h00000754;  wr_data_rom[  469]='h00001188;
    rd_cycle[  470] = 1'b0;  wr_cycle[  470] = 1'b1;  addr_rom[  470]='h00000758;  wr_data_rom[  470]='h000018b4;
    rd_cycle[  471] = 1'b0;  wr_cycle[  471] = 1'b1;  addr_rom[  471]='h0000075c;  wr_data_rom[  471]='h00001117;
    rd_cycle[  472] = 1'b0;  wr_cycle[  472] = 1'b1;  addr_rom[  472]='h00000760;  wr_data_rom[  472]='h0000166c;
    rd_cycle[  473] = 1'b0;  wr_cycle[  473] = 1'b1;  addr_rom[  473]='h00000764;  wr_data_rom[  473]='h00000107;
    rd_cycle[  474] = 1'b0;  wr_cycle[  474] = 1'b1;  addr_rom[  474]='h00000768;  wr_data_rom[  474]='h00001de2;
    rd_cycle[  475] = 1'b0;  wr_cycle[  475] = 1'b1;  addr_rom[  475]='h0000076c;  wr_data_rom[  475]='h00001498;
    rd_cycle[  476] = 1'b0;  wr_cycle[  476] = 1'b1;  addr_rom[  476]='h00000770;  wr_data_rom[  476]='h0000185e;
    rd_cycle[  477] = 1'b0;  wr_cycle[  477] = 1'b1;  addr_rom[  477]='h00000774;  wr_data_rom[  477]='h00001b6d;
    rd_cycle[  478] = 1'b0;  wr_cycle[  478] = 1'b1;  addr_rom[  478]='h00000778;  wr_data_rom[  478]='h00000281;
    rd_cycle[  479] = 1'b0;  wr_cycle[  479] = 1'b1;  addr_rom[  479]='h0000077c;  wr_data_rom[  479]='h000003e9;
    rd_cycle[  480] = 1'b0;  wr_cycle[  480] = 1'b1;  addr_rom[  480]='h00000780;  wr_data_rom[  480]='h0000087e;
    rd_cycle[  481] = 1'b0;  wr_cycle[  481] = 1'b1;  addr_rom[  481]='h00000784;  wr_data_rom[  481]='h000000b1;
    rd_cycle[  482] = 1'b0;  wr_cycle[  482] = 1'b1;  addr_rom[  482]='h00000788;  wr_data_rom[  482]='h00000df1;
    rd_cycle[  483] = 1'b0;  wr_cycle[  483] = 1'b1;  addr_rom[  483]='h0000078c;  wr_data_rom[  483]='h00000ef7;
    rd_cycle[  484] = 1'b0;  wr_cycle[  484] = 1'b1;  addr_rom[  484]='h00000790;  wr_data_rom[  484]='h00000877;
    rd_cycle[  485] = 1'b0;  wr_cycle[  485] = 1'b1;  addr_rom[  485]='h00000794;  wr_data_rom[  485]='h00001363;
    rd_cycle[  486] = 1'b0;  wr_cycle[  486] = 1'b1;  addr_rom[  486]='h00000798;  wr_data_rom[  486]='h00000db0;
    rd_cycle[  487] = 1'b0;  wr_cycle[  487] = 1'b1;  addr_rom[  487]='h0000079c;  wr_data_rom[  487]='h000019fb;
    rd_cycle[  488] = 1'b0;  wr_cycle[  488] = 1'b1;  addr_rom[  488]='h000007a0;  wr_data_rom[  488]='h00001020;
    rd_cycle[  489] = 1'b0;  wr_cycle[  489] = 1'b1;  addr_rom[  489]='h000007a4;  wr_data_rom[  489]='h00000d22;
    rd_cycle[  490] = 1'b0;  wr_cycle[  490] = 1'b1;  addr_rom[  490]='h000007a8;  wr_data_rom[  490]='h0000069b;
    rd_cycle[  491] = 1'b0;  wr_cycle[  491] = 1'b1;  addr_rom[  491]='h000007ac;  wr_data_rom[  491]='h000001fb;
    rd_cycle[  492] = 1'b0;  wr_cycle[  492] = 1'b1;  addr_rom[  492]='h000007b0;  wr_data_rom[  492]='h00001678;
    rd_cycle[  493] = 1'b0;  wr_cycle[  493] = 1'b1;  addr_rom[  493]='h000007b4;  wr_data_rom[  493]='h00001c31;
    rd_cycle[  494] = 1'b0;  wr_cycle[  494] = 1'b1;  addr_rom[  494]='h000007b8;  wr_data_rom[  494]='h00001154;
    rd_cycle[  495] = 1'b0;  wr_cycle[  495] = 1'b1;  addr_rom[  495]='h000007bc;  wr_data_rom[  495]='h00001d24;
    rd_cycle[  496] = 1'b0;  wr_cycle[  496] = 1'b1;  addr_rom[  496]='h000007c0;  wr_data_rom[  496]='h00000b5a;
    rd_cycle[  497] = 1'b0;  wr_cycle[  497] = 1'b1;  addr_rom[  497]='h000007c4;  wr_data_rom[  497]='h00001dbd;
    rd_cycle[  498] = 1'b0;  wr_cycle[  498] = 1'b1;  addr_rom[  498]='h000007c8;  wr_data_rom[  498]='h00001065;
    rd_cycle[  499] = 1'b0;  wr_cycle[  499] = 1'b1;  addr_rom[  499]='h000007cc;  wr_data_rom[  499]='h0000185d;
    rd_cycle[  500] = 1'b0;  wr_cycle[  500] = 1'b1;  addr_rom[  500]='h000007d0;  wr_data_rom[  500]='h00000f32;
    rd_cycle[  501] = 1'b0;  wr_cycle[  501] = 1'b1;  addr_rom[  501]='h000007d4;  wr_data_rom[  501]='h0000072b;
    rd_cycle[  502] = 1'b0;  wr_cycle[  502] = 1'b1;  addr_rom[  502]='h000007d8;  wr_data_rom[  502]='h00000630;
    rd_cycle[  503] = 1'b0;  wr_cycle[  503] = 1'b1;  addr_rom[  503]='h000007dc;  wr_data_rom[  503]='h0000091d;
    rd_cycle[  504] = 1'b0;  wr_cycle[  504] = 1'b1;  addr_rom[  504]='h000007e0;  wr_data_rom[  504]='h00000f63;
    rd_cycle[  505] = 1'b0;  wr_cycle[  505] = 1'b1;  addr_rom[  505]='h000007e4;  wr_data_rom[  505]='h00001d2d;
    rd_cycle[  506] = 1'b0;  wr_cycle[  506] = 1'b1;  addr_rom[  506]='h000007e8;  wr_data_rom[  506]='h00000b8b;
    rd_cycle[  507] = 1'b0;  wr_cycle[  507] = 1'b1;  addr_rom[  507]='h000007ec;  wr_data_rom[  507]='h00000785;
    rd_cycle[  508] = 1'b0;  wr_cycle[  508] = 1'b1;  addr_rom[  508]='h000007f0;  wr_data_rom[  508]='h0000154e;
    rd_cycle[  509] = 1'b0;  wr_cycle[  509] = 1'b1;  addr_rom[  509]='h000007f4;  wr_data_rom[  509]='h000000ec;
    rd_cycle[  510] = 1'b0;  wr_cycle[  510] = 1'b1;  addr_rom[  510]='h000007f8;  wr_data_rom[  510]='h000005f9;
    rd_cycle[  511] = 1'b0;  wr_cycle[  511] = 1'b1;  addr_rom[  511]='h000007fc;  wr_data_rom[  511]='h000007e1;
    rd_cycle[  512] = 1'b0;  wr_cycle[  512] = 1'b1;  addr_rom[  512]='h00000800;  wr_data_rom[  512]='h00001d2a;
    rd_cycle[  513] = 1'b0;  wr_cycle[  513] = 1'b1;  addr_rom[  513]='h00000804;  wr_data_rom[  513]='h00000cad;
    rd_cycle[  514] = 1'b0;  wr_cycle[  514] = 1'b1;  addr_rom[  514]='h00000808;  wr_data_rom[  514]='h00001435;
    rd_cycle[  515] = 1'b0;  wr_cycle[  515] = 1'b1;  addr_rom[  515]='h0000080c;  wr_data_rom[  515]='h00000256;
    rd_cycle[  516] = 1'b0;  wr_cycle[  516] = 1'b1;  addr_rom[  516]='h00000810;  wr_data_rom[  516]='h00001866;
    rd_cycle[  517] = 1'b0;  wr_cycle[  517] = 1'b1;  addr_rom[  517]='h00000814;  wr_data_rom[  517]='h00000e5b;
    rd_cycle[  518] = 1'b0;  wr_cycle[  518] = 1'b1;  addr_rom[  518]='h00000818;  wr_data_rom[  518]='h0000085c;
    rd_cycle[  519] = 1'b0;  wr_cycle[  519] = 1'b1;  addr_rom[  519]='h0000081c;  wr_data_rom[  519]='h00000320;
    rd_cycle[  520] = 1'b0;  wr_cycle[  520] = 1'b1;  addr_rom[  520]='h00000820;  wr_data_rom[  520]='h00001e62;
    rd_cycle[  521] = 1'b0;  wr_cycle[  521] = 1'b1;  addr_rom[  521]='h00000824;  wr_data_rom[  521]='h00000fe1;
    rd_cycle[  522] = 1'b0;  wr_cycle[  522] = 1'b1;  addr_rom[  522]='h00000828;  wr_data_rom[  522]='h000000d7;
    rd_cycle[  523] = 1'b0;  wr_cycle[  523] = 1'b1;  addr_rom[  523]='h0000082c;  wr_data_rom[  523]='h0000104e;
    rd_cycle[  524] = 1'b0;  wr_cycle[  524] = 1'b1;  addr_rom[  524]='h00000830;  wr_data_rom[  524]='h00000a30;
    rd_cycle[  525] = 1'b0;  wr_cycle[  525] = 1'b1;  addr_rom[  525]='h00000834;  wr_data_rom[  525]='h000001f0;
    rd_cycle[  526] = 1'b0;  wr_cycle[  526] = 1'b1;  addr_rom[  526]='h00000838;  wr_data_rom[  526]='h000002c2;
    rd_cycle[  527] = 1'b0;  wr_cycle[  527] = 1'b1;  addr_rom[  527]='h0000083c;  wr_data_rom[  527]='h00001f21;
    rd_cycle[  528] = 1'b0;  wr_cycle[  528] = 1'b1;  addr_rom[  528]='h00000840;  wr_data_rom[  528]='h00000572;
    rd_cycle[  529] = 1'b0;  wr_cycle[  529] = 1'b1;  addr_rom[  529]='h00000844;  wr_data_rom[  529]='h0000136e;
    rd_cycle[  530] = 1'b0;  wr_cycle[  530] = 1'b1;  addr_rom[  530]='h00000848;  wr_data_rom[  530]='h00000355;
    rd_cycle[  531] = 1'b0;  wr_cycle[  531] = 1'b1;  addr_rom[  531]='h0000084c;  wr_data_rom[  531]='h00001dfa;
    rd_cycle[  532] = 1'b0;  wr_cycle[  532] = 1'b1;  addr_rom[  532]='h00000850;  wr_data_rom[  532]='h000008b9;
    rd_cycle[  533] = 1'b0;  wr_cycle[  533] = 1'b1;  addr_rom[  533]='h00000854;  wr_data_rom[  533]='h00000fd7;
    rd_cycle[  534] = 1'b0;  wr_cycle[  534] = 1'b1;  addr_rom[  534]='h00000858;  wr_data_rom[  534]='h000005a3;
    rd_cycle[  535] = 1'b0;  wr_cycle[  535] = 1'b1;  addr_rom[  535]='h0000085c;  wr_data_rom[  535]='h00000a90;
    rd_cycle[  536] = 1'b0;  wr_cycle[  536] = 1'b1;  addr_rom[  536]='h00000860;  wr_data_rom[  536]='h00000051;
    rd_cycle[  537] = 1'b0;  wr_cycle[  537] = 1'b1;  addr_rom[  537]='h00000864;  wr_data_rom[  537]='h00001516;
    rd_cycle[  538] = 1'b0;  wr_cycle[  538] = 1'b1;  addr_rom[  538]='h00000868;  wr_data_rom[  538]='h000003cd;
    rd_cycle[  539] = 1'b0;  wr_cycle[  539] = 1'b1;  addr_rom[  539]='h0000086c;  wr_data_rom[  539]='h000009bb;
    rd_cycle[  540] = 1'b0;  wr_cycle[  540] = 1'b1;  addr_rom[  540]='h00000870;  wr_data_rom[  540]='h00001731;
    rd_cycle[  541] = 1'b0;  wr_cycle[  541] = 1'b1;  addr_rom[  541]='h00000874;  wr_data_rom[  541]='h00001d02;
    rd_cycle[  542] = 1'b0;  wr_cycle[  542] = 1'b1;  addr_rom[  542]='h00000878;  wr_data_rom[  542]='h00001bac;
    rd_cycle[  543] = 1'b0;  wr_cycle[  543] = 1'b1;  addr_rom[  543]='h0000087c;  wr_data_rom[  543]='h000011fe;
    rd_cycle[  544] = 1'b0;  wr_cycle[  544] = 1'b1;  addr_rom[  544]='h00000880;  wr_data_rom[  544]='h00000491;
    rd_cycle[  545] = 1'b0;  wr_cycle[  545] = 1'b1;  addr_rom[  545]='h00000884;  wr_data_rom[  545]='h000009b9;
    rd_cycle[  546] = 1'b0;  wr_cycle[  546] = 1'b1;  addr_rom[  546]='h00000888;  wr_data_rom[  546]='h00000249;
    rd_cycle[  547] = 1'b0;  wr_cycle[  547] = 1'b1;  addr_rom[  547]='h0000088c;  wr_data_rom[  547]='h00001b9d;
    rd_cycle[  548] = 1'b0;  wr_cycle[  548] = 1'b1;  addr_rom[  548]='h00000890;  wr_data_rom[  548]='h00000f4d;
    rd_cycle[  549] = 1'b0;  wr_cycle[  549] = 1'b1;  addr_rom[  549]='h00000894;  wr_data_rom[  549]='h00000a16;
    rd_cycle[  550] = 1'b0;  wr_cycle[  550] = 1'b1;  addr_rom[  550]='h00000898;  wr_data_rom[  550]='h000014e6;
    rd_cycle[  551] = 1'b0;  wr_cycle[  551] = 1'b1;  addr_rom[  551]='h0000089c;  wr_data_rom[  551]='h00000894;
    rd_cycle[  552] = 1'b0;  wr_cycle[  552] = 1'b1;  addr_rom[  552]='h000008a0;  wr_data_rom[  552]='h00000c4c;
    rd_cycle[  553] = 1'b0;  wr_cycle[  553] = 1'b1;  addr_rom[  553]='h000008a4;  wr_data_rom[  553]='h0000120a;
    rd_cycle[  554] = 1'b0;  wr_cycle[  554] = 1'b1;  addr_rom[  554]='h000008a8;  wr_data_rom[  554]='h000011f9;
    rd_cycle[  555] = 1'b0;  wr_cycle[  555] = 1'b1;  addr_rom[  555]='h000008ac;  wr_data_rom[  555]='h00001bdf;
    rd_cycle[  556] = 1'b0;  wr_cycle[  556] = 1'b1;  addr_rom[  556]='h000008b0;  wr_data_rom[  556]='h000016fc;
    rd_cycle[  557] = 1'b0;  wr_cycle[  557] = 1'b1;  addr_rom[  557]='h000008b4;  wr_data_rom[  557]='h0000047d;
    rd_cycle[  558] = 1'b0;  wr_cycle[  558] = 1'b1;  addr_rom[  558]='h000008b8;  wr_data_rom[  558]='h0000197c;
    rd_cycle[  559] = 1'b0;  wr_cycle[  559] = 1'b1;  addr_rom[  559]='h000008bc;  wr_data_rom[  559]='h00000405;
    rd_cycle[  560] = 1'b0;  wr_cycle[  560] = 1'b1;  addr_rom[  560]='h000008c0;  wr_data_rom[  560]='h000004ba;
    rd_cycle[  561] = 1'b0;  wr_cycle[  561] = 1'b1;  addr_rom[  561]='h000008c4;  wr_data_rom[  561]='h00000198;
    rd_cycle[  562] = 1'b0;  wr_cycle[  562] = 1'b1;  addr_rom[  562]='h000008c8;  wr_data_rom[  562]='h00001471;
    rd_cycle[  563] = 1'b0;  wr_cycle[  563] = 1'b1;  addr_rom[  563]='h000008cc;  wr_data_rom[  563]='h00000e4f;
    rd_cycle[  564] = 1'b0;  wr_cycle[  564] = 1'b1;  addr_rom[  564]='h000008d0;  wr_data_rom[  564]='h000012a5;
    rd_cycle[  565] = 1'b0;  wr_cycle[  565] = 1'b1;  addr_rom[  565]='h000008d4;  wr_data_rom[  565]='h00000ddb;
    rd_cycle[  566] = 1'b0;  wr_cycle[  566] = 1'b1;  addr_rom[  566]='h000008d8;  wr_data_rom[  566]='h00001e9e;
    rd_cycle[  567] = 1'b0;  wr_cycle[  567] = 1'b1;  addr_rom[  567]='h000008dc;  wr_data_rom[  567]='h000003e8;
    rd_cycle[  568] = 1'b0;  wr_cycle[  568] = 1'b1;  addr_rom[  568]='h000008e0;  wr_data_rom[  568]='h00000db1;
    rd_cycle[  569] = 1'b0;  wr_cycle[  569] = 1'b1;  addr_rom[  569]='h000008e4;  wr_data_rom[  569]='h0000137a;
    rd_cycle[  570] = 1'b0;  wr_cycle[  570] = 1'b1;  addr_rom[  570]='h000008e8;  wr_data_rom[  570]='h000011ea;
    rd_cycle[  571] = 1'b0;  wr_cycle[  571] = 1'b1;  addr_rom[  571]='h000008ec;  wr_data_rom[  571]='h00000afe;
    rd_cycle[  572] = 1'b0;  wr_cycle[  572] = 1'b1;  addr_rom[  572]='h000008f0;  wr_data_rom[  572]='h000015c2;
    rd_cycle[  573] = 1'b0;  wr_cycle[  573] = 1'b1;  addr_rom[  573]='h000008f4;  wr_data_rom[  573]='h000019f9;
    rd_cycle[  574] = 1'b0;  wr_cycle[  574] = 1'b1;  addr_rom[  574]='h000008f8;  wr_data_rom[  574]='h000018ec;
    rd_cycle[  575] = 1'b0;  wr_cycle[  575] = 1'b1;  addr_rom[  575]='h000008fc;  wr_data_rom[  575]='h000014f2;
    rd_cycle[  576] = 1'b0;  wr_cycle[  576] = 1'b1;  addr_rom[  576]='h00000900;  wr_data_rom[  576]='h00001b2b;
    rd_cycle[  577] = 1'b0;  wr_cycle[  577] = 1'b1;  addr_rom[  577]='h00000904;  wr_data_rom[  577]='h00001b17;
    rd_cycle[  578] = 1'b0;  wr_cycle[  578] = 1'b1;  addr_rom[  578]='h00000908;  wr_data_rom[  578]='h00000270;
    rd_cycle[  579] = 1'b0;  wr_cycle[  579] = 1'b1;  addr_rom[  579]='h0000090c;  wr_data_rom[  579]='h00001800;
    rd_cycle[  580] = 1'b0;  wr_cycle[  580] = 1'b1;  addr_rom[  580]='h00000910;  wr_data_rom[  580]='h000000b7;
    rd_cycle[  581] = 1'b0;  wr_cycle[  581] = 1'b1;  addr_rom[  581]='h00000914;  wr_data_rom[  581]='h00000280;
    rd_cycle[  582] = 1'b0;  wr_cycle[  582] = 1'b1;  addr_rom[  582]='h00000918;  wr_data_rom[  582]='h00000603;
    rd_cycle[  583] = 1'b0;  wr_cycle[  583] = 1'b1;  addr_rom[  583]='h0000091c;  wr_data_rom[  583]='h00000d86;
    rd_cycle[  584] = 1'b0;  wr_cycle[  584] = 1'b1;  addr_rom[  584]='h00000920;  wr_data_rom[  584]='h0000160c;
    rd_cycle[  585] = 1'b0;  wr_cycle[  585] = 1'b1;  addr_rom[  585]='h00000924;  wr_data_rom[  585]='h00001d93;
    rd_cycle[  586] = 1'b0;  wr_cycle[  586] = 1'b1;  addr_rom[  586]='h00000928;  wr_data_rom[  586]='h0000121c;
    rd_cycle[  587] = 1'b0;  wr_cycle[  587] = 1'b1;  addr_rom[  587]='h0000092c;  wr_data_rom[  587]='h00000edd;
    rd_cycle[  588] = 1'b0;  wr_cycle[  588] = 1'b1;  addr_rom[  588]='h00000930;  wr_data_rom[  588]='h0000024d;
    rd_cycle[  589] = 1'b0;  wr_cycle[  589] = 1'b1;  addr_rom[  589]='h00000934;  wr_data_rom[  589]='h0000000d;
    rd_cycle[  590] = 1'b0;  wr_cycle[  590] = 1'b1;  addr_rom[  590]='h00000938;  wr_data_rom[  590]='h000004d3;
    rd_cycle[  591] = 1'b0;  wr_cycle[  591] = 1'b1;  addr_rom[  591]='h0000093c;  wr_data_rom[  591]='h00001493;
    rd_cycle[  592] = 1'b0;  wr_cycle[  592] = 1'b1;  addr_rom[  592]='h00000940;  wr_data_rom[  592]='h00000279;
    rd_cycle[  593] = 1'b0;  wr_cycle[  593] = 1'b1;  addr_rom[  593]='h00000944;  wr_data_rom[  593]='h0000161e;
    rd_cycle[  594] = 1'b0;  wr_cycle[  594] = 1'b1;  addr_rom[  594]='h00000948;  wr_data_rom[  594]='h00000409;
    rd_cycle[  595] = 1'b0;  wr_cycle[  595] = 1'b1;  addr_rom[  595]='h0000094c;  wr_data_rom[  595]='h00001c3b;
    rd_cycle[  596] = 1'b0;  wr_cycle[  596] = 1'b1;  addr_rom[  596]='h00000950;  wr_data_rom[  596]='h00001d9a;
    rd_cycle[  597] = 1'b0;  wr_cycle[  597] = 1'b1;  addr_rom[  597]='h00000954;  wr_data_rom[  597]='h00001c14;
    rd_cycle[  598] = 1'b0;  wr_cycle[  598] = 1'b1;  addr_rom[  598]='h00000958;  wr_data_rom[  598]='h00001d9d;
    rd_cycle[  599] = 1'b0;  wr_cycle[  599] = 1'b1;  addr_rom[  599]='h0000095c;  wr_data_rom[  599]='h00000b52;
    rd_cycle[  600] = 1'b0;  wr_cycle[  600] = 1'b1;  addr_rom[  600]='h00000960;  wr_data_rom[  600]='h00001bf4;
    rd_cycle[  601] = 1'b0;  wr_cycle[  601] = 1'b1;  addr_rom[  601]='h00000964;  wr_data_rom[  601]='h00001e73;
    rd_cycle[  602] = 1'b0;  wr_cycle[  602] = 1'b1;  addr_rom[  602]='h00000968;  wr_data_rom[  602]='h000012e4;
    rd_cycle[  603] = 1'b0;  wr_cycle[  603] = 1'b1;  addr_rom[  603]='h0000096c;  wr_data_rom[  603]='h000014e4;
    rd_cycle[  604] = 1'b0;  wr_cycle[  604] = 1'b1;  addr_rom[  604]='h00000970;  wr_data_rom[  604]='h00001b93;
    rd_cycle[  605] = 1'b0;  wr_cycle[  605] = 1'b1;  addr_rom[  605]='h00000974;  wr_data_rom[  605]='h00001b69;
    rd_cycle[  606] = 1'b0;  wr_cycle[  606] = 1'b1;  addr_rom[  606]='h00000978;  wr_data_rom[  606]='h00001e3a;
    rd_cycle[  607] = 1'b0;  wr_cycle[  607] = 1'b1;  addr_rom[  607]='h0000097c;  wr_data_rom[  607]='h000002da;
    rd_cycle[  608] = 1'b0;  wr_cycle[  608] = 1'b1;  addr_rom[  608]='h00000980;  wr_data_rom[  608]='h00001663;
    rd_cycle[  609] = 1'b0;  wr_cycle[  609] = 1'b1;  addr_rom[  609]='h00000984;  wr_data_rom[  609]='h0000189d;
    rd_cycle[  610] = 1'b0;  wr_cycle[  610] = 1'b1;  addr_rom[  610]='h00000988;  wr_data_rom[  610]='h00000a0c;
    rd_cycle[  611] = 1'b0;  wr_cycle[  611] = 1'b1;  addr_rom[  611]='h0000098c;  wr_data_rom[  611]='h000016bb;
    rd_cycle[  612] = 1'b0;  wr_cycle[  612] = 1'b1;  addr_rom[  612]='h00000990;  wr_data_rom[  612]='h00001bd2;
    rd_cycle[  613] = 1'b0;  wr_cycle[  613] = 1'b1;  addr_rom[  613]='h00000994;  wr_data_rom[  613]='h0000076f;
    rd_cycle[  614] = 1'b0;  wr_cycle[  614] = 1'b1;  addr_rom[  614]='h00000998;  wr_data_rom[  614]='h0000057b;
    rd_cycle[  615] = 1'b0;  wr_cycle[  615] = 1'b1;  addr_rom[  615]='h0000099c;  wr_data_rom[  615]='h00000829;
    rd_cycle[  616] = 1'b0;  wr_cycle[  616] = 1'b1;  addr_rom[  616]='h000009a0;  wr_data_rom[  616]='h00000340;
    rd_cycle[  617] = 1'b0;  wr_cycle[  617] = 1'b1;  addr_rom[  617]='h000009a4;  wr_data_rom[  617]='h00000f2d;
    rd_cycle[  618] = 1'b0;  wr_cycle[  618] = 1'b1;  addr_rom[  618]='h000009a8;  wr_data_rom[  618]='h0000030e;
    rd_cycle[  619] = 1'b0;  wr_cycle[  619] = 1'b1;  addr_rom[  619]='h000009ac;  wr_data_rom[  619]='h00000dc3;
    rd_cycle[  620] = 1'b0;  wr_cycle[  620] = 1'b1;  addr_rom[  620]='h000009b0;  wr_data_rom[  620]='h000016f2;
    rd_cycle[  621] = 1'b0;  wr_cycle[  621] = 1'b1;  addr_rom[  621]='h000009b4;  wr_data_rom[  621]='h00000cf7;
    rd_cycle[  622] = 1'b0;  wr_cycle[  622] = 1'b1;  addr_rom[  622]='h000009b8;  wr_data_rom[  622]='h00000c0d;
    rd_cycle[  623] = 1'b0;  wr_cycle[  623] = 1'b1;  addr_rom[  623]='h000009bc;  wr_data_rom[  623]='h00000c59;
    rd_cycle[  624] = 1'b0;  wr_cycle[  624] = 1'b1;  addr_rom[  624]='h000009c0;  wr_data_rom[  624]='h00000d7e;
    rd_cycle[  625] = 1'b0;  wr_cycle[  625] = 1'b1;  addr_rom[  625]='h000009c4;  wr_data_rom[  625]='h00000f50;
    rd_cycle[  626] = 1'b0;  wr_cycle[  626] = 1'b1;  addr_rom[  626]='h000009c8;  wr_data_rom[  626]='h0000199f;
    rd_cycle[  627] = 1'b0;  wr_cycle[  627] = 1'b1;  addr_rom[  627]='h000009cc;  wr_data_rom[  627]='h00000f03;
    rd_cycle[  628] = 1'b0;  wr_cycle[  628] = 1'b1;  addr_rom[  628]='h000009d0;  wr_data_rom[  628]='h00000d85;
    rd_cycle[  629] = 1'b0;  wr_cycle[  629] = 1'b1;  addr_rom[  629]='h000009d4;  wr_data_rom[  629]='h00000a68;
    rd_cycle[  630] = 1'b0;  wr_cycle[  630] = 1'b1;  addr_rom[  630]='h000009d8;  wr_data_rom[  630]='h0000111d;
    rd_cycle[  631] = 1'b0;  wr_cycle[  631] = 1'b1;  addr_rom[  631]='h000009dc;  wr_data_rom[  631]='h00001338;
    rd_cycle[  632] = 1'b0;  wr_cycle[  632] = 1'b1;  addr_rom[  632]='h000009e0;  wr_data_rom[  632]='h0000045b;
    rd_cycle[  633] = 1'b0;  wr_cycle[  633] = 1'b1;  addr_rom[  633]='h000009e4;  wr_data_rom[  633]='h00000aa0;
    rd_cycle[  634] = 1'b0;  wr_cycle[  634] = 1'b1;  addr_rom[  634]='h000009e8;  wr_data_rom[  634]='h00000b4d;
    rd_cycle[  635] = 1'b0;  wr_cycle[  635] = 1'b1;  addr_rom[  635]='h000009ec;  wr_data_rom[  635]='h00001613;
    rd_cycle[  636] = 1'b0;  wr_cycle[  636] = 1'b1;  addr_rom[  636]='h000009f0;  wr_data_rom[  636]='h00000367;
    rd_cycle[  637] = 1'b0;  wr_cycle[  637] = 1'b1;  addr_rom[  637]='h000009f4;  wr_data_rom[  637]='h00000c30;
    rd_cycle[  638] = 1'b0;  wr_cycle[  638] = 1'b1;  addr_rom[  638]='h000009f8;  wr_data_rom[  638]='h000004e9;
    rd_cycle[  639] = 1'b0;  wr_cycle[  639] = 1'b1;  addr_rom[  639]='h000009fc;  wr_data_rom[  639]='h0000183c;
    rd_cycle[  640] = 1'b0;  wr_cycle[  640] = 1'b1;  addr_rom[  640]='h00000a00;  wr_data_rom[  640]='h00001275;
    rd_cycle[  641] = 1'b0;  wr_cycle[  641] = 1'b1;  addr_rom[  641]='h00000a04;  wr_data_rom[  641]='h000005c7;
    rd_cycle[  642] = 1'b0;  wr_cycle[  642] = 1'b1;  addr_rom[  642]='h00000a08;  wr_data_rom[  642]='h00001c95;
    rd_cycle[  643] = 1'b0;  wr_cycle[  643] = 1'b1;  addr_rom[  643]='h00000a0c;  wr_data_rom[  643]='h000009b1;
    rd_cycle[  644] = 1'b0;  wr_cycle[  644] = 1'b1;  addr_rom[  644]='h00000a10;  wr_data_rom[  644]='h0000006e;
    rd_cycle[  645] = 1'b0;  wr_cycle[  645] = 1'b1;  addr_rom[  645]='h00000a14;  wr_data_rom[  645]='h00001c12;
    rd_cycle[  646] = 1'b0;  wr_cycle[  646] = 1'b1;  addr_rom[  646]='h00000a18;  wr_data_rom[  646]='h000011b3;
    rd_cycle[  647] = 1'b0;  wr_cycle[  647] = 1'b1;  addr_rom[  647]='h00000a1c;  wr_data_rom[  647]='h00001ef4;
    rd_cycle[  648] = 1'b0;  wr_cycle[  648] = 1'b1;  addr_rom[  648]='h00000a20;  wr_data_rom[  648]='h00000a4d;
    rd_cycle[  649] = 1'b0;  wr_cycle[  649] = 1'b1;  addr_rom[  649]='h00000a24;  wr_data_rom[  649]='h00001de7;
    rd_cycle[  650] = 1'b0;  wr_cycle[  650] = 1'b1;  addr_rom[  650]='h00000a28;  wr_data_rom[  650]='h0000125a;
    rd_cycle[  651] = 1'b0;  wr_cycle[  651] = 1'b1;  addr_rom[  651]='h00000a2c;  wr_data_rom[  651]='h0000173c;
    rd_cycle[  652] = 1'b0;  wr_cycle[  652] = 1'b1;  addr_rom[  652]='h00000a30;  wr_data_rom[  652]='h00000f01;
    rd_cycle[  653] = 1'b0;  wr_cycle[  653] = 1'b1;  addr_rom[  653]='h00000a34;  wr_data_rom[  653]='h00000ff9;
    rd_cycle[  654] = 1'b0;  wr_cycle[  654] = 1'b1;  addr_rom[  654]='h00000a38;  wr_data_rom[  654]='h00001a54;
    rd_cycle[  655] = 1'b0;  wr_cycle[  655] = 1'b1;  addr_rom[  655]='h00000a3c;  wr_data_rom[  655]='h00001158;
    rd_cycle[  656] = 1'b0;  wr_cycle[  656] = 1'b1;  addr_rom[  656]='h00000a40;  wr_data_rom[  656]='h0000188e;
    rd_cycle[  657] = 1'b0;  wr_cycle[  657] = 1'b1;  addr_rom[  657]='h00000a44;  wr_data_rom[  657]='h000015ad;
    rd_cycle[  658] = 1'b0;  wr_cycle[  658] = 1'b1;  addr_rom[  658]='h00000a48;  wr_data_rom[  658]='h00000b08;
    rd_cycle[  659] = 1'b0;  wr_cycle[  659] = 1'b1;  addr_rom[  659]='h00000a4c;  wr_data_rom[  659]='h00001469;
    rd_cycle[  660] = 1'b0;  wr_cycle[  660] = 1'b1;  addr_rom[  660]='h00000a50;  wr_data_rom[  660]='h00001672;
    rd_cycle[  661] = 1'b0;  wr_cycle[  661] = 1'b1;  addr_rom[  661]='h00000a54;  wr_data_rom[  661]='h00001340;
    rd_cycle[  662] = 1'b0;  wr_cycle[  662] = 1'b1;  addr_rom[  662]='h00000a58;  wr_data_rom[  662]='h0000087c;
    rd_cycle[  663] = 1'b0;  wr_cycle[  663] = 1'b1;  addr_rom[  663]='h00000a5c;  wr_data_rom[  663]='h000011ff;
    rd_cycle[  664] = 1'b0;  wr_cycle[  664] = 1'b1;  addr_rom[  664]='h00000a60;  wr_data_rom[  664]='h00000089;
    rd_cycle[  665] = 1'b0;  wr_cycle[  665] = 1'b1;  addr_rom[  665]='h00000a64;  wr_data_rom[  665]='h000000fe;
    rd_cycle[  666] = 1'b0;  wr_cycle[  666] = 1'b1;  addr_rom[  666]='h00000a68;  wr_data_rom[  666]='h00000bc9;
    rd_cycle[  667] = 1'b0;  wr_cycle[  667] = 1'b1;  addr_rom[  667]='h00000a6c;  wr_data_rom[  667]='h000001cb;
    rd_cycle[  668] = 1'b0;  wr_cycle[  668] = 1'b1;  addr_rom[  668]='h00000a70;  wr_data_rom[  668]='h000003d7;
    rd_cycle[  669] = 1'b0;  wr_cycle[  669] = 1'b1;  addr_rom[  669]='h00000a74;  wr_data_rom[  669]='h00001852;
    rd_cycle[  670] = 1'b0;  wr_cycle[  670] = 1'b1;  addr_rom[  670]='h00000a78;  wr_data_rom[  670]='h000013af;
    rd_cycle[  671] = 1'b0;  wr_cycle[  671] = 1'b1;  addr_rom[  671]='h00000a7c;  wr_data_rom[  671]='h00000cac;
    rd_cycle[  672] = 1'b0;  wr_cycle[  672] = 1'b1;  addr_rom[  672]='h00000a80;  wr_data_rom[  672]='h00001755;
    rd_cycle[  673] = 1'b0;  wr_cycle[  673] = 1'b1;  addr_rom[  673]='h00000a84;  wr_data_rom[  673]='h0000087f;
    rd_cycle[  674] = 1'b0;  wr_cycle[  674] = 1'b1;  addr_rom[  674]='h00000a88;  wr_data_rom[  674]='h00001320;
    rd_cycle[  675] = 1'b0;  wr_cycle[  675] = 1'b1;  addr_rom[  675]='h00000a8c;  wr_data_rom[  675]='h0000090f;
    rd_cycle[  676] = 1'b0;  wr_cycle[  676] = 1'b1;  addr_rom[  676]='h00000a90;  wr_data_rom[  676]='h00000e23;
    rd_cycle[  677] = 1'b0;  wr_cycle[  677] = 1'b1;  addr_rom[  677]='h00000a94;  wr_data_rom[  677]='h00000a1d;
    rd_cycle[  678] = 1'b0;  wr_cycle[  678] = 1'b1;  addr_rom[  678]='h00000a98;  wr_data_rom[  678]='h0000102f;
    rd_cycle[  679] = 1'b0;  wr_cycle[  679] = 1'b1;  addr_rom[  679]='h00000a9c;  wr_data_rom[  679]='h000016e9;
    rd_cycle[  680] = 1'b0;  wr_cycle[  680] = 1'b1;  addr_rom[  680]='h00000aa0;  wr_data_rom[  680]='h00000928;
    rd_cycle[  681] = 1'b0;  wr_cycle[  681] = 1'b1;  addr_rom[  681]='h00000aa4;  wr_data_rom[  681]='h00000de0;
    rd_cycle[  682] = 1'b0;  wr_cycle[  682] = 1'b1;  addr_rom[  682]='h00000aa8;  wr_data_rom[  682]='h00001e8b;
    rd_cycle[  683] = 1'b0;  wr_cycle[  683] = 1'b1;  addr_rom[  683]='h00000aac;  wr_data_rom[  683]='h000011d3;
    rd_cycle[  684] = 1'b0;  wr_cycle[  684] = 1'b1;  addr_rom[  684]='h00000ab0;  wr_data_rom[  684]='h00001116;
    rd_cycle[  685] = 1'b0;  wr_cycle[  685] = 1'b1;  addr_rom[  685]='h00000ab4;  wr_data_rom[  685]='h00001e00;
    rd_cycle[  686] = 1'b0;  wr_cycle[  686] = 1'b1;  addr_rom[  686]='h00000ab8;  wr_data_rom[  686]='h00001897;
    rd_cycle[  687] = 1'b0;  wr_cycle[  687] = 1'b1;  addr_rom[  687]='h00000abc;  wr_data_rom[  687]='h00001f2d;
    rd_cycle[  688] = 1'b0;  wr_cycle[  688] = 1'b1;  addr_rom[  688]='h00000ac0;  wr_data_rom[  688]='h00000a02;
    rd_cycle[  689] = 1'b0;  wr_cycle[  689] = 1'b1;  addr_rom[  689]='h00000ac4;  wr_data_rom[  689]='h00000360;
    rd_cycle[  690] = 1'b0;  wr_cycle[  690] = 1'b1;  addr_rom[  690]='h00000ac8;  wr_data_rom[  690]='h00001391;
    rd_cycle[  691] = 1'b0;  wr_cycle[  691] = 1'b1;  addr_rom[  691]='h00000acc;  wr_data_rom[  691]='h00001e63;
    rd_cycle[  692] = 1'b0;  wr_cycle[  692] = 1'b1;  addr_rom[  692]='h00000ad0;  wr_data_rom[  692]='h00000517;
    rd_cycle[  693] = 1'b0;  wr_cycle[  693] = 1'b1;  addr_rom[  693]='h00000ad4;  wr_data_rom[  693]='h000001b3;
    rd_cycle[  694] = 1'b0;  wr_cycle[  694] = 1'b1;  addr_rom[  694]='h00000ad8;  wr_data_rom[  694]='h0000053e;
    rd_cycle[  695] = 1'b0;  wr_cycle[  695] = 1'b1;  addr_rom[  695]='h00000adc;  wr_data_rom[  695]='h00001d4a;
    rd_cycle[  696] = 1'b0;  wr_cycle[  696] = 1'b1;  addr_rom[  696]='h00000ae0;  wr_data_rom[  696]='h00000326;
    rd_cycle[  697] = 1'b0;  wr_cycle[  697] = 1'b1;  addr_rom[  697]='h00000ae4;  wr_data_rom[  697]='h00000b74;
    rd_cycle[  698] = 1'b0;  wr_cycle[  698] = 1'b1;  addr_rom[  698]='h00000ae8;  wr_data_rom[  698]='h00000446;
    rd_cycle[  699] = 1'b0;  wr_cycle[  699] = 1'b1;  addr_rom[  699]='h00000aec;  wr_data_rom[  699]='h0000028f;
    rd_cycle[  700] = 1'b0;  wr_cycle[  700] = 1'b1;  addr_rom[  700]='h00000af0;  wr_data_rom[  700]='h000019e8;
    rd_cycle[  701] = 1'b0;  wr_cycle[  701] = 1'b1;  addr_rom[  701]='h00000af4;  wr_data_rom[  701]='h00000674;
    rd_cycle[  702] = 1'b0;  wr_cycle[  702] = 1'b1;  addr_rom[  702]='h00000af8;  wr_data_rom[  702]='h0000141e;
    rd_cycle[  703] = 1'b0;  wr_cycle[  703] = 1'b1;  addr_rom[  703]='h00000afc;  wr_data_rom[  703]='h00000316;
    rd_cycle[  704] = 1'b0;  wr_cycle[  704] = 1'b1;  addr_rom[  704]='h00000b00;  wr_data_rom[  704]='h00001de9;
    rd_cycle[  705] = 1'b0;  wr_cycle[  705] = 1'b1;  addr_rom[  705]='h00000b04;  wr_data_rom[  705]='h00000000;
    rd_cycle[  706] = 1'b0;  wr_cycle[  706] = 1'b1;  addr_rom[  706]='h00000b08;  wr_data_rom[  706]='h00001a6b;
    rd_cycle[  707] = 1'b0;  wr_cycle[  707] = 1'b1;  addr_rom[  707]='h00000b0c;  wr_data_rom[  707]='h000000be;
    rd_cycle[  708] = 1'b0;  wr_cycle[  708] = 1'b1;  addr_rom[  708]='h00000b10;  wr_data_rom[  708]='h00000a29;
    rd_cycle[  709] = 1'b0;  wr_cycle[  709] = 1'b1;  addr_rom[  709]='h00000b14;  wr_data_rom[  709]='h00000f1e;
    rd_cycle[  710] = 1'b0;  wr_cycle[  710] = 1'b1;  addr_rom[  710]='h00000b18;  wr_data_rom[  710]='h000016ab;
    rd_cycle[  711] = 1'b0;  wr_cycle[  711] = 1'b1;  addr_rom[  711]='h00000b1c;  wr_data_rom[  711]='h00001754;
    rd_cycle[  712] = 1'b0;  wr_cycle[  712] = 1'b1;  addr_rom[  712]='h00000b20;  wr_data_rom[  712]='h00001301;
    rd_cycle[  713] = 1'b0;  wr_cycle[  713] = 1'b1;  addr_rom[  713]='h00000b24;  wr_data_rom[  713]='h00000243;
    rd_cycle[  714] = 1'b0;  wr_cycle[  714] = 1'b1;  addr_rom[  714]='h00000b28;  wr_data_rom[  714]='h00001584;
    rd_cycle[  715] = 1'b0;  wr_cycle[  715] = 1'b1;  addr_rom[  715]='h00000b2c;  wr_data_rom[  715]='h00000c40;
    rd_cycle[  716] = 1'b0;  wr_cycle[  716] = 1'b1;  addr_rom[  716]='h00000b30;  wr_data_rom[  716]='h00000308;
    rd_cycle[  717] = 1'b0;  wr_cycle[  717] = 1'b1;  addr_rom[  717]='h00000b34;  wr_data_rom[  717]='h00000365;
    rd_cycle[  718] = 1'b0;  wr_cycle[  718] = 1'b1;  addr_rom[  718]='h00000b38;  wr_data_rom[  718]='h0000106a;
    rd_cycle[  719] = 1'b0;  wr_cycle[  719] = 1'b1;  addr_rom[  719]='h00000b3c;  wr_data_rom[  719]='h000004d7;
    rd_cycle[  720] = 1'b0;  wr_cycle[  720] = 1'b1;  addr_rom[  720]='h00000b40;  wr_data_rom[  720]='h00000595;
    rd_cycle[  721] = 1'b0;  wr_cycle[  721] = 1'b1;  addr_rom[  721]='h00000b44;  wr_data_rom[  721]='h00001441;
    rd_cycle[  722] = 1'b0;  wr_cycle[  722] = 1'b1;  addr_rom[  722]='h00000b48;  wr_data_rom[  722]='h00000a8a;
    rd_cycle[  723] = 1'b0;  wr_cycle[  723] = 1'b1;  addr_rom[  723]='h00000b4c;  wr_data_rom[  723]='h00001ca5;
    rd_cycle[  724] = 1'b0;  wr_cycle[  724] = 1'b1;  addr_rom[  724]='h00000b50;  wr_data_rom[  724]='h0000076c;
    rd_cycle[  725] = 1'b0;  wr_cycle[  725] = 1'b1;  addr_rom[  725]='h00000b54;  wr_data_rom[  725]='h00001464;
    rd_cycle[  726] = 1'b0;  wr_cycle[  726] = 1'b1;  addr_rom[  726]='h00000b58;  wr_data_rom[  726]='h00000faf;
    rd_cycle[  727] = 1'b0;  wr_cycle[  727] = 1'b1;  addr_rom[  727]='h00000b5c;  wr_data_rom[  727]='h000004cc;
    rd_cycle[  728] = 1'b0;  wr_cycle[  728] = 1'b1;  addr_rom[  728]='h00000b60;  wr_data_rom[  728]='h00000e66;
    rd_cycle[  729] = 1'b0;  wr_cycle[  729] = 1'b1;  addr_rom[  729]='h00000b64;  wr_data_rom[  729]='h000013b9;
    rd_cycle[  730] = 1'b0;  wr_cycle[  730] = 1'b1;  addr_rom[  730]='h00000b68;  wr_data_rom[  730]='h00000fbe;
    rd_cycle[  731] = 1'b0;  wr_cycle[  731] = 1'b1;  addr_rom[  731]='h00000b6c;  wr_data_rom[  731]='h0000024b;
    rd_cycle[  732] = 1'b0;  wr_cycle[  732] = 1'b1;  addr_rom[  732]='h00000b70;  wr_data_rom[  732]='h000010bf;
    rd_cycle[  733] = 1'b0;  wr_cycle[  733] = 1'b1;  addr_rom[  733]='h00000b74;  wr_data_rom[  733]='h0000050c;
    rd_cycle[  734] = 1'b0;  wr_cycle[  734] = 1'b1;  addr_rom[  734]='h00000b78;  wr_data_rom[  734]='h000005ef;
    rd_cycle[  735] = 1'b0;  wr_cycle[  735] = 1'b1;  addr_rom[  735]='h00000b7c;  wr_data_rom[  735]='h00000d85;
    rd_cycle[  736] = 1'b0;  wr_cycle[  736] = 1'b1;  addr_rom[  736]='h00000b80;  wr_data_rom[  736]='h000011f3;
    rd_cycle[  737] = 1'b0;  wr_cycle[  737] = 1'b1;  addr_rom[  737]='h00000b84;  wr_data_rom[  737]='h000013be;
    rd_cycle[  738] = 1'b0;  wr_cycle[  738] = 1'b1;  addr_rom[  738]='h00000b88;  wr_data_rom[  738]='h00001c3a;
    rd_cycle[  739] = 1'b0;  wr_cycle[  739] = 1'b1;  addr_rom[  739]='h00000b8c;  wr_data_rom[  739]='h00001e38;
    rd_cycle[  740] = 1'b0;  wr_cycle[  740] = 1'b1;  addr_rom[  740]='h00000b90;  wr_data_rom[  740]='h00000aaa;
    rd_cycle[  741] = 1'b0;  wr_cycle[  741] = 1'b1;  addr_rom[  741]='h00000b94;  wr_data_rom[  741]='h000016b6;
    rd_cycle[  742] = 1'b0;  wr_cycle[  742] = 1'b1;  addr_rom[  742]='h00000b98;  wr_data_rom[  742]='h00000162;
    rd_cycle[  743] = 1'b0;  wr_cycle[  743] = 1'b1;  addr_rom[  743]='h00000b9c;  wr_data_rom[  743]='h00000f01;
    rd_cycle[  744] = 1'b0;  wr_cycle[  744] = 1'b1;  addr_rom[  744]='h00000ba0;  wr_data_rom[  744]='h00001d47;
    rd_cycle[  745] = 1'b0;  wr_cycle[  745] = 1'b1;  addr_rom[  745]='h00000ba4;  wr_data_rom[  745]='h0000014b;
    rd_cycle[  746] = 1'b0;  wr_cycle[  746] = 1'b1;  addr_rom[  746]='h00000ba8;  wr_data_rom[  746]='h00001a54;
    rd_cycle[  747] = 1'b0;  wr_cycle[  747] = 1'b1;  addr_rom[  747]='h00000bac;  wr_data_rom[  747]='h000001d2;
    rd_cycle[  748] = 1'b0;  wr_cycle[  748] = 1'b1;  addr_rom[  748]='h00000bb0;  wr_data_rom[  748]='h00001ba1;
    rd_cycle[  749] = 1'b0;  wr_cycle[  749] = 1'b1;  addr_rom[  749]='h00000bb4;  wr_data_rom[  749]='h0000160f;
    rd_cycle[  750] = 1'b0;  wr_cycle[  750] = 1'b1;  addr_rom[  750]='h00000bb8;  wr_data_rom[  750]='h000009b0;
    rd_cycle[  751] = 1'b0;  wr_cycle[  751] = 1'b1;  addr_rom[  751]='h00000bbc;  wr_data_rom[  751]='h00000c2c;
    rd_cycle[  752] = 1'b0;  wr_cycle[  752] = 1'b1;  addr_rom[  752]='h00000bc0;  wr_data_rom[  752]='h000008f6;
    rd_cycle[  753] = 1'b0;  wr_cycle[  753] = 1'b1;  addr_rom[  753]='h00000bc4;  wr_data_rom[  753]='h0000029e;
    rd_cycle[  754] = 1'b0;  wr_cycle[  754] = 1'b1;  addr_rom[  754]='h00000bc8;  wr_data_rom[  754]='h00000ac4;
    rd_cycle[  755] = 1'b0;  wr_cycle[  755] = 1'b1;  addr_rom[  755]='h00000bcc;  wr_data_rom[  755]='h00001478;
    rd_cycle[  756] = 1'b0;  wr_cycle[  756] = 1'b1;  addr_rom[  756]='h00000bd0;  wr_data_rom[  756]='h000000c2;
    rd_cycle[  757] = 1'b0;  wr_cycle[  757] = 1'b1;  addr_rom[  757]='h00000bd4;  wr_data_rom[  757]='h00000a8f;
    rd_cycle[  758] = 1'b0;  wr_cycle[  758] = 1'b1;  addr_rom[  758]='h00000bd8;  wr_data_rom[  758]='h0000063e;
    rd_cycle[  759] = 1'b0;  wr_cycle[  759] = 1'b1;  addr_rom[  759]='h00000bdc;  wr_data_rom[  759]='h00000e83;
    rd_cycle[  760] = 1'b0;  wr_cycle[  760] = 1'b1;  addr_rom[  760]='h00000be0;  wr_data_rom[  760]='h000008f6;
    rd_cycle[  761] = 1'b0;  wr_cycle[  761] = 1'b1;  addr_rom[  761]='h00000be4;  wr_data_rom[  761]='h000018ad;
    rd_cycle[  762] = 1'b0;  wr_cycle[  762] = 1'b1;  addr_rom[  762]='h00000be8;  wr_data_rom[  762]='h00001749;
    rd_cycle[  763] = 1'b0;  wr_cycle[  763] = 1'b1;  addr_rom[  763]='h00000bec;  wr_data_rom[  763]='h0000163f;
    rd_cycle[  764] = 1'b0;  wr_cycle[  764] = 1'b1;  addr_rom[  764]='h00000bf0;  wr_data_rom[  764]='h00000df3;
    rd_cycle[  765] = 1'b0;  wr_cycle[  765] = 1'b1;  addr_rom[  765]='h00000bf4;  wr_data_rom[  765]='h000011fd;
    rd_cycle[  766] = 1'b0;  wr_cycle[  766] = 1'b1;  addr_rom[  766]='h00000bf8;  wr_data_rom[  766]='h00001d45;
    rd_cycle[  767] = 1'b0;  wr_cycle[  767] = 1'b1;  addr_rom[  767]='h00000bfc;  wr_data_rom[  767]='h00001790;
    rd_cycle[  768] = 1'b0;  wr_cycle[  768] = 1'b1;  addr_rom[  768]='h00000c00;  wr_data_rom[  768]='h00001913;
    rd_cycle[  769] = 1'b0;  wr_cycle[  769] = 1'b1;  addr_rom[  769]='h00000c04;  wr_data_rom[  769]='h00000fa9;
    rd_cycle[  770] = 1'b0;  wr_cycle[  770] = 1'b1;  addr_rom[  770]='h00000c08;  wr_data_rom[  770]='h000015d8;
    rd_cycle[  771] = 1'b0;  wr_cycle[  771] = 1'b1;  addr_rom[  771]='h00000c0c;  wr_data_rom[  771]='h00000f1c;
    rd_cycle[  772] = 1'b0;  wr_cycle[  772] = 1'b1;  addr_rom[  772]='h00000c10;  wr_data_rom[  772]='h0000016a;
    rd_cycle[  773] = 1'b0;  wr_cycle[  773] = 1'b1;  addr_rom[  773]='h00000c14;  wr_data_rom[  773]='h000010a9;
    rd_cycle[  774] = 1'b0;  wr_cycle[  774] = 1'b1;  addr_rom[  774]='h00000c18;  wr_data_rom[  774]='h00001441;
    rd_cycle[  775] = 1'b0;  wr_cycle[  775] = 1'b1;  addr_rom[  775]='h00000c1c;  wr_data_rom[  775]='h000012fe;
    rd_cycle[  776] = 1'b0;  wr_cycle[  776] = 1'b1;  addr_rom[  776]='h00000c20;  wr_data_rom[  776]='h000001fa;
    rd_cycle[  777] = 1'b0;  wr_cycle[  777] = 1'b1;  addr_rom[  777]='h00000c24;  wr_data_rom[  777]='h0000044d;
    rd_cycle[  778] = 1'b0;  wr_cycle[  778] = 1'b1;  addr_rom[  778]='h00000c28;  wr_data_rom[  778]='h00000a5e;
    rd_cycle[  779] = 1'b0;  wr_cycle[  779] = 1'b1;  addr_rom[  779]='h00000c2c;  wr_data_rom[  779]='h000004f9;
    rd_cycle[  780] = 1'b0;  wr_cycle[  780] = 1'b1;  addr_rom[  780]='h00000c30;  wr_data_rom[  780]='h0000184c;
    rd_cycle[  781] = 1'b0;  wr_cycle[  781] = 1'b1;  addr_rom[  781]='h00000c34;  wr_data_rom[  781]='h00000c20;
    rd_cycle[  782] = 1'b0;  wr_cycle[  782] = 1'b1;  addr_rom[  782]='h00000c38;  wr_data_rom[  782]='h0000097d;
    rd_cycle[  783] = 1'b0;  wr_cycle[  783] = 1'b1;  addr_rom[  783]='h00000c3c;  wr_data_rom[  783]='h00001b06;
    rd_cycle[  784] = 1'b0;  wr_cycle[  784] = 1'b1;  addr_rom[  784]='h00000c40;  wr_data_rom[  784]='h00001c5b;
    rd_cycle[  785] = 1'b0;  wr_cycle[  785] = 1'b1;  addr_rom[  785]='h00000c44;  wr_data_rom[  785]='h00001217;
    rd_cycle[  786] = 1'b0;  wr_cycle[  786] = 1'b1;  addr_rom[  786]='h00000c48;  wr_data_rom[  786]='h00000176;
    rd_cycle[  787] = 1'b0;  wr_cycle[  787] = 1'b1;  addr_rom[  787]='h00000c4c;  wr_data_rom[  787]='h00001829;
    rd_cycle[  788] = 1'b0;  wr_cycle[  788] = 1'b1;  addr_rom[  788]='h00000c50;  wr_data_rom[  788]='h000016d3;
    rd_cycle[  789] = 1'b0;  wr_cycle[  789] = 1'b1;  addr_rom[  789]='h00000c54;  wr_data_rom[  789]='h00000d1d;
    rd_cycle[  790] = 1'b0;  wr_cycle[  790] = 1'b1;  addr_rom[  790]='h00000c58;  wr_data_rom[  790]='h000008a9;
    rd_cycle[  791] = 1'b0;  wr_cycle[  791] = 1'b1;  addr_rom[  791]='h00000c5c;  wr_data_rom[  791]='h00001c5b;
    rd_cycle[  792] = 1'b0;  wr_cycle[  792] = 1'b1;  addr_rom[  792]='h00000c60;  wr_data_rom[  792]='h000004f5;
    rd_cycle[  793] = 1'b0;  wr_cycle[  793] = 1'b1;  addr_rom[  793]='h00000c64;  wr_data_rom[  793]='h00001d65;
    rd_cycle[  794] = 1'b0;  wr_cycle[  794] = 1'b1;  addr_rom[  794]='h00000c68;  wr_data_rom[  794]='h00001e7a;
    rd_cycle[  795] = 1'b0;  wr_cycle[  795] = 1'b1;  addr_rom[  795]='h00000c6c;  wr_data_rom[  795]='h00000103;
    rd_cycle[  796] = 1'b0;  wr_cycle[  796] = 1'b1;  addr_rom[  796]='h00000c70;  wr_data_rom[  796]='h0000011c;
    rd_cycle[  797] = 1'b0;  wr_cycle[  797] = 1'b1;  addr_rom[  797]='h00000c74;  wr_data_rom[  797]='h0000196b;
    rd_cycle[  798] = 1'b0;  wr_cycle[  798] = 1'b1;  addr_rom[  798]='h00000c78;  wr_data_rom[  798]='h000007af;
    rd_cycle[  799] = 1'b0;  wr_cycle[  799] = 1'b1;  addr_rom[  799]='h00000c7c;  wr_data_rom[  799]='h000014c1;
    rd_cycle[  800] = 1'b0;  wr_cycle[  800] = 1'b1;  addr_rom[  800]='h00000c80;  wr_data_rom[  800]='h00001307;
    rd_cycle[  801] = 1'b0;  wr_cycle[  801] = 1'b1;  addr_rom[  801]='h00000c84;  wr_data_rom[  801]='h000007fc;
    rd_cycle[  802] = 1'b0;  wr_cycle[  802] = 1'b1;  addr_rom[  802]='h00000c88;  wr_data_rom[  802]='h00001902;
    rd_cycle[  803] = 1'b0;  wr_cycle[  803] = 1'b1;  addr_rom[  803]='h00000c8c;  wr_data_rom[  803]='h000019b3;
    rd_cycle[  804] = 1'b0;  wr_cycle[  804] = 1'b1;  addr_rom[  804]='h00000c90;  wr_data_rom[  804]='h000006dd;
    rd_cycle[  805] = 1'b0;  wr_cycle[  805] = 1'b1;  addr_rom[  805]='h00000c94;  wr_data_rom[  805]='h000013ea;
    rd_cycle[  806] = 1'b0;  wr_cycle[  806] = 1'b1;  addr_rom[  806]='h00000c98;  wr_data_rom[  806]='h00001be8;
    rd_cycle[  807] = 1'b0;  wr_cycle[  807] = 1'b1;  addr_rom[  807]='h00000c9c;  wr_data_rom[  807]='h000011f7;
    rd_cycle[  808] = 1'b0;  wr_cycle[  808] = 1'b1;  addr_rom[  808]='h00000ca0;  wr_data_rom[  808]='h00000aad;
    rd_cycle[  809] = 1'b0;  wr_cycle[  809] = 1'b1;  addr_rom[  809]='h00000ca4;  wr_data_rom[  809]='h000018c8;
    rd_cycle[  810] = 1'b0;  wr_cycle[  810] = 1'b1;  addr_rom[  810]='h00000ca8;  wr_data_rom[  810]='h00001730;
    rd_cycle[  811] = 1'b0;  wr_cycle[  811] = 1'b1;  addr_rom[  811]='h00000cac;  wr_data_rom[  811]='h00000dcb;
    rd_cycle[  812] = 1'b0;  wr_cycle[  812] = 1'b1;  addr_rom[  812]='h00000cb0;  wr_data_rom[  812]='h000014f9;
    rd_cycle[  813] = 1'b0;  wr_cycle[  813] = 1'b1;  addr_rom[  813]='h00000cb4;  wr_data_rom[  813]='h00000961;
    rd_cycle[  814] = 1'b0;  wr_cycle[  814] = 1'b1;  addr_rom[  814]='h00000cb8;  wr_data_rom[  814]='h00000b4a;
    rd_cycle[  815] = 1'b0;  wr_cycle[  815] = 1'b1;  addr_rom[  815]='h00000cbc;  wr_data_rom[  815]='h00000eca;
    rd_cycle[  816] = 1'b0;  wr_cycle[  816] = 1'b1;  addr_rom[  816]='h00000cc0;  wr_data_rom[  816]='h000011cd;
    rd_cycle[  817] = 1'b0;  wr_cycle[  817] = 1'b1;  addr_rom[  817]='h00000cc4;  wr_data_rom[  817]='h00000a6f;
    rd_cycle[  818] = 1'b0;  wr_cycle[  818] = 1'b1;  addr_rom[  818]='h00000cc8;  wr_data_rom[  818]='h00000c31;
    rd_cycle[  819] = 1'b0;  wr_cycle[  819] = 1'b1;  addr_rom[  819]='h00000ccc;  wr_data_rom[  819]='h00000ca0;
    rd_cycle[  820] = 1'b0;  wr_cycle[  820] = 1'b1;  addr_rom[  820]='h00000cd0;  wr_data_rom[  820]='h000002ee;
    rd_cycle[  821] = 1'b0;  wr_cycle[  821] = 1'b1;  addr_rom[  821]='h00000cd4;  wr_data_rom[  821]='h00000173;
    rd_cycle[  822] = 1'b0;  wr_cycle[  822] = 1'b1;  addr_rom[  822]='h00000cd8;  wr_data_rom[  822]='h00000b5d;
    rd_cycle[  823] = 1'b0;  wr_cycle[  823] = 1'b1;  addr_rom[  823]='h00000cdc;  wr_data_rom[  823]='h000005ef;
    rd_cycle[  824] = 1'b0;  wr_cycle[  824] = 1'b1;  addr_rom[  824]='h00000ce0;  wr_data_rom[  824]='h00000a8b;
    rd_cycle[  825] = 1'b0;  wr_cycle[  825] = 1'b1;  addr_rom[  825]='h00000ce4;  wr_data_rom[  825]='h000008ca;
    rd_cycle[  826] = 1'b0;  wr_cycle[  826] = 1'b1;  addr_rom[  826]='h00000ce8;  wr_data_rom[  826]='h00000b7c;
    rd_cycle[  827] = 1'b0;  wr_cycle[  827] = 1'b1;  addr_rom[  827]='h00000cec;  wr_data_rom[  827]='h0000134e;
    rd_cycle[  828] = 1'b0;  wr_cycle[  828] = 1'b1;  addr_rom[  828]='h00000cf0;  wr_data_rom[  828]='h00001acc;
    rd_cycle[  829] = 1'b0;  wr_cycle[  829] = 1'b1;  addr_rom[  829]='h00000cf4;  wr_data_rom[  829]='h00001ab2;
    rd_cycle[  830] = 1'b0;  wr_cycle[  830] = 1'b1;  addr_rom[  830]='h00000cf8;  wr_data_rom[  830]='h00001da1;
    rd_cycle[  831] = 1'b0;  wr_cycle[  831] = 1'b1;  addr_rom[  831]='h00000cfc;  wr_data_rom[  831]='h000001ff;
    rd_cycle[  832] = 1'b0;  wr_cycle[  832] = 1'b1;  addr_rom[  832]='h00000d00;  wr_data_rom[  832]='h000002b5;
    rd_cycle[  833] = 1'b0;  wr_cycle[  833] = 1'b1;  addr_rom[  833]='h00000d04;  wr_data_rom[  833]='h000014df;
    rd_cycle[  834] = 1'b0;  wr_cycle[  834] = 1'b1;  addr_rom[  834]='h00000d08;  wr_data_rom[  834]='h00000d7e;
    rd_cycle[  835] = 1'b0;  wr_cycle[  835] = 1'b1;  addr_rom[  835]='h00000d0c;  wr_data_rom[  835]='h0000090e;
    rd_cycle[  836] = 1'b0;  wr_cycle[  836] = 1'b1;  addr_rom[  836]='h00000d10;  wr_data_rom[  836]='h00000bb5;
    rd_cycle[  837] = 1'b0;  wr_cycle[  837] = 1'b1;  addr_rom[  837]='h00000d14;  wr_data_rom[  837]='h000010fb;
    rd_cycle[  838] = 1'b0;  wr_cycle[  838] = 1'b1;  addr_rom[  838]='h00000d18;  wr_data_rom[  838]='h0000191a;
    rd_cycle[  839] = 1'b0;  wr_cycle[  839] = 1'b1;  addr_rom[  839]='h00000d1c;  wr_data_rom[  839]='h000014f2;
    rd_cycle[  840] = 1'b0;  wr_cycle[  840] = 1'b1;  addr_rom[  840]='h00000d20;  wr_data_rom[  840]='h0000084d;
    rd_cycle[  841] = 1'b0;  wr_cycle[  841] = 1'b1;  addr_rom[  841]='h00000d24;  wr_data_rom[  841]='h000010a0;
    rd_cycle[  842] = 1'b0;  wr_cycle[  842] = 1'b1;  addr_rom[  842]='h00000d28;  wr_data_rom[  842]='h0000174c;
    rd_cycle[  843] = 1'b0;  wr_cycle[  843] = 1'b1;  addr_rom[  843]='h00000d2c;  wr_data_rom[  843]='h0000142e;
    rd_cycle[  844] = 1'b0;  wr_cycle[  844] = 1'b1;  addr_rom[  844]='h00000d30;  wr_data_rom[  844]='h00000bbf;
    rd_cycle[  845] = 1'b0;  wr_cycle[  845] = 1'b1;  addr_rom[  845]='h00000d34;  wr_data_rom[  845]='h000019fa;
    rd_cycle[  846] = 1'b0;  wr_cycle[  846] = 1'b1;  addr_rom[  846]='h00000d38;  wr_data_rom[  846]='h00001b77;
    rd_cycle[  847] = 1'b0;  wr_cycle[  847] = 1'b1;  addr_rom[  847]='h00000d3c;  wr_data_rom[  847]='h000010dd;
    rd_cycle[  848] = 1'b0;  wr_cycle[  848] = 1'b1;  addr_rom[  848]='h00000d40;  wr_data_rom[  848]='h000002ec;
    rd_cycle[  849] = 1'b0;  wr_cycle[  849] = 1'b1;  addr_rom[  849]='h00000d44;  wr_data_rom[  849]='h00000d2b;
    rd_cycle[  850] = 1'b0;  wr_cycle[  850] = 1'b1;  addr_rom[  850]='h00000d48;  wr_data_rom[  850]='h00001b42;
    rd_cycle[  851] = 1'b0;  wr_cycle[  851] = 1'b1;  addr_rom[  851]='h00000d4c;  wr_data_rom[  851]='h00000a55;
    rd_cycle[  852] = 1'b0;  wr_cycle[  852] = 1'b1;  addr_rom[  852]='h00000d50;  wr_data_rom[  852]='h00001ba6;
    rd_cycle[  853] = 1'b0;  wr_cycle[  853] = 1'b1;  addr_rom[  853]='h00000d54;  wr_data_rom[  853]='h00001eed;
    rd_cycle[  854] = 1'b0;  wr_cycle[  854] = 1'b1;  addr_rom[  854]='h00000d58;  wr_data_rom[  854]='h0000161c;
    rd_cycle[  855] = 1'b0;  wr_cycle[  855] = 1'b1;  addr_rom[  855]='h00000d5c;  wr_data_rom[  855]='h00001c7a;
    rd_cycle[  856] = 1'b0;  wr_cycle[  856] = 1'b1;  addr_rom[  856]='h00000d60;  wr_data_rom[  856]='h00001445;
    rd_cycle[  857] = 1'b0;  wr_cycle[  857] = 1'b1;  addr_rom[  857]='h00000d64;  wr_data_rom[  857]='h0000084f;
    rd_cycle[  858] = 1'b0;  wr_cycle[  858] = 1'b1;  addr_rom[  858]='h00000d68;  wr_data_rom[  858]='h00001bdc;
    rd_cycle[  859] = 1'b0;  wr_cycle[  859] = 1'b1;  addr_rom[  859]='h00000d6c;  wr_data_rom[  859]='h000000e6;
    rd_cycle[  860] = 1'b0;  wr_cycle[  860] = 1'b1;  addr_rom[  860]='h00000d70;  wr_data_rom[  860]='h00001426;
    rd_cycle[  861] = 1'b0;  wr_cycle[  861] = 1'b1;  addr_rom[  861]='h00000d74;  wr_data_rom[  861]='h0000092c;
    rd_cycle[  862] = 1'b0;  wr_cycle[  862] = 1'b1;  addr_rom[  862]='h00000d78;  wr_data_rom[  862]='h00001d01;
    rd_cycle[  863] = 1'b0;  wr_cycle[  863] = 1'b1;  addr_rom[  863]='h00000d7c;  wr_data_rom[  863]='h00000e2a;
    rd_cycle[  864] = 1'b0;  wr_cycle[  864] = 1'b1;  addr_rom[  864]='h00000d80;  wr_data_rom[  864]='h00000ecd;
    rd_cycle[  865] = 1'b0;  wr_cycle[  865] = 1'b1;  addr_rom[  865]='h00000d84;  wr_data_rom[  865]='h00001a27;
    rd_cycle[  866] = 1'b0;  wr_cycle[  866] = 1'b1;  addr_rom[  866]='h00000d88;  wr_data_rom[  866]='h000016b8;
    rd_cycle[  867] = 1'b0;  wr_cycle[  867] = 1'b1;  addr_rom[  867]='h00000d8c;  wr_data_rom[  867]='h0000079a;
    rd_cycle[  868] = 1'b0;  wr_cycle[  868] = 1'b1;  addr_rom[  868]='h00000d90;  wr_data_rom[  868]='h00000fb2;
    rd_cycle[  869] = 1'b0;  wr_cycle[  869] = 1'b1;  addr_rom[  869]='h00000d94;  wr_data_rom[  869]='h0000106b;
    rd_cycle[  870] = 1'b0;  wr_cycle[  870] = 1'b1;  addr_rom[  870]='h00000d98;  wr_data_rom[  870]='h000000c8;
    rd_cycle[  871] = 1'b0;  wr_cycle[  871] = 1'b1;  addr_rom[  871]='h00000d9c;  wr_data_rom[  871]='h0000074f;
    rd_cycle[  872] = 1'b0;  wr_cycle[  872] = 1'b1;  addr_rom[  872]='h00000da0;  wr_data_rom[  872]='h00001a61;
    rd_cycle[  873] = 1'b0;  wr_cycle[  873] = 1'b1;  addr_rom[  873]='h00000da4;  wr_data_rom[  873]='h0000137d;
    rd_cycle[  874] = 1'b0;  wr_cycle[  874] = 1'b1;  addr_rom[  874]='h00000da8;  wr_data_rom[  874]='h0000093a;
    rd_cycle[  875] = 1'b0;  wr_cycle[  875] = 1'b1;  addr_rom[  875]='h00000dac;  wr_data_rom[  875]='h00001438;
    rd_cycle[  876] = 1'b0;  wr_cycle[  876] = 1'b1;  addr_rom[  876]='h00000db0;  wr_data_rom[  876]='h00001a11;
    rd_cycle[  877] = 1'b0;  wr_cycle[  877] = 1'b1;  addr_rom[  877]='h00000db4;  wr_data_rom[  877]='h00001a11;
    rd_cycle[  878] = 1'b0;  wr_cycle[  878] = 1'b1;  addr_rom[  878]='h00000db8;  wr_data_rom[  878]='h00000291;
    rd_cycle[  879] = 1'b0;  wr_cycle[  879] = 1'b1;  addr_rom[  879]='h00000dbc;  wr_data_rom[  879]='h000010c0;
    rd_cycle[  880] = 1'b0;  wr_cycle[  880] = 1'b1;  addr_rom[  880]='h00000dc0;  wr_data_rom[  880]='h00000429;
    rd_cycle[  881] = 1'b0;  wr_cycle[  881] = 1'b1;  addr_rom[  881]='h00000dc4;  wr_data_rom[  881]='h0000097b;
    rd_cycle[  882] = 1'b0;  wr_cycle[  882] = 1'b1;  addr_rom[  882]='h00000dc8;  wr_data_rom[  882]='h00000bec;
    rd_cycle[  883] = 1'b0;  wr_cycle[  883] = 1'b1;  addr_rom[  883]='h00000dcc;  wr_data_rom[  883]='h00001586;
    rd_cycle[  884] = 1'b0;  wr_cycle[  884] = 1'b1;  addr_rom[  884]='h00000dd0;  wr_data_rom[  884]='h00000200;
    rd_cycle[  885] = 1'b0;  wr_cycle[  885] = 1'b1;  addr_rom[  885]='h00000dd4;  wr_data_rom[  885]='h00001214;
    rd_cycle[  886] = 1'b0;  wr_cycle[  886] = 1'b1;  addr_rom[  886]='h00000dd8;  wr_data_rom[  886]='h00000c2f;
    rd_cycle[  887] = 1'b0;  wr_cycle[  887] = 1'b1;  addr_rom[  887]='h00000ddc;  wr_data_rom[  887]='h0000100d;
    rd_cycle[  888] = 1'b0;  wr_cycle[  888] = 1'b1;  addr_rom[  888]='h00000de0;  wr_data_rom[  888]='h000007d9;
    rd_cycle[  889] = 1'b0;  wr_cycle[  889] = 1'b1;  addr_rom[  889]='h00000de4;  wr_data_rom[  889]='h00000763;
    rd_cycle[  890] = 1'b0;  wr_cycle[  890] = 1'b1;  addr_rom[  890]='h00000de8;  wr_data_rom[  890]='h00001592;
    rd_cycle[  891] = 1'b0;  wr_cycle[  891] = 1'b1;  addr_rom[  891]='h00000dec;  wr_data_rom[  891]='h00001ce6;
    rd_cycle[  892] = 1'b0;  wr_cycle[  892] = 1'b1;  addr_rom[  892]='h00000df0;  wr_data_rom[  892]='h00000356;
    rd_cycle[  893] = 1'b0;  wr_cycle[  893] = 1'b1;  addr_rom[  893]='h00000df4;  wr_data_rom[  893]='h000010cb;
    rd_cycle[  894] = 1'b0;  wr_cycle[  894] = 1'b1;  addr_rom[  894]='h00000df8;  wr_data_rom[  894]='h00001a93;
    rd_cycle[  895] = 1'b0;  wr_cycle[  895] = 1'b1;  addr_rom[  895]='h00000dfc;  wr_data_rom[  895]='h00001d65;
    rd_cycle[  896] = 1'b0;  wr_cycle[  896] = 1'b1;  addr_rom[  896]='h00000e00;  wr_data_rom[  896]='h000013c5;
    rd_cycle[  897] = 1'b0;  wr_cycle[  897] = 1'b1;  addr_rom[  897]='h00000e04;  wr_data_rom[  897]='h00001d39;
    rd_cycle[  898] = 1'b0;  wr_cycle[  898] = 1'b1;  addr_rom[  898]='h00000e08;  wr_data_rom[  898]='h00000884;
    rd_cycle[  899] = 1'b0;  wr_cycle[  899] = 1'b1;  addr_rom[  899]='h00000e0c;  wr_data_rom[  899]='h00000cce;
    rd_cycle[  900] = 1'b0;  wr_cycle[  900] = 1'b1;  addr_rom[  900]='h00000e10;  wr_data_rom[  900]='h0000005c;
    rd_cycle[  901] = 1'b0;  wr_cycle[  901] = 1'b1;  addr_rom[  901]='h00000e14;  wr_data_rom[  901]='h00000910;
    rd_cycle[  902] = 1'b0;  wr_cycle[  902] = 1'b1;  addr_rom[  902]='h00000e18;  wr_data_rom[  902]='h000012c4;
    rd_cycle[  903] = 1'b0;  wr_cycle[  903] = 1'b1;  addr_rom[  903]='h00000e1c;  wr_data_rom[  903]='h00000b42;
    rd_cycle[  904] = 1'b0;  wr_cycle[  904] = 1'b1;  addr_rom[  904]='h00000e20;  wr_data_rom[  904]='h000000aa;
    rd_cycle[  905] = 1'b0;  wr_cycle[  905] = 1'b1;  addr_rom[  905]='h00000e24;  wr_data_rom[  905]='h00001802;
    rd_cycle[  906] = 1'b0;  wr_cycle[  906] = 1'b1;  addr_rom[  906]='h00000e28;  wr_data_rom[  906]='h00000237;
    rd_cycle[  907] = 1'b0;  wr_cycle[  907] = 1'b1;  addr_rom[  907]='h00000e2c;  wr_data_rom[  907]='h000016ce;
    rd_cycle[  908] = 1'b0;  wr_cycle[  908] = 1'b1;  addr_rom[  908]='h00000e30;  wr_data_rom[  908]='h000006e0;
    rd_cycle[  909] = 1'b0;  wr_cycle[  909] = 1'b1;  addr_rom[  909]='h00000e34;  wr_data_rom[  909]='h0000143e;
    rd_cycle[  910] = 1'b0;  wr_cycle[  910] = 1'b1;  addr_rom[  910]='h00000e38;  wr_data_rom[  910]='h00001bc1;
    rd_cycle[  911] = 1'b0;  wr_cycle[  911] = 1'b1;  addr_rom[  911]='h00000e3c;  wr_data_rom[  911]='h000002f4;
    rd_cycle[  912] = 1'b0;  wr_cycle[  912] = 1'b1;  addr_rom[  912]='h00000e40;  wr_data_rom[  912]='h000002c2;
    rd_cycle[  913] = 1'b0;  wr_cycle[  913] = 1'b1;  addr_rom[  913]='h00000e44;  wr_data_rom[  913]='h00000992;
    rd_cycle[  914] = 1'b0;  wr_cycle[  914] = 1'b1;  addr_rom[  914]='h00000e48;  wr_data_rom[  914]='h00001267;
    rd_cycle[  915] = 1'b0;  wr_cycle[  915] = 1'b1;  addr_rom[  915]='h00000e4c;  wr_data_rom[  915]='h00000497;
    rd_cycle[  916] = 1'b0;  wr_cycle[  916] = 1'b1;  addr_rom[  916]='h00000e50;  wr_data_rom[  916]='h000005e6;
    rd_cycle[  917] = 1'b0;  wr_cycle[  917] = 1'b1;  addr_rom[  917]='h00000e54;  wr_data_rom[  917]='h0000096e;
    rd_cycle[  918] = 1'b0;  wr_cycle[  918] = 1'b1;  addr_rom[  918]='h00000e58;  wr_data_rom[  918]='h000013fd;
    rd_cycle[  919] = 1'b0;  wr_cycle[  919] = 1'b1;  addr_rom[  919]='h00000e5c;  wr_data_rom[  919]='h000002a1;
    rd_cycle[  920] = 1'b0;  wr_cycle[  920] = 1'b1;  addr_rom[  920]='h00000e60;  wr_data_rom[  920]='h00001700;
    rd_cycle[  921] = 1'b0;  wr_cycle[  921] = 1'b1;  addr_rom[  921]='h00000e64;  wr_data_rom[  921]='h000018e9;
    rd_cycle[  922] = 1'b0;  wr_cycle[  922] = 1'b1;  addr_rom[  922]='h00000e68;  wr_data_rom[  922]='h000008fe;
    rd_cycle[  923] = 1'b0;  wr_cycle[  923] = 1'b1;  addr_rom[  923]='h00000e6c;  wr_data_rom[  923]='h00001e9b;
    rd_cycle[  924] = 1'b0;  wr_cycle[  924] = 1'b1;  addr_rom[  924]='h00000e70;  wr_data_rom[  924]='h000002bc;
    rd_cycle[  925] = 1'b0;  wr_cycle[  925] = 1'b1;  addr_rom[  925]='h00000e74;  wr_data_rom[  925]='h000014a0;
    rd_cycle[  926] = 1'b0;  wr_cycle[  926] = 1'b1;  addr_rom[  926]='h00000e78;  wr_data_rom[  926]='h000001a4;
    rd_cycle[  927] = 1'b0;  wr_cycle[  927] = 1'b1;  addr_rom[  927]='h00000e7c;  wr_data_rom[  927]='h00000536;
    rd_cycle[  928] = 1'b0;  wr_cycle[  928] = 1'b1;  addr_rom[  928]='h00000e80;  wr_data_rom[  928]='h00000322;
    rd_cycle[  929] = 1'b0;  wr_cycle[  929] = 1'b1;  addr_rom[  929]='h00000e84;  wr_data_rom[  929]='h00001294;
    rd_cycle[  930] = 1'b0;  wr_cycle[  930] = 1'b1;  addr_rom[  930]='h00000e88;  wr_data_rom[  930]='h00000b0d;
    rd_cycle[  931] = 1'b0;  wr_cycle[  931] = 1'b1;  addr_rom[  931]='h00000e8c;  wr_data_rom[  931]='h00000ed7;
    rd_cycle[  932] = 1'b0;  wr_cycle[  932] = 1'b1;  addr_rom[  932]='h00000e90;  wr_data_rom[  932]='h00000e42;
    rd_cycle[  933] = 1'b0;  wr_cycle[  933] = 1'b1;  addr_rom[  933]='h00000e94;  wr_data_rom[  933]='h00000a07;
    rd_cycle[  934] = 1'b0;  wr_cycle[  934] = 1'b1;  addr_rom[  934]='h00000e98;  wr_data_rom[  934]='h00001459;
    rd_cycle[  935] = 1'b0;  wr_cycle[  935] = 1'b1;  addr_rom[  935]='h00000e9c;  wr_data_rom[  935]='h0000057e;
    rd_cycle[  936] = 1'b0;  wr_cycle[  936] = 1'b1;  addr_rom[  936]='h00000ea0;  wr_data_rom[  936]='h00000031;
    rd_cycle[  937] = 1'b0;  wr_cycle[  937] = 1'b1;  addr_rom[  937]='h00000ea4;  wr_data_rom[  937]='h0000101e;
    rd_cycle[  938] = 1'b0;  wr_cycle[  938] = 1'b1;  addr_rom[  938]='h00000ea8;  wr_data_rom[  938]='h000011dd;
    rd_cycle[  939] = 1'b0;  wr_cycle[  939] = 1'b1;  addr_rom[  939]='h00000eac;  wr_data_rom[  939]='h00001093;
    rd_cycle[  940] = 1'b0;  wr_cycle[  940] = 1'b1;  addr_rom[  940]='h00000eb0;  wr_data_rom[  940]='h0000004e;
    rd_cycle[  941] = 1'b0;  wr_cycle[  941] = 1'b1;  addr_rom[  941]='h00000eb4;  wr_data_rom[  941]='h000013d0;
    rd_cycle[  942] = 1'b0;  wr_cycle[  942] = 1'b1;  addr_rom[  942]='h00000eb8;  wr_data_rom[  942]='h000010b7;
    rd_cycle[  943] = 1'b0;  wr_cycle[  943] = 1'b1;  addr_rom[  943]='h00000ebc;  wr_data_rom[  943]='h00000ff8;
    rd_cycle[  944] = 1'b0;  wr_cycle[  944] = 1'b1;  addr_rom[  944]='h00000ec0;  wr_data_rom[  944]='h00000277;
    rd_cycle[  945] = 1'b0;  wr_cycle[  945] = 1'b1;  addr_rom[  945]='h00000ec4;  wr_data_rom[  945]='h0000040d;
    rd_cycle[  946] = 1'b0;  wr_cycle[  946] = 1'b1;  addr_rom[  946]='h00000ec8;  wr_data_rom[  946]='h0000019c;
    rd_cycle[  947] = 1'b0;  wr_cycle[  947] = 1'b1;  addr_rom[  947]='h00000ecc;  wr_data_rom[  947]='h00001552;
    rd_cycle[  948] = 1'b0;  wr_cycle[  948] = 1'b1;  addr_rom[  948]='h00000ed0;  wr_data_rom[  948]='h00001400;
    rd_cycle[  949] = 1'b0;  wr_cycle[  949] = 1'b1;  addr_rom[  949]='h00000ed4;  wr_data_rom[  949]='h00000623;
    rd_cycle[  950] = 1'b0;  wr_cycle[  950] = 1'b1;  addr_rom[  950]='h00000ed8;  wr_data_rom[  950]='h00000151;
    rd_cycle[  951] = 1'b0;  wr_cycle[  951] = 1'b1;  addr_rom[  951]='h00000edc;  wr_data_rom[  951]='h00000921;
    rd_cycle[  952] = 1'b0;  wr_cycle[  952] = 1'b1;  addr_rom[  952]='h00000ee0;  wr_data_rom[  952]='h00001a90;
    rd_cycle[  953] = 1'b0;  wr_cycle[  953] = 1'b1;  addr_rom[  953]='h00000ee4;  wr_data_rom[  953]='h00001082;
    rd_cycle[  954] = 1'b0;  wr_cycle[  954] = 1'b1;  addr_rom[  954]='h00000ee8;  wr_data_rom[  954]='h00001caf;
    rd_cycle[  955] = 1'b0;  wr_cycle[  955] = 1'b1;  addr_rom[  955]='h00000eec;  wr_data_rom[  955]='h000007ca;
    rd_cycle[  956] = 1'b0;  wr_cycle[  956] = 1'b1;  addr_rom[  956]='h00000ef0;  wr_data_rom[  956]='h00001c95;
    rd_cycle[  957] = 1'b0;  wr_cycle[  957] = 1'b1;  addr_rom[  957]='h00000ef4;  wr_data_rom[  957]='h00001a03;
    rd_cycle[  958] = 1'b0;  wr_cycle[  958] = 1'b1;  addr_rom[  958]='h00000ef8;  wr_data_rom[  958]='h0000187e;
    rd_cycle[  959] = 1'b0;  wr_cycle[  959] = 1'b1;  addr_rom[  959]='h00000efc;  wr_data_rom[  959]='h00000443;
    rd_cycle[  960] = 1'b0;  wr_cycle[  960] = 1'b1;  addr_rom[  960]='h00000f00;  wr_data_rom[  960]='h000019fa;
    rd_cycle[  961] = 1'b0;  wr_cycle[  961] = 1'b1;  addr_rom[  961]='h00000f04;  wr_data_rom[  961]='h00001d9f;
    rd_cycle[  962] = 1'b0;  wr_cycle[  962] = 1'b1;  addr_rom[  962]='h00000f08;  wr_data_rom[  962]='h00000c40;
    rd_cycle[  963] = 1'b0;  wr_cycle[  963] = 1'b1;  addr_rom[  963]='h00000f0c;  wr_data_rom[  963]='h00001904;
    rd_cycle[  964] = 1'b0;  wr_cycle[  964] = 1'b1;  addr_rom[  964]='h00000f10;  wr_data_rom[  964]='h0000144b;
    rd_cycle[  965] = 1'b0;  wr_cycle[  965] = 1'b1;  addr_rom[  965]='h00000f14;  wr_data_rom[  965]='h00000f7b;
    rd_cycle[  966] = 1'b0;  wr_cycle[  966] = 1'b1;  addr_rom[  966]='h00000f18;  wr_data_rom[  966]='h000019a0;
    rd_cycle[  967] = 1'b0;  wr_cycle[  967] = 1'b1;  addr_rom[  967]='h00000f1c;  wr_data_rom[  967]='h0000017f;
    rd_cycle[  968] = 1'b0;  wr_cycle[  968] = 1'b1;  addr_rom[  968]='h00000f20;  wr_data_rom[  968]='h0000024a;
    rd_cycle[  969] = 1'b0;  wr_cycle[  969] = 1'b1;  addr_rom[  969]='h00000f24;  wr_data_rom[  969]='h0000070b;
    rd_cycle[  970] = 1'b0;  wr_cycle[  970] = 1'b1;  addr_rom[  970]='h00000f28;  wr_data_rom[  970]='h00001a7b;
    rd_cycle[  971] = 1'b0;  wr_cycle[  971] = 1'b1;  addr_rom[  971]='h00000f2c;  wr_data_rom[  971]='h0000055c;
    rd_cycle[  972] = 1'b0;  wr_cycle[  972] = 1'b1;  addr_rom[  972]='h00000f30;  wr_data_rom[  972]='h00000afa;
    rd_cycle[  973] = 1'b0;  wr_cycle[  973] = 1'b1;  addr_rom[  973]='h00000f34;  wr_data_rom[  973]='h0000055a;
    rd_cycle[  974] = 1'b0;  wr_cycle[  974] = 1'b1;  addr_rom[  974]='h00000f38;  wr_data_rom[  974]='h00000edb;
    rd_cycle[  975] = 1'b0;  wr_cycle[  975] = 1'b1;  addr_rom[  975]='h00000f3c;  wr_data_rom[  975]='h00000441;
    rd_cycle[  976] = 1'b0;  wr_cycle[  976] = 1'b1;  addr_rom[  976]='h00000f40;  wr_data_rom[  976]='h00000231;
    rd_cycle[  977] = 1'b0;  wr_cycle[  977] = 1'b1;  addr_rom[  977]='h00000f44;  wr_data_rom[  977]='h000010e0;
    rd_cycle[  978] = 1'b0;  wr_cycle[  978] = 1'b1;  addr_rom[  978]='h00000f48;  wr_data_rom[  978]='h000004b3;
    rd_cycle[  979] = 1'b0;  wr_cycle[  979] = 1'b1;  addr_rom[  979]='h00000f4c;  wr_data_rom[  979]='h000007d0;
    rd_cycle[  980] = 1'b0;  wr_cycle[  980] = 1'b1;  addr_rom[  980]='h00000f50;  wr_data_rom[  980]='h00000dec;
    rd_cycle[  981] = 1'b0;  wr_cycle[  981] = 1'b1;  addr_rom[  981]='h00000f54;  wr_data_rom[  981]='h00000b53;
    rd_cycle[  982] = 1'b0;  wr_cycle[  982] = 1'b1;  addr_rom[  982]='h00000f58;  wr_data_rom[  982]='h000019d5;
    rd_cycle[  983] = 1'b0;  wr_cycle[  983] = 1'b1;  addr_rom[  983]='h00000f5c;  wr_data_rom[  983]='h00000ed2;
    rd_cycle[  984] = 1'b0;  wr_cycle[  984] = 1'b1;  addr_rom[  984]='h00000f60;  wr_data_rom[  984]='h00000c06;
    rd_cycle[  985] = 1'b0;  wr_cycle[  985] = 1'b1;  addr_rom[  985]='h00000f64;  wr_data_rom[  985]='h00001362;
    rd_cycle[  986] = 1'b0;  wr_cycle[  986] = 1'b1;  addr_rom[  986]='h00000f68;  wr_data_rom[  986]='h00000ea5;
    rd_cycle[  987] = 1'b0;  wr_cycle[  987] = 1'b1;  addr_rom[  987]='h00000f6c;  wr_data_rom[  987]='h000018c9;
    rd_cycle[  988] = 1'b0;  wr_cycle[  988] = 1'b1;  addr_rom[  988]='h00000f70;  wr_data_rom[  988]='h00001893;
    rd_cycle[  989] = 1'b0;  wr_cycle[  989] = 1'b1;  addr_rom[  989]='h00000f74;  wr_data_rom[  989]='h00001a3d;
    rd_cycle[  990] = 1'b0;  wr_cycle[  990] = 1'b1;  addr_rom[  990]='h00000f78;  wr_data_rom[  990]='h00001ac5;
    rd_cycle[  991] = 1'b0;  wr_cycle[  991] = 1'b1;  addr_rom[  991]='h00000f7c;  wr_data_rom[  991]='h000018a7;
    rd_cycle[  992] = 1'b0;  wr_cycle[  992] = 1'b1;  addr_rom[  992]='h00000f80;  wr_data_rom[  992]='h00001734;
    rd_cycle[  993] = 1'b0;  wr_cycle[  993] = 1'b1;  addr_rom[  993]='h00000f84;  wr_data_rom[  993]='h000009d5;
    rd_cycle[  994] = 1'b0;  wr_cycle[  994] = 1'b1;  addr_rom[  994]='h00000f88;  wr_data_rom[  994]='h000016a3;
    rd_cycle[  995] = 1'b0;  wr_cycle[  995] = 1'b1;  addr_rom[  995]='h00000f8c;  wr_data_rom[  995]='h000002df;
    rd_cycle[  996] = 1'b0;  wr_cycle[  996] = 1'b1;  addr_rom[  996]='h00000f90;  wr_data_rom[  996]='h00001991;
    rd_cycle[  997] = 1'b0;  wr_cycle[  997] = 1'b1;  addr_rom[  997]='h00000f94;  wr_data_rom[  997]='h00001e59;
    rd_cycle[  998] = 1'b0;  wr_cycle[  998] = 1'b1;  addr_rom[  998]='h00000f98;  wr_data_rom[  998]='h00001724;
    rd_cycle[  999] = 1'b0;  wr_cycle[  999] = 1'b1;  addr_rom[  999]='h00000f9c;  wr_data_rom[  999]='h000017de;
    rd_cycle[ 1000] = 1'b0;  wr_cycle[ 1000] = 1'b1;  addr_rom[ 1000]='h00000fa0;  wr_data_rom[ 1000]='h00001525;
    rd_cycle[ 1001] = 1'b0;  wr_cycle[ 1001] = 1'b1;  addr_rom[ 1001]='h00000fa4;  wr_data_rom[ 1001]='h00001c99;
    rd_cycle[ 1002] = 1'b0;  wr_cycle[ 1002] = 1'b1;  addr_rom[ 1002]='h00000fa8;  wr_data_rom[ 1002]='h00001603;
    rd_cycle[ 1003] = 1'b0;  wr_cycle[ 1003] = 1'b1;  addr_rom[ 1003]='h00000fac;  wr_data_rom[ 1003]='h0000142f;
    rd_cycle[ 1004] = 1'b0;  wr_cycle[ 1004] = 1'b1;  addr_rom[ 1004]='h00000fb0;  wr_data_rom[ 1004]='h00000894;
    rd_cycle[ 1005] = 1'b0;  wr_cycle[ 1005] = 1'b1;  addr_rom[ 1005]='h00000fb4;  wr_data_rom[ 1005]='h00001604;
    rd_cycle[ 1006] = 1'b0;  wr_cycle[ 1006] = 1'b1;  addr_rom[ 1006]='h00000fb8;  wr_data_rom[ 1006]='h0000180e;
    rd_cycle[ 1007] = 1'b0;  wr_cycle[ 1007] = 1'b1;  addr_rom[ 1007]='h00000fbc;  wr_data_rom[ 1007]='h00000984;
    rd_cycle[ 1008] = 1'b0;  wr_cycle[ 1008] = 1'b1;  addr_rom[ 1008]='h00000fc0;  wr_data_rom[ 1008]='h00000a99;
    rd_cycle[ 1009] = 1'b0;  wr_cycle[ 1009] = 1'b1;  addr_rom[ 1009]='h00000fc4;  wr_data_rom[ 1009]='h00001506;
    rd_cycle[ 1010] = 1'b0;  wr_cycle[ 1010] = 1'b1;  addr_rom[ 1010]='h00000fc8;  wr_data_rom[ 1010]='h00000047;
    rd_cycle[ 1011] = 1'b0;  wr_cycle[ 1011] = 1'b1;  addr_rom[ 1011]='h00000fcc;  wr_data_rom[ 1011]='h0000156e;
    rd_cycle[ 1012] = 1'b0;  wr_cycle[ 1012] = 1'b1;  addr_rom[ 1012]='h00000fd0;  wr_data_rom[ 1012]='h00001158;
    rd_cycle[ 1013] = 1'b0;  wr_cycle[ 1013] = 1'b1;  addr_rom[ 1013]='h00000fd4;  wr_data_rom[ 1013]='h00001b1f;
    rd_cycle[ 1014] = 1'b0;  wr_cycle[ 1014] = 1'b1;  addr_rom[ 1014]='h00000fd8;  wr_data_rom[ 1014]='h00001437;
    rd_cycle[ 1015] = 1'b0;  wr_cycle[ 1015] = 1'b1;  addr_rom[ 1015]='h00000fdc;  wr_data_rom[ 1015]='h00001a29;
    rd_cycle[ 1016] = 1'b0;  wr_cycle[ 1016] = 1'b1;  addr_rom[ 1016]='h00000fe0;  wr_data_rom[ 1016]='h00000558;
    rd_cycle[ 1017] = 1'b0;  wr_cycle[ 1017] = 1'b1;  addr_rom[ 1017]='h00000fe4;  wr_data_rom[ 1017]='h000017f0;
    rd_cycle[ 1018] = 1'b0;  wr_cycle[ 1018] = 1'b1;  addr_rom[ 1018]='h00000fe8;  wr_data_rom[ 1018]='h00000b28;
    rd_cycle[ 1019] = 1'b0;  wr_cycle[ 1019] = 1'b1;  addr_rom[ 1019]='h00000fec;  wr_data_rom[ 1019]='h0000033e;
    rd_cycle[ 1020] = 1'b0;  wr_cycle[ 1020] = 1'b1;  addr_rom[ 1020]='h00000ff0;  wr_data_rom[ 1020]='h000007c0;
    rd_cycle[ 1021] = 1'b0;  wr_cycle[ 1021] = 1'b1;  addr_rom[ 1021]='h00000ff4;  wr_data_rom[ 1021]='h000012da;
    rd_cycle[ 1022] = 1'b0;  wr_cycle[ 1022] = 1'b1;  addr_rom[ 1022]='h00000ff8;  wr_data_rom[ 1022]='h00001b4f;
    rd_cycle[ 1023] = 1'b0;  wr_cycle[ 1023] = 1'b1;  addr_rom[ 1023]='h00000ffc;  wr_data_rom[ 1023]='h000004a1;
    rd_cycle[ 1024] = 1'b0;  wr_cycle[ 1024] = 1'b1;  addr_rom[ 1024]='h00001000;  wr_data_rom[ 1024]='h00001c47;
    rd_cycle[ 1025] = 1'b0;  wr_cycle[ 1025] = 1'b1;  addr_rom[ 1025]='h00001004;  wr_data_rom[ 1025]='h00001007;
    rd_cycle[ 1026] = 1'b0;  wr_cycle[ 1026] = 1'b1;  addr_rom[ 1026]='h00001008;  wr_data_rom[ 1026]='h00000dc1;
    rd_cycle[ 1027] = 1'b0;  wr_cycle[ 1027] = 1'b1;  addr_rom[ 1027]='h0000100c;  wr_data_rom[ 1027]='h00001903;
    rd_cycle[ 1028] = 1'b0;  wr_cycle[ 1028] = 1'b1;  addr_rom[ 1028]='h00001010;  wr_data_rom[ 1028]='h0000106c;
    rd_cycle[ 1029] = 1'b0;  wr_cycle[ 1029] = 1'b1;  addr_rom[ 1029]='h00001014;  wr_data_rom[ 1029]='h00001d92;
    rd_cycle[ 1030] = 1'b0;  wr_cycle[ 1030] = 1'b1;  addr_rom[ 1030]='h00001018;  wr_data_rom[ 1030]='h00001577;
    rd_cycle[ 1031] = 1'b0;  wr_cycle[ 1031] = 1'b1;  addr_rom[ 1031]='h0000101c;  wr_data_rom[ 1031]='h00000e93;
    rd_cycle[ 1032] = 1'b0;  wr_cycle[ 1032] = 1'b1;  addr_rom[ 1032]='h00001020;  wr_data_rom[ 1032]='h000017cd;
    rd_cycle[ 1033] = 1'b0;  wr_cycle[ 1033] = 1'b1;  addr_rom[ 1033]='h00001024;  wr_data_rom[ 1033]='h00000579;
    rd_cycle[ 1034] = 1'b0;  wr_cycle[ 1034] = 1'b1;  addr_rom[ 1034]='h00001028;  wr_data_rom[ 1034]='h0000140b;
    rd_cycle[ 1035] = 1'b0;  wr_cycle[ 1035] = 1'b1;  addr_rom[ 1035]='h0000102c;  wr_data_rom[ 1035]='h00000020;
    rd_cycle[ 1036] = 1'b0;  wr_cycle[ 1036] = 1'b1;  addr_rom[ 1036]='h00001030;  wr_data_rom[ 1036]='h0000098c;
    rd_cycle[ 1037] = 1'b0;  wr_cycle[ 1037] = 1'b1;  addr_rom[ 1037]='h00001034;  wr_data_rom[ 1037]='h00000529;
    rd_cycle[ 1038] = 1'b0;  wr_cycle[ 1038] = 1'b1;  addr_rom[ 1038]='h00001038;  wr_data_rom[ 1038]='h00000879;
    rd_cycle[ 1039] = 1'b0;  wr_cycle[ 1039] = 1'b1;  addr_rom[ 1039]='h0000103c;  wr_data_rom[ 1039]='h00001999;
    rd_cycle[ 1040] = 1'b0;  wr_cycle[ 1040] = 1'b1;  addr_rom[ 1040]='h00001040;  wr_data_rom[ 1040]='h00001d09;
    rd_cycle[ 1041] = 1'b0;  wr_cycle[ 1041] = 1'b1;  addr_rom[ 1041]='h00001044;  wr_data_rom[ 1041]='h000017fc;
    rd_cycle[ 1042] = 1'b0;  wr_cycle[ 1042] = 1'b1;  addr_rom[ 1042]='h00001048;  wr_data_rom[ 1042]='h0000199f;
    rd_cycle[ 1043] = 1'b0;  wr_cycle[ 1043] = 1'b1;  addr_rom[ 1043]='h0000104c;  wr_data_rom[ 1043]='h00000658;
    rd_cycle[ 1044] = 1'b0;  wr_cycle[ 1044] = 1'b1;  addr_rom[ 1044]='h00001050;  wr_data_rom[ 1044]='h00001e67;
    rd_cycle[ 1045] = 1'b0;  wr_cycle[ 1045] = 1'b1;  addr_rom[ 1045]='h00001054;  wr_data_rom[ 1045]='h00000af6;
    rd_cycle[ 1046] = 1'b0;  wr_cycle[ 1046] = 1'b1;  addr_rom[ 1046]='h00001058;  wr_data_rom[ 1046]='h00000605;
    rd_cycle[ 1047] = 1'b0;  wr_cycle[ 1047] = 1'b1;  addr_rom[ 1047]='h0000105c;  wr_data_rom[ 1047]='h00001914;
    rd_cycle[ 1048] = 1'b0;  wr_cycle[ 1048] = 1'b1;  addr_rom[ 1048]='h00001060;  wr_data_rom[ 1048]='h00001e7e;
    rd_cycle[ 1049] = 1'b0;  wr_cycle[ 1049] = 1'b1;  addr_rom[ 1049]='h00001064;  wr_data_rom[ 1049]='h0000069d;
    rd_cycle[ 1050] = 1'b0;  wr_cycle[ 1050] = 1'b1;  addr_rom[ 1050]='h00001068;  wr_data_rom[ 1050]='h00001072;
    rd_cycle[ 1051] = 1'b0;  wr_cycle[ 1051] = 1'b1;  addr_rom[ 1051]='h0000106c;  wr_data_rom[ 1051]='h000005ed;
    rd_cycle[ 1052] = 1'b0;  wr_cycle[ 1052] = 1'b1;  addr_rom[ 1052]='h00001070;  wr_data_rom[ 1052]='h00000e1b;
    rd_cycle[ 1053] = 1'b0;  wr_cycle[ 1053] = 1'b1;  addr_rom[ 1053]='h00001074;  wr_data_rom[ 1053]='h00001276;
    rd_cycle[ 1054] = 1'b0;  wr_cycle[ 1054] = 1'b1;  addr_rom[ 1054]='h00001078;  wr_data_rom[ 1054]='h00000a16;
    rd_cycle[ 1055] = 1'b0;  wr_cycle[ 1055] = 1'b1;  addr_rom[ 1055]='h0000107c;  wr_data_rom[ 1055]='h000018f7;
    rd_cycle[ 1056] = 1'b0;  wr_cycle[ 1056] = 1'b1;  addr_rom[ 1056]='h00001080;  wr_data_rom[ 1056]='h00000508;
    rd_cycle[ 1057] = 1'b0;  wr_cycle[ 1057] = 1'b1;  addr_rom[ 1057]='h00001084;  wr_data_rom[ 1057]='h0000130c;
    rd_cycle[ 1058] = 1'b0;  wr_cycle[ 1058] = 1'b1;  addr_rom[ 1058]='h00001088;  wr_data_rom[ 1058]='h00001304;
    rd_cycle[ 1059] = 1'b0;  wr_cycle[ 1059] = 1'b1;  addr_rom[ 1059]='h0000108c;  wr_data_rom[ 1059]='h00000837;
    rd_cycle[ 1060] = 1'b0;  wr_cycle[ 1060] = 1'b1;  addr_rom[ 1060]='h00001090;  wr_data_rom[ 1060]='h00001909;
    rd_cycle[ 1061] = 1'b0;  wr_cycle[ 1061] = 1'b1;  addr_rom[ 1061]='h00001094;  wr_data_rom[ 1061]='h000011e9;
    rd_cycle[ 1062] = 1'b0;  wr_cycle[ 1062] = 1'b1;  addr_rom[ 1062]='h00001098;  wr_data_rom[ 1062]='h00000956;
    rd_cycle[ 1063] = 1'b0;  wr_cycle[ 1063] = 1'b1;  addr_rom[ 1063]='h0000109c;  wr_data_rom[ 1063]='h00001745;
    rd_cycle[ 1064] = 1'b0;  wr_cycle[ 1064] = 1'b1;  addr_rom[ 1064]='h000010a0;  wr_data_rom[ 1064]='h0000017a;
    rd_cycle[ 1065] = 1'b0;  wr_cycle[ 1065] = 1'b1;  addr_rom[ 1065]='h000010a4;  wr_data_rom[ 1065]='h00000bdf;
    rd_cycle[ 1066] = 1'b0;  wr_cycle[ 1066] = 1'b1;  addr_rom[ 1066]='h000010a8;  wr_data_rom[ 1066]='h000005ef;
    rd_cycle[ 1067] = 1'b0;  wr_cycle[ 1067] = 1'b1;  addr_rom[ 1067]='h000010ac;  wr_data_rom[ 1067]='h00000a4c;
    rd_cycle[ 1068] = 1'b0;  wr_cycle[ 1068] = 1'b1;  addr_rom[ 1068]='h000010b0;  wr_data_rom[ 1068]='h00001cc5;
    rd_cycle[ 1069] = 1'b0;  wr_cycle[ 1069] = 1'b1;  addr_rom[ 1069]='h000010b4;  wr_data_rom[ 1069]='h000003da;
    rd_cycle[ 1070] = 1'b0;  wr_cycle[ 1070] = 1'b1;  addr_rom[ 1070]='h000010b8;  wr_data_rom[ 1070]='h00001ea4;
    rd_cycle[ 1071] = 1'b0;  wr_cycle[ 1071] = 1'b1;  addr_rom[ 1071]='h000010bc;  wr_data_rom[ 1071]='h00000de3;
    rd_cycle[ 1072] = 1'b0;  wr_cycle[ 1072] = 1'b1;  addr_rom[ 1072]='h000010c0;  wr_data_rom[ 1072]='h00000b66;
    rd_cycle[ 1073] = 1'b0;  wr_cycle[ 1073] = 1'b1;  addr_rom[ 1073]='h000010c4;  wr_data_rom[ 1073]='h0000005e;
    rd_cycle[ 1074] = 1'b0;  wr_cycle[ 1074] = 1'b1;  addr_rom[ 1074]='h000010c8;  wr_data_rom[ 1074]='h00000bd6;
    rd_cycle[ 1075] = 1'b0;  wr_cycle[ 1075] = 1'b1;  addr_rom[ 1075]='h000010cc;  wr_data_rom[ 1075]='h000006ca;
    rd_cycle[ 1076] = 1'b0;  wr_cycle[ 1076] = 1'b1;  addr_rom[ 1076]='h000010d0;  wr_data_rom[ 1076]='h000000b0;
    rd_cycle[ 1077] = 1'b0;  wr_cycle[ 1077] = 1'b1;  addr_rom[ 1077]='h000010d4;  wr_data_rom[ 1077]='h00001ea9;
    rd_cycle[ 1078] = 1'b0;  wr_cycle[ 1078] = 1'b1;  addr_rom[ 1078]='h000010d8;  wr_data_rom[ 1078]='h00001b59;
    rd_cycle[ 1079] = 1'b0;  wr_cycle[ 1079] = 1'b1;  addr_rom[ 1079]='h000010dc;  wr_data_rom[ 1079]='h00001197;
    rd_cycle[ 1080] = 1'b0;  wr_cycle[ 1080] = 1'b1;  addr_rom[ 1080]='h000010e0;  wr_data_rom[ 1080]='h000012ec;
    rd_cycle[ 1081] = 1'b0;  wr_cycle[ 1081] = 1'b1;  addr_rom[ 1081]='h000010e4;  wr_data_rom[ 1081]='h000019b8;
    rd_cycle[ 1082] = 1'b0;  wr_cycle[ 1082] = 1'b1;  addr_rom[ 1082]='h000010e8;  wr_data_rom[ 1082]='h00000ec3;
    rd_cycle[ 1083] = 1'b0;  wr_cycle[ 1083] = 1'b1;  addr_rom[ 1083]='h000010ec;  wr_data_rom[ 1083]='h0000083d;
    rd_cycle[ 1084] = 1'b0;  wr_cycle[ 1084] = 1'b1;  addr_rom[ 1084]='h000010f0;  wr_data_rom[ 1084]='h00000d11;
    rd_cycle[ 1085] = 1'b0;  wr_cycle[ 1085] = 1'b1;  addr_rom[ 1085]='h000010f4;  wr_data_rom[ 1085]='h0000064d;
    rd_cycle[ 1086] = 1'b0;  wr_cycle[ 1086] = 1'b1;  addr_rom[ 1086]='h000010f8;  wr_data_rom[ 1086]='h000004b3;
    rd_cycle[ 1087] = 1'b0;  wr_cycle[ 1087] = 1'b1;  addr_rom[ 1087]='h000010fc;  wr_data_rom[ 1087]='h0000196a;
    rd_cycle[ 1088] = 1'b0;  wr_cycle[ 1088] = 1'b1;  addr_rom[ 1088]='h00001100;  wr_data_rom[ 1088]='h00000512;
    rd_cycle[ 1089] = 1'b0;  wr_cycle[ 1089] = 1'b1;  addr_rom[ 1089]='h00001104;  wr_data_rom[ 1089]='h00000077;
    rd_cycle[ 1090] = 1'b0;  wr_cycle[ 1090] = 1'b1;  addr_rom[ 1090]='h00001108;  wr_data_rom[ 1090]='h000002cc;
    rd_cycle[ 1091] = 1'b0;  wr_cycle[ 1091] = 1'b1;  addr_rom[ 1091]='h0000110c;  wr_data_rom[ 1091]='h00001da4;
    rd_cycle[ 1092] = 1'b0;  wr_cycle[ 1092] = 1'b1;  addr_rom[ 1092]='h00001110;  wr_data_rom[ 1092]='h00000440;
    rd_cycle[ 1093] = 1'b0;  wr_cycle[ 1093] = 1'b1;  addr_rom[ 1093]='h00001114;  wr_data_rom[ 1093]='h00000f18;
    rd_cycle[ 1094] = 1'b0;  wr_cycle[ 1094] = 1'b1;  addr_rom[ 1094]='h00001118;  wr_data_rom[ 1094]='h0000056f;
    rd_cycle[ 1095] = 1'b0;  wr_cycle[ 1095] = 1'b1;  addr_rom[ 1095]='h0000111c;  wr_data_rom[ 1095]='h00000bed;
    rd_cycle[ 1096] = 1'b0;  wr_cycle[ 1096] = 1'b1;  addr_rom[ 1096]='h00001120;  wr_data_rom[ 1096]='h00000f86;
    rd_cycle[ 1097] = 1'b0;  wr_cycle[ 1097] = 1'b1;  addr_rom[ 1097]='h00001124;  wr_data_rom[ 1097]='h000018b4;
    rd_cycle[ 1098] = 1'b0;  wr_cycle[ 1098] = 1'b1;  addr_rom[ 1098]='h00001128;  wr_data_rom[ 1098]='h00000434;
    rd_cycle[ 1099] = 1'b0;  wr_cycle[ 1099] = 1'b1;  addr_rom[ 1099]='h0000112c;  wr_data_rom[ 1099]='h00001b52;
    rd_cycle[ 1100] = 1'b0;  wr_cycle[ 1100] = 1'b1;  addr_rom[ 1100]='h00001130;  wr_data_rom[ 1100]='h000016f6;
    rd_cycle[ 1101] = 1'b0;  wr_cycle[ 1101] = 1'b1;  addr_rom[ 1101]='h00001134;  wr_data_rom[ 1101]='h000001ca;
    rd_cycle[ 1102] = 1'b0;  wr_cycle[ 1102] = 1'b1;  addr_rom[ 1102]='h00001138;  wr_data_rom[ 1102]='h00001f01;
    rd_cycle[ 1103] = 1'b0;  wr_cycle[ 1103] = 1'b1;  addr_rom[ 1103]='h0000113c;  wr_data_rom[ 1103]='h00001cf2;
    rd_cycle[ 1104] = 1'b0;  wr_cycle[ 1104] = 1'b1;  addr_rom[ 1104]='h00001140;  wr_data_rom[ 1104]='h00000a36;
    rd_cycle[ 1105] = 1'b0;  wr_cycle[ 1105] = 1'b1;  addr_rom[ 1105]='h00001144;  wr_data_rom[ 1105]='h000016b4;
    rd_cycle[ 1106] = 1'b0;  wr_cycle[ 1106] = 1'b1;  addr_rom[ 1106]='h00001148;  wr_data_rom[ 1106]='h00000b11;
    rd_cycle[ 1107] = 1'b0;  wr_cycle[ 1107] = 1'b1;  addr_rom[ 1107]='h0000114c;  wr_data_rom[ 1107]='h00001472;
    rd_cycle[ 1108] = 1'b0;  wr_cycle[ 1108] = 1'b1;  addr_rom[ 1108]='h00001150;  wr_data_rom[ 1108]='h000010ee;
    rd_cycle[ 1109] = 1'b0;  wr_cycle[ 1109] = 1'b1;  addr_rom[ 1109]='h00001154;  wr_data_rom[ 1109]='h0000141b;
    rd_cycle[ 1110] = 1'b0;  wr_cycle[ 1110] = 1'b1;  addr_rom[ 1110]='h00001158;  wr_data_rom[ 1110]='h0000156d;
    rd_cycle[ 1111] = 1'b0;  wr_cycle[ 1111] = 1'b1;  addr_rom[ 1111]='h0000115c;  wr_data_rom[ 1111]='h00000078;
    rd_cycle[ 1112] = 1'b0;  wr_cycle[ 1112] = 1'b1;  addr_rom[ 1112]='h00001160;  wr_data_rom[ 1112]='h00001b8b;
    rd_cycle[ 1113] = 1'b0;  wr_cycle[ 1113] = 1'b1;  addr_rom[ 1113]='h00001164;  wr_data_rom[ 1113]='h0000173e;
    rd_cycle[ 1114] = 1'b0;  wr_cycle[ 1114] = 1'b1;  addr_rom[ 1114]='h00001168;  wr_data_rom[ 1114]='h000013d3;
    rd_cycle[ 1115] = 1'b0;  wr_cycle[ 1115] = 1'b1;  addr_rom[ 1115]='h0000116c;  wr_data_rom[ 1115]='h00001b9b;
    rd_cycle[ 1116] = 1'b0;  wr_cycle[ 1116] = 1'b1;  addr_rom[ 1116]='h00001170;  wr_data_rom[ 1116]='h00000552;
    rd_cycle[ 1117] = 1'b0;  wr_cycle[ 1117] = 1'b1;  addr_rom[ 1117]='h00001174;  wr_data_rom[ 1117]='h000010f2;
    rd_cycle[ 1118] = 1'b0;  wr_cycle[ 1118] = 1'b1;  addr_rom[ 1118]='h00001178;  wr_data_rom[ 1118]='h0000118e;
    rd_cycle[ 1119] = 1'b0;  wr_cycle[ 1119] = 1'b1;  addr_rom[ 1119]='h0000117c;  wr_data_rom[ 1119]='h00000b38;
    rd_cycle[ 1120] = 1'b0;  wr_cycle[ 1120] = 1'b1;  addr_rom[ 1120]='h00001180;  wr_data_rom[ 1120]='h00000aa5;
    rd_cycle[ 1121] = 1'b0;  wr_cycle[ 1121] = 1'b1;  addr_rom[ 1121]='h00001184;  wr_data_rom[ 1121]='h00001a8d;
    rd_cycle[ 1122] = 1'b0;  wr_cycle[ 1122] = 1'b1;  addr_rom[ 1122]='h00001188;  wr_data_rom[ 1122]='h00000c79;
    rd_cycle[ 1123] = 1'b0;  wr_cycle[ 1123] = 1'b1;  addr_rom[ 1123]='h0000118c;  wr_data_rom[ 1123]='h00000136;
    rd_cycle[ 1124] = 1'b0;  wr_cycle[ 1124] = 1'b1;  addr_rom[ 1124]='h00001190;  wr_data_rom[ 1124]='h0000074c;
    rd_cycle[ 1125] = 1'b0;  wr_cycle[ 1125] = 1'b1;  addr_rom[ 1125]='h00001194;  wr_data_rom[ 1125]='h00000cf0;
    rd_cycle[ 1126] = 1'b0;  wr_cycle[ 1126] = 1'b1;  addr_rom[ 1126]='h00001198;  wr_data_rom[ 1126]='h0000023b;
    rd_cycle[ 1127] = 1'b0;  wr_cycle[ 1127] = 1'b1;  addr_rom[ 1127]='h0000119c;  wr_data_rom[ 1127]='h00000645;
    rd_cycle[ 1128] = 1'b0;  wr_cycle[ 1128] = 1'b1;  addr_rom[ 1128]='h000011a0;  wr_data_rom[ 1128]='h00001244;
    rd_cycle[ 1129] = 1'b0;  wr_cycle[ 1129] = 1'b1;  addr_rom[ 1129]='h000011a4;  wr_data_rom[ 1129]='h00001bf7;
    rd_cycle[ 1130] = 1'b0;  wr_cycle[ 1130] = 1'b1;  addr_rom[ 1130]='h000011a8;  wr_data_rom[ 1130]='h00000ece;
    rd_cycle[ 1131] = 1'b0;  wr_cycle[ 1131] = 1'b1;  addr_rom[ 1131]='h000011ac;  wr_data_rom[ 1131]='h00000eb8;
    rd_cycle[ 1132] = 1'b0;  wr_cycle[ 1132] = 1'b1;  addr_rom[ 1132]='h000011b0;  wr_data_rom[ 1132]='h0000081c;
    rd_cycle[ 1133] = 1'b0;  wr_cycle[ 1133] = 1'b1;  addr_rom[ 1133]='h000011b4;  wr_data_rom[ 1133]='h00001448;
    rd_cycle[ 1134] = 1'b0;  wr_cycle[ 1134] = 1'b1;  addr_rom[ 1134]='h000011b8;  wr_data_rom[ 1134]='h00000e9c;
    rd_cycle[ 1135] = 1'b0;  wr_cycle[ 1135] = 1'b1;  addr_rom[ 1135]='h000011bc;  wr_data_rom[ 1135]='h000009b5;
    rd_cycle[ 1136] = 1'b0;  wr_cycle[ 1136] = 1'b1;  addr_rom[ 1136]='h000011c0;  wr_data_rom[ 1136]='h00000501;
    rd_cycle[ 1137] = 1'b0;  wr_cycle[ 1137] = 1'b1;  addr_rom[ 1137]='h000011c4;  wr_data_rom[ 1137]='h00001099;
    rd_cycle[ 1138] = 1'b0;  wr_cycle[ 1138] = 1'b1;  addr_rom[ 1138]='h000011c8;  wr_data_rom[ 1138]='h000019c0;
    rd_cycle[ 1139] = 1'b0;  wr_cycle[ 1139] = 1'b1;  addr_rom[ 1139]='h000011cc;  wr_data_rom[ 1139]='h000019cb;
    rd_cycle[ 1140] = 1'b0;  wr_cycle[ 1140] = 1'b1;  addr_rom[ 1140]='h000011d0;  wr_data_rom[ 1140]='h00000ff1;
    rd_cycle[ 1141] = 1'b0;  wr_cycle[ 1141] = 1'b1;  addr_rom[ 1141]='h000011d4;  wr_data_rom[ 1141]='h00001375;
    rd_cycle[ 1142] = 1'b0;  wr_cycle[ 1142] = 1'b1;  addr_rom[ 1142]='h000011d8;  wr_data_rom[ 1142]='h00000893;
    rd_cycle[ 1143] = 1'b0;  wr_cycle[ 1143] = 1'b1;  addr_rom[ 1143]='h000011dc;  wr_data_rom[ 1143]='h00000ffd;
    rd_cycle[ 1144] = 1'b0;  wr_cycle[ 1144] = 1'b1;  addr_rom[ 1144]='h000011e0;  wr_data_rom[ 1144]='h00001d0b;
    rd_cycle[ 1145] = 1'b0;  wr_cycle[ 1145] = 1'b1;  addr_rom[ 1145]='h000011e4;  wr_data_rom[ 1145]='h00000303;
    rd_cycle[ 1146] = 1'b0;  wr_cycle[ 1146] = 1'b1;  addr_rom[ 1146]='h000011e8;  wr_data_rom[ 1146]='h00001645;
    rd_cycle[ 1147] = 1'b0;  wr_cycle[ 1147] = 1'b1;  addr_rom[ 1147]='h000011ec;  wr_data_rom[ 1147]='h000019ec;
    rd_cycle[ 1148] = 1'b0;  wr_cycle[ 1148] = 1'b1;  addr_rom[ 1148]='h000011f0;  wr_data_rom[ 1148]='h00000776;
    rd_cycle[ 1149] = 1'b0;  wr_cycle[ 1149] = 1'b1;  addr_rom[ 1149]='h000011f4;  wr_data_rom[ 1149]='h00001688;
    rd_cycle[ 1150] = 1'b0;  wr_cycle[ 1150] = 1'b1;  addr_rom[ 1150]='h000011f8;  wr_data_rom[ 1150]='h00000eae;
    rd_cycle[ 1151] = 1'b0;  wr_cycle[ 1151] = 1'b1;  addr_rom[ 1151]='h000011fc;  wr_data_rom[ 1151]='h000006ee;
    rd_cycle[ 1152] = 1'b0;  wr_cycle[ 1152] = 1'b1;  addr_rom[ 1152]='h00001200;  wr_data_rom[ 1152]='h0000063a;
    rd_cycle[ 1153] = 1'b0;  wr_cycle[ 1153] = 1'b1;  addr_rom[ 1153]='h00001204;  wr_data_rom[ 1153]='h00000bc0;
    rd_cycle[ 1154] = 1'b0;  wr_cycle[ 1154] = 1'b1;  addr_rom[ 1154]='h00001208;  wr_data_rom[ 1154]='h00001033;
    rd_cycle[ 1155] = 1'b0;  wr_cycle[ 1155] = 1'b1;  addr_rom[ 1155]='h0000120c;  wr_data_rom[ 1155]='h00001c5d;
    rd_cycle[ 1156] = 1'b0;  wr_cycle[ 1156] = 1'b1;  addr_rom[ 1156]='h00001210;  wr_data_rom[ 1156]='h000011a2;
    rd_cycle[ 1157] = 1'b0;  wr_cycle[ 1157] = 1'b1;  addr_rom[ 1157]='h00001214;  wr_data_rom[ 1157]='h0000048b;
    rd_cycle[ 1158] = 1'b0;  wr_cycle[ 1158] = 1'b1;  addr_rom[ 1158]='h00001218;  wr_data_rom[ 1158]='h00001b31;
    rd_cycle[ 1159] = 1'b0;  wr_cycle[ 1159] = 1'b1;  addr_rom[ 1159]='h0000121c;  wr_data_rom[ 1159]='h0000058a;
    rd_cycle[ 1160] = 1'b0;  wr_cycle[ 1160] = 1'b1;  addr_rom[ 1160]='h00001220;  wr_data_rom[ 1160]='h00001e72;
    rd_cycle[ 1161] = 1'b0;  wr_cycle[ 1161] = 1'b1;  addr_rom[ 1161]='h00001224;  wr_data_rom[ 1161]='h000007c1;
    rd_cycle[ 1162] = 1'b0;  wr_cycle[ 1162] = 1'b1;  addr_rom[ 1162]='h00001228;  wr_data_rom[ 1162]='h00001d9f;
    rd_cycle[ 1163] = 1'b0;  wr_cycle[ 1163] = 1'b1;  addr_rom[ 1163]='h0000122c;  wr_data_rom[ 1163]='h0000188f;
    rd_cycle[ 1164] = 1'b0;  wr_cycle[ 1164] = 1'b1;  addr_rom[ 1164]='h00001230;  wr_data_rom[ 1164]='h00001712;
    rd_cycle[ 1165] = 1'b0;  wr_cycle[ 1165] = 1'b1;  addr_rom[ 1165]='h00001234;  wr_data_rom[ 1165]='h00001b92;
    rd_cycle[ 1166] = 1'b0;  wr_cycle[ 1166] = 1'b1;  addr_rom[ 1166]='h00001238;  wr_data_rom[ 1166]='h00000e08;
    rd_cycle[ 1167] = 1'b0;  wr_cycle[ 1167] = 1'b1;  addr_rom[ 1167]='h0000123c;  wr_data_rom[ 1167]='h00000931;
    rd_cycle[ 1168] = 1'b0;  wr_cycle[ 1168] = 1'b1;  addr_rom[ 1168]='h00001240;  wr_data_rom[ 1168]='h0000171b;
    rd_cycle[ 1169] = 1'b0;  wr_cycle[ 1169] = 1'b1;  addr_rom[ 1169]='h00001244;  wr_data_rom[ 1169]='h00000c72;
    rd_cycle[ 1170] = 1'b0;  wr_cycle[ 1170] = 1'b1;  addr_rom[ 1170]='h00001248;  wr_data_rom[ 1170]='h0000156a;
    rd_cycle[ 1171] = 1'b0;  wr_cycle[ 1171] = 1'b1;  addr_rom[ 1171]='h0000124c;  wr_data_rom[ 1171]='h000005af;
    rd_cycle[ 1172] = 1'b0;  wr_cycle[ 1172] = 1'b1;  addr_rom[ 1172]='h00001250;  wr_data_rom[ 1172]='h00001004;
    rd_cycle[ 1173] = 1'b0;  wr_cycle[ 1173] = 1'b1;  addr_rom[ 1173]='h00001254;  wr_data_rom[ 1173]='h0000166f;
    rd_cycle[ 1174] = 1'b0;  wr_cycle[ 1174] = 1'b1;  addr_rom[ 1174]='h00001258;  wr_data_rom[ 1174]='h00001f25;
    rd_cycle[ 1175] = 1'b0;  wr_cycle[ 1175] = 1'b1;  addr_rom[ 1175]='h0000125c;  wr_data_rom[ 1175]='h000010e3;
    rd_cycle[ 1176] = 1'b0;  wr_cycle[ 1176] = 1'b1;  addr_rom[ 1176]='h00001260;  wr_data_rom[ 1176]='h00001376;
    rd_cycle[ 1177] = 1'b0;  wr_cycle[ 1177] = 1'b1;  addr_rom[ 1177]='h00001264;  wr_data_rom[ 1177]='h00000171;
    rd_cycle[ 1178] = 1'b0;  wr_cycle[ 1178] = 1'b1;  addr_rom[ 1178]='h00001268;  wr_data_rom[ 1178]='h00000640;
    rd_cycle[ 1179] = 1'b0;  wr_cycle[ 1179] = 1'b1;  addr_rom[ 1179]='h0000126c;  wr_data_rom[ 1179]='h0000016b;
    rd_cycle[ 1180] = 1'b0;  wr_cycle[ 1180] = 1'b1;  addr_rom[ 1180]='h00001270;  wr_data_rom[ 1180]='h00000b02;
    rd_cycle[ 1181] = 1'b0;  wr_cycle[ 1181] = 1'b1;  addr_rom[ 1181]='h00001274;  wr_data_rom[ 1181]='h00000eef;
    rd_cycle[ 1182] = 1'b0;  wr_cycle[ 1182] = 1'b1;  addr_rom[ 1182]='h00001278;  wr_data_rom[ 1182]='h00001cbb;
    rd_cycle[ 1183] = 1'b0;  wr_cycle[ 1183] = 1'b1;  addr_rom[ 1183]='h0000127c;  wr_data_rom[ 1183]='h000019ca;
    rd_cycle[ 1184] = 1'b0;  wr_cycle[ 1184] = 1'b1;  addr_rom[ 1184]='h00001280;  wr_data_rom[ 1184]='h00000629;
    rd_cycle[ 1185] = 1'b0;  wr_cycle[ 1185] = 1'b1;  addr_rom[ 1185]='h00001284;  wr_data_rom[ 1185]='h00001347;
    rd_cycle[ 1186] = 1'b0;  wr_cycle[ 1186] = 1'b1;  addr_rom[ 1186]='h00001288;  wr_data_rom[ 1186]='h00001797;
    rd_cycle[ 1187] = 1'b0;  wr_cycle[ 1187] = 1'b1;  addr_rom[ 1187]='h0000128c;  wr_data_rom[ 1187]='h00000f7b;
    rd_cycle[ 1188] = 1'b0;  wr_cycle[ 1188] = 1'b1;  addr_rom[ 1188]='h00001290;  wr_data_rom[ 1188]='h0000052f;
    rd_cycle[ 1189] = 1'b0;  wr_cycle[ 1189] = 1'b1;  addr_rom[ 1189]='h00001294;  wr_data_rom[ 1189]='h00000c86;
    rd_cycle[ 1190] = 1'b0;  wr_cycle[ 1190] = 1'b1;  addr_rom[ 1190]='h00001298;  wr_data_rom[ 1190]='h00000113;
    rd_cycle[ 1191] = 1'b0;  wr_cycle[ 1191] = 1'b1;  addr_rom[ 1191]='h0000129c;  wr_data_rom[ 1191]='h00000299;
    rd_cycle[ 1192] = 1'b0;  wr_cycle[ 1192] = 1'b1;  addr_rom[ 1192]='h000012a0;  wr_data_rom[ 1192]='h00000766;
    rd_cycle[ 1193] = 1'b0;  wr_cycle[ 1193] = 1'b1;  addr_rom[ 1193]='h000012a4;  wr_data_rom[ 1193]='h00000b13;
    rd_cycle[ 1194] = 1'b0;  wr_cycle[ 1194] = 1'b1;  addr_rom[ 1194]='h000012a8;  wr_data_rom[ 1194]='h0000101a;
    rd_cycle[ 1195] = 1'b0;  wr_cycle[ 1195] = 1'b1;  addr_rom[ 1195]='h000012ac;  wr_data_rom[ 1195]='h000013c5;
    rd_cycle[ 1196] = 1'b0;  wr_cycle[ 1196] = 1'b1;  addr_rom[ 1196]='h000012b0;  wr_data_rom[ 1196]='h000016de;
    rd_cycle[ 1197] = 1'b0;  wr_cycle[ 1197] = 1'b1;  addr_rom[ 1197]='h000012b4;  wr_data_rom[ 1197]='h0000058c;
    rd_cycle[ 1198] = 1'b0;  wr_cycle[ 1198] = 1'b1;  addr_rom[ 1198]='h000012b8;  wr_data_rom[ 1198]='h0000158d;
    rd_cycle[ 1199] = 1'b0;  wr_cycle[ 1199] = 1'b1;  addr_rom[ 1199]='h000012bc;  wr_data_rom[ 1199]='h0000064f;
    rd_cycle[ 1200] = 1'b0;  wr_cycle[ 1200] = 1'b1;  addr_rom[ 1200]='h000012c0;  wr_data_rom[ 1200]='h00001523;
    rd_cycle[ 1201] = 1'b0;  wr_cycle[ 1201] = 1'b1;  addr_rom[ 1201]='h000012c4;  wr_data_rom[ 1201]='h000018e4;
    rd_cycle[ 1202] = 1'b0;  wr_cycle[ 1202] = 1'b1;  addr_rom[ 1202]='h000012c8;  wr_data_rom[ 1202]='h00001689;
    rd_cycle[ 1203] = 1'b0;  wr_cycle[ 1203] = 1'b1;  addr_rom[ 1203]='h000012cc;  wr_data_rom[ 1203]='h00000fec;
    rd_cycle[ 1204] = 1'b0;  wr_cycle[ 1204] = 1'b1;  addr_rom[ 1204]='h000012d0;  wr_data_rom[ 1204]='h000005c1;
    rd_cycle[ 1205] = 1'b0;  wr_cycle[ 1205] = 1'b1;  addr_rom[ 1205]='h000012d4;  wr_data_rom[ 1205]='h0000059e;
    rd_cycle[ 1206] = 1'b0;  wr_cycle[ 1206] = 1'b1;  addr_rom[ 1206]='h000012d8;  wr_data_rom[ 1206]='h00000ba9;
    rd_cycle[ 1207] = 1'b0;  wr_cycle[ 1207] = 1'b1;  addr_rom[ 1207]='h000012dc;  wr_data_rom[ 1207]='h0000060a;
    rd_cycle[ 1208] = 1'b0;  wr_cycle[ 1208] = 1'b1;  addr_rom[ 1208]='h000012e0;  wr_data_rom[ 1208]='h000017ae;
    rd_cycle[ 1209] = 1'b0;  wr_cycle[ 1209] = 1'b1;  addr_rom[ 1209]='h000012e4;  wr_data_rom[ 1209]='h0000132b;
    rd_cycle[ 1210] = 1'b0;  wr_cycle[ 1210] = 1'b1;  addr_rom[ 1210]='h000012e8;  wr_data_rom[ 1210]='h00000e73;
    rd_cycle[ 1211] = 1'b0;  wr_cycle[ 1211] = 1'b1;  addr_rom[ 1211]='h000012ec;  wr_data_rom[ 1211]='h000009d0;
    rd_cycle[ 1212] = 1'b0;  wr_cycle[ 1212] = 1'b1;  addr_rom[ 1212]='h000012f0;  wr_data_rom[ 1212]='h00000683;
    rd_cycle[ 1213] = 1'b0;  wr_cycle[ 1213] = 1'b1;  addr_rom[ 1213]='h000012f4;  wr_data_rom[ 1213]='h00000bc7;
    rd_cycle[ 1214] = 1'b0;  wr_cycle[ 1214] = 1'b1;  addr_rom[ 1214]='h000012f8;  wr_data_rom[ 1214]='h00001768;
    rd_cycle[ 1215] = 1'b0;  wr_cycle[ 1215] = 1'b1;  addr_rom[ 1215]='h000012fc;  wr_data_rom[ 1215]='h000013f0;
    rd_cycle[ 1216] = 1'b0;  wr_cycle[ 1216] = 1'b1;  addr_rom[ 1216]='h00001300;  wr_data_rom[ 1216]='h00001491;
    rd_cycle[ 1217] = 1'b0;  wr_cycle[ 1217] = 1'b1;  addr_rom[ 1217]='h00001304;  wr_data_rom[ 1217]='h00000722;
    rd_cycle[ 1218] = 1'b0;  wr_cycle[ 1218] = 1'b1;  addr_rom[ 1218]='h00001308;  wr_data_rom[ 1218]='h00001b70;
    rd_cycle[ 1219] = 1'b0;  wr_cycle[ 1219] = 1'b1;  addr_rom[ 1219]='h0000130c;  wr_data_rom[ 1219]='h00001232;
    rd_cycle[ 1220] = 1'b0;  wr_cycle[ 1220] = 1'b1;  addr_rom[ 1220]='h00001310;  wr_data_rom[ 1220]='h0000072e;
    rd_cycle[ 1221] = 1'b0;  wr_cycle[ 1221] = 1'b1;  addr_rom[ 1221]='h00001314;  wr_data_rom[ 1221]='h00000539;
    rd_cycle[ 1222] = 1'b0;  wr_cycle[ 1222] = 1'b1;  addr_rom[ 1222]='h00001318;  wr_data_rom[ 1222]='h00001b26;
    rd_cycle[ 1223] = 1'b0;  wr_cycle[ 1223] = 1'b1;  addr_rom[ 1223]='h0000131c;  wr_data_rom[ 1223]='h00001c4c;
    rd_cycle[ 1224] = 1'b0;  wr_cycle[ 1224] = 1'b1;  addr_rom[ 1224]='h00001320;  wr_data_rom[ 1224]='h00001e0c;
    rd_cycle[ 1225] = 1'b0;  wr_cycle[ 1225] = 1'b1;  addr_rom[ 1225]='h00001324;  wr_data_rom[ 1225]='h0000085f;
    rd_cycle[ 1226] = 1'b0;  wr_cycle[ 1226] = 1'b1;  addr_rom[ 1226]='h00001328;  wr_data_rom[ 1226]='h00001265;
    rd_cycle[ 1227] = 1'b0;  wr_cycle[ 1227] = 1'b1;  addr_rom[ 1227]='h0000132c;  wr_data_rom[ 1227]='h00000cc5;
    rd_cycle[ 1228] = 1'b0;  wr_cycle[ 1228] = 1'b1;  addr_rom[ 1228]='h00001330;  wr_data_rom[ 1228]='h00000e61;
    rd_cycle[ 1229] = 1'b0;  wr_cycle[ 1229] = 1'b1;  addr_rom[ 1229]='h00001334;  wr_data_rom[ 1229]='h000014a1;
    rd_cycle[ 1230] = 1'b0;  wr_cycle[ 1230] = 1'b1;  addr_rom[ 1230]='h00001338;  wr_data_rom[ 1230]='h00001c32;
    rd_cycle[ 1231] = 1'b0;  wr_cycle[ 1231] = 1'b1;  addr_rom[ 1231]='h0000133c;  wr_data_rom[ 1231]='h0000002f;
    rd_cycle[ 1232] = 1'b0;  wr_cycle[ 1232] = 1'b1;  addr_rom[ 1232]='h00001340;  wr_data_rom[ 1232]='h000006d8;
    rd_cycle[ 1233] = 1'b0;  wr_cycle[ 1233] = 1'b1;  addr_rom[ 1233]='h00001344;  wr_data_rom[ 1233]='h0000014b;
    rd_cycle[ 1234] = 1'b0;  wr_cycle[ 1234] = 1'b1;  addr_rom[ 1234]='h00001348;  wr_data_rom[ 1234]='h00000bec;
    rd_cycle[ 1235] = 1'b0;  wr_cycle[ 1235] = 1'b1;  addr_rom[ 1235]='h0000134c;  wr_data_rom[ 1235]='h000005a0;
    rd_cycle[ 1236] = 1'b0;  wr_cycle[ 1236] = 1'b1;  addr_rom[ 1236]='h00001350;  wr_data_rom[ 1236]='h0000057a;
    rd_cycle[ 1237] = 1'b0;  wr_cycle[ 1237] = 1'b1;  addr_rom[ 1237]='h00001354;  wr_data_rom[ 1237]='h0000115b;
    rd_cycle[ 1238] = 1'b0;  wr_cycle[ 1238] = 1'b1;  addr_rom[ 1238]='h00001358;  wr_data_rom[ 1238]='h00000108;
    rd_cycle[ 1239] = 1'b0;  wr_cycle[ 1239] = 1'b1;  addr_rom[ 1239]='h0000135c;  wr_data_rom[ 1239]='h000013e0;
    rd_cycle[ 1240] = 1'b0;  wr_cycle[ 1240] = 1'b1;  addr_rom[ 1240]='h00001360;  wr_data_rom[ 1240]='h00001200;
    rd_cycle[ 1241] = 1'b0;  wr_cycle[ 1241] = 1'b1;  addr_rom[ 1241]='h00001364;  wr_data_rom[ 1241]='h00001960;
    rd_cycle[ 1242] = 1'b0;  wr_cycle[ 1242] = 1'b1;  addr_rom[ 1242]='h00001368;  wr_data_rom[ 1242]='h000011e5;
    rd_cycle[ 1243] = 1'b0;  wr_cycle[ 1243] = 1'b1;  addr_rom[ 1243]='h0000136c;  wr_data_rom[ 1243]='h0000020e;
    rd_cycle[ 1244] = 1'b0;  wr_cycle[ 1244] = 1'b1;  addr_rom[ 1244]='h00001370;  wr_data_rom[ 1244]='h00001e4d;
    rd_cycle[ 1245] = 1'b0;  wr_cycle[ 1245] = 1'b1;  addr_rom[ 1245]='h00001374;  wr_data_rom[ 1245]='h00001c15;
    rd_cycle[ 1246] = 1'b0;  wr_cycle[ 1246] = 1'b1;  addr_rom[ 1246]='h00001378;  wr_data_rom[ 1246]='h00001887;
    rd_cycle[ 1247] = 1'b0;  wr_cycle[ 1247] = 1'b1;  addr_rom[ 1247]='h0000137c;  wr_data_rom[ 1247]='h000007ef;
    rd_cycle[ 1248] = 1'b0;  wr_cycle[ 1248] = 1'b1;  addr_rom[ 1248]='h00001380;  wr_data_rom[ 1248]='h0000044e;
    rd_cycle[ 1249] = 1'b0;  wr_cycle[ 1249] = 1'b1;  addr_rom[ 1249]='h00001384;  wr_data_rom[ 1249]='h000000fa;
    rd_cycle[ 1250] = 1'b0;  wr_cycle[ 1250] = 1'b1;  addr_rom[ 1250]='h00001388;  wr_data_rom[ 1250]='h00000c8d;
    rd_cycle[ 1251] = 1'b0;  wr_cycle[ 1251] = 1'b1;  addr_rom[ 1251]='h0000138c;  wr_data_rom[ 1251]='h00001db9;
    rd_cycle[ 1252] = 1'b0;  wr_cycle[ 1252] = 1'b1;  addr_rom[ 1252]='h00001390;  wr_data_rom[ 1252]='h0000144e;
    rd_cycle[ 1253] = 1'b0;  wr_cycle[ 1253] = 1'b1;  addr_rom[ 1253]='h00001394;  wr_data_rom[ 1253]='h000003de;
    rd_cycle[ 1254] = 1'b0;  wr_cycle[ 1254] = 1'b1;  addr_rom[ 1254]='h00001398;  wr_data_rom[ 1254]='h00000e35;
    rd_cycle[ 1255] = 1'b0;  wr_cycle[ 1255] = 1'b1;  addr_rom[ 1255]='h0000139c;  wr_data_rom[ 1255]='h0000010e;
    rd_cycle[ 1256] = 1'b0;  wr_cycle[ 1256] = 1'b1;  addr_rom[ 1256]='h000013a0;  wr_data_rom[ 1256]='h00001edc;
    rd_cycle[ 1257] = 1'b0;  wr_cycle[ 1257] = 1'b1;  addr_rom[ 1257]='h000013a4;  wr_data_rom[ 1257]='h00001ca8;
    rd_cycle[ 1258] = 1'b0;  wr_cycle[ 1258] = 1'b1;  addr_rom[ 1258]='h000013a8;  wr_data_rom[ 1258]='h000000f7;
    rd_cycle[ 1259] = 1'b0;  wr_cycle[ 1259] = 1'b1;  addr_rom[ 1259]='h000013ac;  wr_data_rom[ 1259]='h0000028b;
    rd_cycle[ 1260] = 1'b0;  wr_cycle[ 1260] = 1'b1;  addr_rom[ 1260]='h000013b0;  wr_data_rom[ 1260]='h000014d0;
    rd_cycle[ 1261] = 1'b0;  wr_cycle[ 1261] = 1'b1;  addr_rom[ 1261]='h000013b4;  wr_data_rom[ 1261]='h0000070d;
    rd_cycle[ 1262] = 1'b0;  wr_cycle[ 1262] = 1'b1;  addr_rom[ 1262]='h000013b8;  wr_data_rom[ 1262]='h00001666;
    rd_cycle[ 1263] = 1'b0;  wr_cycle[ 1263] = 1'b1;  addr_rom[ 1263]='h000013bc;  wr_data_rom[ 1263]='h00000bb2;
    rd_cycle[ 1264] = 1'b0;  wr_cycle[ 1264] = 1'b1;  addr_rom[ 1264]='h000013c0;  wr_data_rom[ 1264]='h00000208;
    rd_cycle[ 1265] = 1'b0;  wr_cycle[ 1265] = 1'b1;  addr_rom[ 1265]='h000013c4;  wr_data_rom[ 1265]='h00000320;
    rd_cycle[ 1266] = 1'b0;  wr_cycle[ 1266] = 1'b1;  addr_rom[ 1266]='h000013c8;  wr_data_rom[ 1266]='h00000424;
    rd_cycle[ 1267] = 1'b0;  wr_cycle[ 1267] = 1'b1;  addr_rom[ 1267]='h000013cc;  wr_data_rom[ 1267]='h00000fa8;
    rd_cycle[ 1268] = 1'b0;  wr_cycle[ 1268] = 1'b1;  addr_rom[ 1268]='h000013d0;  wr_data_rom[ 1268]='h00001575;
    rd_cycle[ 1269] = 1'b0;  wr_cycle[ 1269] = 1'b1;  addr_rom[ 1269]='h000013d4;  wr_data_rom[ 1269]='h00001349;
    rd_cycle[ 1270] = 1'b0;  wr_cycle[ 1270] = 1'b1;  addr_rom[ 1270]='h000013d8;  wr_data_rom[ 1270]='h00000921;
    rd_cycle[ 1271] = 1'b0;  wr_cycle[ 1271] = 1'b1;  addr_rom[ 1271]='h000013dc;  wr_data_rom[ 1271]='h00000598;
    rd_cycle[ 1272] = 1'b0;  wr_cycle[ 1272] = 1'b1;  addr_rom[ 1272]='h000013e0;  wr_data_rom[ 1272]='h00000d6c;
    rd_cycle[ 1273] = 1'b0;  wr_cycle[ 1273] = 1'b1;  addr_rom[ 1273]='h000013e4;  wr_data_rom[ 1273]='h00000a15;
    rd_cycle[ 1274] = 1'b0;  wr_cycle[ 1274] = 1'b1;  addr_rom[ 1274]='h000013e8;  wr_data_rom[ 1274]='h00000a59;
    rd_cycle[ 1275] = 1'b0;  wr_cycle[ 1275] = 1'b1;  addr_rom[ 1275]='h000013ec;  wr_data_rom[ 1275]='h000002bf;
    rd_cycle[ 1276] = 1'b0;  wr_cycle[ 1276] = 1'b1;  addr_rom[ 1276]='h000013f0;  wr_data_rom[ 1276]='h00000400;
    rd_cycle[ 1277] = 1'b0;  wr_cycle[ 1277] = 1'b1;  addr_rom[ 1277]='h000013f4;  wr_data_rom[ 1277]='h000013e2;
    rd_cycle[ 1278] = 1'b0;  wr_cycle[ 1278] = 1'b1;  addr_rom[ 1278]='h000013f8;  wr_data_rom[ 1278]='h000018fd;
    rd_cycle[ 1279] = 1'b0;  wr_cycle[ 1279] = 1'b1;  addr_rom[ 1279]='h000013fc;  wr_data_rom[ 1279]='h00001a17;
    rd_cycle[ 1280] = 1'b0;  wr_cycle[ 1280] = 1'b1;  addr_rom[ 1280]='h00001400;  wr_data_rom[ 1280]='h000001dc;
    rd_cycle[ 1281] = 1'b0;  wr_cycle[ 1281] = 1'b1;  addr_rom[ 1281]='h00001404;  wr_data_rom[ 1281]='h0000001f;
    rd_cycle[ 1282] = 1'b0;  wr_cycle[ 1282] = 1'b1;  addr_rom[ 1282]='h00001408;  wr_data_rom[ 1282]='h00001bba;
    rd_cycle[ 1283] = 1'b0;  wr_cycle[ 1283] = 1'b1;  addr_rom[ 1283]='h0000140c;  wr_data_rom[ 1283]='h00001020;
    rd_cycle[ 1284] = 1'b0;  wr_cycle[ 1284] = 1'b1;  addr_rom[ 1284]='h00001410;  wr_data_rom[ 1284]='h0000130d;
    rd_cycle[ 1285] = 1'b0;  wr_cycle[ 1285] = 1'b1;  addr_rom[ 1285]='h00001414;  wr_data_rom[ 1285]='h00000b1e;
    rd_cycle[ 1286] = 1'b0;  wr_cycle[ 1286] = 1'b1;  addr_rom[ 1286]='h00001418;  wr_data_rom[ 1286]='h000004bc;
    rd_cycle[ 1287] = 1'b0;  wr_cycle[ 1287] = 1'b1;  addr_rom[ 1287]='h0000141c;  wr_data_rom[ 1287]='h00000f98;
    rd_cycle[ 1288] = 1'b0;  wr_cycle[ 1288] = 1'b1;  addr_rom[ 1288]='h00001420;  wr_data_rom[ 1288]='h00000e6c;
    rd_cycle[ 1289] = 1'b0;  wr_cycle[ 1289] = 1'b1;  addr_rom[ 1289]='h00001424;  wr_data_rom[ 1289]='h00000a5d;
    rd_cycle[ 1290] = 1'b0;  wr_cycle[ 1290] = 1'b1;  addr_rom[ 1290]='h00001428;  wr_data_rom[ 1290]='h00001a99;
    rd_cycle[ 1291] = 1'b0;  wr_cycle[ 1291] = 1'b1;  addr_rom[ 1291]='h0000142c;  wr_data_rom[ 1291]='h000017f9;
    rd_cycle[ 1292] = 1'b0;  wr_cycle[ 1292] = 1'b1;  addr_rom[ 1292]='h00001430;  wr_data_rom[ 1292]='h00000b68;
    rd_cycle[ 1293] = 1'b0;  wr_cycle[ 1293] = 1'b1;  addr_rom[ 1293]='h00001434;  wr_data_rom[ 1293]='h00000767;
    rd_cycle[ 1294] = 1'b0;  wr_cycle[ 1294] = 1'b1;  addr_rom[ 1294]='h00001438;  wr_data_rom[ 1294]='h00001784;
    rd_cycle[ 1295] = 1'b0;  wr_cycle[ 1295] = 1'b1;  addr_rom[ 1295]='h0000143c;  wr_data_rom[ 1295]='h00001c79;
    rd_cycle[ 1296] = 1'b0;  wr_cycle[ 1296] = 1'b1;  addr_rom[ 1296]='h00001440;  wr_data_rom[ 1296]='h00001a4d;
    rd_cycle[ 1297] = 1'b0;  wr_cycle[ 1297] = 1'b1;  addr_rom[ 1297]='h00001444;  wr_data_rom[ 1297]='h00000e6b;
    rd_cycle[ 1298] = 1'b0;  wr_cycle[ 1298] = 1'b1;  addr_rom[ 1298]='h00001448;  wr_data_rom[ 1298]='h00000587;
    rd_cycle[ 1299] = 1'b0;  wr_cycle[ 1299] = 1'b1;  addr_rom[ 1299]='h0000144c;  wr_data_rom[ 1299]='h00000667;
    rd_cycle[ 1300] = 1'b0;  wr_cycle[ 1300] = 1'b1;  addr_rom[ 1300]='h00001450;  wr_data_rom[ 1300]='h000019f6;
    rd_cycle[ 1301] = 1'b0;  wr_cycle[ 1301] = 1'b1;  addr_rom[ 1301]='h00001454;  wr_data_rom[ 1301]='h000015a5;
    rd_cycle[ 1302] = 1'b0;  wr_cycle[ 1302] = 1'b1;  addr_rom[ 1302]='h00001458;  wr_data_rom[ 1302]='h000013e7;
    rd_cycle[ 1303] = 1'b0;  wr_cycle[ 1303] = 1'b1;  addr_rom[ 1303]='h0000145c;  wr_data_rom[ 1303]='h00001d69;
    rd_cycle[ 1304] = 1'b0;  wr_cycle[ 1304] = 1'b1;  addr_rom[ 1304]='h00001460;  wr_data_rom[ 1304]='h000005f5;
    rd_cycle[ 1305] = 1'b0;  wr_cycle[ 1305] = 1'b1;  addr_rom[ 1305]='h00001464;  wr_data_rom[ 1305]='h000009b1;
    rd_cycle[ 1306] = 1'b0;  wr_cycle[ 1306] = 1'b1;  addr_rom[ 1306]='h00001468;  wr_data_rom[ 1306]='h00001884;
    rd_cycle[ 1307] = 1'b0;  wr_cycle[ 1307] = 1'b1;  addr_rom[ 1307]='h0000146c;  wr_data_rom[ 1307]='h00000b55;
    rd_cycle[ 1308] = 1'b0;  wr_cycle[ 1308] = 1'b1;  addr_rom[ 1308]='h00001470;  wr_data_rom[ 1308]='h00001dd5;
    rd_cycle[ 1309] = 1'b0;  wr_cycle[ 1309] = 1'b1;  addr_rom[ 1309]='h00001474;  wr_data_rom[ 1309]='h00001efc;
    rd_cycle[ 1310] = 1'b0;  wr_cycle[ 1310] = 1'b1;  addr_rom[ 1310]='h00001478;  wr_data_rom[ 1310]='h00001d60;
    rd_cycle[ 1311] = 1'b0;  wr_cycle[ 1311] = 1'b1;  addr_rom[ 1311]='h0000147c;  wr_data_rom[ 1311]='h0000032f;
    rd_cycle[ 1312] = 1'b0;  wr_cycle[ 1312] = 1'b1;  addr_rom[ 1312]='h00001480;  wr_data_rom[ 1312]='h00000cb5;
    rd_cycle[ 1313] = 1'b0;  wr_cycle[ 1313] = 1'b1;  addr_rom[ 1313]='h00001484;  wr_data_rom[ 1313]='h0000109a;
    rd_cycle[ 1314] = 1'b0;  wr_cycle[ 1314] = 1'b1;  addr_rom[ 1314]='h00001488;  wr_data_rom[ 1314]='h0000123b;
    rd_cycle[ 1315] = 1'b0;  wr_cycle[ 1315] = 1'b1;  addr_rom[ 1315]='h0000148c;  wr_data_rom[ 1315]='h00001db0;
    rd_cycle[ 1316] = 1'b0;  wr_cycle[ 1316] = 1'b1;  addr_rom[ 1316]='h00001490;  wr_data_rom[ 1316]='h000013a2;
    rd_cycle[ 1317] = 1'b0;  wr_cycle[ 1317] = 1'b1;  addr_rom[ 1317]='h00001494;  wr_data_rom[ 1317]='h00000c19;
    rd_cycle[ 1318] = 1'b0;  wr_cycle[ 1318] = 1'b1;  addr_rom[ 1318]='h00001498;  wr_data_rom[ 1318]='h000009b5;
    rd_cycle[ 1319] = 1'b0;  wr_cycle[ 1319] = 1'b1;  addr_rom[ 1319]='h0000149c;  wr_data_rom[ 1319]='h00001a9f;
    rd_cycle[ 1320] = 1'b0;  wr_cycle[ 1320] = 1'b1;  addr_rom[ 1320]='h000014a0;  wr_data_rom[ 1320]='h000010cc;
    rd_cycle[ 1321] = 1'b0;  wr_cycle[ 1321] = 1'b1;  addr_rom[ 1321]='h000014a4;  wr_data_rom[ 1321]='h00000e2b;
    rd_cycle[ 1322] = 1'b0;  wr_cycle[ 1322] = 1'b1;  addr_rom[ 1322]='h000014a8;  wr_data_rom[ 1322]='h0000127c;
    rd_cycle[ 1323] = 1'b0;  wr_cycle[ 1323] = 1'b1;  addr_rom[ 1323]='h000014ac;  wr_data_rom[ 1323]='h000016ef;
    rd_cycle[ 1324] = 1'b0;  wr_cycle[ 1324] = 1'b1;  addr_rom[ 1324]='h000014b0;  wr_data_rom[ 1324]='h00000f08;
    rd_cycle[ 1325] = 1'b0;  wr_cycle[ 1325] = 1'b1;  addr_rom[ 1325]='h000014b4;  wr_data_rom[ 1325]='h000002c4;
    rd_cycle[ 1326] = 1'b0;  wr_cycle[ 1326] = 1'b1;  addr_rom[ 1326]='h000014b8;  wr_data_rom[ 1326]='h000017c4;
    rd_cycle[ 1327] = 1'b0;  wr_cycle[ 1327] = 1'b1;  addr_rom[ 1327]='h000014bc;  wr_data_rom[ 1327]='h00001bcb;
    rd_cycle[ 1328] = 1'b0;  wr_cycle[ 1328] = 1'b1;  addr_rom[ 1328]='h000014c0;  wr_data_rom[ 1328]='h00000521;
    rd_cycle[ 1329] = 1'b0;  wr_cycle[ 1329] = 1'b1;  addr_rom[ 1329]='h000014c4;  wr_data_rom[ 1329]='h000013a7;
    rd_cycle[ 1330] = 1'b0;  wr_cycle[ 1330] = 1'b1;  addr_rom[ 1330]='h000014c8;  wr_data_rom[ 1330]='h000006a8;
    rd_cycle[ 1331] = 1'b0;  wr_cycle[ 1331] = 1'b1;  addr_rom[ 1331]='h000014cc;  wr_data_rom[ 1331]='h00000473;
    rd_cycle[ 1332] = 1'b0;  wr_cycle[ 1332] = 1'b1;  addr_rom[ 1332]='h000014d0;  wr_data_rom[ 1332]='h00001416;
    rd_cycle[ 1333] = 1'b0;  wr_cycle[ 1333] = 1'b1;  addr_rom[ 1333]='h000014d4;  wr_data_rom[ 1333]='h00000cc8;
    rd_cycle[ 1334] = 1'b0;  wr_cycle[ 1334] = 1'b1;  addr_rom[ 1334]='h000014d8;  wr_data_rom[ 1334]='h00001d71;
    rd_cycle[ 1335] = 1'b0;  wr_cycle[ 1335] = 1'b1;  addr_rom[ 1335]='h000014dc;  wr_data_rom[ 1335]='h00001228;
    rd_cycle[ 1336] = 1'b0;  wr_cycle[ 1336] = 1'b1;  addr_rom[ 1336]='h000014e0;  wr_data_rom[ 1336]='h000010d2;
    rd_cycle[ 1337] = 1'b0;  wr_cycle[ 1337] = 1'b1;  addr_rom[ 1337]='h000014e4;  wr_data_rom[ 1337]='h00001070;
    rd_cycle[ 1338] = 1'b0;  wr_cycle[ 1338] = 1'b1;  addr_rom[ 1338]='h000014e8;  wr_data_rom[ 1338]='h00000ef2;
    rd_cycle[ 1339] = 1'b0;  wr_cycle[ 1339] = 1'b1;  addr_rom[ 1339]='h000014ec;  wr_data_rom[ 1339]='h000002f1;
    rd_cycle[ 1340] = 1'b0;  wr_cycle[ 1340] = 1'b1;  addr_rom[ 1340]='h000014f0;  wr_data_rom[ 1340]='h00001977;
    rd_cycle[ 1341] = 1'b0;  wr_cycle[ 1341] = 1'b1;  addr_rom[ 1341]='h000014f4;  wr_data_rom[ 1341]='h00000d41;
    rd_cycle[ 1342] = 1'b0;  wr_cycle[ 1342] = 1'b1;  addr_rom[ 1342]='h000014f8;  wr_data_rom[ 1342]='h00001ac1;
    rd_cycle[ 1343] = 1'b0;  wr_cycle[ 1343] = 1'b1;  addr_rom[ 1343]='h000014fc;  wr_data_rom[ 1343]='h00000a1f;
    rd_cycle[ 1344] = 1'b0;  wr_cycle[ 1344] = 1'b1;  addr_rom[ 1344]='h00001500;  wr_data_rom[ 1344]='h00001afa;
    rd_cycle[ 1345] = 1'b0;  wr_cycle[ 1345] = 1'b1;  addr_rom[ 1345]='h00001504;  wr_data_rom[ 1345]='h00001a04;
    rd_cycle[ 1346] = 1'b0;  wr_cycle[ 1346] = 1'b1;  addr_rom[ 1346]='h00001508;  wr_data_rom[ 1346]='h000017d2;
    rd_cycle[ 1347] = 1'b0;  wr_cycle[ 1347] = 1'b1;  addr_rom[ 1347]='h0000150c;  wr_data_rom[ 1347]='h0000133f;
    rd_cycle[ 1348] = 1'b0;  wr_cycle[ 1348] = 1'b1;  addr_rom[ 1348]='h00001510;  wr_data_rom[ 1348]='h00000a7a;
    rd_cycle[ 1349] = 1'b0;  wr_cycle[ 1349] = 1'b1;  addr_rom[ 1349]='h00001514;  wr_data_rom[ 1349]='h00001651;
    rd_cycle[ 1350] = 1'b0;  wr_cycle[ 1350] = 1'b1;  addr_rom[ 1350]='h00001518;  wr_data_rom[ 1350]='h000013e3;
    rd_cycle[ 1351] = 1'b0;  wr_cycle[ 1351] = 1'b1;  addr_rom[ 1351]='h0000151c;  wr_data_rom[ 1351]='h00000bf6;
    rd_cycle[ 1352] = 1'b0;  wr_cycle[ 1352] = 1'b1;  addr_rom[ 1352]='h00001520;  wr_data_rom[ 1352]='h000008fc;
    rd_cycle[ 1353] = 1'b0;  wr_cycle[ 1353] = 1'b1;  addr_rom[ 1353]='h00001524;  wr_data_rom[ 1353]='h00000293;
    rd_cycle[ 1354] = 1'b0;  wr_cycle[ 1354] = 1'b1;  addr_rom[ 1354]='h00001528;  wr_data_rom[ 1354]='h000013df;
    rd_cycle[ 1355] = 1'b0;  wr_cycle[ 1355] = 1'b1;  addr_rom[ 1355]='h0000152c;  wr_data_rom[ 1355]='h00001b39;
    rd_cycle[ 1356] = 1'b0;  wr_cycle[ 1356] = 1'b1;  addr_rom[ 1356]='h00001530;  wr_data_rom[ 1356]='h00000fbb;
    rd_cycle[ 1357] = 1'b0;  wr_cycle[ 1357] = 1'b1;  addr_rom[ 1357]='h00001534;  wr_data_rom[ 1357]='h0000151e;
    rd_cycle[ 1358] = 1'b0;  wr_cycle[ 1358] = 1'b1;  addr_rom[ 1358]='h00001538;  wr_data_rom[ 1358]='h000018b9;
    rd_cycle[ 1359] = 1'b0;  wr_cycle[ 1359] = 1'b1;  addr_rom[ 1359]='h0000153c;  wr_data_rom[ 1359]='h00000f1e;
    rd_cycle[ 1360] = 1'b0;  wr_cycle[ 1360] = 1'b1;  addr_rom[ 1360]='h00001540;  wr_data_rom[ 1360]='h000013f5;
    rd_cycle[ 1361] = 1'b0;  wr_cycle[ 1361] = 1'b1;  addr_rom[ 1361]='h00001544;  wr_data_rom[ 1361]='h00000862;
    rd_cycle[ 1362] = 1'b0;  wr_cycle[ 1362] = 1'b1;  addr_rom[ 1362]='h00001548;  wr_data_rom[ 1362]='h00000327;
    rd_cycle[ 1363] = 1'b0;  wr_cycle[ 1363] = 1'b1;  addr_rom[ 1363]='h0000154c;  wr_data_rom[ 1363]='h00000de9;
    rd_cycle[ 1364] = 1'b0;  wr_cycle[ 1364] = 1'b1;  addr_rom[ 1364]='h00001550;  wr_data_rom[ 1364]='h00001152;
    rd_cycle[ 1365] = 1'b0;  wr_cycle[ 1365] = 1'b1;  addr_rom[ 1365]='h00001554;  wr_data_rom[ 1365]='h000002a2;
    rd_cycle[ 1366] = 1'b0;  wr_cycle[ 1366] = 1'b1;  addr_rom[ 1366]='h00001558;  wr_data_rom[ 1366]='h00000bc5;
    rd_cycle[ 1367] = 1'b0;  wr_cycle[ 1367] = 1'b1;  addr_rom[ 1367]='h0000155c;  wr_data_rom[ 1367]='h00000b77;
    rd_cycle[ 1368] = 1'b0;  wr_cycle[ 1368] = 1'b1;  addr_rom[ 1368]='h00001560;  wr_data_rom[ 1368]='h0000187a;
    rd_cycle[ 1369] = 1'b0;  wr_cycle[ 1369] = 1'b1;  addr_rom[ 1369]='h00001564;  wr_data_rom[ 1369]='h00001102;
    rd_cycle[ 1370] = 1'b0;  wr_cycle[ 1370] = 1'b1;  addr_rom[ 1370]='h00001568;  wr_data_rom[ 1370]='h000005bf;
    rd_cycle[ 1371] = 1'b0;  wr_cycle[ 1371] = 1'b1;  addr_rom[ 1371]='h0000156c;  wr_data_rom[ 1371]='h00000373;
    rd_cycle[ 1372] = 1'b0;  wr_cycle[ 1372] = 1'b1;  addr_rom[ 1372]='h00001570;  wr_data_rom[ 1372]='h00001c1e;
    rd_cycle[ 1373] = 1'b0;  wr_cycle[ 1373] = 1'b1;  addr_rom[ 1373]='h00001574;  wr_data_rom[ 1373]='h00000090;
    rd_cycle[ 1374] = 1'b0;  wr_cycle[ 1374] = 1'b1;  addr_rom[ 1374]='h00001578;  wr_data_rom[ 1374]='h000004bf;
    rd_cycle[ 1375] = 1'b0;  wr_cycle[ 1375] = 1'b1;  addr_rom[ 1375]='h0000157c;  wr_data_rom[ 1375]='h00000b2f;
    rd_cycle[ 1376] = 1'b0;  wr_cycle[ 1376] = 1'b1;  addr_rom[ 1376]='h00001580;  wr_data_rom[ 1376]='h00000296;
    rd_cycle[ 1377] = 1'b0;  wr_cycle[ 1377] = 1'b1;  addr_rom[ 1377]='h00001584;  wr_data_rom[ 1377]='h000010e1;
    rd_cycle[ 1378] = 1'b0;  wr_cycle[ 1378] = 1'b1;  addr_rom[ 1378]='h00001588;  wr_data_rom[ 1378]='h00001b94;
    rd_cycle[ 1379] = 1'b0;  wr_cycle[ 1379] = 1'b1;  addr_rom[ 1379]='h0000158c;  wr_data_rom[ 1379]='h00001677;
    rd_cycle[ 1380] = 1'b0;  wr_cycle[ 1380] = 1'b1;  addr_rom[ 1380]='h00001590;  wr_data_rom[ 1380]='h000013b0;
    rd_cycle[ 1381] = 1'b0;  wr_cycle[ 1381] = 1'b1;  addr_rom[ 1381]='h00001594;  wr_data_rom[ 1381]='h0000008a;
    rd_cycle[ 1382] = 1'b0;  wr_cycle[ 1382] = 1'b1;  addr_rom[ 1382]='h00001598;  wr_data_rom[ 1382]='h000000be;
    rd_cycle[ 1383] = 1'b0;  wr_cycle[ 1383] = 1'b1;  addr_rom[ 1383]='h0000159c;  wr_data_rom[ 1383]='h0000026b;
    rd_cycle[ 1384] = 1'b0;  wr_cycle[ 1384] = 1'b1;  addr_rom[ 1384]='h000015a0;  wr_data_rom[ 1384]='h00000a19;
    rd_cycle[ 1385] = 1'b0;  wr_cycle[ 1385] = 1'b1;  addr_rom[ 1385]='h000015a4;  wr_data_rom[ 1385]='h00001c9e;
    rd_cycle[ 1386] = 1'b0;  wr_cycle[ 1386] = 1'b1;  addr_rom[ 1386]='h000015a8;  wr_data_rom[ 1386]='h00001250;
    rd_cycle[ 1387] = 1'b0;  wr_cycle[ 1387] = 1'b1;  addr_rom[ 1387]='h000015ac;  wr_data_rom[ 1387]='h00001e63;
    rd_cycle[ 1388] = 1'b0;  wr_cycle[ 1388] = 1'b1;  addr_rom[ 1388]='h000015b0;  wr_data_rom[ 1388]='h0000001a;
    rd_cycle[ 1389] = 1'b0;  wr_cycle[ 1389] = 1'b1;  addr_rom[ 1389]='h000015b4;  wr_data_rom[ 1389]='h00001349;
    rd_cycle[ 1390] = 1'b0;  wr_cycle[ 1390] = 1'b1;  addr_rom[ 1390]='h000015b8;  wr_data_rom[ 1390]='h000017cc;
    rd_cycle[ 1391] = 1'b0;  wr_cycle[ 1391] = 1'b1;  addr_rom[ 1391]='h000015bc;  wr_data_rom[ 1391]='h000003f7;
    rd_cycle[ 1392] = 1'b0;  wr_cycle[ 1392] = 1'b1;  addr_rom[ 1392]='h000015c0;  wr_data_rom[ 1392]='h0000035c;
    rd_cycle[ 1393] = 1'b0;  wr_cycle[ 1393] = 1'b1;  addr_rom[ 1393]='h000015c4;  wr_data_rom[ 1393]='h000018ae;
    rd_cycle[ 1394] = 1'b0;  wr_cycle[ 1394] = 1'b1;  addr_rom[ 1394]='h000015c8;  wr_data_rom[ 1394]='h0000143e;
    rd_cycle[ 1395] = 1'b0;  wr_cycle[ 1395] = 1'b1;  addr_rom[ 1395]='h000015cc;  wr_data_rom[ 1395]='h0000167b;
    rd_cycle[ 1396] = 1'b0;  wr_cycle[ 1396] = 1'b1;  addr_rom[ 1396]='h000015d0;  wr_data_rom[ 1396]='h0000109d;
    rd_cycle[ 1397] = 1'b0;  wr_cycle[ 1397] = 1'b1;  addr_rom[ 1397]='h000015d4;  wr_data_rom[ 1397]='h00000188;
    rd_cycle[ 1398] = 1'b0;  wr_cycle[ 1398] = 1'b1;  addr_rom[ 1398]='h000015d8;  wr_data_rom[ 1398]='h00000411;
    rd_cycle[ 1399] = 1'b0;  wr_cycle[ 1399] = 1'b1;  addr_rom[ 1399]='h000015dc;  wr_data_rom[ 1399]='h00000d0b;
    rd_cycle[ 1400] = 1'b0;  wr_cycle[ 1400] = 1'b1;  addr_rom[ 1400]='h000015e0;  wr_data_rom[ 1400]='h00000862;
    rd_cycle[ 1401] = 1'b0;  wr_cycle[ 1401] = 1'b1;  addr_rom[ 1401]='h000015e4;  wr_data_rom[ 1401]='h000008bb;
    rd_cycle[ 1402] = 1'b0;  wr_cycle[ 1402] = 1'b1;  addr_rom[ 1402]='h000015e8;  wr_data_rom[ 1402]='h00001723;
    rd_cycle[ 1403] = 1'b0;  wr_cycle[ 1403] = 1'b1;  addr_rom[ 1403]='h000015ec;  wr_data_rom[ 1403]='h00001068;
    rd_cycle[ 1404] = 1'b0;  wr_cycle[ 1404] = 1'b1;  addr_rom[ 1404]='h000015f0;  wr_data_rom[ 1404]='h00000913;
    rd_cycle[ 1405] = 1'b0;  wr_cycle[ 1405] = 1'b1;  addr_rom[ 1405]='h000015f4;  wr_data_rom[ 1405]='h00000983;
    rd_cycle[ 1406] = 1'b0;  wr_cycle[ 1406] = 1'b1;  addr_rom[ 1406]='h000015f8;  wr_data_rom[ 1406]='h00001122;
    rd_cycle[ 1407] = 1'b0;  wr_cycle[ 1407] = 1'b1;  addr_rom[ 1407]='h000015fc;  wr_data_rom[ 1407]='h0000010c;
    rd_cycle[ 1408] = 1'b0;  wr_cycle[ 1408] = 1'b1;  addr_rom[ 1408]='h00001600;  wr_data_rom[ 1408]='h000000cf;
    rd_cycle[ 1409] = 1'b0;  wr_cycle[ 1409] = 1'b1;  addr_rom[ 1409]='h00001604;  wr_data_rom[ 1409]='h000005ae;
    rd_cycle[ 1410] = 1'b0;  wr_cycle[ 1410] = 1'b1;  addr_rom[ 1410]='h00001608;  wr_data_rom[ 1410]='h00000a45;
    rd_cycle[ 1411] = 1'b0;  wr_cycle[ 1411] = 1'b1;  addr_rom[ 1411]='h0000160c;  wr_data_rom[ 1411]='h00000f49;
    rd_cycle[ 1412] = 1'b0;  wr_cycle[ 1412] = 1'b1;  addr_rom[ 1412]='h00001610;  wr_data_rom[ 1412]='h00001a36;
    rd_cycle[ 1413] = 1'b0;  wr_cycle[ 1413] = 1'b1;  addr_rom[ 1413]='h00001614;  wr_data_rom[ 1413]='h000016c4;
    rd_cycle[ 1414] = 1'b0;  wr_cycle[ 1414] = 1'b1;  addr_rom[ 1414]='h00001618;  wr_data_rom[ 1414]='h000006ea;
    rd_cycle[ 1415] = 1'b0;  wr_cycle[ 1415] = 1'b1;  addr_rom[ 1415]='h0000161c;  wr_data_rom[ 1415]='h000000d5;
    rd_cycle[ 1416] = 1'b0;  wr_cycle[ 1416] = 1'b1;  addr_rom[ 1416]='h00001620;  wr_data_rom[ 1416]='h00000e70;
    rd_cycle[ 1417] = 1'b0;  wr_cycle[ 1417] = 1'b1;  addr_rom[ 1417]='h00001624;  wr_data_rom[ 1417]='h000016db;
    rd_cycle[ 1418] = 1'b0;  wr_cycle[ 1418] = 1'b1;  addr_rom[ 1418]='h00001628;  wr_data_rom[ 1418]='h00001047;
    rd_cycle[ 1419] = 1'b0;  wr_cycle[ 1419] = 1'b1;  addr_rom[ 1419]='h0000162c;  wr_data_rom[ 1419]='h00000f1c;
    rd_cycle[ 1420] = 1'b0;  wr_cycle[ 1420] = 1'b1;  addr_rom[ 1420]='h00001630;  wr_data_rom[ 1420]='h00000f5f;
    rd_cycle[ 1421] = 1'b0;  wr_cycle[ 1421] = 1'b1;  addr_rom[ 1421]='h00001634;  wr_data_rom[ 1421]='h00001a56;
    rd_cycle[ 1422] = 1'b0;  wr_cycle[ 1422] = 1'b1;  addr_rom[ 1422]='h00001638;  wr_data_rom[ 1422]='h00000a0b;
    rd_cycle[ 1423] = 1'b0;  wr_cycle[ 1423] = 1'b1;  addr_rom[ 1423]='h0000163c;  wr_data_rom[ 1423]='h0000195c;
    rd_cycle[ 1424] = 1'b0;  wr_cycle[ 1424] = 1'b1;  addr_rom[ 1424]='h00001640;  wr_data_rom[ 1424]='h000016cf;
    rd_cycle[ 1425] = 1'b0;  wr_cycle[ 1425] = 1'b1;  addr_rom[ 1425]='h00001644;  wr_data_rom[ 1425]='h00001450;
    rd_cycle[ 1426] = 1'b0;  wr_cycle[ 1426] = 1'b1;  addr_rom[ 1426]='h00001648;  wr_data_rom[ 1426]='h00000533;
    rd_cycle[ 1427] = 1'b0;  wr_cycle[ 1427] = 1'b1;  addr_rom[ 1427]='h0000164c;  wr_data_rom[ 1427]='h00000065;
    rd_cycle[ 1428] = 1'b0;  wr_cycle[ 1428] = 1'b1;  addr_rom[ 1428]='h00001650;  wr_data_rom[ 1428]='h000001cf;
    rd_cycle[ 1429] = 1'b0;  wr_cycle[ 1429] = 1'b1;  addr_rom[ 1429]='h00001654;  wr_data_rom[ 1429]='h000014f4;
    rd_cycle[ 1430] = 1'b0;  wr_cycle[ 1430] = 1'b1;  addr_rom[ 1430]='h00001658;  wr_data_rom[ 1430]='h00000926;
    rd_cycle[ 1431] = 1'b0;  wr_cycle[ 1431] = 1'b1;  addr_rom[ 1431]='h0000165c;  wr_data_rom[ 1431]='h00001289;
    rd_cycle[ 1432] = 1'b0;  wr_cycle[ 1432] = 1'b1;  addr_rom[ 1432]='h00001660;  wr_data_rom[ 1432]='h00000ffa;
    rd_cycle[ 1433] = 1'b0;  wr_cycle[ 1433] = 1'b1;  addr_rom[ 1433]='h00001664;  wr_data_rom[ 1433]='h00001a1e;
    rd_cycle[ 1434] = 1'b0;  wr_cycle[ 1434] = 1'b1;  addr_rom[ 1434]='h00001668;  wr_data_rom[ 1434]='h00000775;
    rd_cycle[ 1435] = 1'b0;  wr_cycle[ 1435] = 1'b1;  addr_rom[ 1435]='h0000166c;  wr_data_rom[ 1435]='h00001ade;
    rd_cycle[ 1436] = 1'b0;  wr_cycle[ 1436] = 1'b1;  addr_rom[ 1436]='h00001670;  wr_data_rom[ 1436]='h00000cee;
    rd_cycle[ 1437] = 1'b0;  wr_cycle[ 1437] = 1'b1;  addr_rom[ 1437]='h00001674;  wr_data_rom[ 1437]='h00000dbf;
    rd_cycle[ 1438] = 1'b0;  wr_cycle[ 1438] = 1'b1;  addr_rom[ 1438]='h00001678;  wr_data_rom[ 1438]='h00000a56;
    rd_cycle[ 1439] = 1'b0;  wr_cycle[ 1439] = 1'b1;  addr_rom[ 1439]='h0000167c;  wr_data_rom[ 1439]='h00001826;
    rd_cycle[ 1440] = 1'b0;  wr_cycle[ 1440] = 1'b1;  addr_rom[ 1440]='h00001680;  wr_data_rom[ 1440]='h000002e3;
    rd_cycle[ 1441] = 1'b0;  wr_cycle[ 1441] = 1'b1;  addr_rom[ 1441]='h00001684;  wr_data_rom[ 1441]='h000002f0;
    rd_cycle[ 1442] = 1'b0;  wr_cycle[ 1442] = 1'b1;  addr_rom[ 1442]='h00001688;  wr_data_rom[ 1442]='h0000101a;
    rd_cycle[ 1443] = 1'b0;  wr_cycle[ 1443] = 1'b1;  addr_rom[ 1443]='h0000168c;  wr_data_rom[ 1443]='h00001ac0;
    rd_cycle[ 1444] = 1'b0;  wr_cycle[ 1444] = 1'b1;  addr_rom[ 1444]='h00001690;  wr_data_rom[ 1444]='h0000151a;
    rd_cycle[ 1445] = 1'b0;  wr_cycle[ 1445] = 1'b1;  addr_rom[ 1445]='h00001694;  wr_data_rom[ 1445]='h00000f1f;
    rd_cycle[ 1446] = 1'b0;  wr_cycle[ 1446] = 1'b1;  addr_rom[ 1446]='h00001698;  wr_data_rom[ 1446]='h000017c0;
    rd_cycle[ 1447] = 1'b0;  wr_cycle[ 1447] = 1'b1;  addr_rom[ 1447]='h0000169c;  wr_data_rom[ 1447]='h00000f19;
    rd_cycle[ 1448] = 1'b0;  wr_cycle[ 1448] = 1'b1;  addr_rom[ 1448]='h000016a0;  wr_data_rom[ 1448]='h000018e8;
    rd_cycle[ 1449] = 1'b0;  wr_cycle[ 1449] = 1'b1;  addr_rom[ 1449]='h000016a4;  wr_data_rom[ 1449]='h00000ddf;
    rd_cycle[ 1450] = 1'b0;  wr_cycle[ 1450] = 1'b1;  addr_rom[ 1450]='h000016a8;  wr_data_rom[ 1450]='h00001077;
    rd_cycle[ 1451] = 1'b0;  wr_cycle[ 1451] = 1'b1;  addr_rom[ 1451]='h000016ac;  wr_data_rom[ 1451]='h00001217;
    rd_cycle[ 1452] = 1'b0;  wr_cycle[ 1452] = 1'b1;  addr_rom[ 1452]='h000016b0;  wr_data_rom[ 1452]='h00001c94;
    rd_cycle[ 1453] = 1'b0;  wr_cycle[ 1453] = 1'b1;  addr_rom[ 1453]='h000016b4;  wr_data_rom[ 1453]='h00001c8a;
    rd_cycle[ 1454] = 1'b0;  wr_cycle[ 1454] = 1'b1;  addr_rom[ 1454]='h000016b8;  wr_data_rom[ 1454]='h00000847;
    rd_cycle[ 1455] = 1'b0;  wr_cycle[ 1455] = 1'b1;  addr_rom[ 1455]='h000016bc;  wr_data_rom[ 1455]='h00001723;
    rd_cycle[ 1456] = 1'b0;  wr_cycle[ 1456] = 1'b1;  addr_rom[ 1456]='h000016c0;  wr_data_rom[ 1456]='h000014af;
    rd_cycle[ 1457] = 1'b0;  wr_cycle[ 1457] = 1'b1;  addr_rom[ 1457]='h000016c4;  wr_data_rom[ 1457]='h000015ea;
    rd_cycle[ 1458] = 1'b0;  wr_cycle[ 1458] = 1'b1;  addr_rom[ 1458]='h000016c8;  wr_data_rom[ 1458]='h00001b8a;
    rd_cycle[ 1459] = 1'b0;  wr_cycle[ 1459] = 1'b1;  addr_rom[ 1459]='h000016cc;  wr_data_rom[ 1459]='h0000117a;
    rd_cycle[ 1460] = 1'b0;  wr_cycle[ 1460] = 1'b1;  addr_rom[ 1460]='h000016d0;  wr_data_rom[ 1460]='h00000342;
    rd_cycle[ 1461] = 1'b0;  wr_cycle[ 1461] = 1'b1;  addr_rom[ 1461]='h000016d4;  wr_data_rom[ 1461]='h00001c71;
    rd_cycle[ 1462] = 1'b0;  wr_cycle[ 1462] = 1'b1;  addr_rom[ 1462]='h000016d8;  wr_data_rom[ 1462]='h00001d1e;
    rd_cycle[ 1463] = 1'b0;  wr_cycle[ 1463] = 1'b1;  addr_rom[ 1463]='h000016dc;  wr_data_rom[ 1463]='h0000005a;
    rd_cycle[ 1464] = 1'b0;  wr_cycle[ 1464] = 1'b1;  addr_rom[ 1464]='h000016e0;  wr_data_rom[ 1464]='h000007f4;
    rd_cycle[ 1465] = 1'b0;  wr_cycle[ 1465] = 1'b1;  addr_rom[ 1465]='h000016e4;  wr_data_rom[ 1465]='h00000d37;
    rd_cycle[ 1466] = 1'b0;  wr_cycle[ 1466] = 1'b1;  addr_rom[ 1466]='h000016e8;  wr_data_rom[ 1466]='h00000576;
    rd_cycle[ 1467] = 1'b0;  wr_cycle[ 1467] = 1'b1;  addr_rom[ 1467]='h000016ec;  wr_data_rom[ 1467]='h00001dc8;
    rd_cycle[ 1468] = 1'b0;  wr_cycle[ 1468] = 1'b1;  addr_rom[ 1468]='h000016f0;  wr_data_rom[ 1468]='h00000754;
    rd_cycle[ 1469] = 1'b0;  wr_cycle[ 1469] = 1'b1;  addr_rom[ 1469]='h000016f4;  wr_data_rom[ 1469]='h000013c2;
    rd_cycle[ 1470] = 1'b0;  wr_cycle[ 1470] = 1'b1;  addr_rom[ 1470]='h000016f8;  wr_data_rom[ 1470]='h00000bb8;
    rd_cycle[ 1471] = 1'b0;  wr_cycle[ 1471] = 1'b1;  addr_rom[ 1471]='h000016fc;  wr_data_rom[ 1471]='h00001623;
    rd_cycle[ 1472] = 1'b0;  wr_cycle[ 1472] = 1'b1;  addr_rom[ 1472]='h00001700;  wr_data_rom[ 1472]='h00001a1f;
    rd_cycle[ 1473] = 1'b0;  wr_cycle[ 1473] = 1'b1;  addr_rom[ 1473]='h00001704;  wr_data_rom[ 1473]='h00001afc;
    rd_cycle[ 1474] = 1'b0;  wr_cycle[ 1474] = 1'b1;  addr_rom[ 1474]='h00001708;  wr_data_rom[ 1474]='h00000477;
    rd_cycle[ 1475] = 1'b0;  wr_cycle[ 1475] = 1'b1;  addr_rom[ 1475]='h0000170c;  wr_data_rom[ 1475]='h00000cda;
    rd_cycle[ 1476] = 1'b0;  wr_cycle[ 1476] = 1'b1;  addr_rom[ 1476]='h00001710;  wr_data_rom[ 1476]='h00000875;
    rd_cycle[ 1477] = 1'b0;  wr_cycle[ 1477] = 1'b1;  addr_rom[ 1477]='h00001714;  wr_data_rom[ 1477]='h00000cf1;
    rd_cycle[ 1478] = 1'b0;  wr_cycle[ 1478] = 1'b1;  addr_rom[ 1478]='h00001718;  wr_data_rom[ 1478]='h00000b3f;
    rd_cycle[ 1479] = 1'b0;  wr_cycle[ 1479] = 1'b1;  addr_rom[ 1479]='h0000171c;  wr_data_rom[ 1479]='h00000085;
    rd_cycle[ 1480] = 1'b0;  wr_cycle[ 1480] = 1'b1;  addr_rom[ 1480]='h00001720;  wr_data_rom[ 1480]='h00001d09;
    rd_cycle[ 1481] = 1'b0;  wr_cycle[ 1481] = 1'b1;  addr_rom[ 1481]='h00001724;  wr_data_rom[ 1481]='h000014fe;
    rd_cycle[ 1482] = 1'b0;  wr_cycle[ 1482] = 1'b1;  addr_rom[ 1482]='h00001728;  wr_data_rom[ 1482]='h00000b06;
    rd_cycle[ 1483] = 1'b0;  wr_cycle[ 1483] = 1'b1;  addr_rom[ 1483]='h0000172c;  wr_data_rom[ 1483]='h00001720;
    rd_cycle[ 1484] = 1'b0;  wr_cycle[ 1484] = 1'b1;  addr_rom[ 1484]='h00001730;  wr_data_rom[ 1484]='h00000bb5;
    rd_cycle[ 1485] = 1'b0;  wr_cycle[ 1485] = 1'b1;  addr_rom[ 1485]='h00001734;  wr_data_rom[ 1485]='h00000892;
    rd_cycle[ 1486] = 1'b0;  wr_cycle[ 1486] = 1'b1;  addr_rom[ 1486]='h00001738;  wr_data_rom[ 1486]='h000008f6;
    rd_cycle[ 1487] = 1'b0;  wr_cycle[ 1487] = 1'b1;  addr_rom[ 1487]='h0000173c;  wr_data_rom[ 1487]='h000012ea;
    rd_cycle[ 1488] = 1'b0;  wr_cycle[ 1488] = 1'b1;  addr_rom[ 1488]='h00001740;  wr_data_rom[ 1488]='h000004e4;
    rd_cycle[ 1489] = 1'b0;  wr_cycle[ 1489] = 1'b1;  addr_rom[ 1489]='h00001744;  wr_data_rom[ 1489]='h00000cb3;
    rd_cycle[ 1490] = 1'b0;  wr_cycle[ 1490] = 1'b1;  addr_rom[ 1490]='h00001748;  wr_data_rom[ 1490]='h000013e7;
    rd_cycle[ 1491] = 1'b0;  wr_cycle[ 1491] = 1'b1;  addr_rom[ 1491]='h0000174c;  wr_data_rom[ 1491]='h00001c93;
    rd_cycle[ 1492] = 1'b0;  wr_cycle[ 1492] = 1'b1;  addr_rom[ 1492]='h00001750;  wr_data_rom[ 1492]='h000019b0;
    rd_cycle[ 1493] = 1'b0;  wr_cycle[ 1493] = 1'b1;  addr_rom[ 1493]='h00001754;  wr_data_rom[ 1493]='h00000ac7;
    rd_cycle[ 1494] = 1'b0;  wr_cycle[ 1494] = 1'b1;  addr_rom[ 1494]='h00001758;  wr_data_rom[ 1494]='h00001eb5;
    rd_cycle[ 1495] = 1'b0;  wr_cycle[ 1495] = 1'b1;  addr_rom[ 1495]='h0000175c;  wr_data_rom[ 1495]='h00000004;
    rd_cycle[ 1496] = 1'b0;  wr_cycle[ 1496] = 1'b1;  addr_rom[ 1496]='h00001760;  wr_data_rom[ 1496]='h00000f52;
    rd_cycle[ 1497] = 1'b0;  wr_cycle[ 1497] = 1'b1;  addr_rom[ 1497]='h00001764;  wr_data_rom[ 1497]='h00001688;
    rd_cycle[ 1498] = 1'b0;  wr_cycle[ 1498] = 1'b1;  addr_rom[ 1498]='h00001768;  wr_data_rom[ 1498]='h00001018;
    rd_cycle[ 1499] = 1'b0;  wr_cycle[ 1499] = 1'b1;  addr_rom[ 1499]='h0000176c;  wr_data_rom[ 1499]='h00000e5b;
    rd_cycle[ 1500] = 1'b0;  wr_cycle[ 1500] = 1'b1;  addr_rom[ 1500]='h00001770;  wr_data_rom[ 1500]='h00000b6a;
    rd_cycle[ 1501] = 1'b0;  wr_cycle[ 1501] = 1'b1;  addr_rom[ 1501]='h00001774;  wr_data_rom[ 1501]='h00001ca1;
    rd_cycle[ 1502] = 1'b0;  wr_cycle[ 1502] = 1'b1;  addr_rom[ 1502]='h00001778;  wr_data_rom[ 1502]='h00000902;
    rd_cycle[ 1503] = 1'b0;  wr_cycle[ 1503] = 1'b1;  addr_rom[ 1503]='h0000177c;  wr_data_rom[ 1503]='h0000151b;
    rd_cycle[ 1504] = 1'b0;  wr_cycle[ 1504] = 1'b1;  addr_rom[ 1504]='h00001780;  wr_data_rom[ 1504]='h0000007f;
    rd_cycle[ 1505] = 1'b0;  wr_cycle[ 1505] = 1'b1;  addr_rom[ 1505]='h00001784;  wr_data_rom[ 1505]='h0000138a;
    rd_cycle[ 1506] = 1'b0;  wr_cycle[ 1506] = 1'b1;  addr_rom[ 1506]='h00001788;  wr_data_rom[ 1506]='h000000b2;
    rd_cycle[ 1507] = 1'b0;  wr_cycle[ 1507] = 1'b1;  addr_rom[ 1507]='h0000178c;  wr_data_rom[ 1507]='h000009b5;
    rd_cycle[ 1508] = 1'b0;  wr_cycle[ 1508] = 1'b1;  addr_rom[ 1508]='h00001790;  wr_data_rom[ 1508]='h00000cd6;
    rd_cycle[ 1509] = 1'b0;  wr_cycle[ 1509] = 1'b1;  addr_rom[ 1509]='h00001794;  wr_data_rom[ 1509]='h00001c8c;
    rd_cycle[ 1510] = 1'b0;  wr_cycle[ 1510] = 1'b1;  addr_rom[ 1510]='h00001798;  wr_data_rom[ 1510]='h00001d6b;
    rd_cycle[ 1511] = 1'b0;  wr_cycle[ 1511] = 1'b1;  addr_rom[ 1511]='h0000179c;  wr_data_rom[ 1511]='h00001b40;
    rd_cycle[ 1512] = 1'b0;  wr_cycle[ 1512] = 1'b1;  addr_rom[ 1512]='h000017a0;  wr_data_rom[ 1512]='h000004a6;
    rd_cycle[ 1513] = 1'b0;  wr_cycle[ 1513] = 1'b1;  addr_rom[ 1513]='h000017a4;  wr_data_rom[ 1513]='h00000252;
    rd_cycle[ 1514] = 1'b0;  wr_cycle[ 1514] = 1'b1;  addr_rom[ 1514]='h000017a8;  wr_data_rom[ 1514]='h000008a7;
    rd_cycle[ 1515] = 1'b0;  wr_cycle[ 1515] = 1'b1;  addr_rom[ 1515]='h000017ac;  wr_data_rom[ 1515]='h00000c5e;
    rd_cycle[ 1516] = 1'b0;  wr_cycle[ 1516] = 1'b1;  addr_rom[ 1516]='h000017b0;  wr_data_rom[ 1516]='h000007ed;
    rd_cycle[ 1517] = 1'b0;  wr_cycle[ 1517] = 1'b1;  addr_rom[ 1517]='h000017b4;  wr_data_rom[ 1517]='h00000abe;
    rd_cycle[ 1518] = 1'b0;  wr_cycle[ 1518] = 1'b1;  addr_rom[ 1518]='h000017b8;  wr_data_rom[ 1518]='h00001314;
    rd_cycle[ 1519] = 1'b0;  wr_cycle[ 1519] = 1'b1;  addr_rom[ 1519]='h000017bc;  wr_data_rom[ 1519]='h0000118d;
    rd_cycle[ 1520] = 1'b0;  wr_cycle[ 1520] = 1'b1;  addr_rom[ 1520]='h000017c0;  wr_data_rom[ 1520]='h00000660;
    rd_cycle[ 1521] = 1'b0;  wr_cycle[ 1521] = 1'b1;  addr_rom[ 1521]='h000017c4;  wr_data_rom[ 1521]='h0000062d;
    rd_cycle[ 1522] = 1'b0;  wr_cycle[ 1522] = 1'b1;  addr_rom[ 1522]='h000017c8;  wr_data_rom[ 1522]='h000009f8;
    rd_cycle[ 1523] = 1'b0;  wr_cycle[ 1523] = 1'b1;  addr_rom[ 1523]='h000017cc;  wr_data_rom[ 1523]='h00001f1f;
    rd_cycle[ 1524] = 1'b0;  wr_cycle[ 1524] = 1'b1;  addr_rom[ 1524]='h000017d0;  wr_data_rom[ 1524]='h000010e2;
    rd_cycle[ 1525] = 1'b0;  wr_cycle[ 1525] = 1'b1;  addr_rom[ 1525]='h000017d4;  wr_data_rom[ 1525]='h00001be9;
    rd_cycle[ 1526] = 1'b0;  wr_cycle[ 1526] = 1'b1;  addr_rom[ 1526]='h000017d8;  wr_data_rom[ 1526]='h0000174b;
    rd_cycle[ 1527] = 1'b0;  wr_cycle[ 1527] = 1'b1;  addr_rom[ 1527]='h000017dc;  wr_data_rom[ 1527]='h000003d5;
    rd_cycle[ 1528] = 1'b0;  wr_cycle[ 1528] = 1'b1;  addr_rom[ 1528]='h000017e0;  wr_data_rom[ 1528]='h00001271;
    rd_cycle[ 1529] = 1'b0;  wr_cycle[ 1529] = 1'b1;  addr_rom[ 1529]='h000017e4;  wr_data_rom[ 1529]='h00000be5;
    rd_cycle[ 1530] = 1'b0;  wr_cycle[ 1530] = 1'b1;  addr_rom[ 1530]='h000017e8;  wr_data_rom[ 1530]='h00000983;
    rd_cycle[ 1531] = 1'b0;  wr_cycle[ 1531] = 1'b1;  addr_rom[ 1531]='h000017ec;  wr_data_rom[ 1531]='h00001b46;
    rd_cycle[ 1532] = 1'b0;  wr_cycle[ 1532] = 1'b1;  addr_rom[ 1532]='h000017f0;  wr_data_rom[ 1532]='h00000da2;
    rd_cycle[ 1533] = 1'b0;  wr_cycle[ 1533] = 1'b1;  addr_rom[ 1533]='h000017f4;  wr_data_rom[ 1533]='h00001033;
    rd_cycle[ 1534] = 1'b0;  wr_cycle[ 1534] = 1'b1;  addr_rom[ 1534]='h000017f8;  wr_data_rom[ 1534]='h00001ae9;
    rd_cycle[ 1535] = 1'b0;  wr_cycle[ 1535] = 1'b1;  addr_rom[ 1535]='h000017fc;  wr_data_rom[ 1535]='h00000afb;
    rd_cycle[ 1536] = 1'b0;  wr_cycle[ 1536] = 1'b1;  addr_rom[ 1536]='h00001800;  wr_data_rom[ 1536]='h00000d54;
    rd_cycle[ 1537] = 1'b0;  wr_cycle[ 1537] = 1'b1;  addr_rom[ 1537]='h00001804;  wr_data_rom[ 1537]='h0000061b;
    rd_cycle[ 1538] = 1'b0;  wr_cycle[ 1538] = 1'b1;  addr_rom[ 1538]='h00001808;  wr_data_rom[ 1538]='h00001bdc;
    rd_cycle[ 1539] = 1'b0;  wr_cycle[ 1539] = 1'b1;  addr_rom[ 1539]='h0000180c;  wr_data_rom[ 1539]='h000019af;
    rd_cycle[ 1540] = 1'b0;  wr_cycle[ 1540] = 1'b1;  addr_rom[ 1540]='h00001810;  wr_data_rom[ 1540]='h000015d2;
    rd_cycle[ 1541] = 1'b0;  wr_cycle[ 1541] = 1'b1;  addr_rom[ 1541]='h00001814;  wr_data_rom[ 1541]='h00000e7c;
    rd_cycle[ 1542] = 1'b0;  wr_cycle[ 1542] = 1'b1;  addr_rom[ 1542]='h00001818;  wr_data_rom[ 1542]='h00000234;
    rd_cycle[ 1543] = 1'b0;  wr_cycle[ 1543] = 1'b1;  addr_rom[ 1543]='h0000181c;  wr_data_rom[ 1543]='h000019e5;
    rd_cycle[ 1544] = 1'b0;  wr_cycle[ 1544] = 1'b1;  addr_rom[ 1544]='h00001820;  wr_data_rom[ 1544]='h00000d0d;
    rd_cycle[ 1545] = 1'b0;  wr_cycle[ 1545] = 1'b1;  addr_rom[ 1545]='h00001824;  wr_data_rom[ 1545]='h0000136f;
    rd_cycle[ 1546] = 1'b0;  wr_cycle[ 1546] = 1'b1;  addr_rom[ 1546]='h00001828;  wr_data_rom[ 1546]='h00000a48;
    rd_cycle[ 1547] = 1'b0;  wr_cycle[ 1547] = 1'b1;  addr_rom[ 1547]='h0000182c;  wr_data_rom[ 1547]='h00001d36;
    rd_cycle[ 1548] = 1'b0;  wr_cycle[ 1548] = 1'b1;  addr_rom[ 1548]='h00001830;  wr_data_rom[ 1548]='h00001a6d;
    rd_cycle[ 1549] = 1'b0;  wr_cycle[ 1549] = 1'b1;  addr_rom[ 1549]='h00001834;  wr_data_rom[ 1549]='h00001b66;
    rd_cycle[ 1550] = 1'b0;  wr_cycle[ 1550] = 1'b1;  addr_rom[ 1550]='h00001838;  wr_data_rom[ 1550]='h000017cb;
    rd_cycle[ 1551] = 1'b0;  wr_cycle[ 1551] = 1'b1;  addr_rom[ 1551]='h0000183c;  wr_data_rom[ 1551]='h00001d29;
    rd_cycle[ 1552] = 1'b0;  wr_cycle[ 1552] = 1'b1;  addr_rom[ 1552]='h00001840;  wr_data_rom[ 1552]='h00001aae;
    rd_cycle[ 1553] = 1'b0;  wr_cycle[ 1553] = 1'b1;  addr_rom[ 1553]='h00001844;  wr_data_rom[ 1553]='h00000797;
    rd_cycle[ 1554] = 1'b0;  wr_cycle[ 1554] = 1'b1;  addr_rom[ 1554]='h00001848;  wr_data_rom[ 1554]='h0000126b;
    rd_cycle[ 1555] = 1'b0;  wr_cycle[ 1555] = 1'b1;  addr_rom[ 1555]='h0000184c;  wr_data_rom[ 1555]='h00001b45;
    rd_cycle[ 1556] = 1'b0;  wr_cycle[ 1556] = 1'b1;  addr_rom[ 1556]='h00001850;  wr_data_rom[ 1556]='h00001879;
    rd_cycle[ 1557] = 1'b0;  wr_cycle[ 1557] = 1'b1;  addr_rom[ 1557]='h00001854;  wr_data_rom[ 1557]='h000014c7;
    rd_cycle[ 1558] = 1'b0;  wr_cycle[ 1558] = 1'b1;  addr_rom[ 1558]='h00001858;  wr_data_rom[ 1558]='h00000f61;
    rd_cycle[ 1559] = 1'b0;  wr_cycle[ 1559] = 1'b1;  addr_rom[ 1559]='h0000185c;  wr_data_rom[ 1559]='h00000845;
    rd_cycle[ 1560] = 1'b0;  wr_cycle[ 1560] = 1'b1;  addr_rom[ 1560]='h00001860;  wr_data_rom[ 1560]='h00000bee;
    rd_cycle[ 1561] = 1'b0;  wr_cycle[ 1561] = 1'b1;  addr_rom[ 1561]='h00001864;  wr_data_rom[ 1561]='h00000153;
    rd_cycle[ 1562] = 1'b0;  wr_cycle[ 1562] = 1'b1;  addr_rom[ 1562]='h00001868;  wr_data_rom[ 1562]='h0000013a;
    rd_cycle[ 1563] = 1'b0;  wr_cycle[ 1563] = 1'b1;  addr_rom[ 1563]='h0000186c;  wr_data_rom[ 1563]='h000009b1;
    rd_cycle[ 1564] = 1'b0;  wr_cycle[ 1564] = 1'b1;  addr_rom[ 1564]='h00001870;  wr_data_rom[ 1564]='h00001e38;
    rd_cycle[ 1565] = 1'b0;  wr_cycle[ 1565] = 1'b1;  addr_rom[ 1565]='h00001874;  wr_data_rom[ 1565]='h00000450;
    rd_cycle[ 1566] = 1'b0;  wr_cycle[ 1566] = 1'b1;  addr_rom[ 1566]='h00001878;  wr_data_rom[ 1566]='h0000181b;
    rd_cycle[ 1567] = 1'b0;  wr_cycle[ 1567] = 1'b1;  addr_rom[ 1567]='h0000187c;  wr_data_rom[ 1567]='h00000698;
    rd_cycle[ 1568] = 1'b0;  wr_cycle[ 1568] = 1'b1;  addr_rom[ 1568]='h00001880;  wr_data_rom[ 1568]='h00001ecf;
    rd_cycle[ 1569] = 1'b0;  wr_cycle[ 1569] = 1'b1;  addr_rom[ 1569]='h00001884;  wr_data_rom[ 1569]='h000000df;
    rd_cycle[ 1570] = 1'b0;  wr_cycle[ 1570] = 1'b1;  addr_rom[ 1570]='h00001888;  wr_data_rom[ 1570]='h00000814;
    rd_cycle[ 1571] = 1'b0;  wr_cycle[ 1571] = 1'b1;  addr_rom[ 1571]='h0000188c;  wr_data_rom[ 1571]='h0000091f;
    rd_cycle[ 1572] = 1'b0;  wr_cycle[ 1572] = 1'b1;  addr_rom[ 1572]='h00001890;  wr_data_rom[ 1572]='h00001a99;
    rd_cycle[ 1573] = 1'b0;  wr_cycle[ 1573] = 1'b1;  addr_rom[ 1573]='h00001894;  wr_data_rom[ 1573]='h00000c1b;
    rd_cycle[ 1574] = 1'b0;  wr_cycle[ 1574] = 1'b1;  addr_rom[ 1574]='h00001898;  wr_data_rom[ 1574]='h000010bf;
    rd_cycle[ 1575] = 1'b0;  wr_cycle[ 1575] = 1'b1;  addr_rom[ 1575]='h0000189c;  wr_data_rom[ 1575]='h00000696;
    rd_cycle[ 1576] = 1'b0;  wr_cycle[ 1576] = 1'b1;  addr_rom[ 1576]='h000018a0;  wr_data_rom[ 1576]='h00000e11;
    rd_cycle[ 1577] = 1'b0;  wr_cycle[ 1577] = 1'b1;  addr_rom[ 1577]='h000018a4;  wr_data_rom[ 1577]='h00001ae9;
    rd_cycle[ 1578] = 1'b0;  wr_cycle[ 1578] = 1'b1;  addr_rom[ 1578]='h000018a8;  wr_data_rom[ 1578]='h00000684;
    rd_cycle[ 1579] = 1'b0;  wr_cycle[ 1579] = 1'b1;  addr_rom[ 1579]='h000018ac;  wr_data_rom[ 1579]='h00000776;
    rd_cycle[ 1580] = 1'b0;  wr_cycle[ 1580] = 1'b1;  addr_rom[ 1580]='h000018b0;  wr_data_rom[ 1580]='h0000176a;
    rd_cycle[ 1581] = 1'b0;  wr_cycle[ 1581] = 1'b1;  addr_rom[ 1581]='h000018b4;  wr_data_rom[ 1581]='h00001532;
    rd_cycle[ 1582] = 1'b0;  wr_cycle[ 1582] = 1'b1;  addr_rom[ 1582]='h000018b8;  wr_data_rom[ 1582]='h00000052;
    rd_cycle[ 1583] = 1'b0;  wr_cycle[ 1583] = 1'b1;  addr_rom[ 1583]='h000018bc;  wr_data_rom[ 1583]='h000016bb;
    rd_cycle[ 1584] = 1'b0;  wr_cycle[ 1584] = 1'b1;  addr_rom[ 1584]='h000018c0;  wr_data_rom[ 1584]='h00000824;
    rd_cycle[ 1585] = 1'b0;  wr_cycle[ 1585] = 1'b1;  addr_rom[ 1585]='h000018c4;  wr_data_rom[ 1585]='h00001272;
    rd_cycle[ 1586] = 1'b0;  wr_cycle[ 1586] = 1'b1;  addr_rom[ 1586]='h000018c8;  wr_data_rom[ 1586]='h00000315;
    rd_cycle[ 1587] = 1'b0;  wr_cycle[ 1587] = 1'b1;  addr_rom[ 1587]='h000018cc;  wr_data_rom[ 1587]='h00000ba7;
    rd_cycle[ 1588] = 1'b0;  wr_cycle[ 1588] = 1'b1;  addr_rom[ 1588]='h000018d0;  wr_data_rom[ 1588]='h0000130b;
    rd_cycle[ 1589] = 1'b0;  wr_cycle[ 1589] = 1'b1;  addr_rom[ 1589]='h000018d4;  wr_data_rom[ 1589]='h00000ca6;
    rd_cycle[ 1590] = 1'b0;  wr_cycle[ 1590] = 1'b1;  addr_rom[ 1590]='h000018d8;  wr_data_rom[ 1590]='h00000fb2;
    rd_cycle[ 1591] = 1'b0;  wr_cycle[ 1591] = 1'b1;  addr_rom[ 1591]='h000018dc;  wr_data_rom[ 1591]='h0000082c;
    rd_cycle[ 1592] = 1'b0;  wr_cycle[ 1592] = 1'b1;  addr_rom[ 1592]='h000018e0;  wr_data_rom[ 1592]='h00000d14;
    rd_cycle[ 1593] = 1'b0;  wr_cycle[ 1593] = 1'b1;  addr_rom[ 1593]='h000018e4;  wr_data_rom[ 1593]='h00000d8e;
    rd_cycle[ 1594] = 1'b0;  wr_cycle[ 1594] = 1'b1;  addr_rom[ 1594]='h000018e8;  wr_data_rom[ 1594]='h00001a85;
    rd_cycle[ 1595] = 1'b0;  wr_cycle[ 1595] = 1'b1;  addr_rom[ 1595]='h000018ec;  wr_data_rom[ 1595]='h000006ac;
    rd_cycle[ 1596] = 1'b0;  wr_cycle[ 1596] = 1'b1;  addr_rom[ 1596]='h000018f0;  wr_data_rom[ 1596]='h00001ee8;
    rd_cycle[ 1597] = 1'b0;  wr_cycle[ 1597] = 1'b1;  addr_rom[ 1597]='h000018f4;  wr_data_rom[ 1597]='h00001a67;
    rd_cycle[ 1598] = 1'b0;  wr_cycle[ 1598] = 1'b1;  addr_rom[ 1598]='h000018f8;  wr_data_rom[ 1598]='h000001c2;
    rd_cycle[ 1599] = 1'b0;  wr_cycle[ 1599] = 1'b1;  addr_rom[ 1599]='h000018fc;  wr_data_rom[ 1599]='h00000ba0;
    rd_cycle[ 1600] = 1'b0;  wr_cycle[ 1600] = 1'b1;  addr_rom[ 1600]='h00001900;  wr_data_rom[ 1600]='h000000c2;
    rd_cycle[ 1601] = 1'b0;  wr_cycle[ 1601] = 1'b1;  addr_rom[ 1601]='h00001904;  wr_data_rom[ 1601]='h00001745;
    rd_cycle[ 1602] = 1'b0;  wr_cycle[ 1602] = 1'b1;  addr_rom[ 1602]='h00001908;  wr_data_rom[ 1602]='h00000378;
    rd_cycle[ 1603] = 1'b0;  wr_cycle[ 1603] = 1'b1;  addr_rom[ 1603]='h0000190c;  wr_data_rom[ 1603]='h00001464;
    rd_cycle[ 1604] = 1'b0;  wr_cycle[ 1604] = 1'b1;  addr_rom[ 1604]='h00001910;  wr_data_rom[ 1604]='h0000099f;
    rd_cycle[ 1605] = 1'b0;  wr_cycle[ 1605] = 1'b1;  addr_rom[ 1605]='h00001914;  wr_data_rom[ 1605]='h00000d6c;
    rd_cycle[ 1606] = 1'b0;  wr_cycle[ 1606] = 1'b1;  addr_rom[ 1606]='h00001918;  wr_data_rom[ 1606]='h00000f0b;
    rd_cycle[ 1607] = 1'b0;  wr_cycle[ 1607] = 1'b1;  addr_rom[ 1607]='h0000191c;  wr_data_rom[ 1607]='h000007e9;
    rd_cycle[ 1608] = 1'b0;  wr_cycle[ 1608] = 1'b1;  addr_rom[ 1608]='h00001920;  wr_data_rom[ 1608]='h00001060;
    rd_cycle[ 1609] = 1'b0;  wr_cycle[ 1609] = 1'b1;  addr_rom[ 1609]='h00001924;  wr_data_rom[ 1609]='h000006d6;
    rd_cycle[ 1610] = 1'b0;  wr_cycle[ 1610] = 1'b1;  addr_rom[ 1610]='h00001928;  wr_data_rom[ 1610]='h00000d3d;
    rd_cycle[ 1611] = 1'b0;  wr_cycle[ 1611] = 1'b1;  addr_rom[ 1611]='h0000192c;  wr_data_rom[ 1611]='h000012ef;
    rd_cycle[ 1612] = 1'b0;  wr_cycle[ 1612] = 1'b1;  addr_rom[ 1612]='h00001930;  wr_data_rom[ 1612]='h00000114;
    rd_cycle[ 1613] = 1'b0;  wr_cycle[ 1613] = 1'b1;  addr_rom[ 1613]='h00001934;  wr_data_rom[ 1613]='h0000156a;
    rd_cycle[ 1614] = 1'b0;  wr_cycle[ 1614] = 1'b1;  addr_rom[ 1614]='h00001938;  wr_data_rom[ 1614]='h0000063e;
    rd_cycle[ 1615] = 1'b0;  wr_cycle[ 1615] = 1'b1;  addr_rom[ 1615]='h0000193c;  wr_data_rom[ 1615]='h000004e8;
    rd_cycle[ 1616] = 1'b0;  wr_cycle[ 1616] = 1'b1;  addr_rom[ 1616]='h00001940;  wr_data_rom[ 1616]='h000012b4;
    rd_cycle[ 1617] = 1'b0;  wr_cycle[ 1617] = 1'b1;  addr_rom[ 1617]='h00001944;  wr_data_rom[ 1617]='h000007db;
    rd_cycle[ 1618] = 1'b0;  wr_cycle[ 1618] = 1'b1;  addr_rom[ 1618]='h00001948;  wr_data_rom[ 1618]='h00000fd9;
    rd_cycle[ 1619] = 1'b0;  wr_cycle[ 1619] = 1'b1;  addr_rom[ 1619]='h0000194c;  wr_data_rom[ 1619]='h00000463;
    rd_cycle[ 1620] = 1'b0;  wr_cycle[ 1620] = 1'b1;  addr_rom[ 1620]='h00001950;  wr_data_rom[ 1620]='h000017f7;
    rd_cycle[ 1621] = 1'b0;  wr_cycle[ 1621] = 1'b1;  addr_rom[ 1621]='h00001954;  wr_data_rom[ 1621]='h000015db;
    rd_cycle[ 1622] = 1'b0;  wr_cycle[ 1622] = 1'b1;  addr_rom[ 1622]='h00001958;  wr_data_rom[ 1622]='h000007fe;
    rd_cycle[ 1623] = 1'b0;  wr_cycle[ 1623] = 1'b1;  addr_rom[ 1623]='h0000195c;  wr_data_rom[ 1623]='h00001b39;
    rd_cycle[ 1624] = 1'b0;  wr_cycle[ 1624] = 1'b1;  addr_rom[ 1624]='h00001960;  wr_data_rom[ 1624]='h00001e2e;
    rd_cycle[ 1625] = 1'b0;  wr_cycle[ 1625] = 1'b1;  addr_rom[ 1625]='h00001964;  wr_data_rom[ 1625]='h000003c2;
    rd_cycle[ 1626] = 1'b0;  wr_cycle[ 1626] = 1'b1;  addr_rom[ 1626]='h00001968;  wr_data_rom[ 1626]='h000008b0;
    rd_cycle[ 1627] = 1'b0;  wr_cycle[ 1627] = 1'b1;  addr_rom[ 1627]='h0000196c;  wr_data_rom[ 1627]='h0000197f;
    rd_cycle[ 1628] = 1'b0;  wr_cycle[ 1628] = 1'b1;  addr_rom[ 1628]='h00001970;  wr_data_rom[ 1628]='h00000436;
    rd_cycle[ 1629] = 1'b0;  wr_cycle[ 1629] = 1'b1;  addr_rom[ 1629]='h00001974;  wr_data_rom[ 1629]='h00001a7c;
    rd_cycle[ 1630] = 1'b0;  wr_cycle[ 1630] = 1'b1;  addr_rom[ 1630]='h00001978;  wr_data_rom[ 1630]='h000011a7;
    rd_cycle[ 1631] = 1'b0;  wr_cycle[ 1631] = 1'b1;  addr_rom[ 1631]='h0000197c;  wr_data_rom[ 1631]='h00000e4b;
    rd_cycle[ 1632] = 1'b0;  wr_cycle[ 1632] = 1'b1;  addr_rom[ 1632]='h00001980;  wr_data_rom[ 1632]='h00000a73;
    rd_cycle[ 1633] = 1'b0;  wr_cycle[ 1633] = 1'b1;  addr_rom[ 1633]='h00001984;  wr_data_rom[ 1633]='h000006e0;
    rd_cycle[ 1634] = 1'b0;  wr_cycle[ 1634] = 1'b1;  addr_rom[ 1634]='h00001988;  wr_data_rom[ 1634]='h000014d2;
    rd_cycle[ 1635] = 1'b0;  wr_cycle[ 1635] = 1'b1;  addr_rom[ 1635]='h0000198c;  wr_data_rom[ 1635]='h000016d4;
    rd_cycle[ 1636] = 1'b0;  wr_cycle[ 1636] = 1'b1;  addr_rom[ 1636]='h00001990;  wr_data_rom[ 1636]='h00000271;
    rd_cycle[ 1637] = 1'b0;  wr_cycle[ 1637] = 1'b1;  addr_rom[ 1637]='h00001994;  wr_data_rom[ 1637]='h00000d2e;
    rd_cycle[ 1638] = 1'b0;  wr_cycle[ 1638] = 1'b1;  addr_rom[ 1638]='h00001998;  wr_data_rom[ 1638]='h00000281;
    rd_cycle[ 1639] = 1'b0;  wr_cycle[ 1639] = 1'b1;  addr_rom[ 1639]='h0000199c;  wr_data_rom[ 1639]='h0000028b;
    rd_cycle[ 1640] = 1'b0;  wr_cycle[ 1640] = 1'b1;  addr_rom[ 1640]='h000019a0;  wr_data_rom[ 1640]='h000002e8;
    rd_cycle[ 1641] = 1'b0;  wr_cycle[ 1641] = 1'b1;  addr_rom[ 1641]='h000019a4;  wr_data_rom[ 1641]='h00001331;
    rd_cycle[ 1642] = 1'b0;  wr_cycle[ 1642] = 1'b1;  addr_rom[ 1642]='h000019a8;  wr_data_rom[ 1642]='h0000185f;
    rd_cycle[ 1643] = 1'b0;  wr_cycle[ 1643] = 1'b1;  addr_rom[ 1643]='h000019ac;  wr_data_rom[ 1643]='h0000178e;
    rd_cycle[ 1644] = 1'b0;  wr_cycle[ 1644] = 1'b1;  addr_rom[ 1644]='h000019b0;  wr_data_rom[ 1644]='h00000741;
    rd_cycle[ 1645] = 1'b0;  wr_cycle[ 1645] = 1'b1;  addr_rom[ 1645]='h000019b4;  wr_data_rom[ 1645]='h0000109b;
    rd_cycle[ 1646] = 1'b0;  wr_cycle[ 1646] = 1'b1;  addr_rom[ 1646]='h000019b8;  wr_data_rom[ 1646]='h00001908;
    rd_cycle[ 1647] = 1'b0;  wr_cycle[ 1647] = 1'b1;  addr_rom[ 1647]='h000019bc;  wr_data_rom[ 1647]='h000010b9;
    rd_cycle[ 1648] = 1'b0;  wr_cycle[ 1648] = 1'b1;  addr_rom[ 1648]='h000019c0;  wr_data_rom[ 1648]='h00001192;
    rd_cycle[ 1649] = 1'b0;  wr_cycle[ 1649] = 1'b1;  addr_rom[ 1649]='h000019c4;  wr_data_rom[ 1649]='h00000a94;
    rd_cycle[ 1650] = 1'b0;  wr_cycle[ 1650] = 1'b1;  addr_rom[ 1650]='h000019c8;  wr_data_rom[ 1650]='h0000041b;
    rd_cycle[ 1651] = 1'b0;  wr_cycle[ 1651] = 1'b1;  addr_rom[ 1651]='h000019cc;  wr_data_rom[ 1651]='h00001e36;
    rd_cycle[ 1652] = 1'b0;  wr_cycle[ 1652] = 1'b1;  addr_rom[ 1652]='h000019d0;  wr_data_rom[ 1652]='h00001e90;
    rd_cycle[ 1653] = 1'b0;  wr_cycle[ 1653] = 1'b1;  addr_rom[ 1653]='h000019d4;  wr_data_rom[ 1653]='h00001866;
    rd_cycle[ 1654] = 1'b0;  wr_cycle[ 1654] = 1'b1;  addr_rom[ 1654]='h000019d8;  wr_data_rom[ 1654]='h00000358;
    rd_cycle[ 1655] = 1'b0;  wr_cycle[ 1655] = 1'b1;  addr_rom[ 1655]='h000019dc;  wr_data_rom[ 1655]='h0000136b;
    rd_cycle[ 1656] = 1'b0;  wr_cycle[ 1656] = 1'b1;  addr_rom[ 1656]='h000019e0;  wr_data_rom[ 1656]='h0000132a;
    rd_cycle[ 1657] = 1'b0;  wr_cycle[ 1657] = 1'b1;  addr_rom[ 1657]='h000019e4;  wr_data_rom[ 1657]='h0000190e;
    rd_cycle[ 1658] = 1'b0;  wr_cycle[ 1658] = 1'b1;  addr_rom[ 1658]='h000019e8;  wr_data_rom[ 1658]='h00000bec;
    rd_cycle[ 1659] = 1'b0;  wr_cycle[ 1659] = 1'b1;  addr_rom[ 1659]='h000019ec;  wr_data_rom[ 1659]='h000018f3;
    rd_cycle[ 1660] = 1'b0;  wr_cycle[ 1660] = 1'b1;  addr_rom[ 1660]='h000019f0;  wr_data_rom[ 1660]='h00001094;
    rd_cycle[ 1661] = 1'b0;  wr_cycle[ 1661] = 1'b1;  addr_rom[ 1661]='h000019f4;  wr_data_rom[ 1661]='h00000691;
    rd_cycle[ 1662] = 1'b0;  wr_cycle[ 1662] = 1'b1;  addr_rom[ 1662]='h000019f8;  wr_data_rom[ 1662]='h00000c3f;
    rd_cycle[ 1663] = 1'b0;  wr_cycle[ 1663] = 1'b1;  addr_rom[ 1663]='h000019fc;  wr_data_rom[ 1663]='h00000013;
    rd_cycle[ 1664] = 1'b0;  wr_cycle[ 1664] = 1'b1;  addr_rom[ 1664]='h00001a00;  wr_data_rom[ 1664]='h00000c82;
    rd_cycle[ 1665] = 1'b0;  wr_cycle[ 1665] = 1'b1;  addr_rom[ 1665]='h00001a04;  wr_data_rom[ 1665]='h00001a07;
    rd_cycle[ 1666] = 1'b0;  wr_cycle[ 1666] = 1'b1;  addr_rom[ 1666]='h00001a08;  wr_data_rom[ 1666]='h000015b6;
    rd_cycle[ 1667] = 1'b0;  wr_cycle[ 1667] = 1'b1;  addr_rom[ 1667]='h00001a0c;  wr_data_rom[ 1667]='h00001edd;
    rd_cycle[ 1668] = 1'b0;  wr_cycle[ 1668] = 1'b1;  addr_rom[ 1668]='h00001a10;  wr_data_rom[ 1668]='h000015f0;
    rd_cycle[ 1669] = 1'b0;  wr_cycle[ 1669] = 1'b1;  addr_rom[ 1669]='h00001a14;  wr_data_rom[ 1669]='h000000be;
    rd_cycle[ 1670] = 1'b0;  wr_cycle[ 1670] = 1'b1;  addr_rom[ 1670]='h00001a18;  wr_data_rom[ 1670]='h00001f16;
    rd_cycle[ 1671] = 1'b0;  wr_cycle[ 1671] = 1'b1;  addr_rom[ 1671]='h00001a1c;  wr_data_rom[ 1671]='h000005f5;
    rd_cycle[ 1672] = 1'b0;  wr_cycle[ 1672] = 1'b1;  addr_rom[ 1672]='h00001a20;  wr_data_rom[ 1672]='h00000fc3;
    rd_cycle[ 1673] = 1'b0;  wr_cycle[ 1673] = 1'b1;  addr_rom[ 1673]='h00001a24;  wr_data_rom[ 1673]='h00000a3c;
    rd_cycle[ 1674] = 1'b0;  wr_cycle[ 1674] = 1'b1;  addr_rom[ 1674]='h00001a28;  wr_data_rom[ 1674]='h000006fc;
    rd_cycle[ 1675] = 1'b0;  wr_cycle[ 1675] = 1'b1;  addr_rom[ 1675]='h00001a2c;  wr_data_rom[ 1675]='h00000a27;
    rd_cycle[ 1676] = 1'b0;  wr_cycle[ 1676] = 1'b1;  addr_rom[ 1676]='h00001a30;  wr_data_rom[ 1676]='h00000644;
    rd_cycle[ 1677] = 1'b0;  wr_cycle[ 1677] = 1'b1;  addr_rom[ 1677]='h00001a34;  wr_data_rom[ 1677]='h00000f12;
    rd_cycle[ 1678] = 1'b0;  wr_cycle[ 1678] = 1'b1;  addr_rom[ 1678]='h00001a38;  wr_data_rom[ 1678]='h00000b48;
    rd_cycle[ 1679] = 1'b0;  wr_cycle[ 1679] = 1'b1;  addr_rom[ 1679]='h00001a3c;  wr_data_rom[ 1679]='h00000df8;
    rd_cycle[ 1680] = 1'b0;  wr_cycle[ 1680] = 1'b1;  addr_rom[ 1680]='h00001a40;  wr_data_rom[ 1680]='h00001eab;
    rd_cycle[ 1681] = 1'b0;  wr_cycle[ 1681] = 1'b1;  addr_rom[ 1681]='h00001a44;  wr_data_rom[ 1681]='h00000529;
    rd_cycle[ 1682] = 1'b0;  wr_cycle[ 1682] = 1'b1;  addr_rom[ 1682]='h00001a48;  wr_data_rom[ 1682]='h00001b57;
    rd_cycle[ 1683] = 1'b0;  wr_cycle[ 1683] = 1'b1;  addr_rom[ 1683]='h00001a4c;  wr_data_rom[ 1683]='h00001457;
    rd_cycle[ 1684] = 1'b0;  wr_cycle[ 1684] = 1'b1;  addr_rom[ 1684]='h00001a50;  wr_data_rom[ 1684]='h00001241;
    rd_cycle[ 1685] = 1'b0;  wr_cycle[ 1685] = 1'b1;  addr_rom[ 1685]='h00001a54;  wr_data_rom[ 1685]='h0000143f;
    rd_cycle[ 1686] = 1'b0;  wr_cycle[ 1686] = 1'b1;  addr_rom[ 1686]='h00001a58;  wr_data_rom[ 1686]='h000005dc;
    rd_cycle[ 1687] = 1'b0;  wr_cycle[ 1687] = 1'b1;  addr_rom[ 1687]='h00001a5c;  wr_data_rom[ 1687]='h000000e1;
    rd_cycle[ 1688] = 1'b0;  wr_cycle[ 1688] = 1'b1;  addr_rom[ 1688]='h00001a60;  wr_data_rom[ 1688]='h00000f6b;
    rd_cycle[ 1689] = 1'b0;  wr_cycle[ 1689] = 1'b1;  addr_rom[ 1689]='h00001a64;  wr_data_rom[ 1689]='h00001909;
    rd_cycle[ 1690] = 1'b0;  wr_cycle[ 1690] = 1'b1;  addr_rom[ 1690]='h00001a68;  wr_data_rom[ 1690]='h00001d32;
    rd_cycle[ 1691] = 1'b0;  wr_cycle[ 1691] = 1'b1;  addr_rom[ 1691]='h00001a6c;  wr_data_rom[ 1691]='h0000136d;
    rd_cycle[ 1692] = 1'b0;  wr_cycle[ 1692] = 1'b1;  addr_rom[ 1692]='h00001a70;  wr_data_rom[ 1692]='h000008e4;
    rd_cycle[ 1693] = 1'b0;  wr_cycle[ 1693] = 1'b1;  addr_rom[ 1693]='h00001a74;  wr_data_rom[ 1693]='h00001ca1;
    rd_cycle[ 1694] = 1'b0;  wr_cycle[ 1694] = 1'b1;  addr_rom[ 1694]='h00001a78;  wr_data_rom[ 1694]='h00000b93;
    rd_cycle[ 1695] = 1'b0;  wr_cycle[ 1695] = 1'b1;  addr_rom[ 1695]='h00001a7c;  wr_data_rom[ 1695]='h00001465;
    rd_cycle[ 1696] = 1'b0;  wr_cycle[ 1696] = 1'b1;  addr_rom[ 1696]='h00001a80;  wr_data_rom[ 1696]='h00000d83;
    rd_cycle[ 1697] = 1'b0;  wr_cycle[ 1697] = 1'b1;  addr_rom[ 1697]='h00001a84;  wr_data_rom[ 1697]='h000007ae;
    rd_cycle[ 1698] = 1'b0;  wr_cycle[ 1698] = 1'b1;  addr_rom[ 1698]='h00001a88;  wr_data_rom[ 1698]='h000004fd;
    rd_cycle[ 1699] = 1'b0;  wr_cycle[ 1699] = 1'b1;  addr_rom[ 1699]='h00001a8c;  wr_data_rom[ 1699]='h000002cd;
    rd_cycle[ 1700] = 1'b0;  wr_cycle[ 1700] = 1'b1;  addr_rom[ 1700]='h00001a90;  wr_data_rom[ 1700]='h00001323;
    rd_cycle[ 1701] = 1'b0;  wr_cycle[ 1701] = 1'b1;  addr_rom[ 1701]='h00001a94;  wr_data_rom[ 1701]='h000019d5;
    rd_cycle[ 1702] = 1'b0;  wr_cycle[ 1702] = 1'b1;  addr_rom[ 1702]='h00001a98;  wr_data_rom[ 1702]='h000003b2;
    rd_cycle[ 1703] = 1'b0;  wr_cycle[ 1703] = 1'b1;  addr_rom[ 1703]='h00001a9c;  wr_data_rom[ 1703]='h0000151d;
    rd_cycle[ 1704] = 1'b0;  wr_cycle[ 1704] = 1'b1;  addr_rom[ 1704]='h00001aa0;  wr_data_rom[ 1704]='h000015fd;
    rd_cycle[ 1705] = 1'b0;  wr_cycle[ 1705] = 1'b1;  addr_rom[ 1705]='h00001aa4;  wr_data_rom[ 1705]='h00001f05;
    rd_cycle[ 1706] = 1'b0;  wr_cycle[ 1706] = 1'b1;  addr_rom[ 1706]='h00001aa8;  wr_data_rom[ 1706]='h00000360;
    rd_cycle[ 1707] = 1'b0;  wr_cycle[ 1707] = 1'b1;  addr_rom[ 1707]='h00001aac;  wr_data_rom[ 1707]='h00000d4b;
    rd_cycle[ 1708] = 1'b0;  wr_cycle[ 1708] = 1'b1;  addr_rom[ 1708]='h00001ab0;  wr_data_rom[ 1708]='h00001d00;
    rd_cycle[ 1709] = 1'b0;  wr_cycle[ 1709] = 1'b1;  addr_rom[ 1709]='h00001ab4;  wr_data_rom[ 1709]='h0000088f;
    rd_cycle[ 1710] = 1'b0;  wr_cycle[ 1710] = 1'b1;  addr_rom[ 1710]='h00001ab8;  wr_data_rom[ 1710]='h00000dd3;
    rd_cycle[ 1711] = 1'b0;  wr_cycle[ 1711] = 1'b1;  addr_rom[ 1711]='h00001abc;  wr_data_rom[ 1711]='h00000456;
    rd_cycle[ 1712] = 1'b0;  wr_cycle[ 1712] = 1'b1;  addr_rom[ 1712]='h00001ac0;  wr_data_rom[ 1712]='h00001952;
    rd_cycle[ 1713] = 1'b0;  wr_cycle[ 1713] = 1'b1;  addr_rom[ 1713]='h00001ac4;  wr_data_rom[ 1713]='h0000123c;
    rd_cycle[ 1714] = 1'b0;  wr_cycle[ 1714] = 1'b1;  addr_rom[ 1714]='h00001ac8;  wr_data_rom[ 1714]='h00001cea;
    rd_cycle[ 1715] = 1'b0;  wr_cycle[ 1715] = 1'b1;  addr_rom[ 1715]='h00001acc;  wr_data_rom[ 1715]='h000015b2;
    rd_cycle[ 1716] = 1'b0;  wr_cycle[ 1716] = 1'b1;  addr_rom[ 1716]='h00001ad0;  wr_data_rom[ 1716]='h00001942;
    rd_cycle[ 1717] = 1'b0;  wr_cycle[ 1717] = 1'b1;  addr_rom[ 1717]='h00001ad4;  wr_data_rom[ 1717]='h00000b94;
    rd_cycle[ 1718] = 1'b0;  wr_cycle[ 1718] = 1'b1;  addr_rom[ 1718]='h00001ad8;  wr_data_rom[ 1718]='h0000061b;
    rd_cycle[ 1719] = 1'b0;  wr_cycle[ 1719] = 1'b1;  addr_rom[ 1719]='h00001adc;  wr_data_rom[ 1719]='h00001890;
    rd_cycle[ 1720] = 1'b0;  wr_cycle[ 1720] = 1'b1;  addr_rom[ 1720]='h00001ae0;  wr_data_rom[ 1720]='h00001806;
    rd_cycle[ 1721] = 1'b0;  wr_cycle[ 1721] = 1'b1;  addr_rom[ 1721]='h00001ae4;  wr_data_rom[ 1721]='h0000199d;
    rd_cycle[ 1722] = 1'b0;  wr_cycle[ 1722] = 1'b1;  addr_rom[ 1722]='h00001ae8;  wr_data_rom[ 1722]='h00001103;
    rd_cycle[ 1723] = 1'b0;  wr_cycle[ 1723] = 1'b1;  addr_rom[ 1723]='h00001aec;  wr_data_rom[ 1723]='h0000070a;
    rd_cycle[ 1724] = 1'b0;  wr_cycle[ 1724] = 1'b1;  addr_rom[ 1724]='h00001af0;  wr_data_rom[ 1724]='h000014c7;
    rd_cycle[ 1725] = 1'b0;  wr_cycle[ 1725] = 1'b1;  addr_rom[ 1725]='h00001af4;  wr_data_rom[ 1725]='h0000022a;
    rd_cycle[ 1726] = 1'b0;  wr_cycle[ 1726] = 1'b1;  addr_rom[ 1726]='h00001af8;  wr_data_rom[ 1726]='h00001ac3;
    rd_cycle[ 1727] = 1'b0;  wr_cycle[ 1727] = 1'b1;  addr_rom[ 1727]='h00001afc;  wr_data_rom[ 1727]='h00001a5b;
    rd_cycle[ 1728] = 1'b0;  wr_cycle[ 1728] = 1'b1;  addr_rom[ 1728]='h00001b00;  wr_data_rom[ 1728]='h000001c5;
    rd_cycle[ 1729] = 1'b0;  wr_cycle[ 1729] = 1'b1;  addr_rom[ 1729]='h00001b04;  wr_data_rom[ 1729]='h00001f05;
    rd_cycle[ 1730] = 1'b0;  wr_cycle[ 1730] = 1'b1;  addr_rom[ 1730]='h00001b08;  wr_data_rom[ 1730]='h00001856;
    rd_cycle[ 1731] = 1'b0;  wr_cycle[ 1731] = 1'b1;  addr_rom[ 1731]='h00001b0c;  wr_data_rom[ 1731]='h00001e22;
    rd_cycle[ 1732] = 1'b0;  wr_cycle[ 1732] = 1'b1;  addr_rom[ 1732]='h00001b10;  wr_data_rom[ 1732]='h0000020f;
    rd_cycle[ 1733] = 1'b0;  wr_cycle[ 1733] = 1'b1;  addr_rom[ 1733]='h00001b14;  wr_data_rom[ 1733]='h000015e5;
    rd_cycle[ 1734] = 1'b0;  wr_cycle[ 1734] = 1'b1;  addr_rom[ 1734]='h00001b18;  wr_data_rom[ 1734]='h00001660;
    rd_cycle[ 1735] = 1'b0;  wr_cycle[ 1735] = 1'b1;  addr_rom[ 1735]='h00001b1c;  wr_data_rom[ 1735]='h00000254;
    rd_cycle[ 1736] = 1'b0;  wr_cycle[ 1736] = 1'b1;  addr_rom[ 1736]='h00001b20;  wr_data_rom[ 1736]='h000013ee;
    rd_cycle[ 1737] = 1'b0;  wr_cycle[ 1737] = 1'b1;  addr_rom[ 1737]='h00001b24;  wr_data_rom[ 1737]='h0000001a;
    rd_cycle[ 1738] = 1'b0;  wr_cycle[ 1738] = 1'b1;  addr_rom[ 1738]='h00001b28;  wr_data_rom[ 1738]='h00001e96;
    rd_cycle[ 1739] = 1'b0;  wr_cycle[ 1739] = 1'b1;  addr_rom[ 1739]='h00001b2c;  wr_data_rom[ 1739]='h000013c2;
    rd_cycle[ 1740] = 1'b0;  wr_cycle[ 1740] = 1'b1;  addr_rom[ 1740]='h00001b30;  wr_data_rom[ 1740]='h00001ae2;
    rd_cycle[ 1741] = 1'b0;  wr_cycle[ 1741] = 1'b1;  addr_rom[ 1741]='h00001b34;  wr_data_rom[ 1741]='h000008b2;
    rd_cycle[ 1742] = 1'b0;  wr_cycle[ 1742] = 1'b1;  addr_rom[ 1742]='h00001b38;  wr_data_rom[ 1742]='h0000049d;
    rd_cycle[ 1743] = 1'b0;  wr_cycle[ 1743] = 1'b1;  addr_rom[ 1743]='h00001b3c;  wr_data_rom[ 1743]='h00001ed0;
    rd_cycle[ 1744] = 1'b0;  wr_cycle[ 1744] = 1'b1;  addr_rom[ 1744]='h00001b40;  wr_data_rom[ 1744]='h000009c1;
    rd_cycle[ 1745] = 1'b0;  wr_cycle[ 1745] = 1'b1;  addr_rom[ 1745]='h00001b44;  wr_data_rom[ 1745]='h00001c10;
    rd_cycle[ 1746] = 1'b0;  wr_cycle[ 1746] = 1'b1;  addr_rom[ 1746]='h00001b48;  wr_data_rom[ 1746]='h0000060b;
    rd_cycle[ 1747] = 1'b0;  wr_cycle[ 1747] = 1'b1;  addr_rom[ 1747]='h00001b4c;  wr_data_rom[ 1747]='h000013cd;
    rd_cycle[ 1748] = 1'b0;  wr_cycle[ 1748] = 1'b1;  addr_rom[ 1748]='h00001b50;  wr_data_rom[ 1748]='h0000052f;
    rd_cycle[ 1749] = 1'b0;  wr_cycle[ 1749] = 1'b1;  addr_rom[ 1749]='h00001b54;  wr_data_rom[ 1749]='h000011cc;
    rd_cycle[ 1750] = 1'b0;  wr_cycle[ 1750] = 1'b1;  addr_rom[ 1750]='h00001b58;  wr_data_rom[ 1750]='h000017b1;
    rd_cycle[ 1751] = 1'b0;  wr_cycle[ 1751] = 1'b1;  addr_rom[ 1751]='h00001b5c;  wr_data_rom[ 1751]='h0000154d;
    rd_cycle[ 1752] = 1'b0;  wr_cycle[ 1752] = 1'b1;  addr_rom[ 1752]='h00001b60;  wr_data_rom[ 1752]='h00001199;
    rd_cycle[ 1753] = 1'b0;  wr_cycle[ 1753] = 1'b1;  addr_rom[ 1753]='h00001b64;  wr_data_rom[ 1753]='h00000e79;
    rd_cycle[ 1754] = 1'b0;  wr_cycle[ 1754] = 1'b1;  addr_rom[ 1754]='h00001b68;  wr_data_rom[ 1754]='h000000e0;
    rd_cycle[ 1755] = 1'b0;  wr_cycle[ 1755] = 1'b1;  addr_rom[ 1755]='h00001b6c;  wr_data_rom[ 1755]='h00000c43;
    rd_cycle[ 1756] = 1'b0;  wr_cycle[ 1756] = 1'b1;  addr_rom[ 1756]='h00001b70;  wr_data_rom[ 1756]='h00001234;
    rd_cycle[ 1757] = 1'b0;  wr_cycle[ 1757] = 1'b1;  addr_rom[ 1757]='h00001b74;  wr_data_rom[ 1757]='h000008aa;
    rd_cycle[ 1758] = 1'b0;  wr_cycle[ 1758] = 1'b1;  addr_rom[ 1758]='h00001b78;  wr_data_rom[ 1758]='h00000eab;
    rd_cycle[ 1759] = 1'b0;  wr_cycle[ 1759] = 1'b1;  addr_rom[ 1759]='h00001b7c;  wr_data_rom[ 1759]='h000012d6;
    rd_cycle[ 1760] = 1'b0;  wr_cycle[ 1760] = 1'b1;  addr_rom[ 1760]='h00001b80;  wr_data_rom[ 1760]='h00001054;
    rd_cycle[ 1761] = 1'b0;  wr_cycle[ 1761] = 1'b1;  addr_rom[ 1761]='h00001b84;  wr_data_rom[ 1761]='h00001c22;
    rd_cycle[ 1762] = 1'b0;  wr_cycle[ 1762] = 1'b1;  addr_rom[ 1762]='h00001b88;  wr_data_rom[ 1762]='h00000855;
    rd_cycle[ 1763] = 1'b0;  wr_cycle[ 1763] = 1'b1;  addr_rom[ 1763]='h00001b8c;  wr_data_rom[ 1763]='h0000105e;
    rd_cycle[ 1764] = 1'b0;  wr_cycle[ 1764] = 1'b1;  addr_rom[ 1764]='h00001b90;  wr_data_rom[ 1764]='h00000267;
    rd_cycle[ 1765] = 1'b0;  wr_cycle[ 1765] = 1'b1;  addr_rom[ 1765]='h00001b94;  wr_data_rom[ 1765]='h0000010b;
    rd_cycle[ 1766] = 1'b0;  wr_cycle[ 1766] = 1'b1;  addr_rom[ 1766]='h00001b98;  wr_data_rom[ 1766]='h0000127d;
    rd_cycle[ 1767] = 1'b0;  wr_cycle[ 1767] = 1'b1;  addr_rom[ 1767]='h00001b9c;  wr_data_rom[ 1767]='h00001b15;
    rd_cycle[ 1768] = 1'b0;  wr_cycle[ 1768] = 1'b1;  addr_rom[ 1768]='h00001ba0;  wr_data_rom[ 1768]='h00000848;
    rd_cycle[ 1769] = 1'b0;  wr_cycle[ 1769] = 1'b1;  addr_rom[ 1769]='h00001ba4;  wr_data_rom[ 1769]='h00000e8b;
    rd_cycle[ 1770] = 1'b0;  wr_cycle[ 1770] = 1'b1;  addr_rom[ 1770]='h00001ba8;  wr_data_rom[ 1770]='h00000e3e;
    rd_cycle[ 1771] = 1'b0;  wr_cycle[ 1771] = 1'b1;  addr_rom[ 1771]='h00001bac;  wr_data_rom[ 1771]='h00000ada;
    rd_cycle[ 1772] = 1'b0;  wr_cycle[ 1772] = 1'b1;  addr_rom[ 1772]='h00001bb0;  wr_data_rom[ 1772]='h000006f3;
    rd_cycle[ 1773] = 1'b0;  wr_cycle[ 1773] = 1'b1;  addr_rom[ 1773]='h00001bb4;  wr_data_rom[ 1773]='h00000010;
    rd_cycle[ 1774] = 1'b0;  wr_cycle[ 1774] = 1'b1;  addr_rom[ 1774]='h00001bb8;  wr_data_rom[ 1774]='h000012dd;
    rd_cycle[ 1775] = 1'b0;  wr_cycle[ 1775] = 1'b1;  addr_rom[ 1775]='h00001bbc;  wr_data_rom[ 1775]='h00000a8b;
    rd_cycle[ 1776] = 1'b0;  wr_cycle[ 1776] = 1'b1;  addr_rom[ 1776]='h00001bc0;  wr_data_rom[ 1776]='h00001193;
    rd_cycle[ 1777] = 1'b0;  wr_cycle[ 1777] = 1'b1;  addr_rom[ 1777]='h00001bc4;  wr_data_rom[ 1777]='h00001ea7;
    rd_cycle[ 1778] = 1'b0;  wr_cycle[ 1778] = 1'b1;  addr_rom[ 1778]='h00001bc8;  wr_data_rom[ 1778]='h0000023e;
    rd_cycle[ 1779] = 1'b0;  wr_cycle[ 1779] = 1'b1;  addr_rom[ 1779]='h00001bcc;  wr_data_rom[ 1779]='h00000e45;
    rd_cycle[ 1780] = 1'b0;  wr_cycle[ 1780] = 1'b1;  addr_rom[ 1780]='h00001bd0;  wr_data_rom[ 1780]='h00001468;
    rd_cycle[ 1781] = 1'b0;  wr_cycle[ 1781] = 1'b1;  addr_rom[ 1781]='h00001bd4;  wr_data_rom[ 1781]='h00001b92;
    rd_cycle[ 1782] = 1'b0;  wr_cycle[ 1782] = 1'b1;  addr_rom[ 1782]='h00001bd8;  wr_data_rom[ 1782]='h00001dac;
    rd_cycle[ 1783] = 1'b0;  wr_cycle[ 1783] = 1'b1;  addr_rom[ 1783]='h00001bdc;  wr_data_rom[ 1783]='h00000bfb;
    rd_cycle[ 1784] = 1'b0;  wr_cycle[ 1784] = 1'b1;  addr_rom[ 1784]='h00001be0;  wr_data_rom[ 1784]='h000013e7;
    rd_cycle[ 1785] = 1'b0;  wr_cycle[ 1785] = 1'b1;  addr_rom[ 1785]='h00001be4;  wr_data_rom[ 1785]='h000015ac;
    rd_cycle[ 1786] = 1'b0;  wr_cycle[ 1786] = 1'b1;  addr_rom[ 1786]='h00001be8;  wr_data_rom[ 1786]='h0000177b;
    rd_cycle[ 1787] = 1'b0;  wr_cycle[ 1787] = 1'b1;  addr_rom[ 1787]='h00001bec;  wr_data_rom[ 1787]='h00000398;
    rd_cycle[ 1788] = 1'b0;  wr_cycle[ 1788] = 1'b1;  addr_rom[ 1788]='h00001bf0;  wr_data_rom[ 1788]='h00001007;
    rd_cycle[ 1789] = 1'b0;  wr_cycle[ 1789] = 1'b1;  addr_rom[ 1789]='h00001bf4;  wr_data_rom[ 1789]='h00001338;
    rd_cycle[ 1790] = 1'b0;  wr_cycle[ 1790] = 1'b1;  addr_rom[ 1790]='h00001bf8;  wr_data_rom[ 1790]='h00001265;
    rd_cycle[ 1791] = 1'b0;  wr_cycle[ 1791] = 1'b1;  addr_rom[ 1791]='h00001bfc;  wr_data_rom[ 1791]='h000011d2;
    rd_cycle[ 1792] = 1'b0;  wr_cycle[ 1792] = 1'b1;  addr_rom[ 1792]='h00001c00;  wr_data_rom[ 1792]='h00000c24;
    rd_cycle[ 1793] = 1'b0;  wr_cycle[ 1793] = 1'b1;  addr_rom[ 1793]='h00001c04;  wr_data_rom[ 1793]='h000009da;
    rd_cycle[ 1794] = 1'b0;  wr_cycle[ 1794] = 1'b1;  addr_rom[ 1794]='h00001c08;  wr_data_rom[ 1794]='h00001576;
    rd_cycle[ 1795] = 1'b0;  wr_cycle[ 1795] = 1'b1;  addr_rom[ 1795]='h00001c0c;  wr_data_rom[ 1795]='h00000d75;
    rd_cycle[ 1796] = 1'b0;  wr_cycle[ 1796] = 1'b1;  addr_rom[ 1796]='h00001c10;  wr_data_rom[ 1796]='h00000cb6;
    rd_cycle[ 1797] = 1'b0;  wr_cycle[ 1797] = 1'b1;  addr_rom[ 1797]='h00001c14;  wr_data_rom[ 1797]='h000004e4;
    rd_cycle[ 1798] = 1'b0;  wr_cycle[ 1798] = 1'b1;  addr_rom[ 1798]='h00001c18;  wr_data_rom[ 1798]='h00001a19;
    rd_cycle[ 1799] = 1'b0;  wr_cycle[ 1799] = 1'b1;  addr_rom[ 1799]='h00001c1c;  wr_data_rom[ 1799]='h00001b17;
    rd_cycle[ 1800] = 1'b0;  wr_cycle[ 1800] = 1'b1;  addr_rom[ 1800]='h00001c20;  wr_data_rom[ 1800]='h00001716;
    rd_cycle[ 1801] = 1'b0;  wr_cycle[ 1801] = 1'b1;  addr_rom[ 1801]='h00001c24;  wr_data_rom[ 1801]='h00001610;
    rd_cycle[ 1802] = 1'b0;  wr_cycle[ 1802] = 1'b1;  addr_rom[ 1802]='h00001c28;  wr_data_rom[ 1802]='h00000cc0;
    rd_cycle[ 1803] = 1'b0;  wr_cycle[ 1803] = 1'b1;  addr_rom[ 1803]='h00001c2c;  wr_data_rom[ 1803]='h0000155d;
    rd_cycle[ 1804] = 1'b0;  wr_cycle[ 1804] = 1'b1;  addr_rom[ 1804]='h00001c30;  wr_data_rom[ 1804]='h000001cc;
    rd_cycle[ 1805] = 1'b0;  wr_cycle[ 1805] = 1'b1;  addr_rom[ 1805]='h00001c34;  wr_data_rom[ 1805]='h0000025e;
    rd_cycle[ 1806] = 1'b0;  wr_cycle[ 1806] = 1'b1;  addr_rom[ 1806]='h00001c38;  wr_data_rom[ 1806]='h0000002c;
    rd_cycle[ 1807] = 1'b0;  wr_cycle[ 1807] = 1'b1;  addr_rom[ 1807]='h00001c3c;  wr_data_rom[ 1807]='h0000191a;
    rd_cycle[ 1808] = 1'b0;  wr_cycle[ 1808] = 1'b1;  addr_rom[ 1808]='h00001c40;  wr_data_rom[ 1808]='h0000095d;
    rd_cycle[ 1809] = 1'b0;  wr_cycle[ 1809] = 1'b1;  addr_rom[ 1809]='h00001c44;  wr_data_rom[ 1809]='h00001caa;
    rd_cycle[ 1810] = 1'b0;  wr_cycle[ 1810] = 1'b1;  addr_rom[ 1810]='h00001c48;  wr_data_rom[ 1810]='h0000072d;
    rd_cycle[ 1811] = 1'b0;  wr_cycle[ 1811] = 1'b1;  addr_rom[ 1811]='h00001c4c;  wr_data_rom[ 1811]='h0000150a;
    rd_cycle[ 1812] = 1'b0;  wr_cycle[ 1812] = 1'b1;  addr_rom[ 1812]='h00001c50;  wr_data_rom[ 1812]='h0000175d;
    rd_cycle[ 1813] = 1'b0;  wr_cycle[ 1813] = 1'b1;  addr_rom[ 1813]='h00001c54;  wr_data_rom[ 1813]='h000001f5;
    rd_cycle[ 1814] = 1'b0;  wr_cycle[ 1814] = 1'b1;  addr_rom[ 1814]='h00001c58;  wr_data_rom[ 1814]='h00000a51;
    rd_cycle[ 1815] = 1'b0;  wr_cycle[ 1815] = 1'b1;  addr_rom[ 1815]='h00001c5c;  wr_data_rom[ 1815]='h00000946;
    rd_cycle[ 1816] = 1'b0;  wr_cycle[ 1816] = 1'b1;  addr_rom[ 1816]='h00001c60;  wr_data_rom[ 1816]='h00001807;
    rd_cycle[ 1817] = 1'b0;  wr_cycle[ 1817] = 1'b1;  addr_rom[ 1817]='h00001c64;  wr_data_rom[ 1817]='h00001e60;
    rd_cycle[ 1818] = 1'b0;  wr_cycle[ 1818] = 1'b1;  addr_rom[ 1818]='h00001c68;  wr_data_rom[ 1818]='h00000452;
    rd_cycle[ 1819] = 1'b0;  wr_cycle[ 1819] = 1'b1;  addr_rom[ 1819]='h00001c6c;  wr_data_rom[ 1819]='h00001ec8;
    rd_cycle[ 1820] = 1'b0;  wr_cycle[ 1820] = 1'b1;  addr_rom[ 1820]='h00001c70;  wr_data_rom[ 1820]='h000015e8;
    rd_cycle[ 1821] = 1'b0;  wr_cycle[ 1821] = 1'b1;  addr_rom[ 1821]='h00001c74;  wr_data_rom[ 1821]='h000000fb;
    rd_cycle[ 1822] = 1'b0;  wr_cycle[ 1822] = 1'b1;  addr_rom[ 1822]='h00001c78;  wr_data_rom[ 1822]='h000005e9;
    rd_cycle[ 1823] = 1'b0;  wr_cycle[ 1823] = 1'b1;  addr_rom[ 1823]='h00001c7c;  wr_data_rom[ 1823]='h000008ed;
    rd_cycle[ 1824] = 1'b0;  wr_cycle[ 1824] = 1'b1;  addr_rom[ 1824]='h00001c80;  wr_data_rom[ 1824]='h00001539;
    rd_cycle[ 1825] = 1'b0;  wr_cycle[ 1825] = 1'b1;  addr_rom[ 1825]='h00001c84;  wr_data_rom[ 1825]='h00001bf3;
    rd_cycle[ 1826] = 1'b0;  wr_cycle[ 1826] = 1'b1;  addr_rom[ 1826]='h00001c88;  wr_data_rom[ 1826]='h00000a43;
    rd_cycle[ 1827] = 1'b0;  wr_cycle[ 1827] = 1'b1;  addr_rom[ 1827]='h00001c8c;  wr_data_rom[ 1827]='h0000001a;
    rd_cycle[ 1828] = 1'b0;  wr_cycle[ 1828] = 1'b1;  addr_rom[ 1828]='h00001c90;  wr_data_rom[ 1828]='h00001d48;
    rd_cycle[ 1829] = 1'b0;  wr_cycle[ 1829] = 1'b1;  addr_rom[ 1829]='h00001c94;  wr_data_rom[ 1829]='h000004b3;
    rd_cycle[ 1830] = 1'b0;  wr_cycle[ 1830] = 1'b1;  addr_rom[ 1830]='h00001c98;  wr_data_rom[ 1830]='h0000101e;
    rd_cycle[ 1831] = 1'b0;  wr_cycle[ 1831] = 1'b1;  addr_rom[ 1831]='h00001c9c;  wr_data_rom[ 1831]='h000005dc;
    rd_cycle[ 1832] = 1'b0;  wr_cycle[ 1832] = 1'b1;  addr_rom[ 1832]='h00001ca0;  wr_data_rom[ 1832]='h000009e0;
    rd_cycle[ 1833] = 1'b0;  wr_cycle[ 1833] = 1'b1;  addr_rom[ 1833]='h00001ca4;  wr_data_rom[ 1833]='h00000eb9;
    rd_cycle[ 1834] = 1'b0;  wr_cycle[ 1834] = 1'b1;  addr_rom[ 1834]='h00001ca8;  wr_data_rom[ 1834]='h000018d1;
    rd_cycle[ 1835] = 1'b0;  wr_cycle[ 1835] = 1'b1;  addr_rom[ 1835]='h00001cac;  wr_data_rom[ 1835]='h00001d27;
    rd_cycle[ 1836] = 1'b0;  wr_cycle[ 1836] = 1'b1;  addr_rom[ 1836]='h00001cb0;  wr_data_rom[ 1836]='h00000e15;
    rd_cycle[ 1837] = 1'b0;  wr_cycle[ 1837] = 1'b1;  addr_rom[ 1837]='h00001cb4;  wr_data_rom[ 1837]='h00001664;
    rd_cycle[ 1838] = 1'b0;  wr_cycle[ 1838] = 1'b1;  addr_rom[ 1838]='h00001cb8;  wr_data_rom[ 1838]='h00000584;
    rd_cycle[ 1839] = 1'b0;  wr_cycle[ 1839] = 1'b1;  addr_rom[ 1839]='h00001cbc;  wr_data_rom[ 1839]='h00000cdb;
    rd_cycle[ 1840] = 1'b0;  wr_cycle[ 1840] = 1'b1;  addr_rom[ 1840]='h00001cc0;  wr_data_rom[ 1840]='h00000905;
    rd_cycle[ 1841] = 1'b0;  wr_cycle[ 1841] = 1'b1;  addr_rom[ 1841]='h00001cc4;  wr_data_rom[ 1841]='h00000e19;
    rd_cycle[ 1842] = 1'b0;  wr_cycle[ 1842] = 1'b1;  addr_rom[ 1842]='h00001cc8;  wr_data_rom[ 1842]='h0000030e;
    rd_cycle[ 1843] = 1'b0;  wr_cycle[ 1843] = 1'b1;  addr_rom[ 1843]='h00001ccc;  wr_data_rom[ 1843]='h00001ac7;
    rd_cycle[ 1844] = 1'b0;  wr_cycle[ 1844] = 1'b1;  addr_rom[ 1844]='h00001cd0;  wr_data_rom[ 1844]='h000018eb;
    rd_cycle[ 1845] = 1'b0;  wr_cycle[ 1845] = 1'b1;  addr_rom[ 1845]='h00001cd4;  wr_data_rom[ 1845]='h00000d9f;
    rd_cycle[ 1846] = 1'b0;  wr_cycle[ 1846] = 1'b1;  addr_rom[ 1846]='h00001cd8;  wr_data_rom[ 1846]='h00000876;
    rd_cycle[ 1847] = 1'b0;  wr_cycle[ 1847] = 1'b1;  addr_rom[ 1847]='h00001cdc;  wr_data_rom[ 1847]='h00001c5b;
    rd_cycle[ 1848] = 1'b0;  wr_cycle[ 1848] = 1'b1;  addr_rom[ 1848]='h00001ce0;  wr_data_rom[ 1848]='h000000f7;
    rd_cycle[ 1849] = 1'b0;  wr_cycle[ 1849] = 1'b1;  addr_rom[ 1849]='h00001ce4;  wr_data_rom[ 1849]='h00001c1b;
    rd_cycle[ 1850] = 1'b0;  wr_cycle[ 1850] = 1'b1;  addr_rom[ 1850]='h00001ce8;  wr_data_rom[ 1850]='h00001f02;
    rd_cycle[ 1851] = 1'b0;  wr_cycle[ 1851] = 1'b1;  addr_rom[ 1851]='h00001cec;  wr_data_rom[ 1851]='h00001e45;
    rd_cycle[ 1852] = 1'b0;  wr_cycle[ 1852] = 1'b1;  addr_rom[ 1852]='h00001cf0;  wr_data_rom[ 1852]='h00001da2;
    rd_cycle[ 1853] = 1'b0;  wr_cycle[ 1853] = 1'b1;  addr_rom[ 1853]='h00001cf4;  wr_data_rom[ 1853]='h0000153f;
    rd_cycle[ 1854] = 1'b0;  wr_cycle[ 1854] = 1'b1;  addr_rom[ 1854]='h00001cf8;  wr_data_rom[ 1854]='h00000ab4;
    rd_cycle[ 1855] = 1'b0;  wr_cycle[ 1855] = 1'b1;  addr_rom[ 1855]='h00001cfc;  wr_data_rom[ 1855]='h000001b3;
    rd_cycle[ 1856] = 1'b0;  wr_cycle[ 1856] = 1'b1;  addr_rom[ 1856]='h00001d00;  wr_data_rom[ 1856]='h000004b5;
    rd_cycle[ 1857] = 1'b0;  wr_cycle[ 1857] = 1'b1;  addr_rom[ 1857]='h00001d04;  wr_data_rom[ 1857]='h00000a46;
    rd_cycle[ 1858] = 1'b0;  wr_cycle[ 1858] = 1'b1;  addr_rom[ 1858]='h00001d08;  wr_data_rom[ 1858]='h00001adc;
    rd_cycle[ 1859] = 1'b0;  wr_cycle[ 1859] = 1'b1;  addr_rom[ 1859]='h00001d0c;  wr_data_rom[ 1859]='h00001878;
    rd_cycle[ 1860] = 1'b0;  wr_cycle[ 1860] = 1'b1;  addr_rom[ 1860]='h00001d10;  wr_data_rom[ 1860]='h00001b2e;
    rd_cycle[ 1861] = 1'b0;  wr_cycle[ 1861] = 1'b1;  addr_rom[ 1861]='h00001d14;  wr_data_rom[ 1861]='h00001335;
    rd_cycle[ 1862] = 1'b0;  wr_cycle[ 1862] = 1'b1;  addr_rom[ 1862]='h00001d18;  wr_data_rom[ 1862]='h00001a6d;
    rd_cycle[ 1863] = 1'b0;  wr_cycle[ 1863] = 1'b1;  addr_rom[ 1863]='h00001d1c;  wr_data_rom[ 1863]='h00001944;
    rd_cycle[ 1864] = 1'b0;  wr_cycle[ 1864] = 1'b1;  addr_rom[ 1864]='h00001d20;  wr_data_rom[ 1864]='h000014da;
    rd_cycle[ 1865] = 1'b0;  wr_cycle[ 1865] = 1'b1;  addr_rom[ 1865]='h00001d24;  wr_data_rom[ 1865]='h00001350;
    rd_cycle[ 1866] = 1'b0;  wr_cycle[ 1866] = 1'b1;  addr_rom[ 1866]='h00001d28;  wr_data_rom[ 1866]='h0000048c;
    rd_cycle[ 1867] = 1'b0;  wr_cycle[ 1867] = 1'b1;  addr_rom[ 1867]='h00001d2c;  wr_data_rom[ 1867]='h00000968;
    rd_cycle[ 1868] = 1'b0;  wr_cycle[ 1868] = 1'b1;  addr_rom[ 1868]='h00001d30;  wr_data_rom[ 1868]='h00000d54;
    rd_cycle[ 1869] = 1'b0;  wr_cycle[ 1869] = 1'b1;  addr_rom[ 1869]='h00001d34;  wr_data_rom[ 1869]='h00000671;
    rd_cycle[ 1870] = 1'b0;  wr_cycle[ 1870] = 1'b1;  addr_rom[ 1870]='h00001d38;  wr_data_rom[ 1870]='h000004b0;
    rd_cycle[ 1871] = 1'b0;  wr_cycle[ 1871] = 1'b1;  addr_rom[ 1871]='h00001d3c;  wr_data_rom[ 1871]='h00000dfc;
    rd_cycle[ 1872] = 1'b0;  wr_cycle[ 1872] = 1'b1;  addr_rom[ 1872]='h00001d40;  wr_data_rom[ 1872]='h00000e9f;
    rd_cycle[ 1873] = 1'b0;  wr_cycle[ 1873] = 1'b1;  addr_rom[ 1873]='h00001d44;  wr_data_rom[ 1873]='h0000103f;
    rd_cycle[ 1874] = 1'b0;  wr_cycle[ 1874] = 1'b1;  addr_rom[ 1874]='h00001d48;  wr_data_rom[ 1874]='h0000178f;
    rd_cycle[ 1875] = 1'b0;  wr_cycle[ 1875] = 1'b1;  addr_rom[ 1875]='h00001d4c;  wr_data_rom[ 1875]='h000012a2;
    rd_cycle[ 1876] = 1'b0;  wr_cycle[ 1876] = 1'b1;  addr_rom[ 1876]='h00001d50;  wr_data_rom[ 1876]='h000006af;
    rd_cycle[ 1877] = 1'b0;  wr_cycle[ 1877] = 1'b1;  addr_rom[ 1877]='h00001d54;  wr_data_rom[ 1877]='h0000048b;
    rd_cycle[ 1878] = 1'b0;  wr_cycle[ 1878] = 1'b1;  addr_rom[ 1878]='h00001d58;  wr_data_rom[ 1878]='h00001690;
    rd_cycle[ 1879] = 1'b0;  wr_cycle[ 1879] = 1'b1;  addr_rom[ 1879]='h00001d5c;  wr_data_rom[ 1879]='h000015c4;
    rd_cycle[ 1880] = 1'b0;  wr_cycle[ 1880] = 1'b1;  addr_rom[ 1880]='h00001d60;  wr_data_rom[ 1880]='h0000037c;
    rd_cycle[ 1881] = 1'b0;  wr_cycle[ 1881] = 1'b1;  addr_rom[ 1881]='h00001d64;  wr_data_rom[ 1881]='h0000057e;
    rd_cycle[ 1882] = 1'b0;  wr_cycle[ 1882] = 1'b1;  addr_rom[ 1882]='h00001d68;  wr_data_rom[ 1882]='h00000950;
    rd_cycle[ 1883] = 1'b0;  wr_cycle[ 1883] = 1'b1;  addr_rom[ 1883]='h00001d6c;  wr_data_rom[ 1883]='h00000334;
    rd_cycle[ 1884] = 1'b0;  wr_cycle[ 1884] = 1'b1;  addr_rom[ 1884]='h00001d70;  wr_data_rom[ 1884]='h000004a9;
    rd_cycle[ 1885] = 1'b0;  wr_cycle[ 1885] = 1'b1;  addr_rom[ 1885]='h00001d74;  wr_data_rom[ 1885]='h00000ba1;
    rd_cycle[ 1886] = 1'b0;  wr_cycle[ 1886] = 1'b1;  addr_rom[ 1886]='h00001d78;  wr_data_rom[ 1886]='h00001b40;
    rd_cycle[ 1887] = 1'b0;  wr_cycle[ 1887] = 1'b1;  addr_rom[ 1887]='h00001d7c;  wr_data_rom[ 1887]='h00000397;
    rd_cycle[ 1888] = 1'b0;  wr_cycle[ 1888] = 1'b1;  addr_rom[ 1888]='h00001d80;  wr_data_rom[ 1888]='h000016ff;
    rd_cycle[ 1889] = 1'b0;  wr_cycle[ 1889] = 1'b1;  addr_rom[ 1889]='h00001d84;  wr_data_rom[ 1889]='h00000d96;
    rd_cycle[ 1890] = 1'b0;  wr_cycle[ 1890] = 1'b1;  addr_rom[ 1890]='h00001d88;  wr_data_rom[ 1890]='h00000917;
    rd_cycle[ 1891] = 1'b0;  wr_cycle[ 1891] = 1'b1;  addr_rom[ 1891]='h00001d8c;  wr_data_rom[ 1891]='h00001e75;
    rd_cycle[ 1892] = 1'b0;  wr_cycle[ 1892] = 1'b1;  addr_rom[ 1892]='h00001d90;  wr_data_rom[ 1892]='h0000134c;
    rd_cycle[ 1893] = 1'b0;  wr_cycle[ 1893] = 1'b1;  addr_rom[ 1893]='h00001d94;  wr_data_rom[ 1893]='h000008b7;
    rd_cycle[ 1894] = 1'b0;  wr_cycle[ 1894] = 1'b1;  addr_rom[ 1894]='h00001d98;  wr_data_rom[ 1894]='h00000498;
    rd_cycle[ 1895] = 1'b0;  wr_cycle[ 1895] = 1'b1;  addr_rom[ 1895]='h00001d9c;  wr_data_rom[ 1895]='h0000069b;
    rd_cycle[ 1896] = 1'b0;  wr_cycle[ 1896] = 1'b1;  addr_rom[ 1896]='h00001da0;  wr_data_rom[ 1896]='h00001c05;
    rd_cycle[ 1897] = 1'b0;  wr_cycle[ 1897] = 1'b1;  addr_rom[ 1897]='h00001da4;  wr_data_rom[ 1897]='h000002ce;
    rd_cycle[ 1898] = 1'b0;  wr_cycle[ 1898] = 1'b1;  addr_rom[ 1898]='h00001da8;  wr_data_rom[ 1898]='h00001172;
    rd_cycle[ 1899] = 1'b0;  wr_cycle[ 1899] = 1'b1;  addr_rom[ 1899]='h00001dac;  wr_data_rom[ 1899]='h000008d7;
    rd_cycle[ 1900] = 1'b0;  wr_cycle[ 1900] = 1'b1;  addr_rom[ 1900]='h00001db0;  wr_data_rom[ 1900]='h00000bce;
    rd_cycle[ 1901] = 1'b0;  wr_cycle[ 1901] = 1'b1;  addr_rom[ 1901]='h00001db4;  wr_data_rom[ 1901]='h00001a22;
    rd_cycle[ 1902] = 1'b0;  wr_cycle[ 1902] = 1'b1;  addr_rom[ 1902]='h00001db8;  wr_data_rom[ 1902]='h000001e9;
    rd_cycle[ 1903] = 1'b0;  wr_cycle[ 1903] = 1'b1;  addr_rom[ 1903]='h00001dbc;  wr_data_rom[ 1903]='h00001849;
    rd_cycle[ 1904] = 1'b0;  wr_cycle[ 1904] = 1'b1;  addr_rom[ 1904]='h00001dc0;  wr_data_rom[ 1904]='h000000f3;
    rd_cycle[ 1905] = 1'b0;  wr_cycle[ 1905] = 1'b1;  addr_rom[ 1905]='h00001dc4;  wr_data_rom[ 1905]='h00000e72;
    rd_cycle[ 1906] = 1'b0;  wr_cycle[ 1906] = 1'b1;  addr_rom[ 1906]='h00001dc8;  wr_data_rom[ 1906]='h00000e29;
    rd_cycle[ 1907] = 1'b0;  wr_cycle[ 1907] = 1'b1;  addr_rom[ 1907]='h00001dcc;  wr_data_rom[ 1907]='h00001215;
    rd_cycle[ 1908] = 1'b0;  wr_cycle[ 1908] = 1'b1;  addr_rom[ 1908]='h00001dd0;  wr_data_rom[ 1908]='h000013fa;
    rd_cycle[ 1909] = 1'b0;  wr_cycle[ 1909] = 1'b1;  addr_rom[ 1909]='h00001dd4;  wr_data_rom[ 1909]='h000004e6;
    rd_cycle[ 1910] = 1'b0;  wr_cycle[ 1910] = 1'b1;  addr_rom[ 1910]='h00001dd8;  wr_data_rom[ 1910]='h00000955;
    rd_cycle[ 1911] = 1'b0;  wr_cycle[ 1911] = 1'b1;  addr_rom[ 1911]='h00001ddc;  wr_data_rom[ 1911]='h00000b4f;
    rd_cycle[ 1912] = 1'b0;  wr_cycle[ 1912] = 1'b1;  addr_rom[ 1912]='h00001de0;  wr_data_rom[ 1912]='h000017dd;
    rd_cycle[ 1913] = 1'b0;  wr_cycle[ 1913] = 1'b1;  addr_rom[ 1913]='h00001de4;  wr_data_rom[ 1913]='h00001375;
    rd_cycle[ 1914] = 1'b0;  wr_cycle[ 1914] = 1'b1;  addr_rom[ 1914]='h00001de8;  wr_data_rom[ 1914]='h00001b61;
    rd_cycle[ 1915] = 1'b0;  wr_cycle[ 1915] = 1'b1;  addr_rom[ 1915]='h00001dec;  wr_data_rom[ 1915]='h00001abd;
    rd_cycle[ 1916] = 1'b0;  wr_cycle[ 1916] = 1'b1;  addr_rom[ 1916]='h00001df0;  wr_data_rom[ 1916]='h00000b60;
    rd_cycle[ 1917] = 1'b0;  wr_cycle[ 1917] = 1'b1;  addr_rom[ 1917]='h00001df4;  wr_data_rom[ 1917]='h0000135b;
    rd_cycle[ 1918] = 1'b0;  wr_cycle[ 1918] = 1'b1;  addr_rom[ 1918]='h00001df8;  wr_data_rom[ 1918]='h00001728;
    rd_cycle[ 1919] = 1'b0;  wr_cycle[ 1919] = 1'b1;  addr_rom[ 1919]='h00001dfc;  wr_data_rom[ 1919]='h000010b6;
    rd_cycle[ 1920] = 1'b0;  wr_cycle[ 1920] = 1'b1;  addr_rom[ 1920]='h00001e00;  wr_data_rom[ 1920]='h00001cef;
    rd_cycle[ 1921] = 1'b0;  wr_cycle[ 1921] = 1'b1;  addr_rom[ 1921]='h00001e04;  wr_data_rom[ 1921]='h000004ae;
    rd_cycle[ 1922] = 1'b0;  wr_cycle[ 1922] = 1'b1;  addr_rom[ 1922]='h00001e08;  wr_data_rom[ 1922]='h00000b6e;
    rd_cycle[ 1923] = 1'b0;  wr_cycle[ 1923] = 1'b1;  addr_rom[ 1923]='h00001e0c;  wr_data_rom[ 1923]='h00001a7c;
    rd_cycle[ 1924] = 1'b0;  wr_cycle[ 1924] = 1'b1;  addr_rom[ 1924]='h00001e10;  wr_data_rom[ 1924]='h0000001a;
    rd_cycle[ 1925] = 1'b0;  wr_cycle[ 1925] = 1'b1;  addr_rom[ 1925]='h00001e14;  wr_data_rom[ 1925]='h0000183d;
    rd_cycle[ 1926] = 1'b0;  wr_cycle[ 1926] = 1'b1;  addr_rom[ 1926]='h00001e18;  wr_data_rom[ 1926]='h00000487;
    rd_cycle[ 1927] = 1'b0;  wr_cycle[ 1927] = 1'b1;  addr_rom[ 1927]='h00001e1c;  wr_data_rom[ 1927]='h00000413;
    rd_cycle[ 1928] = 1'b0;  wr_cycle[ 1928] = 1'b1;  addr_rom[ 1928]='h00001e20;  wr_data_rom[ 1928]='h000001ec;
    rd_cycle[ 1929] = 1'b0;  wr_cycle[ 1929] = 1'b1;  addr_rom[ 1929]='h00001e24;  wr_data_rom[ 1929]='h00000fc4;
    rd_cycle[ 1930] = 1'b0;  wr_cycle[ 1930] = 1'b1;  addr_rom[ 1930]='h00001e28;  wr_data_rom[ 1930]='h00000b40;
    rd_cycle[ 1931] = 1'b0;  wr_cycle[ 1931] = 1'b1;  addr_rom[ 1931]='h00001e2c;  wr_data_rom[ 1931]='h000007b5;
    rd_cycle[ 1932] = 1'b0;  wr_cycle[ 1932] = 1'b1;  addr_rom[ 1932]='h00001e30;  wr_data_rom[ 1932]='h000000bc;
    rd_cycle[ 1933] = 1'b0;  wr_cycle[ 1933] = 1'b1;  addr_rom[ 1933]='h00001e34;  wr_data_rom[ 1933]='h00000169;
    rd_cycle[ 1934] = 1'b0;  wr_cycle[ 1934] = 1'b1;  addr_rom[ 1934]='h00001e38;  wr_data_rom[ 1934]='h00001d27;
    rd_cycle[ 1935] = 1'b0;  wr_cycle[ 1935] = 1'b1;  addr_rom[ 1935]='h00001e3c;  wr_data_rom[ 1935]='h00000a51;
    rd_cycle[ 1936] = 1'b0;  wr_cycle[ 1936] = 1'b1;  addr_rom[ 1936]='h00001e40;  wr_data_rom[ 1936]='h00000c1b;
    rd_cycle[ 1937] = 1'b0;  wr_cycle[ 1937] = 1'b1;  addr_rom[ 1937]='h00001e44;  wr_data_rom[ 1937]='h000016d0;
    rd_cycle[ 1938] = 1'b0;  wr_cycle[ 1938] = 1'b1;  addr_rom[ 1938]='h00001e48;  wr_data_rom[ 1938]='h00001dda;
    rd_cycle[ 1939] = 1'b0;  wr_cycle[ 1939] = 1'b1;  addr_rom[ 1939]='h00001e4c;  wr_data_rom[ 1939]='h00000411;
    rd_cycle[ 1940] = 1'b0;  wr_cycle[ 1940] = 1'b1;  addr_rom[ 1940]='h00001e50;  wr_data_rom[ 1940]='h00001d0f;
    rd_cycle[ 1941] = 1'b0;  wr_cycle[ 1941] = 1'b1;  addr_rom[ 1941]='h00001e54;  wr_data_rom[ 1941]='h00001acd;
    rd_cycle[ 1942] = 1'b0;  wr_cycle[ 1942] = 1'b1;  addr_rom[ 1942]='h00001e58;  wr_data_rom[ 1942]='h00001d41;
    rd_cycle[ 1943] = 1'b0;  wr_cycle[ 1943] = 1'b1;  addr_rom[ 1943]='h00001e5c;  wr_data_rom[ 1943]='h000011a5;
    rd_cycle[ 1944] = 1'b0;  wr_cycle[ 1944] = 1'b1;  addr_rom[ 1944]='h00001e60;  wr_data_rom[ 1944]='h000015bb;
    rd_cycle[ 1945] = 1'b0;  wr_cycle[ 1945] = 1'b1;  addr_rom[ 1945]='h00001e64;  wr_data_rom[ 1945]='h000005e3;
    rd_cycle[ 1946] = 1'b0;  wr_cycle[ 1946] = 1'b1;  addr_rom[ 1946]='h00001e68;  wr_data_rom[ 1946]='h00001bf9;
    rd_cycle[ 1947] = 1'b0;  wr_cycle[ 1947] = 1'b1;  addr_rom[ 1947]='h00001e6c;  wr_data_rom[ 1947]='h000015ca;
    rd_cycle[ 1948] = 1'b0;  wr_cycle[ 1948] = 1'b1;  addr_rom[ 1948]='h00001e70;  wr_data_rom[ 1948]='h00001072;
    rd_cycle[ 1949] = 1'b0;  wr_cycle[ 1949] = 1'b1;  addr_rom[ 1949]='h00001e74;  wr_data_rom[ 1949]='h00000b28;
    rd_cycle[ 1950] = 1'b0;  wr_cycle[ 1950] = 1'b1;  addr_rom[ 1950]='h00001e78;  wr_data_rom[ 1950]='h00000ab8;
    rd_cycle[ 1951] = 1'b0;  wr_cycle[ 1951] = 1'b1;  addr_rom[ 1951]='h00001e7c;  wr_data_rom[ 1951]='h00000714;
    rd_cycle[ 1952] = 1'b0;  wr_cycle[ 1952] = 1'b1;  addr_rom[ 1952]='h00001e80;  wr_data_rom[ 1952]='h000019ac;
    rd_cycle[ 1953] = 1'b0;  wr_cycle[ 1953] = 1'b1;  addr_rom[ 1953]='h00001e84;  wr_data_rom[ 1953]='h00001805;
    rd_cycle[ 1954] = 1'b0;  wr_cycle[ 1954] = 1'b1;  addr_rom[ 1954]='h00001e88;  wr_data_rom[ 1954]='h0000020e;
    rd_cycle[ 1955] = 1'b0;  wr_cycle[ 1955] = 1'b1;  addr_rom[ 1955]='h00001e8c;  wr_data_rom[ 1955]='h00000746;
    rd_cycle[ 1956] = 1'b0;  wr_cycle[ 1956] = 1'b1;  addr_rom[ 1956]='h00001e90;  wr_data_rom[ 1956]='h00001c6f;
    rd_cycle[ 1957] = 1'b0;  wr_cycle[ 1957] = 1'b1;  addr_rom[ 1957]='h00001e94;  wr_data_rom[ 1957]='h000003af;
    rd_cycle[ 1958] = 1'b0;  wr_cycle[ 1958] = 1'b1;  addr_rom[ 1958]='h00001e98;  wr_data_rom[ 1958]='h000013ee;
    rd_cycle[ 1959] = 1'b0;  wr_cycle[ 1959] = 1'b1;  addr_rom[ 1959]='h00001e9c;  wr_data_rom[ 1959]='h000019ed;
    rd_cycle[ 1960] = 1'b0;  wr_cycle[ 1960] = 1'b1;  addr_rom[ 1960]='h00001ea0;  wr_data_rom[ 1960]='h00001a04;
    rd_cycle[ 1961] = 1'b0;  wr_cycle[ 1961] = 1'b1;  addr_rom[ 1961]='h00001ea4;  wr_data_rom[ 1961]='h00000962;
    rd_cycle[ 1962] = 1'b0;  wr_cycle[ 1962] = 1'b1;  addr_rom[ 1962]='h00001ea8;  wr_data_rom[ 1962]='h000006a9;
    rd_cycle[ 1963] = 1'b0;  wr_cycle[ 1963] = 1'b1;  addr_rom[ 1963]='h00001eac;  wr_data_rom[ 1963]='h00001941;
    rd_cycle[ 1964] = 1'b0;  wr_cycle[ 1964] = 1'b1;  addr_rom[ 1964]='h00001eb0;  wr_data_rom[ 1964]='h000000a1;
    rd_cycle[ 1965] = 1'b0;  wr_cycle[ 1965] = 1'b1;  addr_rom[ 1965]='h00001eb4;  wr_data_rom[ 1965]='h00001d58;
    rd_cycle[ 1966] = 1'b0;  wr_cycle[ 1966] = 1'b1;  addr_rom[ 1966]='h00001eb8;  wr_data_rom[ 1966]='h00000884;
    rd_cycle[ 1967] = 1'b0;  wr_cycle[ 1967] = 1'b1;  addr_rom[ 1967]='h00001ebc;  wr_data_rom[ 1967]='h0000144e;
    rd_cycle[ 1968] = 1'b0;  wr_cycle[ 1968] = 1'b1;  addr_rom[ 1968]='h00001ec0;  wr_data_rom[ 1968]='h00000e7d;
    rd_cycle[ 1969] = 1'b0;  wr_cycle[ 1969] = 1'b1;  addr_rom[ 1969]='h00001ec4;  wr_data_rom[ 1969]='h00000161;
    rd_cycle[ 1970] = 1'b0;  wr_cycle[ 1970] = 1'b1;  addr_rom[ 1970]='h00001ec8;  wr_data_rom[ 1970]='h00001488;
    rd_cycle[ 1971] = 1'b0;  wr_cycle[ 1971] = 1'b1;  addr_rom[ 1971]='h00001ecc;  wr_data_rom[ 1971]='h00000be8;
    rd_cycle[ 1972] = 1'b0;  wr_cycle[ 1972] = 1'b1;  addr_rom[ 1972]='h00001ed0;  wr_data_rom[ 1972]='h000015d3;
    rd_cycle[ 1973] = 1'b0;  wr_cycle[ 1973] = 1'b1;  addr_rom[ 1973]='h00001ed4;  wr_data_rom[ 1973]='h000008c1;
    rd_cycle[ 1974] = 1'b0;  wr_cycle[ 1974] = 1'b1;  addr_rom[ 1974]='h00001ed8;  wr_data_rom[ 1974]='h00001997;
    rd_cycle[ 1975] = 1'b0;  wr_cycle[ 1975] = 1'b1;  addr_rom[ 1975]='h00001edc;  wr_data_rom[ 1975]='h00001820;
    rd_cycle[ 1976] = 1'b0;  wr_cycle[ 1976] = 1'b1;  addr_rom[ 1976]='h00001ee0;  wr_data_rom[ 1976]='h00001340;
    rd_cycle[ 1977] = 1'b0;  wr_cycle[ 1977] = 1'b1;  addr_rom[ 1977]='h00001ee4;  wr_data_rom[ 1977]='h00000459;
    rd_cycle[ 1978] = 1'b0;  wr_cycle[ 1978] = 1'b1;  addr_rom[ 1978]='h00001ee8;  wr_data_rom[ 1978]='h00000579;
    rd_cycle[ 1979] = 1'b0;  wr_cycle[ 1979] = 1'b1;  addr_rom[ 1979]='h00001eec;  wr_data_rom[ 1979]='h0000197f;
    rd_cycle[ 1980] = 1'b0;  wr_cycle[ 1980] = 1'b1;  addr_rom[ 1980]='h00001ef0;  wr_data_rom[ 1980]='h00000207;
    rd_cycle[ 1981] = 1'b0;  wr_cycle[ 1981] = 1'b1;  addr_rom[ 1981]='h00001ef4;  wr_data_rom[ 1981]='h00001a6a;
    rd_cycle[ 1982] = 1'b0;  wr_cycle[ 1982] = 1'b1;  addr_rom[ 1982]='h00001ef8;  wr_data_rom[ 1982]='h000003df;
    rd_cycle[ 1983] = 1'b0;  wr_cycle[ 1983] = 1'b1;  addr_rom[ 1983]='h00001efc;  wr_data_rom[ 1983]='h000015d0;
    rd_cycle[ 1984] = 1'b0;  wr_cycle[ 1984] = 1'b1;  addr_rom[ 1984]='h00001f00;  wr_data_rom[ 1984]='h000010f3;
    rd_cycle[ 1985] = 1'b0;  wr_cycle[ 1985] = 1'b1;  addr_rom[ 1985]='h00001f04;  wr_data_rom[ 1985]='h0000056a;
    rd_cycle[ 1986] = 1'b0;  wr_cycle[ 1986] = 1'b1;  addr_rom[ 1986]='h00001f08;  wr_data_rom[ 1986]='h000019fd;
    rd_cycle[ 1987] = 1'b0;  wr_cycle[ 1987] = 1'b1;  addr_rom[ 1987]='h00001f0c;  wr_data_rom[ 1987]='h00001b6d;
    rd_cycle[ 1988] = 1'b0;  wr_cycle[ 1988] = 1'b1;  addr_rom[ 1988]='h00001f10;  wr_data_rom[ 1988]='h00001629;
    rd_cycle[ 1989] = 1'b0;  wr_cycle[ 1989] = 1'b1;  addr_rom[ 1989]='h00001f14;  wr_data_rom[ 1989]='h00001171;
    rd_cycle[ 1990] = 1'b0;  wr_cycle[ 1990] = 1'b1;  addr_rom[ 1990]='h00001f18;  wr_data_rom[ 1990]='h00000bae;
    rd_cycle[ 1991] = 1'b0;  wr_cycle[ 1991] = 1'b1;  addr_rom[ 1991]='h00001f1c;  wr_data_rom[ 1991]='h00000900;
    rd_cycle[ 1992] = 1'b0;  wr_cycle[ 1992] = 1'b1;  addr_rom[ 1992]='h00001f20;  wr_data_rom[ 1992]='h0000070c;
    rd_cycle[ 1993] = 1'b0;  wr_cycle[ 1993] = 1'b1;  addr_rom[ 1993]='h00001f24;  wr_data_rom[ 1993]='h00000036;
    rd_cycle[ 1994] = 1'b0;  wr_cycle[ 1994] = 1'b1;  addr_rom[ 1994]='h00001f28;  wr_data_rom[ 1994]='h000012cd;
    rd_cycle[ 1995] = 1'b0;  wr_cycle[ 1995] = 1'b1;  addr_rom[ 1995]='h00001f2c;  wr_data_rom[ 1995]='h000006cd;
    rd_cycle[ 1996] = 1'b0;  wr_cycle[ 1996] = 1'b1;  addr_rom[ 1996]='h00001f30;  wr_data_rom[ 1996]='h0000045f;
    rd_cycle[ 1997] = 1'b0;  wr_cycle[ 1997] = 1'b1;  addr_rom[ 1997]='h00001f34;  wr_data_rom[ 1997]='h000006c7;
    rd_cycle[ 1998] = 1'b0;  wr_cycle[ 1998] = 1'b1;  addr_rom[ 1998]='h00001f38;  wr_data_rom[ 1998]='h0000065f;
    rd_cycle[ 1999] = 1'b0;  wr_cycle[ 1999] = 1'b1;  addr_rom[ 1999]='h00001f3c;  wr_data_rom[ 1999]='h00001148;
    // 6000 random read and write cycles
    rd_cycle[ 2000] = 1'b1;  wr_cycle[ 2000] = 1'b0;  addr_rom[ 2000]='h000005b8;  wr_data_rom[ 2000]='h00000000;
    rd_cycle[ 2001] = 1'b1;  wr_cycle[ 2001] = 1'b0;  addr_rom[ 2001]='h00000d48;  wr_data_rom[ 2001]='h00000000;
    rd_cycle[ 2002] = 1'b1;  wr_cycle[ 2002] = 1'b0;  addr_rom[ 2002]='h00000694;  wr_data_rom[ 2002]='h00000000;
    rd_cycle[ 2003] = 1'b0;  wr_cycle[ 2003] = 1'b1;  addr_rom[ 2003]='h0000130c;  wr_data_rom[ 2003]='h000006ea;
    rd_cycle[ 2004] = 1'b0;  wr_cycle[ 2004] = 1'b1;  addr_rom[ 2004]='h00001bfc;  wr_data_rom[ 2004]='h00000a64;
    rd_cycle[ 2005] = 1'b1;  wr_cycle[ 2005] = 1'b0;  addr_rom[ 2005]='h00000438;  wr_data_rom[ 2005]='h00000000;
    rd_cycle[ 2006] = 1'b1;  wr_cycle[ 2006] = 1'b0;  addr_rom[ 2006]='h00000fa8;  wr_data_rom[ 2006]='h00000000;
    rd_cycle[ 2007] = 1'b0;  wr_cycle[ 2007] = 1'b1;  addr_rom[ 2007]='h0000036c;  wr_data_rom[ 2007]='h00001890;
    rd_cycle[ 2008] = 1'b0;  wr_cycle[ 2008] = 1'b1;  addr_rom[ 2008]='h000010e8;  wr_data_rom[ 2008]='h0000036e;
    rd_cycle[ 2009] = 1'b0;  wr_cycle[ 2009] = 1'b1;  addr_rom[ 2009]='h00000824;  wr_data_rom[ 2009]='h00000f42;
    rd_cycle[ 2010] = 1'b1;  wr_cycle[ 2010] = 1'b0;  addr_rom[ 2010]='h00001e34;  wr_data_rom[ 2010]='h00000000;
    rd_cycle[ 2011] = 1'b1;  wr_cycle[ 2011] = 1'b0;  addr_rom[ 2011]='h00000208;  wr_data_rom[ 2011]='h00000000;
    rd_cycle[ 2012] = 1'b1;  wr_cycle[ 2012] = 1'b0;  addr_rom[ 2012]='h000003fc;  wr_data_rom[ 2012]='h00000000;
    rd_cycle[ 2013] = 1'b0;  wr_cycle[ 2013] = 1'b1;  addr_rom[ 2013]='h000001e0;  wr_data_rom[ 2013]='h000001d1;
    rd_cycle[ 2014] = 1'b1;  wr_cycle[ 2014] = 1'b0;  addr_rom[ 2014]='h00000b64;  wr_data_rom[ 2014]='h00000000;
    rd_cycle[ 2015] = 1'b1;  wr_cycle[ 2015] = 1'b0;  addr_rom[ 2015]='h000006bc;  wr_data_rom[ 2015]='h00000000;
    rd_cycle[ 2016] = 1'b0;  wr_cycle[ 2016] = 1'b1;  addr_rom[ 2016]='h00001c80;  wr_data_rom[ 2016]='h00000c22;
    rd_cycle[ 2017] = 1'b1;  wr_cycle[ 2017] = 1'b0;  addr_rom[ 2017]='h00001848;  wr_data_rom[ 2017]='h00000000;
    rd_cycle[ 2018] = 1'b0;  wr_cycle[ 2018] = 1'b1;  addr_rom[ 2018]='h00000ae0;  wr_data_rom[ 2018]='h00000d5a;
    rd_cycle[ 2019] = 1'b1;  wr_cycle[ 2019] = 1'b0;  addr_rom[ 2019]='h0000014c;  wr_data_rom[ 2019]='h00000000;
    rd_cycle[ 2020] = 1'b1;  wr_cycle[ 2020] = 1'b0;  addr_rom[ 2020]='h00000cf4;  wr_data_rom[ 2020]='h00000000;
    rd_cycle[ 2021] = 1'b0;  wr_cycle[ 2021] = 1'b1;  addr_rom[ 2021]='h000019a4;  wr_data_rom[ 2021]='h000001df;
    rd_cycle[ 2022] = 1'b0;  wr_cycle[ 2022] = 1'b1;  addr_rom[ 2022]='h00000ba8;  wr_data_rom[ 2022]='h000008b0;
    rd_cycle[ 2023] = 1'b1;  wr_cycle[ 2023] = 1'b0;  addr_rom[ 2023]='h00000f44;  wr_data_rom[ 2023]='h00000000;
    rd_cycle[ 2024] = 1'b0;  wr_cycle[ 2024] = 1'b1;  addr_rom[ 2024]='h000016f4;  wr_data_rom[ 2024]='h00000f58;
    rd_cycle[ 2025] = 1'b0;  wr_cycle[ 2025] = 1'b1;  addr_rom[ 2025]='h00000168;  wr_data_rom[ 2025]='h000004da;
    rd_cycle[ 2026] = 1'b1;  wr_cycle[ 2026] = 1'b0;  addr_rom[ 2026]='h00000558;  wr_data_rom[ 2026]='h00000000;
    rd_cycle[ 2027] = 1'b0;  wr_cycle[ 2027] = 1'b1;  addr_rom[ 2027]='h00001d34;  wr_data_rom[ 2027]='h00000204;
    rd_cycle[ 2028] = 1'b1;  wr_cycle[ 2028] = 1'b0;  addr_rom[ 2028]='h000003b0;  wr_data_rom[ 2028]='h00000000;
    rd_cycle[ 2029] = 1'b0;  wr_cycle[ 2029] = 1'b1;  addr_rom[ 2029]='h00001e08;  wr_data_rom[ 2029]='h00000d2d;
    rd_cycle[ 2030] = 1'b1;  wr_cycle[ 2030] = 1'b0;  addr_rom[ 2030]='h000004b4;  wr_data_rom[ 2030]='h00000000;
    rd_cycle[ 2031] = 1'b1;  wr_cycle[ 2031] = 1'b0;  addr_rom[ 2031]='h00000598;  wr_data_rom[ 2031]='h00000000;
    rd_cycle[ 2032] = 1'b0;  wr_cycle[ 2032] = 1'b1;  addr_rom[ 2032]='h00001bd0;  wr_data_rom[ 2032]='h0000161d;
    rd_cycle[ 2033] = 1'b1;  wr_cycle[ 2033] = 1'b0;  addr_rom[ 2033]='h00000a10;  wr_data_rom[ 2033]='h00000000;
    rd_cycle[ 2034] = 1'b1;  wr_cycle[ 2034] = 1'b0;  addr_rom[ 2034]='h00000e6c;  wr_data_rom[ 2034]='h00000000;
    rd_cycle[ 2035] = 1'b0;  wr_cycle[ 2035] = 1'b1;  addr_rom[ 2035]='h000012d8;  wr_data_rom[ 2035]='h000009a8;
    rd_cycle[ 2036] = 1'b0;  wr_cycle[ 2036] = 1'b1;  addr_rom[ 2036]='h00001d18;  wr_data_rom[ 2036]='h000001de;
    rd_cycle[ 2037] = 1'b0;  wr_cycle[ 2037] = 1'b1;  addr_rom[ 2037]='h00001028;  wr_data_rom[ 2037]='h000016af;
    rd_cycle[ 2038] = 1'b0;  wr_cycle[ 2038] = 1'b1;  addr_rom[ 2038]='h00000090;  wr_data_rom[ 2038]='h000000f0;
    rd_cycle[ 2039] = 1'b1;  wr_cycle[ 2039] = 1'b0;  addr_rom[ 2039]='h00001848;  wr_data_rom[ 2039]='h00000000;
    rd_cycle[ 2040] = 1'b1;  wr_cycle[ 2040] = 1'b0;  addr_rom[ 2040]='h0000058c;  wr_data_rom[ 2040]='h00000000;
    rd_cycle[ 2041] = 1'b1;  wr_cycle[ 2041] = 1'b0;  addr_rom[ 2041]='h0000095c;  wr_data_rom[ 2041]='h00000000;
    rd_cycle[ 2042] = 1'b0;  wr_cycle[ 2042] = 1'b1;  addr_rom[ 2042]='h00001f24;  wr_data_rom[ 2042]='h000017d6;
    rd_cycle[ 2043] = 1'b0;  wr_cycle[ 2043] = 1'b1;  addr_rom[ 2043]='h00000f4c;  wr_data_rom[ 2043]='h0000112b;
    rd_cycle[ 2044] = 1'b1;  wr_cycle[ 2044] = 1'b0;  addr_rom[ 2044]='h00000970;  wr_data_rom[ 2044]='h00000000;
    rd_cycle[ 2045] = 1'b1;  wr_cycle[ 2045] = 1'b0;  addr_rom[ 2045]='h00001e9c;  wr_data_rom[ 2045]='h00000000;
    rd_cycle[ 2046] = 1'b0;  wr_cycle[ 2046] = 1'b1;  addr_rom[ 2046]='h00000c60;  wr_data_rom[ 2046]='h00001938;
    rd_cycle[ 2047] = 1'b1;  wr_cycle[ 2047] = 1'b0;  addr_rom[ 2047]='h00000ae8;  wr_data_rom[ 2047]='h00000000;
    rd_cycle[ 2048] = 1'b0;  wr_cycle[ 2048] = 1'b1;  addr_rom[ 2048]='h0000125c;  wr_data_rom[ 2048]='h0000171d;
    rd_cycle[ 2049] = 1'b1;  wr_cycle[ 2049] = 1'b0;  addr_rom[ 2049]='h00000c38;  wr_data_rom[ 2049]='h00000000;
    rd_cycle[ 2050] = 1'b0;  wr_cycle[ 2050] = 1'b1;  addr_rom[ 2050]='h000014a4;  wr_data_rom[ 2050]='h00001474;
    rd_cycle[ 2051] = 1'b0;  wr_cycle[ 2051] = 1'b1;  addr_rom[ 2051]='h00001b6c;  wr_data_rom[ 2051]='h00000753;
    rd_cycle[ 2052] = 1'b1;  wr_cycle[ 2052] = 1'b0;  addr_rom[ 2052]='h00000b14;  wr_data_rom[ 2052]='h00000000;
    rd_cycle[ 2053] = 1'b0;  wr_cycle[ 2053] = 1'b1;  addr_rom[ 2053]='h00000228;  wr_data_rom[ 2053]='h00000bc1;
    rd_cycle[ 2054] = 1'b1;  wr_cycle[ 2054] = 1'b0;  addr_rom[ 2054]='h00001738;  wr_data_rom[ 2054]='h00000000;
    rd_cycle[ 2055] = 1'b1;  wr_cycle[ 2055] = 1'b0;  addr_rom[ 2055]='h00000800;  wr_data_rom[ 2055]='h00000000;
    rd_cycle[ 2056] = 1'b0;  wr_cycle[ 2056] = 1'b1;  addr_rom[ 2056]='h00000b08;  wr_data_rom[ 2056]='h00000a6e;
    rd_cycle[ 2057] = 1'b1;  wr_cycle[ 2057] = 1'b0;  addr_rom[ 2057]='h000007e8;  wr_data_rom[ 2057]='h00000000;
    rd_cycle[ 2058] = 1'b0;  wr_cycle[ 2058] = 1'b1;  addr_rom[ 2058]='h00000b94;  wr_data_rom[ 2058]='h00001e7a;
    rd_cycle[ 2059] = 1'b0;  wr_cycle[ 2059] = 1'b1;  addr_rom[ 2059]='h0000095c;  wr_data_rom[ 2059]='h000009d7;
    rd_cycle[ 2060] = 1'b1;  wr_cycle[ 2060] = 1'b0;  addr_rom[ 2060]='h0000017c;  wr_data_rom[ 2060]='h00000000;
    rd_cycle[ 2061] = 1'b0;  wr_cycle[ 2061] = 1'b1;  addr_rom[ 2061]='h000012f4;  wr_data_rom[ 2061]='h00001ee8;
    rd_cycle[ 2062] = 1'b1;  wr_cycle[ 2062] = 1'b0;  addr_rom[ 2062]='h00001844;  wr_data_rom[ 2062]='h00000000;
    rd_cycle[ 2063] = 1'b0;  wr_cycle[ 2063] = 1'b1;  addr_rom[ 2063]='h00001588;  wr_data_rom[ 2063]='h00000888;
    rd_cycle[ 2064] = 1'b0;  wr_cycle[ 2064] = 1'b1;  addr_rom[ 2064]='h0000060c;  wr_data_rom[ 2064]='h0000039b;
    rd_cycle[ 2065] = 1'b0;  wr_cycle[ 2065] = 1'b1;  addr_rom[ 2065]='h00000a9c;  wr_data_rom[ 2065]='h000012d0;
    rd_cycle[ 2066] = 1'b1;  wr_cycle[ 2066] = 1'b0;  addr_rom[ 2066]='h00000904;  wr_data_rom[ 2066]='h00000000;
    rd_cycle[ 2067] = 1'b0;  wr_cycle[ 2067] = 1'b1;  addr_rom[ 2067]='h000011f4;  wr_data_rom[ 2067]='h00001d3b;
    rd_cycle[ 2068] = 1'b1;  wr_cycle[ 2068] = 1'b0;  addr_rom[ 2068]='h00000450;  wr_data_rom[ 2068]='h00000000;
    rd_cycle[ 2069] = 1'b1;  wr_cycle[ 2069] = 1'b0;  addr_rom[ 2069]='h000011b4;  wr_data_rom[ 2069]='h00000000;
    rd_cycle[ 2070] = 1'b1;  wr_cycle[ 2070] = 1'b0;  addr_rom[ 2070]='h00000ec4;  wr_data_rom[ 2070]='h00000000;
    rd_cycle[ 2071] = 1'b0;  wr_cycle[ 2071] = 1'b1;  addr_rom[ 2071]='h0000198c;  wr_data_rom[ 2071]='h0000085b;
    rd_cycle[ 2072] = 1'b0;  wr_cycle[ 2072] = 1'b1;  addr_rom[ 2072]='h000000f4;  wr_data_rom[ 2072]='h000004aa;
    rd_cycle[ 2073] = 1'b0;  wr_cycle[ 2073] = 1'b1;  addr_rom[ 2073]='h00000d28;  wr_data_rom[ 2073]='h00001a70;
    rd_cycle[ 2074] = 1'b1;  wr_cycle[ 2074] = 1'b0;  addr_rom[ 2074]='h00001d74;  wr_data_rom[ 2074]='h00000000;
    rd_cycle[ 2075] = 1'b0;  wr_cycle[ 2075] = 1'b1;  addr_rom[ 2075]='h000016dc;  wr_data_rom[ 2075]='h00001472;
    rd_cycle[ 2076] = 1'b0;  wr_cycle[ 2076] = 1'b1;  addr_rom[ 2076]='h00000db4;  wr_data_rom[ 2076]='h00000b0a;
    rd_cycle[ 2077] = 1'b1;  wr_cycle[ 2077] = 1'b0;  addr_rom[ 2077]='h0000151c;  wr_data_rom[ 2077]='h00000000;
    rd_cycle[ 2078] = 1'b1;  wr_cycle[ 2078] = 1'b0;  addr_rom[ 2078]='h000002b4;  wr_data_rom[ 2078]='h00000000;
    rd_cycle[ 2079] = 1'b0;  wr_cycle[ 2079] = 1'b1;  addr_rom[ 2079]='h00000e1c;  wr_data_rom[ 2079]='h00000c96;
    rd_cycle[ 2080] = 1'b1;  wr_cycle[ 2080] = 1'b0;  addr_rom[ 2080]='h00000490;  wr_data_rom[ 2080]='h00000000;
    rd_cycle[ 2081] = 1'b1;  wr_cycle[ 2081] = 1'b0;  addr_rom[ 2081]='h00001e70;  wr_data_rom[ 2081]='h00000000;
    rd_cycle[ 2082] = 1'b0;  wr_cycle[ 2082] = 1'b1;  addr_rom[ 2082]='h00000818;  wr_data_rom[ 2082]='h00001c30;
    rd_cycle[ 2083] = 1'b0;  wr_cycle[ 2083] = 1'b1;  addr_rom[ 2083]='h000014dc;  wr_data_rom[ 2083]='h00001004;
    rd_cycle[ 2084] = 1'b0;  wr_cycle[ 2084] = 1'b1;  addr_rom[ 2084]='h00001870;  wr_data_rom[ 2084]='h00001c16;
    rd_cycle[ 2085] = 1'b0;  wr_cycle[ 2085] = 1'b1;  addr_rom[ 2085]='h000005cc;  wr_data_rom[ 2085]='h00000cd8;
    rd_cycle[ 2086] = 1'b1;  wr_cycle[ 2086] = 1'b0;  addr_rom[ 2086]='h000015ac;  wr_data_rom[ 2086]='h00000000;
    rd_cycle[ 2087] = 1'b1;  wr_cycle[ 2087] = 1'b0;  addr_rom[ 2087]='h00001c9c;  wr_data_rom[ 2087]='h00000000;
    rd_cycle[ 2088] = 1'b0;  wr_cycle[ 2088] = 1'b1;  addr_rom[ 2088]='h0000103c;  wr_data_rom[ 2088]='h000000de;
    rd_cycle[ 2089] = 1'b1;  wr_cycle[ 2089] = 1'b0;  addr_rom[ 2089]='h00000484;  wr_data_rom[ 2089]='h00000000;
    rd_cycle[ 2090] = 1'b0;  wr_cycle[ 2090] = 1'b1;  addr_rom[ 2090]='h00001440;  wr_data_rom[ 2090]='h00001691;
    rd_cycle[ 2091] = 1'b1;  wr_cycle[ 2091] = 1'b0;  addr_rom[ 2091]='h0000106c;  wr_data_rom[ 2091]='h00000000;
    rd_cycle[ 2092] = 1'b0;  wr_cycle[ 2092] = 1'b1;  addr_rom[ 2092]='h00000294;  wr_data_rom[ 2092]='h000005e3;
    rd_cycle[ 2093] = 1'b0;  wr_cycle[ 2093] = 1'b1;  addr_rom[ 2093]='h00001f00;  wr_data_rom[ 2093]='h00001e05;
    rd_cycle[ 2094] = 1'b0;  wr_cycle[ 2094] = 1'b1;  addr_rom[ 2094]='h000002fc;  wr_data_rom[ 2094]='h00000ccf;
    rd_cycle[ 2095] = 1'b1;  wr_cycle[ 2095] = 1'b0;  addr_rom[ 2095]='h0000111c;  wr_data_rom[ 2095]='h00000000;
    rd_cycle[ 2096] = 1'b0;  wr_cycle[ 2096] = 1'b1;  addr_rom[ 2096]='h00000fd4;  wr_data_rom[ 2096]='h000019e5;
    rd_cycle[ 2097] = 1'b1;  wr_cycle[ 2097] = 1'b0;  addr_rom[ 2097]='h00001120;  wr_data_rom[ 2097]='h00000000;
    rd_cycle[ 2098] = 1'b1;  wr_cycle[ 2098] = 1'b0;  addr_rom[ 2098]='h00001eac;  wr_data_rom[ 2098]='h00000000;
    rd_cycle[ 2099] = 1'b0;  wr_cycle[ 2099] = 1'b1;  addr_rom[ 2099]='h00000afc;  wr_data_rom[ 2099]='h0000063f;
    rd_cycle[ 2100] = 1'b0;  wr_cycle[ 2100] = 1'b1;  addr_rom[ 2100]='h00001148;  wr_data_rom[ 2100]='h0000004a;
    rd_cycle[ 2101] = 1'b1;  wr_cycle[ 2101] = 1'b0;  addr_rom[ 2101]='h00000250;  wr_data_rom[ 2101]='h00000000;
    rd_cycle[ 2102] = 1'b1;  wr_cycle[ 2102] = 1'b0;  addr_rom[ 2102]='h00000a5c;  wr_data_rom[ 2102]='h00000000;
    rd_cycle[ 2103] = 1'b0;  wr_cycle[ 2103] = 1'b1;  addr_rom[ 2103]='h0000049c;  wr_data_rom[ 2103]='h00000c50;
    rd_cycle[ 2104] = 1'b0;  wr_cycle[ 2104] = 1'b1;  addr_rom[ 2104]='h00001b24;  wr_data_rom[ 2104]='h000012f4;
    rd_cycle[ 2105] = 1'b1;  wr_cycle[ 2105] = 1'b0;  addr_rom[ 2105]='h00000a38;  wr_data_rom[ 2105]='h00000000;
    rd_cycle[ 2106] = 1'b1;  wr_cycle[ 2106] = 1'b0;  addr_rom[ 2106]='h00000964;  wr_data_rom[ 2106]='h00000000;
    rd_cycle[ 2107] = 1'b0;  wr_cycle[ 2107] = 1'b1;  addr_rom[ 2107]='h00000cf4;  wr_data_rom[ 2107]='h00000425;
    rd_cycle[ 2108] = 1'b0;  wr_cycle[ 2108] = 1'b1;  addr_rom[ 2108]='h0000126c;  wr_data_rom[ 2108]='h0000157c;
    rd_cycle[ 2109] = 1'b1;  wr_cycle[ 2109] = 1'b0;  addr_rom[ 2109]='h00001b74;  wr_data_rom[ 2109]='h00000000;
    rd_cycle[ 2110] = 1'b0;  wr_cycle[ 2110] = 1'b1;  addr_rom[ 2110]='h00001f38;  wr_data_rom[ 2110]='h000015d9;
    rd_cycle[ 2111] = 1'b0;  wr_cycle[ 2111] = 1'b1;  addr_rom[ 2111]='h00001d64;  wr_data_rom[ 2111]='h00001794;
    rd_cycle[ 2112] = 1'b0;  wr_cycle[ 2112] = 1'b1;  addr_rom[ 2112]='h0000134c;  wr_data_rom[ 2112]='h00000d5a;
    rd_cycle[ 2113] = 1'b1;  wr_cycle[ 2113] = 1'b0;  addr_rom[ 2113]='h00001c24;  wr_data_rom[ 2113]='h00000000;
    rd_cycle[ 2114] = 1'b1;  wr_cycle[ 2114] = 1'b0;  addr_rom[ 2114]='h00000ed8;  wr_data_rom[ 2114]='h00000000;
    rd_cycle[ 2115] = 1'b0;  wr_cycle[ 2115] = 1'b1;  addr_rom[ 2115]='h00001c60;  wr_data_rom[ 2115]='h00001629;
    rd_cycle[ 2116] = 1'b1;  wr_cycle[ 2116] = 1'b0;  addr_rom[ 2116]='h000004e8;  wr_data_rom[ 2116]='h00000000;
    rd_cycle[ 2117] = 1'b0;  wr_cycle[ 2117] = 1'b1;  addr_rom[ 2117]='h00001e50;  wr_data_rom[ 2117]='h000008c9;
    rd_cycle[ 2118] = 1'b0;  wr_cycle[ 2118] = 1'b1;  addr_rom[ 2118]='h00000298;  wr_data_rom[ 2118]='h00000274;
    rd_cycle[ 2119] = 1'b0;  wr_cycle[ 2119] = 1'b1;  addr_rom[ 2119]='h0000138c;  wr_data_rom[ 2119]='h00001ef0;
    rd_cycle[ 2120] = 1'b0;  wr_cycle[ 2120] = 1'b1;  addr_rom[ 2120]='h00000ea8;  wr_data_rom[ 2120]='h0000029b;
    rd_cycle[ 2121] = 1'b1;  wr_cycle[ 2121] = 1'b0;  addr_rom[ 2121]='h00001408;  wr_data_rom[ 2121]='h00000000;
    rd_cycle[ 2122] = 1'b1;  wr_cycle[ 2122] = 1'b0;  addr_rom[ 2122]='h000001b8;  wr_data_rom[ 2122]='h00000000;
    rd_cycle[ 2123] = 1'b0;  wr_cycle[ 2123] = 1'b1;  addr_rom[ 2123]='h000013e4;  wr_data_rom[ 2123]='h00000d45;
    rd_cycle[ 2124] = 1'b1;  wr_cycle[ 2124] = 1'b0;  addr_rom[ 2124]='h00000684;  wr_data_rom[ 2124]='h00000000;
    rd_cycle[ 2125] = 1'b1;  wr_cycle[ 2125] = 1'b0;  addr_rom[ 2125]='h00001d64;  wr_data_rom[ 2125]='h00000000;
    rd_cycle[ 2126] = 1'b0;  wr_cycle[ 2126] = 1'b1;  addr_rom[ 2126]='h00000e4c;  wr_data_rom[ 2126]='h00001271;
    rd_cycle[ 2127] = 1'b1;  wr_cycle[ 2127] = 1'b0;  addr_rom[ 2127]='h00000cc0;  wr_data_rom[ 2127]='h00000000;
    rd_cycle[ 2128] = 1'b1;  wr_cycle[ 2128] = 1'b0;  addr_rom[ 2128]='h0000032c;  wr_data_rom[ 2128]='h00000000;
    rd_cycle[ 2129] = 1'b0;  wr_cycle[ 2129] = 1'b1;  addr_rom[ 2129]='h0000003c;  wr_data_rom[ 2129]='h00000e13;
    rd_cycle[ 2130] = 1'b1;  wr_cycle[ 2130] = 1'b0;  addr_rom[ 2130]='h00001558;  wr_data_rom[ 2130]='h00000000;
    rd_cycle[ 2131] = 1'b1;  wr_cycle[ 2131] = 1'b0;  addr_rom[ 2131]='h000005c4;  wr_data_rom[ 2131]='h00000000;
    rd_cycle[ 2132] = 1'b1;  wr_cycle[ 2132] = 1'b0;  addr_rom[ 2132]='h00001ed4;  wr_data_rom[ 2132]='h00000000;
    rd_cycle[ 2133] = 1'b1;  wr_cycle[ 2133] = 1'b0;  addr_rom[ 2133]='h00000cdc;  wr_data_rom[ 2133]='h00000000;
    rd_cycle[ 2134] = 1'b1;  wr_cycle[ 2134] = 1'b0;  addr_rom[ 2134]='h00001658;  wr_data_rom[ 2134]='h00000000;
    rd_cycle[ 2135] = 1'b1;  wr_cycle[ 2135] = 1'b0;  addr_rom[ 2135]='h00001700;  wr_data_rom[ 2135]='h00000000;
    rd_cycle[ 2136] = 1'b0;  wr_cycle[ 2136] = 1'b1;  addr_rom[ 2136]='h000004e0;  wr_data_rom[ 2136]='h00001847;
    rd_cycle[ 2137] = 1'b0;  wr_cycle[ 2137] = 1'b1;  addr_rom[ 2137]='h00000688;  wr_data_rom[ 2137]='h0000153d;
    rd_cycle[ 2138] = 1'b0;  wr_cycle[ 2138] = 1'b1;  addr_rom[ 2138]='h0000154c;  wr_data_rom[ 2138]='h0000061f;
    rd_cycle[ 2139] = 1'b1;  wr_cycle[ 2139] = 1'b0;  addr_rom[ 2139]='h00001668;  wr_data_rom[ 2139]='h00000000;
    rd_cycle[ 2140] = 1'b1;  wr_cycle[ 2140] = 1'b0;  addr_rom[ 2140]='h00000040;  wr_data_rom[ 2140]='h00000000;
    rd_cycle[ 2141] = 1'b1;  wr_cycle[ 2141] = 1'b0;  addr_rom[ 2141]='h00000d64;  wr_data_rom[ 2141]='h00000000;
    rd_cycle[ 2142] = 1'b1;  wr_cycle[ 2142] = 1'b0;  addr_rom[ 2142]='h00001e84;  wr_data_rom[ 2142]='h00000000;
    rd_cycle[ 2143] = 1'b1;  wr_cycle[ 2143] = 1'b0;  addr_rom[ 2143]='h000017f0;  wr_data_rom[ 2143]='h00000000;
    rd_cycle[ 2144] = 1'b1;  wr_cycle[ 2144] = 1'b0;  addr_rom[ 2144]='h00000f80;  wr_data_rom[ 2144]='h00000000;
    rd_cycle[ 2145] = 1'b1;  wr_cycle[ 2145] = 1'b0;  addr_rom[ 2145]='h000016a8;  wr_data_rom[ 2145]='h00000000;
    rd_cycle[ 2146] = 1'b1;  wr_cycle[ 2146] = 1'b0;  addr_rom[ 2146]='h0000001c;  wr_data_rom[ 2146]='h00000000;
    rd_cycle[ 2147] = 1'b1;  wr_cycle[ 2147] = 1'b0;  addr_rom[ 2147]='h000000f8;  wr_data_rom[ 2147]='h00000000;
    rd_cycle[ 2148] = 1'b0;  wr_cycle[ 2148] = 1'b1;  addr_rom[ 2148]='h000004a8;  wr_data_rom[ 2148]='h00001c7a;
    rd_cycle[ 2149] = 1'b1;  wr_cycle[ 2149] = 1'b0;  addr_rom[ 2149]='h00001520;  wr_data_rom[ 2149]='h00000000;
    rd_cycle[ 2150] = 1'b0;  wr_cycle[ 2150] = 1'b1;  addr_rom[ 2150]='h00000730;  wr_data_rom[ 2150]='h00001e69;
    rd_cycle[ 2151] = 1'b1;  wr_cycle[ 2151] = 1'b0;  addr_rom[ 2151]='h000002c4;  wr_data_rom[ 2151]='h00000000;
    rd_cycle[ 2152] = 1'b1;  wr_cycle[ 2152] = 1'b0;  addr_rom[ 2152]='h00001988;  wr_data_rom[ 2152]='h00000000;
    rd_cycle[ 2153] = 1'b1;  wr_cycle[ 2153] = 1'b0;  addr_rom[ 2153]='h0000060c;  wr_data_rom[ 2153]='h00000000;
    rd_cycle[ 2154] = 1'b1;  wr_cycle[ 2154] = 1'b0;  addr_rom[ 2154]='h000015ac;  wr_data_rom[ 2154]='h00000000;
    rd_cycle[ 2155] = 1'b0;  wr_cycle[ 2155] = 1'b1;  addr_rom[ 2155]='h00000764;  wr_data_rom[ 2155]='h00001dfb;
    rd_cycle[ 2156] = 1'b0;  wr_cycle[ 2156] = 1'b1;  addr_rom[ 2156]='h00001e10;  wr_data_rom[ 2156]='h00000dd8;
    rd_cycle[ 2157] = 1'b0;  wr_cycle[ 2157] = 1'b1;  addr_rom[ 2157]='h00001998;  wr_data_rom[ 2157]='h00000c97;
    rd_cycle[ 2158] = 1'b1;  wr_cycle[ 2158] = 1'b0;  addr_rom[ 2158]='h00000d90;  wr_data_rom[ 2158]='h00000000;
    rd_cycle[ 2159] = 1'b0;  wr_cycle[ 2159] = 1'b1;  addr_rom[ 2159]='h00001f38;  wr_data_rom[ 2159]='h000008f1;
    rd_cycle[ 2160] = 1'b0;  wr_cycle[ 2160] = 1'b1;  addr_rom[ 2160]='h0000104c;  wr_data_rom[ 2160]='h000001bf;
    rd_cycle[ 2161] = 1'b0;  wr_cycle[ 2161] = 1'b1;  addr_rom[ 2161]='h00001848;  wr_data_rom[ 2161]='h000017be;
    rd_cycle[ 2162] = 1'b0;  wr_cycle[ 2162] = 1'b1;  addr_rom[ 2162]='h00000128;  wr_data_rom[ 2162]='h0000047f;
    rd_cycle[ 2163] = 1'b1;  wr_cycle[ 2163] = 1'b0;  addr_rom[ 2163]='h00001910;  wr_data_rom[ 2163]='h00000000;
    rd_cycle[ 2164] = 1'b1;  wr_cycle[ 2164] = 1'b0;  addr_rom[ 2164]='h00001bb4;  wr_data_rom[ 2164]='h00000000;
    rd_cycle[ 2165] = 1'b0;  wr_cycle[ 2165] = 1'b1;  addr_rom[ 2165]='h00001d68;  wr_data_rom[ 2165]='h000003c7;
    rd_cycle[ 2166] = 1'b0;  wr_cycle[ 2166] = 1'b1;  addr_rom[ 2166]='h000005e8;  wr_data_rom[ 2166]='h00000de7;
    rd_cycle[ 2167] = 1'b1;  wr_cycle[ 2167] = 1'b0;  addr_rom[ 2167]='h00001674;  wr_data_rom[ 2167]='h00000000;
    rd_cycle[ 2168] = 1'b1;  wr_cycle[ 2168] = 1'b0;  addr_rom[ 2168]='h00000600;  wr_data_rom[ 2168]='h00000000;
    rd_cycle[ 2169] = 1'b1;  wr_cycle[ 2169] = 1'b0;  addr_rom[ 2169]='h0000060c;  wr_data_rom[ 2169]='h00000000;
    rd_cycle[ 2170] = 1'b1;  wr_cycle[ 2170] = 1'b0;  addr_rom[ 2170]='h00000690;  wr_data_rom[ 2170]='h00000000;
    rd_cycle[ 2171] = 1'b1;  wr_cycle[ 2171] = 1'b0;  addr_rom[ 2171]='h00000fd8;  wr_data_rom[ 2171]='h00000000;
    rd_cycle[ 2172] = 1'b1;  wr_cycle[ 2172] = 1'b0;  addr_rom[ 2172]='h00001cd4;  wr_data_rom[ 2172]='h00000000;
    rd_cycle[ 2173] = 1'b0;  wr_cycle[ 2173] = 1'b1;  addr_rom[ 2173]='h00001864;  wr_data_rom[ 2173]='h00001c22;
    rd_cycle[ 2174] = 1'b0;  wr_cycle[ 2174] = 1'b1;  addr_rom[ 2174]='h00001ec4;  wr_data_rom[ 2174]='h00000911;
    rd_cycle[ 2175] = 1'b0;  wr_cycle[ 2175] = 1'b1;  addr_rom[ 2175]='h00000fc8;  wr_data_rom[ 2175]='h000015f1;
    rd_cycle[ 2176] = 1'b0;  wr_cycle[ 2176] = 1'b1;  addr_rom[ 2176]='h00000e08;  wr_data_rom[ 2176]='h00000e50;
    rd_cycle[ 2177] = 1'b0;  wr_cycle[ 2177] = 1'b1;  addr_rom[ 2177]='h00000f64;  wr_data_rom[ 2177]='h00001234;
    rd_cycle[ 2178] = 1'b1;  wr_cycle[ 2178] = 1'b0;  addr_rom[ 2178]='h00000f8c;  wr_data_rom[ 2178]='h00000000;
    rd_cycle[ 2179] = 1'b1;  wr_cycle[ 2179] = 1'b0;  addr_rom[ 2179]='h00001ae8;  wr_data_rom[ 2179]='h00000000;
    rd_cycle[ 2180] = 1'b1;  wr_cycle[ 2180] = 1'b0;  addr_rom[ 2180]='h00000ed4;  wr_data_rom[ 2180]='h00000000;
    rd_cycle[ 2181] = 1'b0;  wr_cycle[ 2181] = 1'b1;  addr_rom[ 2181]='h000003d0;  wr_data_rom[ 2181]='h00000041;
    rd_cycle[ 2182] = 1'b0;  wr_cycle[ 2182] = 1'b1;  addr_rom[ 2182]='h00000e94;  wr_data_rom[ 2182]='h00000a7a;
    rd_cycle[ 2183] = 1'b0;  wr_cycle[ 2183] = 1'b1;  addr_rom[ 2183]='h00000540;  wr_data_rom[ 2183]='h00001662;
    rd_cycle[ 2184] = 1'b1;  wr_cycle[ 2184] = 1'b0;  addr_rom[ 2184]='h00000c7c;  wr_data_rom[ 2184]='h00000000;
    rd_cycle[ 2185] = 1'b0;  wr_cycle[ 2185] = 1'b1;  addr_rom[ 2185]='h00001570;  wr_data_rom[ 2185]='h00000d67;
    rd_cycle[ 2186] = 1'b0;  wr_cycle[ 2186] = 1'b1;  addr_rom[ 2186]='h00000f0c;  wr_data_rom[ 2186]='h00000779;
    rd_cycle[ 2187] = 1'b1;  wr_cycle[ 2187] = 1'b0;  addr_rom[ 2187]='h00001064;  wr_data_rom[ 2187]='h00000000;
    rd_cycle[ 2188] = 1'b1;  wr_cycle[ 2188] = 1'b0;  addr_rom[ 2188]='h000004ac;  wr_data_rom[ 2188]='h00000000;
    rd_cycle[ 2189] = 1'b0;  wr_cycle[ 2189] = 1'b1;  addr_rom[ 2189]='h00001540;  wr_data_rom[ 2189]='h00000910;
    rd_cycle[ 2190] = 1'b0;  wr_cycle[ 2190] = 1'b1;  addr_rom[ 2190]='h00001ae4;  wr_data_rom[ 2190]='h0000026b;
    rd_cycle[ 2191] = 1'b0;  wr_cycle[ 2191] = 1'b1;  addr_rom[ 2191]='h00001434;  wr_data_rom[ 2191]='h00001cb3;
    rd_cycle[ 2192] = 1'b1;  wr_cycle[ 2192] = 1'b0;  addr_rom[ 2192]='h000012b0;  wr_data_rom[ 2192]='h00000000;
    rd_cycle[ 2193] = 1'b1;  wr_cycle[ 2193] = 1'b0;  addr_rom[ 2193]='h00000e30;  wr_data_rom[ 2193]='h00000000;
    rd_cycle[ 2194] = 1'b1;  wr_cycle[ 2194] = 1'b0;  addr_rom[ 2194]='h00000f38;  wr_data_rom[ 2194]='h00000000;
    rd_cycle[ 2195] = 1'b0;  wr_cycle[ 2195] = 1'b1;  addr_rom[ 2195]='h00001290;  wr_data_rom[ 2195]='h00000f14;
    rd_cycle[ 2196] = 1'b1;  wr_cycle[ 2196] = 1'b0;  addr_rom[ 2196]='h00001000;  wr_data_rom[ 2196]='h00000000;
    rd_cycle[ 2197] = 1'b1;  wr_cycle[ 2197] = 1'b0;  addr_rom[ 2197]='h00001340;  wr_data_rom[ 2197]='h00000000;
    rd_cycle[ 2198] = 1'b0;  wr_cycle[ 2198] = 1'b1;  addr_rom[ 2198]='h00001868;  wr_data_rom[ 2198]='h00001569;
    rd_cycle[ 2199] = 1'b1;  wr_cycle[ 2199] = 1'b0;  addr_rom[ 2199]='h000005fc;  wr_data_rom[ 2199]='h00000000;
    rd_cycle[ 2200] = 1'b0;  wr_cycle[ 2200] = 1'b1;  addr_rom[ 2200]='h0000193c;  wr_data_rom[ 2200]='h00001f15;
    rd_cycle[ 2201] = 1'b1;  wr_cycle[ 2201] = 1'b0;  addr_rom[ 2201]='h00001940;  wr_data_rom[ 2201]='h00000000;
    rd_cycle[ 2202] = 1'b1;  wr_cycle[ 2202] = 1'b0;  addr_rom[ 2202]='h0000096c;  wr_data_rom[ 2202]='h00000000;
    rd_cycle[ 2203] = 1'b0;  wr_cycle[ 2203] = 1'b1;  addr_rom[ 2203]='h00001a74;  wr_data_rom[ 2203]='h00001f2e;
    rd_cycle[ 2204] = 1'b0;  wr_cycle[ 2204] = 1'b1;  addr_rom[ 2204]='h00000368;  wr_data_rom[ 2204]='h00001d6f;
    rd_cycle[ 2205] = 1'b1;  wr_cycle[ 2205] = 1'b0;  addr_rom[ 2205]='h00000094;  wr_data_rom[ 2205]='h00000000;
    rd_cycle[ 2206] = 1'b1;  wr_cycle[ 2206] = 1'b0;  addr_rom[ 2206]='h000015c4;  wr_data_rom[ 2206]='h00000000;
    rd_cycle[ 2207] = 1'b0;  wr_cycle[ 2207] = 1'b1;  addr_rom[ 2207]='h00001ee8;  wr_data_rom[ 2207]='h00000d9e;
    rd_cycle[ 2208] = 1'b1;  wr_cycle[ 2208] = 1'b0;  addr_rom[ 2208]='h00000fc0;  wr_data_rom[ 2208]='h00000000;
    rd_cycle[ 2209] = 1'b0;  wr_cycle[ 2209] = 1'b1;  addr_rom[ 2209]='h00000f48;  wr_data_rom[ 2209]='h000019dc;
    rd_cycle[ 2210] = 1'b0;  wr_cycle[ 2210] = 1'b1;  addr_rom[ 2210]='h000009d8;  wr_data_rom[ 2210]='h0000018e;
    rd_cycle[ 2211] = 1'b1;  wr_cycle[ 2211] = 1'b0;  addr_rom[ 2211]='h00000d1c;  wr_data_rom[ 2211]='h00000000;
    rd_cycle[ 2212] = 1'b1;  wr_cycle[ 2212] = 1'b0;  addr_rom[ 2212]='h00000020;  wr_data_rom[ 2212]='h00000000;
    rd_cycle[ 2213] = 1'b0;  wr_cycle[ 2213] = 1'b1;  addr_rom[ 2213]='h00001240;  wr_data_rom[ 2213]='h00000fd2;
    rd_cycle[ 2214] = 1'b0;  wr_cycle[ 2214] = 1'b1;  addr_rom[ 2214]='h00000dac;  wr_data_rom[ 2214]='h00001ebe;
    rd_cycle[ 2215] = 1'b1;  wr_cycle[ 2215] = 1'b0;  addr_rom[ 2215]='h00000ef0;  wr_data_rom[ 2215]='h00000000;
    rd_cycle[ 2216] = 1'b0;  wr_cycle[ 2216] = 1'b1;  addr_rom[ 2216]='h000001dc;  wr_data_rom[ 2216]='h000003c9;
    rd_cycle[ 2217] = 1'b1;  wr_cycle[ 2217] = 1'b0;  addr_rom[ 2217]='h00001978;  wr_data_rom[ 2217]='h00000000;
    rd_cycle[ 2218] = 1'b1;  wr_cycle[ 2218] = 1'b0;  addr_rom[ 2218]='h00000234;  wr_data_rom[ 2218]='h00000000;
    rd_cycle[ 2219] = 1'b1;  wr_cycle[ 2219] = 1'b0;  addr_rom[ 2219]='h00000074;  wr_data_rom[ 2219]='h00000000;
    rd_cycle[ 2220] = 1'b0;  wr_cycle[ 2220] = 1'b1;  addr_rom[ 2220]='h00000f00;  wr_data_rom[ 2220]='h000014ad;
    rd_cycle[ 2221] = 1'b1;  wr_cycle[ 2221] = 1'b0;  addr_rom[ 2221]='h00000a50;  wr_data_rom[ 2221]='h00000000;
    rd_cycle[ 2222] = 1'b1;  wr_cycle[ 2222] = 1'b0;  addr_rom[ 2222]='h0000103c;  wr_data_rom[ 2222]='h00000000;
    rd_cycle[ 2223] = 1'b0;  wr_cycle[ 2223] = 1'b1;  addr_rom[ 2223]='h00001188;  wr_data_rom[ 2223]='h0000005a;
    rd_cycle[ 2224] = 1'b0;  wr_cycle[ 2224] = 1'b1;  addr_rom[ 2224]='h000008c8;  wr_data_rom[ 2224]='h0000058b;
    rd_cycle[ 2225] = 1'b1;  wr_cycle[ 2225] = 1'b0;  addr_rom[ 2225]='h00000274;  wr_data_rom[ 2225]='h00000000;
    rd_cycle[ 2226] = 1'b1;  wr_cycle[ 2226] = 1'b0;  addr_rom[ 2226]='h00001e60;  wr_data_rom[ 2226]='h00000000;
    rd_cycle[ 2227] = 1'b0;  wr_cycle[ 2227] = 1'b1;  addr_rom[ 2227]='h00000608;  wr_data_rom[ 2227]='h000010e3;
    rd_cycle[ 2228] = 1'b0;  wr_cycle[ 2228] = 1'b1;  addr_rom[ 2228]='h00001720;  wr_data_rom[ 2228]='h00000cee;
    rd_cycle[ 2229] = 1'b1;  wr_cycle[ 2229] = 1'b0;  addr_rom[ 2229]='h00001ac8;  wr_data_rom[ 2229]='h00000000;
    rd_cycle[ 2230] = 1'b0;  wr_cycle[ 2230] = 1'b1;  addr_rom[ 2230]='h00001988;  wr_data_rom[ 2230]='h00001ee5;
    rd_cycle[ 2231] = 1'b0;  wr_cycle[ 2231] = 1'b1;  addr_rom[ 2231]='h00000c70;  wr_data_rom[ 2231]='h0000123d;
    rd_cycle[ 2232] = 1'b0;  wr_cycle[ 2232] = 1'b1;  addr_rom[ 2232]='h00001f34;  wr_data_rom[ 2232]='h000009c1;
    rd_cycle[ 2233] = 1'b1;  wr_cycle[ 2233] = 1'b0;  addr_rom[ 2233]='h00001698;  wr_data_rom[ 2233]='h00000000;
    rd_cycle[ 2234] = 1'b1;  wr_cycle[ 2234] = 1'b0;  addr_rom[ 2234]='h00001970;  wr_data_rom[ 2234]='h00000000;
    rd_cycle[ 2235] = 1'b1;  wr_cycle[ 2235] = 1'b0;  addr_rom[ 2235]='h000014c0;  wr_data_rom[ 2235]='h00000000;
    rd_cycle[ 2236] = 1'b0;  wr_cycle[ 2236] = 1'b1;  addr_rom[ 2236]='h00001d84;  wr_data_rom[ 2236]='h0000169c;
    rd_cycle[ 2237] = 1'b1;  wr_cycle[ 2237] = 1'b0;  addr_rom[ 2237]='h00001c6c;  wr_data_rom[ 2237]='h00000000;
    rd_cycle[ 2238] = 1'b1;  wr_cycle[ 2238] = 1'b0;  addr_rom[ 2238]='h000009cc;  wr_data_rom[ 2238]='h00000000;
    rd_cycle[ 2239] = 1'b1;  wr_cycle[ 2239] = 1'b0;  addr_rom[ 2239]='h00001554;  wr_data_rom[ 2239]='h00000000;
    rd_cycle[ 2240] = 1'b1;  wr_cycle[ 2240] = 1'b0;  addr_rom[ 2240]='h0000119c;  wr_data_rom[ 2240]='h00000000;
    rd_cycle[ 2241] = 1'b0;  wr_cycle[ 2241] = 1'b1;  addr_rom[ 2241]='h00001800;  wr_data_rom[ 2241]='h000014a3;
    rd_cycle[ 2242] = 1'b1;  wr_cycle[ 2242] = 1'b0;  addr_rom[ 2242]='h00000094;  wr_data_rom[ 2242]='h00000000;
    rd_cycle[ 2243] = 1'b1;  wr_cycle[ 2243] = 1'b0;  addr_rom[ 2243]='h00001888;  wr_data_rom[ 2243]='h00000000;
    rd_cycle[ 2244] = 1'b1;  wr_cycle[ 2244] = 1'b0;  addr_rom[ 2244]='h000010ac;  wr_data_rom[ 2244]='h00000000;
    rd_cycle[ 2245] = 1'b1;  wr_cycle[ 2245] = 1'b0;  addr_rom[ 2245]='h0000173c;  wr_data_rom[ 2245]='h00000000;
    rd_cycle[ 2246] = 1'b1;  wr_cycle[ 2246] = 1'b0;  addr_rom[ 2246]='h000011a4;  wr_data_rom[ 2246]='h00000000;
    rd_cycle[ 2247] = 1'b0;  wr_cycle[ 2247] = 1'b1;  addr_rom[ 2247]='h00001ee0;  wr_data_rom[ 2247]='h00001550;
    rd_cycle[ 2248] = 1'b1;  wr_cycle[ 2248] = 1'b0;  addr_rom[ 2248]='h00000a14;  wr_data_rom[ 2248]='h00000000;
    rd_cycle[ 2249] = 1'b0;  wr_cycle[ 2249] = 1'b1;  addr_rom[ 2249]='h00001458;  wr_data_rom[ 2249]='h00000b84;
    rd_cycle[ 2250] = 1'b0;  wr_cycle[ 2250] = 1'b1;  addr_rom[ 2250]='h0000163c;  wr_data_rom[ 2250]='h000010cf;
    rd_cycle[ 2251] = 1'b1;  wr_cycle[ 2251] = 1'b0;  addr_rom[ 2251]='h0000186c;  wr_data_rom[ 2251]='h00000000;
    rd_cycle[ 2252] = 1'b1;  wr_cycle[ 2252] = 1'b0;  addr_rom[ 2252]='h00000ff0;  wr_data_rom[ 2252]='h00000000;
    rd_cycle[ 2253] = 1'b0;  wr_cycle[ 2253] = 1'b1;  addr_rom[ 2253]='h000014cc;  wr_data_rom[ 2253]='h000010be;
    rd_cycle[ 2254] = 1'b1;  wr_cycle[ 2254] = 1'b0;  addr_rom[ 2254]='h00001b34;  wr_data_rom[ 2254]='h00000000;
    rd_cycle[ 2255] = 1'b0;  wr_cycle[ 2255] = 1'b1;  addr_rom[ 2255]='h00001bc4;  wr_data_rom[ 2255]='h00001dfc;
    rd_cycle[ 2256] = 1'b0;  wr_cycle[ 2256] = 1'b1;  addr_rom[ 2256]='h00000a6c;  wr_data_rom[ 2256]='h00000c75;
    rd_cycle[ 2257] = 1'b0;  wr_cycle[ 2257] = 1'b1;  addr_rom[ 2257]='h00000dac;  wr_data_rom[ 2257]='h0000104a;
    rd_cycle[ 2258] = 1'b0;  wr_cycle[ 2258] = 1'b1;  addr_rom[ 2258]='h00001d08;  wr_data_rom[ 2258]='h00001c2b;
    rd_cycle[ 2259] = 1'b1;  wr_cycle[ 2259] = 1'b0;  addr_rom[ 2259]='h000002dc;  wr_data_rom[ 2259]='h00000000;
    rd_cycle[ 2260] = 1'b1;  wr_cycle[ 2260] = 1'b0;  addr_rom[ 2260]='h00001e94;  wr_data_rom[ 2260]='h00000000;
    rd_cycle[ 2261] = 1'b0;  wr_cycle[ 2261] = 1'b1;  addr_rom[ 2261]='h00000ab4;  wr_data_rom[ 2261]='h000007c8;
    rd_cycle[ 2262] = 1'b1;  wr_cycle[ 2262] = 1'b0;  addr_rom[ 2262]='h00000774;  wr_data_rom[ 2262]='h00000000;
    rd_cycle[ 2263] = 1'b0;  wr_cycle[ 2263] = 1'b1;  addr_rom[ 2263]='h00000744;  wr_data_rom[ 2263]='h00001345;
    rd_cycle[ 2264] = 1'b0;  wr_cycle[ 2264] = 1'b1;  addr_rom[ 2264]='h000011b8;  wr_data_rom[ 2264]='h0000113e;
    rd_cycle[ 2265] = 1'b1;  wr_cycle[ 2265] = 1'b0;  addr_rom[ 2265]='h000009d0;  wr_data_rom[ 2265]='h00000000;
    rd_cycle[ 2266] = 1'b0;  wr_cycle[ 2266] = 1'b1;  addr_rom[ 2266]='h00001c4c;  wr_data_rom[ 2266]='h00000817;
    rd_cycle[ 2267] = 1'b0;  wr_cycle[ 2267] = 1'b1;  addr_rom[ 2267]='h00001384;  wr_data_rom[ 2267]='h000007fe;
    rd_cycle[ 2268] = 1'b0;  wr_cycle[ 2268] = 1'b1;  addr_rom[ 2268]='h00001178;  wr_data_rom[ 2268]='h000009d9;
    rd_cycle[ 2269] = 1'b1;  wr_cycle[ 2269] = 1'b0;  addr_rom[ 2269]='h00001798;  wr_data_rom[ 2269]='h00000000;
    rd_cycle[ 2270] = 1'b1;  wr_cycle[ 2270] = 1'b0;  addr_rom[ 2270]='h00000ae4;  wr_data_rom[ 2270]='h00000000;
    rd_cycle[ 2271] = 1'b0;  wr_cycle[ 2271] = 1'b1;  addr_rom[ 2271]='h00000394;  wr_data_rom[ 2271]='h000012fb;
    rd_cycle[ 2272] = 1'b1;  wr_cycle[ 2272] = 1'b0;  addr_rom[ 2272]='h000003f4;  wr_data_rom[ 2272]='h00000000;
    rd_cycle[ 2273] = 1'b0;  wr_cycle[ 2273] = 1'b1;  addr_rom[ 2273]='h000012a0;  wr_data_rom[ 2273]='h00001f05;
    rd_cycle[ 2274] = 1'b0;  wr_cycle[ 2274] = 1'b1;  addr_rom[ 2274]='h000004a4;  wr_data_rom[ 2274]='h0000149b;
    rd_cycle[ 2275] = 1'b0;  wr_cycle[ 2275] = 1'b1;  addr_rom[ 2275]='h00001278;  wr_data_rom[ 2275]='h00001c09;
    rd_cycle[ 2276] = 1'b0;  wr_cycle[ 2276] = 1'b1;  addr_rom[ 2276]='h00000e74;  wr_data_rom[ 2276]='h00000d9b;
    rd_cycle[ 2277] = 1'b0;  wr_cycle[ 2277] = 1'b1;  addr_rom[ 2277]='h0000120c;  wr_data_rom[ 2277]='h00000538;
    rd_cycle[ 2278] = 1'b1;  wr_cycle[ 2278] = 1'b0;  addr_rom[ 2278]='h00000f5c;  wr_data_rom[ 2278]='h00000000;
    rd_cycle[ 2279] = 1'b1;  wr_cycle[ 2279] = 1'b0;  addr_rom[ 2279]='h00001098;  wr_data_rom[ 2279]='h00000000;
    rd_cycle[ 2280] = 1'b0;  wr_cycle[ 2280] = 1'b1;  addr_rom[ 2280]='h00001668;  wr_data_rom[ 2280]='h00001442;
    rd_cycle[ 2281] = 1'b0;  wr_cycle[ 2281] = 1'b1;  addr_rom[ 2281]='h000000dc;  wr_data_rom[ 2281]='h00001e6f;
    rd_cycle[ 2282] = 1'b0;  wr_cycle[ 2282] = 1'b1;  addr_rom[ 2282]='h00001e74;  wr_data_rom[ 2282]='h00001a3b;
    rd_cycle[ 2283] = 1'b1;  wr_cycle[ 2283] = 1'b0;  addr_rom[ 2283]='h00001504;  wr_data_rom[ 2283]='h00000000;
    rd_cycle[ 2284] = 1'b1;  wr_cycle[ 2284] = 1'b0;  addr_rom[ 2284]='h00000060;  wr_data_rom[ 2284]='h00000000;
    rd_cycle[ 2285] = 1'b1;  wr_cycle[ 2285] = 1'b0;  addr_rom[ 2285]='h00000e8c;  wr_data_rom[ 2285]='h00000000;
    rd_cycle[ 2286] = 1'b0;  wr_cycle[ 2286] = 1'b1;  addr_rom[ 2286]='h00001478;  wr_data_rom[ 2286]='h00000e51;
    rd_cycle[ 2287] = 1'b1;  wr_cycle[ 2287] = 1'b0;  addr_rom[ 2287]='h000013e8;  wr_data_rom[ 2287]='h00000000;
    rd_cycle[ 2288] = 1'b0;  wr_cycle[ 2288] = 1'b1;  addr_rom[ 2288]='h00001998;  wr_data_rom[ 2288]='h00000189;
    rd_cycle[ 2289] = 1'b0;  wr_cycle[ 2289] = 1'b1;  addr_rom[ 2289]='h0000165c;  wr_data_rom[ 2289]='h00000180;
    rd_cycle[ 2290] = 1'b1;  wr_cycle[ 2290] = 1'b0;  addr_rom[ 2290]='h00001090;  wr_data_rom[ 2290]='h00000000;
    rd_cycle[ 2291] = 1'b1;  wr_cycle[ 2291] = 1'b0;  addr_rom[ 2291]='h000007b4;  wr_data_rom[ 2291]='h00000000;
    rd_cycle[ 2292] = 1'b1;  wr_cycle[ 2292] = 1'b0;  addr_rom[ 2292]='h000017d4;  wr_data_rom[ 2292]='h00000000;
    rd_cycle[ 2293] = 1'b0;  wr_cycle[ 2293] = 1'b1;  addr_rom[ 2293]='h00000f40;  wr_data_rom[ 2293]='h00001a20;
    rd_cycle[ 2294] = 1'b0;  wr_cycle[ 2294] = 1'b1;  addr_rom[ 2294]='h00001bc4;  wr_data_rom[ 2294]='h000001f1;
    rd_cycle[ 2295] = 1'b0;  wr_cycle[ 2295] = 1'b1;  addr_rom[ 2295]='h00001c8c;  wr_data_rom[ 2295]='h00000759;
    rd_cycle[ 2296] = 1'b0;  wr_cycle[ 2296] = 1'b1;  addr_rom[ 2296]='h00001070;  wr_data_rom[ 2296]='h000013a7;
    rd_cycle[ 2297] = 1'b0;  wr_cycle[ 2297] = 1'b1;  addr_rom[ 2297]='h00001860;  wr_data_rom[ 2297]='h000005c4;
    rd_cycle[ 2298] = 1'b1;  wr_cycle[ 2298] = 1'b0;  addr_rom[ 2298]='h00001450;  wr_data_rom[ 2298]='h00000000;
    rd_cycle[ 2299] = 1'b0;  wr_cycle[ 2299] = 1'b1;  addr_rom[ 2299]='h000004a4;  wr_data_rom[ 2299]='h00001431;
    rd_cycle[ 2300] = 1'b0;  wr_cycle[ 2300] = 1'b1;  addr_rom[ 2300]='h00001cb8;  wr_data_rom[ 2300]='h000019f1;
    rd_cycle[ 2301] = 1'b0;  wr_cycle[ 2301] = 1'b1;  addr_rom[ 2301]='h00000084;  wr_data_rom[ 2301]='h00000ec3;
    rd_cycle[ 2302] = 1'b1;  wr_cycle[ 2302] = 1'b0;  addr_rom[ 2302]='h00001258;  wr_data_rom[ 2302]='h00000000;
    rd_cycle[ 2303] = 1'b1;  wr_cycle[ 2303] = 1'b0;  addr_rom[ 2303]='h00000ef8;  wr_data_rom[ 2303]='h00000000;
    rd_cycle[ 2304] = 1'b0;  wr_cycle[ 2304] = 1'b1;  addr_rom[ 2304]='h00000474;  wr_data_rom[ 2304]='h000001ca;
    rd_cycle[ 2305] = 1'b0;  wr_cycle[ 2305] = 1'b1;  addr_rom[ 2305]='h00001dac;  wr_data_rom[ 2305]='h000005b6;
    rd_cycle[ 2306] = 1'b0;  wr_cycle[ 2306] = 1'b1;  addr_rom[ 2306]='h00000950;  wr_data_rom[ 2306]='h00000482;
    rd_cycle[ 2307] = 1'b0;  wr_cycle[ 2307] = 1'b1;  addr_rom[ 2307]='h00001764;  wr_data_rom[ 2307]='h00000079;
    rd_cycle[ 2308] = 1'b1;  wr_cycle[ 2308] = 1'b0;  addr_rom[ 2308]='h00001374;  wr_data_rom[ 2308]='h00000000;
    rd_cycle[ 2309] = 1'b0;  wr_cycle[ 2309] = 1'b1;  addr_rom[ 2309]='h00000a58;  wr_data_rom[ 2309]='h0000060a;
    rd_cycle[ 2310] = 1'b1;  wr_cycle[ 2310] = 1'b0;  addr_rom[ 2310]='h00001d1c;  wr_data_rom[ 2310]='h00000000;
    rd_cycle[ 2311] = 1'b1;  wr_cycle[ 2311] = 1'b0;  addr_rom[ 2311]='h000013d4;  wr_data_rom[ 2311]='h00000000;
    rd_cycle[ 2312] = 1'b0;  wr_cycle[ 2312] = 1'b1;  addr_rom[ 2312]='h0000028c;  wr_data_rom[ 2312]='h00000da7;
    rd_cycle[ 2313] = 1'b0;  wr_cycle[ 2313] = 1'b1;  addr_rom[ 2313]='h00001a7c;  wr_data_rom[ 2313]='h00000d8f;
    rd_cycle[ 2314] = 1'b0;  wr_cycle[ 2314] = 1'b1;  addr_rom[ 2314]='h00000dcc;  wr_data_rom[ 2314]='h000008eb;
    rd_cycle[ 2315] = 1'b1;  wr_cycle[ 2315] = 1'b0;  addr_rom[ 2315]='h00001a8c;  wr_data_rom[ 2315]='h00000000;
    rd_cycle[ 2316] = 1'b0;  wr_cycle[ 2316] = 1'b1;  addr_rom[ 2316]='h0000058c;  wr_data_rom[ 2316]='h00001a21;
    rd_cycle[ 2317] = 1'b1;  wr_cycle[ 2317] = 1'b0;  addr_rom[ 2317]='h00000120;  wr_data_rom[ 2317]='h00000000;
    rd_cycle[ 2318] = 1'b1;  wr_cycle[ 2318] = 1'b0;  addr_rom[ 2318]='h0000018c;  wr_data_rom[ 2318]='h00000000;
    rd_cycle[ 2319] = 1'b0;  wr_cycle[ 2319] = 1'b1;  addr_rom[ 2319]='h00001810;  wr_data_rom[ 2319]='h000004c7;
    rd_cycle[ 2320] = 1'b1;  wr_cycle[ 2320] = 1'b0;  addr_rom[ 2320]='h00001ca4;  wr_data_rom[ 2320]='h00000000;
    rd_cycle[ 2321] = 1'b0;  wr_cycle[ 2321] = 1'b1;  addr_rom[ 2321]='h0000159c;  wr_data_rom[ 2321]='h00001e70;
    rd_cycle[ 2322] = 1'b1;  wr_cycle[ 2322] = 1'b0;  addr_rom[ 2322]='h00000ebc;  wr_data_rom[ 2322]='h00000000;
    rd_cycle[ 2323] = 1'b1;  wr_cycle[ 2323] = 1'b0;  addr_rom[ 2323]='h00000b58;  wr_data_rom[ 2323]='h00000000;
    rd_cycle[ 2324] = 1'b1;  wr_cycle[ 2324] = 1'b0;  addr_rom[ 2324]='h000000a0;  wr_data_rom[ 2324]='h00000000;
    rd_cycle[ 2325] = 1'b1;  wr_cycle[ 2325] = 1'b0;  addr_rom[ 2325]='h000010a8;  wr_data_rom[ 2325]='h00000000;
    rd_cycle[ 2326] = 1'b0;  wr_cycle[ 2326] = 1'b1;  addr_rom[ 2326]='h000001e4;  wr_data_rom[ 2326]='h000011f3;
    rd_cycle[ 2327] = 1'b1;  wr_cycle[ 2327] = 1'b0;  addr_rom[ 2327]='h00001378;  wr_data_rom[ 2327]='h00000000;
    rd_cycle[ 2328] = 1'b1;  wr_cycle[ 2328] = 1'b0;  addr_rom[ 2328]='h00000fec;  wr_data_rom[ 2328]='h00000000;
    rd_cycle[ 2329] = 1'b1;  wr_cycle[ 2329] = 1'b0;  addr_rom[ 2329]='h0000009c;  wr_data_rom[ 2329]='h00000000;
    rd_cycle[ 2330] = 1'b0;  wr_cycle[ 2330] = 1'b1;  addr_rom[ 2330]='h000009f4;  wr_data_rom[ 2330]='h00000801;
    rd_cycle[ 2331] = 1'b0;  wr_cycle[ 2331] = 1'b1;  addr_rom[ 2331]='h00000d64;  wr_data_rom[ 2331]='h00000109;
    rd_cycle[ 2332] = 1'b0;  wr_cycle[ 2332] = 1'b1;  addr_rom[ 2332]='h00000e98;  wr_data_rom[ 2332]='h00000e8a;
    rd_cycle[ 2333] = 1'b1;  wr_cycle[ 2333] = 1'b0;  addr_rom[ 2333]='h00000e34;  wr_data_rom[ 2333]='h00000000;
    rd_cycle[ 2334] = 1'b1;  wr_cycle[ 2334] = 1'b0;  addr_rom[ 2334]='h00001b98;  wr_data_rom[ 2334]='h00000000;
    rd_cycle[ 2335] = 1'b1;  wr_cycle[ 2335] = 1'b0;  addr_rom[ 2335]='h00001a74;  wr_data_rom[ 2335]='h00000000;
    rd_cycle[ 2336] = 1'b0;  wr_cycle[ 2336] = 1'b1;  addr_rom[ 2336]='h000008c8;  wr_data_rom[ 2336]='h00001730;
    rd_cycle[ 2337] = 1'b0;  wr_cycle[ 2337] = 1'b1;  addr_rom[ 2337]='h00001600;  wr_data_rom[ 2337]='h00001718;
    rd_cycle[ 2338] = 1'b0;  wr_cycle[ 2338] = 1'b1;  addr_rom[ 2338]='h00001464;  wr_data_rom[ 2338]='h000006f5;
    rd_cycle[ 2339] = 1'b1;  wr_cycle[ 2339] = 1'b0;  addr_rom[ 2339]='h00001d4c;  wr_data_rom[ 2339]='h00000000;
    rd_cycle[ 2340] = 1'b1;  wr_cycle[ 2340] = 1'b0;  addr_rom[ 2340]='h00000e50;  wr_data_rom[ 2340]='h00000000;
    rd_cycle[ 2341] = 1'b1;  wr_cycle[ 2341] = 1'b0;  addr_rom[ 2341]='h000009b8;  wr_data_rom[ 2341]='h00000000;
    rd_cycle[ 2342] = 1'b1;  wr_cycle[ 2342] = 1'b0;  addr_rom[ 2342]='h00000a68;  wr_data_rom[ 2342]='h00000000;
    rd_cycle[ 2343] = 1'b1;  wr_cycle[ 2343] = 1'b0;  addr_rom[ 2343]='h00000ca8;  wr_data_rom[ 2343]='h00000000;
    rd_cycle[ 2344] = 1'b0;  wr_cycle[ 2344] = 1'b1;  addr_rom[ 2344]='h000005f4;  wr_data_rom[ 2344]='h000005d3;
    rd_cycle[ 2345] = 1'b0;  wr_cycle[ 2345] = 1'b1;  addr_rom[ 2345]='h00000e44;  wr_data_rom[ 2345]='h00000a4a;
    rd_cycle[ 2346] = 1'b0;  wr_cycle[ 2346] = 1'b1;  addr_rom[ 2346]='h000015c4;  wr_data_rom[ 2346]='h00000981;
    rd_cycle[ 2347] = 1'b1;  wr_cycle[ 2347] = 1'b0;  addr_rom[ 2347]='h00000ba8;  wr_data_rom[ 2347]='h00000000;
    rd_cycle[ 2348] = 1'b0;  wr_cycle[ 2348] = 1'b1;  addr_rom[ 2348]='h00001698;  wr_data_rom[ 2348]='h00001c4f;
    rd_cycle[ 2349] = 1'b0;  wr_cycle[ 2349] = 1'b1;  addr_rom[ 2349]='h00000fd0;  wr_data_rom[ 2349]='h00001f37;
    rd_cycle[ 2350] = 1'b0;  wr_cycle[ 2350] = 1'b1;  addr_rom[ 2350]='h00000d4c;  wr_data_rom[ 2350]='h000018fb;
    rd_cycle[ 2351] = 1'b1;  wr_cycle[ 2351] = 1'b0;  addr_rom[ 2351]='h00001770;  wr_data_rom[ 2351]='h00000000;
    rd_cycle[ 2352] = 1'b1;  wr_cycle[ 2352] = 1'b0;  addr_rom[ 2352]='h00001ec0;  wr_data_rom[ 2352]='h00000000;
    rd_cycle[ 2353] = 1'b0;  wr_cycle[ 2353] = 1'b1;  addr_rom[ 2353]='h00001aec;  wr_data_rom[ 2353]='h000005df;
    rd_cycle[ 2354] = 1'b1;  wr_cycle[ 2354] = 1'b0;  addr_rom[ 2354]='h00000fe0;  wr_data_rom[ 2354]='h00000000;
    rd_cycle[ 2355] = 1'b0;  wr_cycle[ 2355] = 1'b1;  addr_rom[ 2355]='h00000b08;  wr_data_rom[ 2355]='h00000910;
    rd_cycle[ 2356] = 1'b0;  wr_cycle[ 2356] = 1'b1;  addr_rom[ 2356]='h00001178;  wr_data_rom[ 2356]='h00001600;
    rd_cycle[ 2357] = 1'b0;  wr_cycle[ 2357] = 1'b1;  addr_rom[ 2357]='h00000230;  wr_data_rom[ 2357]='h00001861;
    rd_cycle[ 2358] = 1'b0;  wr_cycle[ 2358] = 1'b1;  addr_rom[ 2358]='h00000b88;  wr_data_rom[ 2358]='h00001690;
    rd_cycle[ 2359] = 1'b1;  wr_cycle[ 2359] = 1'b0;  addr_rom[ 2359]='h000009bc;  wr_data_rom[ 2359]='h00000000;
    rd_cycle[ 2360] = 1'b0;  wr_cycle[ 2360] = 1'b1;  addr_rom[ 2360]='h00001e90;  wr_data_rom[ 2360]='h00001b1e;
    rd_cycle[ 2361] = 1'b0;  wr_cycle[ 2361] = 1'b1;  addr_rom[ 2361]='h00000630;  wr_data_rom[ 2361]='h00000405;
    rd_cycle[ 2362] = 1'b1;  wr_cycle[ 2362] = 1'b0;  addr_rom[ 2362]='h00001dc4;  wr_data_rom[ 2362]='h00000000;
    rd_cycle[ 2363] = 1'b1;  wr_cycle[ 2363] = 1'b0;  addr_rom[ 2363]='h00000014;  wr_data_rom[ 2363]='h00000000;
    rd_cycle[ 2364] = 1'b1;  wr_cycle[ 2364] = 1'b0;  addr_rom[ 2364]='h000004d8;  wr_data_rom[ 2364]='h00000000;
    rd_cycle[ 2365] = 1'b1;  wr_cycle[ 2365] = 1'b0;  addr_rom[ 2365]='h00000c20;  wr_data_rom[ 2365]='h00000000;
    rd_cycle[ 2366] = 1'b1;  wr_cycle[ 2366] = 1'b0;  addr_rom[ 2366]='h000011ec;  wr_data_rom[ 2366]='h00000000;
    rd_cycle[ 2367] = 1'b1;  wr_cycle[ 2367] = 1'b0;  addr_rom[ 2367]='h000006c0;  wr_data_rom[ 2367]='h00000000;
    rd_cycle[ 2368] = 1'b0;  wr_cycle[ 2368] = 1'b1;  addr_rom[ 2368]='h00001e58;  wr_data_rom[ 2368]='h000000e2;
    rd_cycle[ 2369] = 1'b0;  wr_cycle[ 2369] = 1'b1;  addr_rom[ 2369]='h00000134;  wr_data_rom[ 2369]='h00001605;
    rd_cycle[ 2370] = 1'b0;  wr_cycle[ 2370] = 1'b1;  addr_rom[ 2370]='h00001d54;  wr_data_rom[ 2370]='h000012a2;
    rd_cycle[ 2371] = 1'b1;  wr_cycle[ 2371] = 1'b0;  addr_rom[ 2371]='h00000e7c;  wr_data_rom[ 2371]='h00000000;
    rd_cycle[ 2372] = 1'b0;  wr_cycle[ 2372] = 1'b1;  addr_rom[ 2372]='h00000b74;  wr_data_rom[ 2372]='h00001be3;
    rd_cycle[ 2373] = 1'b1;  wr_cycle[ 2373] = 1'b0;  addr_rom[ 2373]='h00000240;  wr_data_rom[ 2373]='h00000000;
    rd_cycle[ 2374] = 1'b0;  wr_cycle[ 2374] = 1'b1;  addr_rom[ 2374]='h00000054;  wr_data_rom[ 2374]='h00000deb;
    rd_cycle[ 2375] = 1'b0;  wr_cycle[ 2375] = 1'b1;  addr_rom[ 2375]='h000009f0;  wr_data_rom[ 2375]='h0000151a;
    rd_cycle[ 2376] = 1'b1;  wr_cycle[ 2376] = 1'b0;  addr_rom[ 2376]='h00001d90;  wr_data_rom[ 2376]='h00000000;
    rd_cycle[ 2377] = 1'b0;  wr_cycle[ 2377] = 1'b1;  addr_rom[ 2377]='h000000e4;  wr_data_rom[ 2377]='h00001c3b;
    rd_cycle[ 2378] = 1'b0;  wr_cycle[ 2378] = 1'b1;  addr_rom[ 2378]='h00001bd0;  wr_data_rom[ 2378]='h000000f9;
    rd_cycle[ 2379] = 1'b0;  wr_cycle[ 2379] = 1'b1;  addr_rom[ 2379]='h0000065c;  wr_data_rom[ 2379]='h000002ce;
    rd_cycle[ 2380] = 1'b1;  wr_cycle[ 2380] = 1'b0;  addr_rom[ 2380]='h00000e78;  wr_data_rom[ 2380]='h00000000;
    rd_cycle[ 2381] = 1'b1;  wr_cycle[ 2381] = 1'b0;  addr_rom[ 2381]='h0000014c;  wr_data_rom[ 2381]='h00000000;
    rd_cycle[ 2382] = 1'b0;  wr_cycle[ 2382] = 1'b1;  addr_rom[ 2382]='h00000200;  wr_data_rom[ 2382]='h00000578;
    rd_cycle[ 2383] = 1'b0;  wr_cycle[ 2383] = 1'b1;  addr_rom[ 2383]='h00001174;  wr_data_rom[ 2383]='h0000141e;
    rd_cycle[ 2384] = 1'b1;  wr_cycle[ 2384] = 1'b0;  addr_rom[ 2384]='h00001d3c;  wr_data_rom[ 2384]='h00000000;
    rd_cycle[ 2385] = 1'b1;  wr_cycle[ 2385] = 1'b0;  addr_rom[ 2385]='h00001074;  wr_data_rom[ 2385]='h00000000;
    rd_cycle[ 2386] = 1'b1;  wr_cycle[ 2386] = 1'b0;  addr_rom[ 2386]='h00000eac;  wr_data_rom[ 2386]='h00000000;
    rd_cycle[ 2387] = 1'b0;  wr_cycle[ 2387] = 1'b1;  addr_rom[ 2387]='h00001574;  wr_data_rom[ 2387]='h00000247;
    rd_cycle[ 2388] = 1'b0;  wr_cycle[ 2388] = 1'b1;  addr_rom[ 2388]='h000007d8;  wr_data_rom[ 2388]='h0000170e;
    rd_cycle[ 2389] = 1'b1;  wr_cycle[ 2389] = 1'b0;  addr_rom[ 2389]='h0000057c;  wr_data_rom[ 2389]='h00000000;
    rd_cycle[ 2390] = 1'b0;  wr_cycle[ 2390] = 1'b1;  addr_rom[ 2390]='h00001434;  wr_data_rom[ 2390]='h000008a3;
    rd_cycle[ 2391] = 1'b1;  wr_cycle[ 2391] = 1'b0;  addr_rom[ 2391]='h00000870;  wr_data_rom[ 2391]='h00000000;
    rd_cycle[ 2392] = 1'b0;  wr_cycle[ 2392] = 1'b1;  addr_rom[ 2392]='h00000370;  wr_data_rom[ 2392]='h00001d17;
    rd_cycle[ 2393] = 1'b0;  wr_cycle[ 2393] = 1'b1;  addr_rom[ 2393]='h00000434;  wr_data_rom[ 2393]='h0000149b;
    rd_cycle[ 2394] = 1'b0;  wr_cycle[ 2394] = 1'b1;  addr_rom[ 2394]='h000019fc;  wr_data_rom[ 2394]='h00000f19;
    rd_cycle[ 2395] = 1'b0;  wr_cycle[ 2395] = 1'b1;  addr_rom[ 2395]='h000003a8;  wr_data_rom[ 2395]='h0000197e;
    rd_cycle[ 2396] = 1'b1;  wr_cycle[ 2396] = 1'b0;  addr_rom[ 2396]='h000000cc;  wr_data_rom[ 2396]='h00000000;
    rd_cycle[ 2397] = 1'b0;  wr_cycle[ 2397] = 1'b1;  addr_rom[ 2397]='h00001500;  wr_data_rom[ 2397]='h000009f8;
    rd_cycle[ 2398] = 1'b1;  wr_cycle[ 2398] = 1'b0;  addr_rom[ 2398]='h0000069c;  wr_data_rom[ 2398]='h00000000;
    rd_cycle[ 2399] = 1'b0;  wr_cycle[ 2399] = 1'b1;  addr_rom[ 2399]='h0000012c;  wr_data_rom[ 2399]='h00000b99;
    rd_cycle[ 2400] = 1'b0;  wr_cycle[ 2400] = 1'b1;  addr_rom[ 2400]='h0000108c;  wr_data_rom[ 2400]='h0000198b;
    rd_cycle[ 2401] = 1'b1;  wr_cycle[ 2401] = 1'b0;  addr_rom[ 2401]='h00000be8;  wr_data_rom[ 2401]='h00000000;
    rd_cycle[ 2402] = 1'b0;  wr_cycle[ 2402] = 1'b1;  addr_rom[ 2402]='h000010fc;  wr_data_rom[ 2402]='h00001852;
    rd_cycle[ 2403] = 1'b1;  wr_cycle[ 2403] = 1'b0;  addr_rom[ 2403]='h00001e94;  wr_data_rom[ 2403]='h00000000;
    rd_cycle[ 2404] = 1'b1;  wr_cycle[ 2404] = 1'b0;  addr_rom[ 2404]='h00001098;  wr_data_rom[ 2404]='h00000000;
    rd_cycle[ 2405] = 1'b0;  wr_cycle[ 2405] = 1'b1;  addr_rom[ 2405]='h00001948;  wr_data_rom[ 2405]='h000016f3;
    rd_cycle[ 2406] = 1'b1;  wr_cycle[ 2406] = 1'b0;  addr_rom[ 2406]='h00001694;  wr_data_rom[ 2406]='h00000000;
    rd_cycle[ 2407] = 1'b1;  wr_cycle[ 2407] = 1'b0;  addr_rom[ 2407]='h000017c0;  wr_data_rom[ 2407]='h00000000;
    rd_cycle[ 2408] = 1'b0;  wr_cycle[ 2408] = 1'b1;  addr_rom[ 2408]='h00001a0c;  wr_data_rom[ 2408]='h000013ea;
    rd_cycle[ 2409] = 1'b0;  wr_cycle[ 2409] = 1'b1;  addr_rom[ 2409]='h0000129c;  wr_data_rom[ 2409]='h00001f0a;
    rd_cycle[ 2410] = 1'b0;  wr_cycle[ 2410] = 1'b1;  addr_rom[ 2410]='h00000d8c;  wr_data_rom[ 2410]='h00001d5b;
    rd_cycle[ 2411] = 1'b1;  wr_cycle[ 2411] = 1'b0;  addr_rom[ 2411]='h000004a4;  wr_data_rom[ 2411]='h00000000;
    rd_cycle[ 2412] = 1'b0;  wr_cycle[ 2412] = 1'b1;  addr_rom[ 2412]='h00000540;  wr_data_rom[ 2412]='h00000b54;
    rd_cycle[ 2413] = 1'b0;  wr_cycle[ 2413] = 1'b1;  addr_rom[ 2413]='h00000ef4;  wr_data_rom[ 2413]='h000003ad;
    rd_cycle[ 2414] = 1'b1;  wr_cycle[ 2414] = 1'b0;  addr_rom[ 2414]='h000002f0;  wr_data_rom[ 2414]='h00000000;
    rd_cycle[ 2415] = 1'b1;  wr_cycle[ 2415] = 1'b0;  addr_rom[ 2415]='h00000cac;  wr_data_rom[ 2415]='h00000000;
    rd_cycle[ 2416] = 1'b0;  wr_cycle[ 2416] = 1'b1;  addr_rom[ 2416]='h00000d98;  wr_data_rom[ 2416]='h00000f07;
    rd_cycle[ 2417] = 1'b0;  wr_cycle[ 2417] = 1'b1;  addr_rom[ 2417]='h00000f90;  wr_data_rom[ 2417]='h00000166;
    rd_cycle[ 2418] = 1'b1;  wr_cycle[ 2418] = 1'b0;  addr_rom[ 2418]='h000007bc;  wr_data_rom[ 2418]='h00000000;
    rd_cycle[ 2419] = 1'b1;  wr_cycle[ 2419] = 1'b0;  addr_rom[ 2419]='h000015c8;  wr_data_rom[ 2419]='h00000000;
    rd_cycle[ 2420] = 1'b1;  wr_cycle[ 2420] = 1'b0;  addr_rom[ 2420]='h000015fc;  wr_data_rom[ 2420]='h00000000;
    rd_cycle[ 2421] = 1'b1;  wr_cycle[ 2421] = 1'b0;  addr_rom[ 2421]='h000005e8;  wr_data_rom[ 2421]='h00000000;
    rd_cycle[ 2422] = 1'b1;  wr_cycle[ 2422] = 1'b0;  addr_rom[ 2422]='h0000106c;  wr_data_rom[ 2422]='h00000000;
    rd_cycle[ 2423] = 1'b0;  wr_cycle[ 2423] = 1'b1;  addr_rom[ 2423]='h00001140;  wr_data_rom[ 2423]='h0000064d;
    rd_cycle[ 2424] = 1'b0;  wr_cycle[ 2424] = 1'b1;  addr_rom[ 2424]='h00001bec;  wr_data_rom[ 2424]='h00000cf2;
    rd_cycle[ 2425] = 1'b1;  wr_cycle[ 2425] = 1'b0;  addr_rom[ 2425]='h00000608;  wr_data_rom[ 2425]='h00000000;
    rd_cycle[ 2426] = 1'b0;  wr_cycle[ 2426] = 1'b1;  addr_rom[ 2426]='h000016f4;  wr_data_rom[ 2426]='h000013e8;
    rd_cycle[ 2427] = 1'b1;  wr_cycle[ 2427] = 1'b0;  addr_rom[ 2427]='h0000005c;  wr_data_rom[ 2427]='h00000000;
    rd_cycle[ 2428] = 1'b0;  wr_cycle[ 2428] = 1'b1;  addr_rom[ 2428]='h00000038;  wr_data_rom[ 2428]='h00000265;
    rd_cycle[ 2429] = 1'b1;  wr_cycle[ 2429] = 1'b0;  addr_rom[ 2429]='h00000fd0;  wr_data_rom[ 2429]='h00000000;
    rd_cycle[ 2430] = 1'b1;  wr_cycle[ 2430] = 1'b0;  addr_rom[ 2430]='h000004e4;  wr_data_rom[ 2430]='h00000000;
    rd_cycle[ 2431] = 1'b1;  wr_cycle[ 2431] = 1'b0;  addr_rom[ 2431]='h00001010;  wr_data_rom[ 2431]='h00000000;
    rd_cycle[ 2432] = 1'b1;  wr_cycle[ 2432] = 1'b0;  addr_rom[ 2432]='h00001c18;  wr_data_rom[ 2432]='h00000000;
    rd_cycle[ 2433] = 1'b1;  wr_cycle[ 2433] = 1'b0;  addr_rom[ 2433]='h00000d48;  wr_data_rom[ 2433]='h00000000;
    rd_cycle[ 2434] = 1'b1;  wr_cycle[ 2434] = 1'b0;  addr_rom[ 2434]='h00001168;  wr_data_rom[ 2434]='h00000000;
    rd_cycle[ 2435] = 1'b0;  wr_cycle[ 2435] = 1'b1;  addr_rom[ 2435]='h00001cd8;  wr_data_rom[ 2435]='h00000a85;
    rd_cycle[ 2436] = 1'b1;  wr_cycle[ 2436] = 1'b0;  addr_rom[ 2436]='h00000518;  wr_data_rom[ 2436]='h00000000;
    rd_cycle[ 2437] = 1'b1;  wr_cycle[ 2437] = 1'b0;  addr_rom[ 2437]='h000019e4;  wr_data_rom[ 2437]='h00000000;
    rd_cycle[ 2438] = 1'b0;  wr_cycle[ 2438] = 1'b1;  addr_rom[ 2438]='h00000c0c;  wr_data_rom[ 2438]='h00001d5b;
    rd_cycle[ 2439] = 1'b0;  wr_cycle[ 2439] = 1'b1;  addr_rom[ 2439]='h000004d8;  wr_data_rom[ 2439]='h00001a24;
    rd_cycle[ 2440] = 1'b1;  wr_cycle[ 2440] = 1'b0;  addr_rom[ 2440]='h00000fc8;  wr_data_rom[ 2440]='h00000000;
    rd_cycle[ 2441] = 1'b0;  wr_cycle[ 2441] = 1'b1;  addr_rom[ 2441]='h000013d8;  wr_data_rom[ 2441]='h00000204;
    rd_cycle[ 2442] = 1'b1;  wr_cycle[ 2442] = 1'b0;  addr_rom[ 2442]='h00000240;  wr_data_rom[ 2442]='h00000000;
    rd_cycle[ 2443] = 1'b0;  wr_cycle[ 2443] = 1'b1;  addr_rom[ 2443]='h000013e0;  wr_data_rom[ 2443]='h00000ce0;
    rd_cycle[ 2444] = 1'b0;  wr_cycle[ 2444] = 1'b1;  addr_rom[ 2444]='h00001180;  wr_data_rom[ 2444]='h00001a92;
    rd_cycle[ 2445] = 1'b1;  wr_cycle[ 2445] = 1'b0;  addr_rom[ 2445]='h00000500;  wr_data_rom[ 2445]='h00000000;
    rd_cycle[ 2446] = 1'b1;  wr_cycle[ 2446] = 1'b0;  addr_rom[ 2446]='h00001064;  wr_data_rom[ 2446]='h00000000;
    rd_cycle[ 2447] = 1'b1;  wr_cycle[ 2447] = 1'b0;  addr_rom[ 2447]='h00000ca0;  wr_data_rom[ 2447]='h00000000;
    rd_cycle[ 2448] = 1'b0;  wr_cycle[ 2448] = 1'b1;  addr_rom[ 2448]='h00001d30;  wr_data_rom[ 2448]='h00001428;
    rd_cycle[ 2449] = 1'b1;  wr_cycle[ 2449] = 1'b0;  addr_rom[ 2449]='h00001084;  wr_data_rom[ 2449]='h00000000;
    rd_cycle[ 2450] = 1'b1;  wr_cycle[ 2450] = 1'b0;  addr_rom[ 2450]='h000012f8;  wr_data_rom[ 2450]='h00000000;
    rd_cycle[ 2451] = 1'b1;  wr_cycle[ 2451] = 1'b0;  addr_rom[ 2451]='h000011e8;  wr_data_rom[ 2451]='h00000000;
    rd_cycle[ 2452] = 1'b0;  wr_cycle[ 2452] = 1'b1;  addr_rom[ 2452]='h000016bc;  wr_data_rom[ 2452]='h00000bd6;
    rd_cycle[ 2453] = 1'b0;  wr_cycle[ 2453] = 1'b1;  addr_rom[ 2453]='h0000087c;  wr_data_rom[ 2453]='h00001f16;
    rd_cycle[ 2454] = 1'b0;  wr_cycle[ 2454] = 1'b1;  addr_rom[ 2454]='h00001a14;  wr_data_rom[ 2454]='h000014a7;
    rd_cycle[ 2455] = 1'b1;  wr_cycle[ 2455] = 1'b0;  addr_rom[ 2455]='h00000408;  wr_data_rom[ 2455]='h00000000;
    rd_cycle[ 2456] = 1'b0;  wr_cycle[ 2456] = 1'b1;  addr_rom[ 2456]='h000018f8;  wr_data_rom[ 2456]='h0000150c;
    rd_cycle[ 2457] = 1'b1;  wr_cycle[ 2457] = 1'b0;  addr_rom[ 2457]='h00001728;  wr_data_rom[ 2457]='h00000000;
    rd_cycle[ 2458] = 1'b1;  wr_cycle[ 2458] = 1'b0;  addr_rom[ 2458]='h00000160;  wr_data_rom[ 2458]='h00000000;
    rd_cycle[ 2459] = 1'b0;  wr_cycle[ 2459] = 1'b1;  addr_rom[ 2459]='h00000aa4;  wr_data_rom[ 2459]='h0000061a;
    rd_cycle[ 2460] = 1'b1;  wr_cycle[ 2460] = 1'b0;  addr_rom[ 2460]='h00000e40;  wr_data_rom[ 2460]='h00000000;
    rd_cycle[ 2461] = 1'b0;  wr_cycle[ 2461] = 1'b1;  addr_rom[ 2461]='h000013c0;  wr_data_rom[ 2461]='h00000b88;
    rd_cycle[ 2462] = 1'b1;  wr_cycle[ 2462] = 1'b0;  addr_rom[ 2462]='h000004d4;  wr_data_rom[ 2462]='h00000000;
    rd_cycle[ 2463] = 1'b0;  wr_cycle[ 2463] = 1'b1;  addr_rom[ 2463]='h000007f8;  wr_data_rom[ 2463]='h000000f3;
    rd_cycle[ 2464] = 1'b0;  wr_cycle[ 2464] = 1'b1;  addr_rom[ 2464]='h00001538;  wr_data_rom[ 2464]='h00000830;
    rd_cycle[ 2465] = 1'b1;  wr_cycle[ 2465] = 1'b0;  addr_rom[ 2465]='h0000025c;  wr_data_rom[ 2465]='h00000000;
    rd_cycle[ 2466] = 1'b1;  wr_cycle[ 2466] = 1'b0;  addr_rom[ 2466]='h00000868;  wr_data_rom[ 2466]='h00000000;
    rd_cycle[ 2467] = 1'b0;  wr_cycle[ 2467] = 1'b1;  addr_rom[ 2467]='h00001b68;  wr_data_rom[ 2467]='h000005a6;
    rd_cycle[ 2468] = 1'b1;  wr_cycle[ 2468] = 1'b0;  addr_rom[ 2468]='h00000ea0;  wr_data_rom[ 2468]='h00000000;
    rd_cycle[ 2469] = 1'b0;  wr_cycle[ 2469] = 1'b1;  addr_rom[ 2469]='h000000e4;  wr_data_rom[ 2469]='h00001147;
    rd_cycle[ 2470] = 1'b0;  wr_cycle[ 2470] = 1'b1;  addr_rom[ 2470]='h00001070;  wr_data_rom[ 2470]='h00000556;
    rd_cycle[ 2471] = 1'b0;  wr_cycle[ 2471] = 1'b1;  addr_rom[ 2471]='h0000070c;  wr_data_rom[ 2471]='h00001e63;
    rd_cycle[ 2472] = 1'b0;  wr_cycle[ 2472] = 1'b1;  addr_rom[ 2472]='h00000ed0;  wr_data_rom[ 2472]='h000018af;
    rd_cycle[ 2473] = 1'b1;  wr_cycle[ 2473] = 1'b0;  addr_rom[ 2473]='h00001b78;  wr_data_rom[ 2473]='h00000000;
    rd_cycle[ 2474] = 1'b1;  wr_cycle[ 2474] = 1'b0;  addr_rom[ 2474]='h00001500;  wr_data_rom[ 2474]='h00000000;
    rd_cycle[ 2475] = 1'b0;  wr_cycle[ 2475] = 1'b1;  addr_rom[ 2475]='h00000f84;  wr_data_rom[ 2475]='h000012ee;
    rd_cycle[ 2476] = 1'b0;  wr_cycle[ 2476] = 1'b1;  addr_rom[ 2476]='h00000ab8;  wr_data_rom[ 2476]='h00000b76;
    rd_cycle[ 2477] = 1'b1;  wr_cycle[ 2477] = 1'b0;  addr_rom[ 2477]='h00000a78;  wr_data_rom[ 2477]='h00000000;
    rd_cycle[ 2478] = 1'b0;  wr_cycle[ 2478] = 1'b1;  addr_rom[ 2478]='h0000035c;  wr_data_rom[ 2478]='h0000158f;
    rd_cycle[ 2479] = 1'b1;  wr_cycle[ 2479] = 1'b0;  addr_rom[ 2479]='h00000b54;  wr_data_rom[ 2479]='h00000000;
    rd_cycle[ 2480] = 1'b1;  wr_cycle[ 2480] = 1'b0;  addr_rom[ 2480]='h00000fe8;  wr_data_rom[ 2480]='h00000000;
    rd_cycle[ 2481] = 1'b0;  wr_cycle[ 2481] = 1'b1;  addr_rom[ 2481]='h0000149c;  wr_data_rom[ 2481]='h00001a2f;
    rd_cycle[ 2482] = 1'b1;  wr_cycle[ 2482] = 1'b0;  addr_rom[ 2482]='h000014fc;  wr_data_rom[ 2482]='h00000000;
    rd_cycle[ 2483] = 1'b0;  wr_cycle[ 2483] = 1'b1;  addr_rom[ 2483]='h00001120;  wr_data_rom[ 2483]='h00001231;
    rd_cycle[ 2484] = 1'b0;  wr_cycle[ 2484] = 1'b1;  addr_rom[ 2484]='h00001b98;  wr_data_rom[ 2484]='h00001261;
    rd_cycle[ 2485] = 1'b0;  wr_cycle[ 2485] = 1'b1;  addr_rom[ 2485]='h00000c5c;  wr_data_rom[ 2485]='h0000139a;
    rd_cycle[ 2486] = 1'b1;  wr_cycle[ 2486] = 1'b0;  addr_rom[ 2486]='h000015e8;  wr_data_rom[ 2486]='h00000000;
    rd_cycle[ 2487] = 1'b0;  wr_cycle[ 2487] = 1'b1;  addr_rom[ 2487]='h00000d94;  wr_data_rom[ 2487]='h0000062f;
    rd_cycle[ 2488] = 1'b1;  wr_cycle[ 2488] = 1'b0;  addr_rom[ 2488]='h000007c0;  wr_data_rom[ 2488]='h00000000;
    rd_cycle[ 2489] = 1'b1;  wr_cycle[ 2489] = 1'b0;  addr_rom[ 2489]='h000002c0;  wr_data_rom[ 2489]='h00000000;
    rd_cycle[ 2490] = 1'b0;  wr_cycle[ 2490] = 1'b1;  addr_rom[ 2490]='h00001700;  wr_data_rom[ 2490]='h00001281;
    rd_cycle[ 2491] = 1'b1;  wr_cycle[ 2491] = 1'b0;  addr_rom[ 2491]='h00000338;  wr_data_rom[ 2491]='h00000000;
    rd_cycle[ 2492] = 1'b0;  wr_cycle[ 2492] = 1'b1;  addr_rom[ 2492]='h00001780;  wr_data_rom[ 2492]='h00000561;
    rd_cycle[ 2493] = 1'b1;  wr_cycle[ 2493] = 1'b0;  addr_rom[ 2493]='h00000150;  wr_data_rom[ 2493]='h00000000;
    rd_cycle[ 2494] = 1'b1;  wr_cycle[ 2494] = 1'b0;  addr_rom[ 2494]='h00001d50;  wr_data_rom[ 2494]='h00000000;
    rd_cycle[ 2495] = 1'b1;  wr_cycle[ 2495] = 1'b0;  addr_rom[ 2495]='h00000cd0;  wr_data_rom[ 2495]='h00000000;
    rd_cycle[ 2496] = 1'b0;  wr_cycle[ 2496] = 1'b1;  addr_rom[ 2496]='h00000d00;  wr_data_rom[ 2496]='h000005fe;
    rd_cycle[ 2497] = 1'b0;  wr_cycle[ 2497] = 1'b1;  addr_rom[ 2497]='h00001e9c;  wr_data_rom[ 2497]='h000016a6;
    rd_cycle[ 2498] = 1'b0;  wr_cycle[ 2498] = 1'b1;  addr_rom[ 2498]='h00000184;  wr_data_rom[ 2498]='h00001e6e;
    rd_cycle[ 2499] = 1'b1;  wr_cycle[ 2499] = 1'b0;  addr_rom[ 2499]='h00000450;  wr_data_rom[ 2499]='h00000000;
    rd_cycle[ 2500] = 1'b1;  wr_cycle[ 2500] = 1'b0;  addr_rom[ 2500]='h00000480;  wr_data_rom[ 2500]='h00000000;
    rd_cycle[ 2501] = 1'b1;  wr_cycle[ 2501] = 1'b0;  addr_rom[ 2501]='h00001a5c;  wr_data_rom[ 2501]='h00000000;
    rd_cycle[ 2502] = 1'b1;  wr_cycle[ 2502] = 1'b0;  addr_rom[ 2502]='h00001b9c;  wr_data_rom[ 2502]='h00000000;
    rd_cycle[ 2503] = 1'b1;  wr_cycle[ 2503] = 1'b0;  addr_rom[ 2503]='h00001f30;  wr_data_rom[ 2503]='h00000000;
    rd_cycle[ 2504] = 1'b1;  wr_cycle[ 2504] = 1'b0;  addr_rom[ 2504]='h0000138c;  wr_data_rom[ 2504]='h00000000;
    rd_cycle[ 2505] = 1'b0;  wr_cycle[ 2505] = 1'b1;  addr_rom[ 2505]='h00000b38;  wr_data_rom[ 2505]='h00000410;
    rd_cycle[ 2506] = 1'b0;  wr_cycle[ 2506] = 1'b1;  addr_rom[ 2506]='h0000030c;  wr_data_rom[ 2506]='h00001bc3;
    rd_cycle[ 2507] = 1'b1;  wr_cycle[ 2507] = 1'b0;  addr_rom[ 2507]='h0000094c;  wr_data_rom[ 2507]='h00000000;
    rd_cycle[ 2508] = 1'b0;  wr_cycle[ 2508] = 1'b1;  addr_rom[ 2508]='h0000178c;  wr_data_rom[ 2508]='h00001452;
    rd_cycle[ 2509] = 1'b0;  wr_cycle[ 2509] = 1'b1;  addr_rom[ 2509]='h000018a0;  wr_data_rom[ 2509]='h000019fc;
    rd_cycle[ 2510] = 1'b0;  wr_cycle[ 2510] = 1'b1;  addr_rom[ 2510]='h00001698;  wr_data_rom[ 2510]='h00001898;
    rd_cycle[ 2511] = 1'b1;  wr_cycle[ 2511] = 1'b0;  addr_rom[ 2511]='h00000c10;  wr_data_rom[ 2511]='h00000000;
    rd_cycle[ 2512] = 1'b0;  wr_cycle[ 2512] = 1'b1;  addr_rom[ 2512]='h000010d0;  wr_data_rom[ 2512]='h00001c1e;
    rd_cycle[ 2513] = 1'b0;  wr_cycle[ 2513] = 1'b1;  addr_rom[ 2513]='h00001b94;  wr_data_rom[ 2513]='h00001dc1;
    rd_cycle[ 2514] = 1'b1;  wr_cycle[ 2514] = 1'b0;  addr_rom[ 2514]='h00000668;  wr_data_rom[ 2514]='h00000000;
    rd_cycle[ 2515] = 1'b1;  wr_cycle[ 2515] = 1'b0;  addr_rom[ 2515]='h000008e4;  wr_data_rom[ 2515]='h00000000;
    rd_cycle[ 2516] = 1'b0;  wr_cycle[ 2516] = 1'b1;  addr_rom[ 2516]='h00001bcc;  wr_data_rom[ 2516]='h00000477;
    rd_cycle[ 2517] = 1'b0;  wr_cycle[ 2517] = 1'b1;  addr_rom[ 2517]='h000005a4;  wr_data_rom[ 2517]='h00000bcc;
    rd_cycle[ 2518] = 1'b0;  wr_cycle[ 2518] = 1'b1;  addr_rom[ 2518]='h000006d4;  wr_data_rom[ 2518]='h000002dd;
    rd_cycle[ 2519] = 1'b0;  wr_cycle[ 2519] = 1'b1;  addr_rom[ 2519]='h00001318;  wr_data_rom[ 2519]='h000003ea;
    rd_cycle[ 2520] = 1'b1;  wr_cycle[ 2520] = 1'b0;  addr_rom[ 2520]='h00001424;  wr_data_rom[ 2520]='h00000000;
    rd_cycle[ 2521] = 1'b1;  wr_cycle[ 2521] = 1'b0;  addr_rom[ 2521]='h00001358;  wr_data_rom[ 2521]='h00000000;
    rd_cycle[ 2522] = 1'b0;  wr_cycle[ 2522] = 1'b1;  addr_rom[ 2522]='h00001770;  wr_data_rom[ 2522]='h000003e2;
    rd_cycle[ 2523] = 1'b1;  wr_cycle[ 2523] = 1'b0;  addr_rom[ 2523]='h00001840;  wr_data_rom[ 2523]='h00000000;
    rd_cycle[ 2524] = 1'b1;  wr_cycle[ 2524] = 1'b0;  addr_rom[ 2524]='h000012f0;  wr_data_rom[ 2524]='h00000000;
    rd_cycle[ 2525] = 1'b0;  wr_cycle[ 2525] = 1'b1;  addr_rom[ 2525]='h00000dc0;  wr_data_rom[ 2525]='h000012d3;
    rd_cycle[ 2526] = 1'b1;  wr_cycle[ 2526] = 1'b0;  addr_rom[ 2526]='h000009e8;  wr_data_rom[ 2526]='h00000000;
    rd_cycle[ 2527] = 1'b1;  wr_cycle[ 2527] = 1'b0;  addr_rom[ 2527]='h0000088c;  wr_data_rom[ 2527]='h00000000;
    rd_cycle[ 2528] = 1'b0;  wr_cycle[ 2528] = 1'b1;  addr_rom[ 2528]='h0000087c;  wr_data_rom[ 2528]='h00001acf;
    rd_cycle[ 2529] = 1'b0;  wr_cycle[ 2529] = 1'b1;  addr_rom[ 2529]='h00001e9c;  wr_data_rom[ 2529]='h00000ca0;
    rd_cycle[ 2530] = 1'b0;  wr_cycle[ 2530] = 1'b1;  addr_rom[ 2530]='h00000524;  wr_data_rom[ 2530]='h0000144a;
    rd_cycle[ 2531] = 1'b1;  wr_cycle[ 2531] = 1'b0;  addr_rom[ 2531]='h00001428;  wr_data_rom[ 2531]='h00000000;
    rd_cycle[ 2532] = 1'b1;  wr_cycle[ 2532] = 1'b0;  addr_rom[ 2532]='h00000cc4;  wr_data_rom[ 2532]='h00000000;
    rd_cycle[ 2533] = 1'b1;  wr_cycle[ 2533] = 1'b0;  addr_rom[ 2533]='h00000ba4;  wr_data_rom[ 2533]='h00000000;
    rd_cycle[ 2534] = 1'b0;  wr_cycle[ 2534] = 1'b1;  addr_rom[ 2534]='h00001490;  wr_data_rom[ 2534]='h0000089d;
    rd_cycle[ 2535] = 1'b0;  wr_cycle[ 2535] = 1'b1;  addr_rom[ 2535]='h00000844;  wr_data_rom[ 2535]='h00001edb;
    rd_cycle[ 2536] = 1'b0;  wr_cycle[ 2536] = 1'b1;  addr_rom[ 2536]='h000016fc;  wr_data_rom[ 2536]='h00000d2e;
    rd_cycle[ 2537] = 1'b1;  wr_cycle[ 2537] = 1'b0;  addr_rom[ 2537]='h00001128;  wr_data_rom[ 2537]='h00000000;
    rd_cycle[ 2538] = 1'b0;  wr_cycle[ 2538] = 1'b1;  addr_rom[ 2538]='h00001e14;  wr_data_rom[ 2538]='h00000de2;
    rd_cycle[ 2539] = 1'b1;  wr_cycle[ 2539] = 1'b0;  addr_rom[ 2539]='h00001be8;  wr_data_rom[ 2539]='h00000000;
    rd_cycle[ 2540] = 1'b0;  wr_cycle[ 2540] = 1'b1;  addr_rom[ 2540]='h00000ccc;  wr_data_rom[ 2540]='h00000569;
    rd_cycle[ 2541] = 1'b0;  wr_cycle[ 2541] = 1'b1;  addr_rom[ 2541]='h00000d3c;  wr_data_rom[ 2541]='h00000906;
    rd_cycle[ 2542] = 1'b0;  wr_cycle[ 2542] = 1'b1;  addr_rom[ 2542]='h000009fc;  wr_data_rom[ 2542]='h000000dd;
    rd_cycle[ 2543] = 1'b1;  wr_cycle[ 2543] = 1'b0;  addr_rom[ 2543]='h000016b4;  wr_data_rom[ 2543]='h00000000;
    rd_cycle[ 2544] = 1'b1;  wr_cycle[ 2544] = 1'b0;  addr_rom[ 2544]='h00000f70;  wr_data_rom[ 2544]='h00000000;
    rd_cycle[ 2545] = 1'b0;  wr_cycle[ 2545] = 1'b1;  addr_rom[ 2545]='h0000040c;  wr_data_rom[ 2545]='h000007ea;
    rd_cycle[ 2546] = 1'b0;  wr_cycle[ 2546] = 1'b1;  addr_rom[ 2546]='h00001ee0;  wr_data_rom[ 2546]='h00000a0e;
    rd_cycle[ 2547] = 1'b1;  wr_cycle[ 2547] = 1'b0;  addr_rom[ 2547]='h00000448;  wr_data_rom[ 2547]='h00000000;
    rd_cycle[ 2548] = 1'b1;  wr_cycle[ 2548] = 1'b0;  addr_rom[ 2548]='h000001ac;  wr_data_rom[ 2548]='h00000000;
    rd_cycle[ 2549] = 1'b1;  wr_cycle[ 2549] = 1'b0;  addr_rom[ 2549]='h000004dc;  wr_data_rom[ 2549]='h00000000;
    rd_cycle[ 2550] = 1'b0;  wr_cycle[ 2550] = 1'b1;  addr_rom[ 2550]='h00000988;  wr_data_rom[ 2550]='h0000089f;
    rd_cycle[ 2551] = 1'b1;  wr_cycle[ 2551] = 1'b0;  addr_rom[ 2551]='h000013f8;  wr_data_rom[ 2551]='h00000000;
    rd_cycle[ 2552] = 1'b0;  wr_cycle[ 2552] = 1'b1;  addr_rom[ 2552]='h000013c0;  wr_data_rom[ 2552]='h00000655;
    rd_cycle[ 2553] = 1'b1;  wr_cycle[ 2553] = 1'b0;  addr_rom[ 2553]='h00001d98;  wr_data_rom[ 2553]='h00000000;
    rd_cycle[ 2554] = 1'b1;  wr_cycle[ 2554] = 1'b0;  addr_rom[ 2554]='h00000134;  wr_data_rom[ 2554]='h00000000;
    rd_cycle[ 2555] = 1'b0;  wr_cycle[ 2555] = 1'b1;  addr_rom[ 2555]='h00001cc0;  wr_data_rom[ 2555]='h00000faa;
    rd_cycle[ 2556] = 1'b0;  wr_cycle[ 2556] = 1'b1;  addr_rom[ 2556]='h0000178c;  wr_data_rom[ 2556]='h00000187;
    rd_cycle[ 2557] = 1'b0;  wr_cycle[ 2557] = 1'b1;  addr_rom[ 2557]='h000001a4;  wr_data_rom[ 2557]='h00000ea2;
    rd_cycle[ 2558] = 1'b1;  wr_cycle[ 2558] = 1'b0;  addr_rom[ 2558]='h00000dcc;  wr_data_rom[ 2558]='h00000000;
    rd_cycle[ 2559] = 1'b1;  wr_cycle[ 2559] = 1'b0;  addr_rom[ 2559]='h00001c38;  wr_data_rom[ 2559]='h00000000;
    rd_cycle[ 2560] = 1'b1;  wr_cycle[ 2560] = 1'b0;  addr_rom[ 2560]='h00001ca4;  wr_data_rom[ 2560]='h00000000;
    rd_cycle[ 2561] = 1'b0;  wr_cycle[ 2561] = 1'b1;  addr_rom[ 2561]='h00001958;  wr_data_rom[ 2561]='h00000b9b;
    rd_cycle[ 2562] = 1'b0;  wr_cycle[ 2562] = 1'b1;  addr_rom[ 2562]='h000009f0;  wr_data_rom[ 2562]='h0000165b;
    rd_cycle[ 2563] = 1'b0;  wr_cycle[ 2563] = 1'b1;  addr_rom[ 2563]='h0000029c;  wr_data_rom[ 2563]='h00001e5b;
    rd_cycle[ 2564] = 1'b1;  wr_cycle[ 2564] = 1'b0;  addr_rom[ 2564]='h00001880;  wr_data_rom[ 2564]='h00000000;
    rd_cycle[ 2565] = 1'b0;  wr_cycle[ 2565] = 1'b1;  addr_rom[ 2565]='h000006cc;  wr_data_rom[ 2565]='h00001cd7;
    rd_cycle[ 2566] = 1'b0;  wr_cycle[ 2566] = 1'b1;  addr_rom[ 2566]='h00000d68;  wr_data_rom[ 2566]='h00001155;
    rd_cycle[ 2567] = 1'b0;  wr_cycle[ 2567] = 1'b1;  addr_rom[ 2567]='h00000f44;  wr_data_rom[ 2567]='h00000af8;
    rd_cycle[ 2568] = 1'b0;  wr_cycle[ 2568] = 1'b1;  addr_rom[ 2568]='h00000aac;  wr_data_rom[ 2568]='h00001f39;
    rd_cycle[ 2569] = 1'b1;  wr_cycle[ 2569] = 1'b0;  addr_rom[ 2569]='h00001b84;  wr_data_rom[ 2569]='h00000000;
    rd_cycle[ 2570] = 1'b1;  wr_cycle[ 2570] = 1'b0;  addr_rom[ 2570]='h00001328;  wr_data_rom[ 2570]='h00000000;
    rd_cycle[ 2571] = 1'b1;  wr_cycle[ 2571] = 1'b0;  addr_rom[ 2571]='h00000f58;  wr_data_rom[ 2571]='h00000000;
    rd_cycle[ 2572] = 1'b1;  wr_cycle[ 2572] = 1'b0;  addr_rom[ 2572]='h00000b18;  wr_data_rom[ 2572]='h00000000;
    rd_cycle[ 2573] = 1'b1;  wr_cycle[ 2573] = 1'b0;  addr_rom[ 2573]='h00000458;  wr_data_rom[ 2573]='h00000000;
    rd_cycle[ 2574] = 1'b1;  wr_cycle[ 2574] = 1'b0;  addr_rom[ 2574]='h00000020;  wr_data_rom[ 2574]='h00000000;
    rd_cycle[ 2575] = 1'b0;  wr_cycle[ 2575] = 1'b1;  addr_rom[ 2575]='h00001874;  wr_data_rom[ 2575]='h00001d7a;
    rd_cycle[ 2576] = 1'b0;  wr_cycle[ 2576] = 1'b1;  addr_rom[ 2576]='h000000f0;  wr_data_rom[ 2576]='h000012de;
    rd_cycle[ 2577] = 1'b0;  wr_cycle[ 2577] = 1'b1;  addr_rom[ 2577]='h00000638;  wr_data_rom[ 2577]='h00001027;
    rd_cycle[ 2578] = 1'b1;  wr_cycle[ 2578] = 1'b0;  addr_rom[ 2578]='h000009ac;  wr_data_rom[ 2578]='h00000000;
    rd_cycle[ 2579] = 1'b1;  wr_cycle[ 2579] = 1'b0;  addr_rom[ 2579]='h00001294;  wr_data_rom[ 2579]='h00000000;
    rd_cycle[ 2580] = 1'b0;  wr_cycle[ 2580] = 1'b1;  addr_rom[ 2580]='h00000d8c;  wr_data_rom[ 2580]='h00001e5a;
    rd_cycle[ 2581] = 1'b1;  wr_cycle[ 2581] = 1'b0;  addr_rom[ 2581]='h0000080c;  wr_data_rom[ 2581]='h00000000;
    rd_cycle[ 2582] = 1'b0;  wr_cycle[ 2582] = 1'b1;  addr_rom[ 2582]='h000005d0;  wr_data_rom[ 2582]='h0000108b;
    rd_cycle[ 2583] = 1'b1;  wr_cycle[ 2583] = 1'b0;  addr_rom[ 2583]='h00000dc8;  wr_data_rom[ 2583]='h00000000;
    rd_cycle[ 2584] = 1'b1;  wr_cycle[ 2584] = 1'b0;  addr_rom[ 2584]='h00001898;  wr_data_rom[ 2584]='h00000000;
    rd_cycle[ 2585] = 1'b0;  wr_cycle[ 2585] = 1'b1;  addr_rom[ 2585]='h000002f8;  wr_data_rom[ 2585]='h00000d91;
    rd_cycle[ 2586] = 1'b0;  wr_cycle[ 2586] = 1'b1;  addr_rom[ 2586]='h000012a8;  wr_data_rom[ 2586]='h00001541;
    rd_cycle[ 2587] = 1'b1;  wr_cycle[ 2587] = 1'b0;  addr_rom[ 2587]='h0000008c;  wr_data_rom[ 2587]='h00000000;
    rd_cycle[ 2588] = 1'b0;  wr_cycle[ 2588] = 1'b1;  addr_rom[ 2588]='h00001c38;  wr_data_rom[ 2588]='h00001df5;
    rd_cycle[ 2589] = 1'b0;  wr_cycle[ 2589] = 1'b1;  addr_rom[ 2589]='h00000c90;  wr_data_rom[ 2589]='h00001a74;
    rd_cycle[ 2590] = 1'b0;  wr_cycle[ 2590] = 1'b1;  addr_rom[ 2590]='h000019dc;  wr_data_rom[ 2590]='h00000fe9;
    rd_cycle[ 2591] = 1'b0;  wr_cycle[ 2591] = 1'b1;  addr_rom[ 2591]='h00001408;  wr_data_rom[ 2591]='h000002a7;
    rd_cycle[ 2592] = 1'b1;  wr_cycle[ 2592] = 1'b0;  addr_rom[ 2592]='h00000058;  wr_data_rom[ 2592]='h00000000;
    rd_cycle[ 2593] = 1'b1;  wr_cycle[ 2593] = 1'b0;  addr_rom[ 2593]='h00001878;  wr_data_rom[ 2593]='h00000000;
    rd_cycle[ 2594] = 1'b1;  wr_cycle[ 2594] = 1'b0;  addr_rom[ 2594]='h00001910;  wr_data_rom[ 2594]='h00000000;
    rd_cycle[ 2595] = 1'b0;  wr_cycle[ 2595] = 1'b1;  addr_rom[ 2595]='h00001c04;  wr_data_rom[ 2595]='h00001d22;
    rd_cycle[ 2596] = 1'b1;  wr_cycle[ 2596] = 1'b0;  addr_rom[ 2596]='h00000ae4;  wr_data_rom[ 2596]='h00000000;
    rd_cycle[ 2597] = 1'b0;  wr_cycle[ 2597] = 1'b1;  addr_rom[ 2597]='h00000a10;  wr_data_rom[ 2597]='h00000fd4;
    rd_cycle[ 2598] = 1'b1;  wr_cycle[ 2598] = 1'b0;  addr_rom[ 2598]='h00001828;  wr_data_rom[ 2598]='h00000000;
    rd_cycle[ 2599] = 1'b1;  wr_cycle[ 2599] = 1'b0;  addr_rom[ 2599]='h000014a8;  wr_data_rom[ 2599]='h00000000;
    rd_cycle[ 2600] = 1'b1;  wr_cycle[ 2600] = 1'b0;  addr_rom[ 2600]='h0000192c;  wr_data_rom[ 2600]='h00000000;
    rd_cycle[ 2601] = 1'b0;  wr_cycle[ 2601] = 1'b1;  addr_rom[ 2601]='h00000984;  wr_data_rom[ 2601]='h00000f0c;
    rd_cycle[ 2602] = 1'b0;  wr_cycle[ 2602] = 1'b1;  addr_rom[ 2602]='h00001a44;  wr_data_rom[ 2602]='h00000a8d;
    rd_cycle[ 2603] = 1'b0;  wr_cycle[ 2603] = 1'b1;  addr_rom[ 2603]='h00001128;  wr_data_rom[ 2603]='h00000fdf;
    rd_cycle[ 2604] = 1'b1;  wr_cycle[ 2604] = 1'b0;  addr_rom[ 2604]='h00001e6c;  wr_data_rom[ 2604]='h00000000;
    rd_cycle[ 2605] = 1'b1;  wr_cycle[ 2605] = 1'b0;  addr_rom[ 2605]='h00001a78;  wr_data_rom[ 2605]='h00000000;
    rd_cycle[ 2606] = 1'b1;  wr_cycle[ 2606] = 1'b0;  addr_rom[ 2606]='h00000580;  wr_data_rom[ 2606]='h00000000;
    rd_cycle[ 2607] = 1'b0;  wr_cycle[ 2607] = 1'b1;  addr_rom[ 2607]='h00000cec;  wr_data_rom[ 2607]='h00000abb;
    rd_cycle[ 2608] = 1'b1;  wr_cycle[ 2608] = 1'b0;  addr_rom[ 2608]='h000013ec;  wr_data_rom[ 2608]='h00000000;
    rd_cycle[ 2609] = 1'b1;  wr_cycle[ 2609] = 1'b0;  addr_rom[ 2609]='h000003cc;  wr_data_rom[ 2609]='h00000000;
    rd_cycle[ 2610] = 1'b1;  wr_cycle[ 2610] = 1'b0;  addr_rom[ 2610]='h00000f54;  wr_data_rom[ 2610]='h00000000;
    rd_cycle[ 2611] = 1'b1;  wr_cycle[ 2611] = 1'b0;  addr_rom[ 2611]='h00001574;  wr_data_rom[ 2611]='h00000000;
    rd_cycle[ 2612] = 1'b0;  wr_cycle[ 2612] = 1'b1;  addr_rom[ 2612]='h00001cf8;  wr_data_rom[ 2612]='h000004d8;
    rd_cycle[ 2613] = 1'b0;  wr_cycle[ 2613] = 1'b1;  addr_rom[ 2613]='h00000e28;  wr_data_rom[ 2613]='h00000a77;
    rd_cycle[ 2614] = 1'b0;  wr_cycle[ 2614] = 1'b1;  addr_rom[ 2614]='h00001094;  wr_data_rom[ 2614]='h000007d4;
    rd_cycle[ 2615] = 1'b0;  wr_cycle[ 2615] = 1'b1;  addr_rom[ 2615]='h000003f8;  wr_data_rom[ 2615]='h000004cf;
    rd_cycle[ 2616] = 1'b0;  wr_cycle[ 2616] = 1'b1;  addr_rom[ 2616]='h00001454;  wr_data_rom[ 2616]='h00000eaa;
    rd_cycle[ 2617] = 1'b1;  wr_cycle[ 2617] = 1'b0;  addr_rom[ 2617]='h00001610;  wr_data_rom[ 2617]='h00000000;
    rd_cycle[ 2618] = 1'b0;  wr_cycle[ 2618] = 1'b1;  addr_rom[ 2618]='h00001460;  wr_data_rom[ 2618]='h0000009f;
    rd_cycle[ 2619] = 1'b0;  wr_cycle[ 2619] = 1'b1;  addr_rom[ 2619]='h00001a10;  wr_data_rom[ 2619]='h00000705;
    rd_cycle[ 2620] = 1'b0;  wr_cycle[ 2620] = 1'b1;  addr_rom[ 2620]='h0000144c;  wr_data_rom[ 2620]='h000000cd;
    rd_cycle[ 2621] = 1'b1;  wr_cycle[ 2621] = 1'b0;  addr_rom[ 2621]='h000010f8;  wr_data_rom[ 2621]='h00000000;
    rd_cycle[ 2622] = 1'b1;  wr_cycle[ 2622] = 1'b0;  addr_rom[ 2622]='h00001454;  wr_data_rom[ 2622]='h00000000;
    rd_cycle[ 2623] = 1'b0;  wr_cycle[ 2623] = 1'b1;  addr_rom[ 2623]='h00001e3c;  wr_data_rom[ 2623]='h00000014;
    rd_cycle[ 2624] = 1'b0;  wr_cycle[ 2624] = 1'b1;  addr_rom[ 2624]='h00000930;  wr_data_rom[ 2624]='h00000f0f;
    rd_cycle[ 2625] = 1'b0;  wr_cycle[ 2625] = 1'b1;  addr_rom[ 2625]='h000010d0;  wr_data_rom[ 2625]='h0000173a;
    rd_cycle[ 2626] = 1'b0;  wr_cycle[ 2626] = 1'b1;  addr_rom[ 2626]='h000019d4;  wr_data_rom[ 2626]='h00001069;
    rd_cycle[ 2627] = 1'b1;  wr_cycle[ 2627] = 1'b0;  addr_rom[ 2627]='h00001500;  wr_data_rom[ 2627]='h00000000;
    rd_cycle[ 2628] = 1'b1;  wr_cycle[ 2628] = 1'b0;  addr_rom[ 2628]='h00001574;  wr_data_rom[ 2628]='h00000000;
    rd_cycle[ 2629] = 1'b0;  wr_cycle[ 2629] = 1'b1;  addr_rom[ 2629]='h00001274;  wr_data_rom[ 2629]='h000017db;
    rd_cycle[ 2630] = 1'b0;  wr_cycle[ 2630] = 1'b1;  addr_rom[ 2630]='h00000f24;  wr_data_rom[ 2630]='h00001c59;
    rd_cycle[ 2631] = 1'b0;  wr_cycle[ 2631] = 1'b1;  addr_rom[ 2631]='h00001144;  wr_data_rom[ 2631]='h00001c6a;
    rd_cycle[ 2632] = 1'b0;  wr_cycle[ 2632] = 1'b1;  addr_rom[ 2632]='h00001944;  wr_data_rom[ 2632]='h00001211;
    rd_cycle[ 2633] = 1'b0;  wr_cycle[ 2633] = 1'b1;  addr_rom[ 2633]='h00001c84;  wr_data_rom[ 2633]='h00001d25;
    rd_cycle[ 2634] = 1'b0;  wr_cycle[ 2634] = 1'b1;  addr_rom[ 2634]='h000003ac;  wr_data_rom[ 2634]='h000015b4;
    rd_cycle[ 2635] = 1'b0;  wr_cycle[ 2635] = 1'b1;  addr_rom[ 2635]='h000008bc;  wr_data_rom[ 2635]='h000016df;
    rd_cycle[ 2636] = 1'b1;  wr_cycle[ 2636] = 1'b0;  addr_rom[ 2636]='h0000085c;  wr_data_rom[ 2636]='h00000000;
    rd_cycle[ 2637] = 1'b1;  wr_cycle[ 2637] = 1'b0;  addr_rom[ 2637]='h00000fb8;  wr_data_rom[ 2637]='h00000000;
    rd_cycle[ 2638] = 1'b0;  wr_cycle[ 2638] = 1'b1;  addr_rom[ 2638]='h00001b98;  wr_data_rom[ 2638]='h00000f23;
    rd_cycle[ 2639] = 1'b0;  wr_cycle[ 2639] = 1'b1;  addr_rom[ 2639]='h000011e8;  wr_data_rom[ 2639]='h00001e38;
    rd_cycle[ 2640] = 1'b0;  wr_cycle[ 2640] = 1'b1;  addr_rom[ 2640]='h00001ce8;  wr_data_rom[ 2640]='h000011ea;
    rd_cycle[ 2641] = 1'b0;  wr_cycle[ 2641] = 1'b1;  addr_rom[ 2641]='h00000690;  wr_data_rom[ 2641]='h00001ba2;
    rd_cycle[ 2642] = 1'b0;  wr_cycle[ 2642] = 1'b1;  addr_rom[ 2642]='h000004f4;  wr_data_rom[ 2642]='h000008f6;
    rd_cycle[ 2643] = 1'b1;  wr_cycle[ 2643] = 1'b0;  addr_rom[ 2643]='h00001e18;  wr_data_rom[ 2643]='h00000000;
    rd_cycle[ 2644] = 1'b0;  wr_cycle[ 2644] = 1'b1;  addr_rom[ 2644]='h000012f4;  wr_data_rom[ 2644]='h00001e76;
    rd_cycle[ 2645] = 1'b1;  wr_cycle[ 2645] = 1'b0;  addr_rom[ 2645]='h0000146c;  wr_data_rom[ 2645]='h00000000;
    rd_cycle[ 2646] = 1'b0;  wr_cycle[ 2646] = 1'b1;  addr_rom[ 2646]='h0000024c;  wr_data_rom[ 2646]='h000018cc;
    rd_cycle[ 2647] = 1'b0;  wr_cycle[ 2647] = 1'b1;  addr_rom[ 2647]='h00001be0;  wr_data_rom[ 2647]='h0000150f;
    rd_cycle[ 2648] = 1'b1;  wr_cycle[ 2648] = 1'b0;  addr_rom[ 2648]='h00001040;  wr_data_rom[ 2648]='h00000000;
    rd_cycle[ 2649] = 1'b1;  wr_cycle[ 2649] = 1'b0;  addr_rom[ 2649]='h00001784;  wr_data_rom[ 2649]='h00000000;
    rd_cycle[ 2650] = 1'b1;  wr_cycle[ 2650] = 1'b0;  addr_rom[ 2650]='h00001e60;  wr_data_rom[ 2650]='h00000000;
    rd_cycle[ 2651] = 1'b1;  wr_cycle[ 2651] = 1'b0;  addr_rom[ 2651]='h00001310;  wr_data_rom[ 2651]='h00000000;
    rd_cycle[ 2652] = 1'b0;  wr_cycle[ 2652] = 1'b1;  addr_rom[ 2652]='h00000e38;  wr_data_rom[ 2652]='h00000c98;
    rd_cycle[ 2653] = 1'b1;  wr_cycle[ 2653] = 1'b0;  addr_rom[ 2653]='h00001024;  wr_data_rom[ 2653]='h00000000;
    rd_cycle[ 2654] = 1'b0;  wr_cycle[ 2654] = 1'b1;  addr_rom[ 2654]='h00000ec0;  wr_data_rom[ 2654]='h0000035d;
    rd_cycle[ 2655] = 1'b1;  wr_cycle[ 2655] = 1'b0;  addr_rom[ 2655]='h000007a0;  wr_data_rom[ 2655]='h00000000;
    rd_cycle[ 2656] = 1'b1;  wr_cycle[ 2656] = 1'b0;  addr_rom[ 2656]='h000005e4;  wr_data_rom[ 2656]='h00000000;
    rd_cycle[ 2657] = 1'b0;  wr_cycle[ 2657] = 1'b1;  addr_rom[ 2657]='h00001060;  wr_data_rom[ 2657]='h000016fb;
    rd_cycle[ 2658] = 1'b1;  wr_cycle[ 2658] = 1'b0;  addr_rom[ 2658]='h00001958;  wr_data_rom[ 2658]='h00000000;
    rd_cycle[ 2659] = 1'b0;  wr_cycle[ 2659] = 1'b1;  addr_rom[ 2659]='h000015a4;  wr_data_rom[ 2659]='h00001c81;
    rd_cycle[ 2660] = 1'b0;  wr_cycle[ 2660] = 1'b1;  addr_rom[ 2660]='h000005e4;  wr_data_rom[ 2660]='h000007c9;
    rd_cycle[ 2661] = 1'b0;  wr_cycle[ 2661] = 1'b1;  addr_rom[ 2661]='h00001034;  wr_data_rom[ 2661]='h00001e9c;
    rd_cycle[ 2662] = 1'b1;  wr_cycle[ 2662] = 1'b0;  addr_rom[ 2662]='h000017d8;  wr_data_rom[ 2662]='h00000000;
    rd_cycle[ 2663] = 1'b1;  wr_cycle[ 2663] = 1'b0;  addr_rom[ 2663]='h00001834;  wr_data_rom[ 2663]='h00000000;
    rd_cycle[ 2664] = 1'b1;  wr_cycle[ 2664] = 1'b0;  addr_rom[ 2664]='h00001048;  wr_data_rom[ 2664]='h00000000;
    rd_cycle[ 2665] = 1'b1;  wr_cycle[ 2665] = 1'b0;  addr_rom[ 2665]='h00000db0;  wr_data_rom[ 2665]='h00000000;
    rd_cycle[ 2666] = 1'b0;  wr_cycle[ 2666] = 1'b1;  addr_rom[ 2666]='h00000bd8;  wr_data_rom[ 2666]='h00001078;
    rd_cycle[ 2667] = 1'b1;  wr_cycle[ 2667] = 1'b0;  addr_rom[ 2667]='h00001a8c;  wr_data_rom[ 2667]='h00000000;
    rd_cycle[ 2668] = 1'b1;  wr_cycle[ 2668] = 1'b0;  addr_rom[ 2668]='h00000d2c;  wr_data_rom[ 2668]='h00000000;
    rd_cycle[ 2669] = 1'b1;  wr_cycle[ 2669] = 1'b0;  addr_rom[ 2669]='h00000c54;  wr_data_rom[ 2669]='h00000000;
    rd_cycle[ 2670] = 1'b1;  wr_cycle[ 2670] = 1'b0;  addr_rom[ 2670]='h000013bc;  wr_data_rom[ 2670]='h00000000;
    rd_cycle[ 2671] = 1'b0;  wr_cycle[ 2671] = 1'b1;  addr_rom[ 2671]='h00001b84;  wr_data_rom[ 2671]='h0000096a;
    rd_cycle[ 2672] = 1'b0;  wr_cycle[ 2672] = 1'b1;  addr_rom[ 2672]='h00000d4c;  wr_data_rom[ 2672]='h0000104e;
    rd_cycle[ 2673] = 1'b0;  wr_cycle[ 2673] = 1'b1;  addr_rom[ 2673]='h000016c0;  wr_data_rom[ 2673]='h00000cde;
    rd_cycle[ 2674] = 1'b1;  wr_cycle[ 2674] = 1'b0;  addr_rom[ 2674]='h0000189c;  wr_data_rom[ 2674]='h00000000;
    rd_cycle[ 2675] = 1'b0;  wr_cycle[ 2675] = 1'b1;  addr_rom[ 2675]='h00001c0c;  wr_data_rom[ 2675]='h00001bf3;
    rd_cycle[ 2676] = 1'b1;  wr_cycle[ 2676] = 1'b0;  addr_rom[ 2676]='h000006bc;  wr_data_rom[ 2676]='h00000000;
    rd_cycle[ 2677] = 1'b1;  wr_cycle[ 2677] = 1'b0;  addr_rom[ 2677]='h000018ec;  wr_data_rom[ 2677]='h00000000;
    rd_cycle[ 2678] = 1'b0;  wr_cycle[ 2678] = 1'b1;  addr_rom[ 2678]='h000002fc;  wr_data_rom[ 2678]='h00001ab1;
    rd_cycle[ 2679] = 1'b1;  wr_cycle[ 2679] = 1'b0;  addr_rom[ 2679]='h000000b4;  wr_data_rom[ 2679]='h00000000;
    rd_cycle[ 2680] = 1'b1;  wr_cycle[ 2680] = 1'b0;  addr_rom[ 2680]='h00000048;  wr_data_rom[ 2680]='h00000000;
    rd_cycle[ 2681] = 1'b0;  wr_cycle[ 2681] = 1'b1;  addr_rom[ 2681]='h00001310;  wr_data_rom[ 2681]='h00001364;
    rd_cycle[ 2682] = 1'b0;  wr_cycle[ 2682] = 1'b1;  addr_rom[ 2682]='h000003f4;  wr_data_rom[ 2682]='h00001902;
    rd_cycle[ 2683] = 1'b1;  wr_cycle[ 2683] = 1'b0;  addr_rom[ 2683]='h00000c88;  wr_data_rom[ 2683]='h00000000;
    rd_cycle[ 2684] = 1'b0;  wr_cycle[ 2684] = 1'b1;  addr_rom[ 2684]='h000007d8;  wr_data_rom[ 2684]='h0000159d;
    rd_cycle[ 2685] = 1'b0;  wr_cycle[ 2685] = 1'b1;  addr_rom[ 2685]='h00001898;  wr_data_rom[ 2685]='h00001e00;
    rd_cycle[ 2686] = 1'b1;  wr_cycle[ 2686] = 1'b0;  addr_rom[ 2686]='h00000ed0;  wr_data_rom[ 2686]='h00000000;
    rd_cycle[ 2687] = 1'b1;  wr_cycle[ 2687] = 1'b0;  addr_rom[ 2687]='h00001c3c;  wr_data_rom[ 2687]='h00000000;
    rd_cycle[ 2688] = 1'b1;  wr_cycle[ 2688] = 1'b0;  addr_rom[ 2688]='h00000ce4;  wr_data_rom[ 2688]='h00000000;
    rd_cycle[ 2689] = 1'b1;  wr_cycle[ 2689] = 1'b0;  addr_rom[ 2689]='h00000dc0;  wr_data_rom[ 2689]='h00000000;
    rd_cycle[ 2690] = 1'b0;  wr_cycle[ 2690] = 1'b1;  addr_rom[ 2690]='h00000304;  wr_data_rom[ 2690]='h00000644;
    rd_cycle[ 2691] = 1'b1;  wr_cycle[ 2691] = 1'b0;  addr_rom[ 2691]='h00001e0c;  wr_data_rom[ 2691]='h00000000;
    rd_cycle[ 2692] = 1'b0;  wr_cycle[ 2692] = 1'b1;  addr_rom[ 2692]='h00001c84;  wr_data_rom[ 2692]='h00000f6c;
    rd_cycle[ 2693] = 1'b0;  wr_cycle[ 2693] = 1'b1;  addr_rom[ 2693]='h00000670;  wr_data_rom[ 2693]='h00001a80;
    rd_cycle[ 2694] = 1'b1;  wr_cycle[ 2694] = 1'b0;  addr_rom[ 2694]='h00001890;  wr_data_rom[ 2694]='h00000000;
    rd_cycle[ 2695] = 1'b0;  wr_cycle[ 2695] = 1'b1;  addr_rom[ 2695]='h00001c74;  wr_data_rom[ 2695]='h00000088;
    rd_cycle[ 2696] = 1'b0;  wr_cycle[ 2696] = 1'b1;  addr_rom[ 2696]='h000011e8;  wr_data_rom[ 2696]='h00001c07;
    rd_cycle[ 2697] = 1'b0;  wr_cycle[ 2697] = 1'b1;  addr_rom[ 2697]='h000008e8;  wr_data_rom[ 2697]='h00000107;
    rd_cycle[ 2698] = 1'b0;  wr_cycle[ 2698] = 1'b1;  addr_rom[ 2698]='h00001c80;  wr_data_rom[ 2698]='h00001dd7;
    rd_cycle[ 2699] = 1'b1;  wr_cycle[ 2699] = 1'b0;  addr_rom[ 2699]='h0000055c;  wr_data_rom[ 2699]='h00000000;
    rd_cycle[ 2700] = 1'b1;  wr_cycle[ 2700] = 1'b0;  addr_rom[ 2700]='h00001c1c;  wr_data_rom[ 2700]='h00000000;
    rd_cycle[ 2701] = 1'b1;  wr_cycle[ 2701] = 1'b0;  addr_rom[ 2701]='h00000a04;  wr_data_rom[ 2701]='h00000000;
    rd_cycle[ 2702] = 1'b0;  wr_cycle[ 2702] = 1'b1;  addr_rom[ 2702]='h000016b4;  wr_data_rom[ 2702]='h00000fad;
    rd_cycle[ 2703] = 1'b0;  wr_cycle[ 2703] = 1'b1;  addr_rom[ 2703]='h00000e6c;  wr_data_rom[ 2703]='h00000ac6;
    rd_cycle[ 2704] = 1'b1;  wr_cycle[ 2704] = 1'b0;  addr_rom[ 2704]='h00000948;  wr_data_rom[ 2704]='h00000000;
    rd_cycle[ 2705] = 1'b0;  wr_cycle[ 2705] = 1'b1;  addr_rom[ 2705]='h00000d38;  wr_data_rom[ 2705]='h00000921;
    rd_cycle[ 2706] = 1'b1;  wr_cycle[ 2706] = 1'b0;  addr_rom[ 2706]='h00001bbc;  wr_data_rom[ 2706]='h00000000;
    rd_cycle[ 2707] = 1'b0;  wr_cycle[ 2707] = 1'b1;  addr_rom[ 2707]='h0000029c;  wr_data_rom[ 2707]='h00000a82;
    rd_cycle[ 2708] = 1'b0;  wr_cycle[ 2708] = 1'b1;  addr_rom[ 2708]='h0000135c;  wr_data_rom[ 2708]='h00001637;
    rd_cycle[ 2709] = 1'b1;  wr_cycle[ 2709] = 1'b0;  addr_rom[ 2709]='h00000dc0;  wr_data_rom[ 2709]='h00000000;
    rd_cycle[ 2710] = 1'b0;  wr_cycle[ 2710] = 1'b1;  addr_rom[ 2710]='h0000029c;  wr_data_rom[ 2710]='h00000fb7;
    rd_cycle[ 2711] = 1'b1;  wr_cycle[ 2711] = 1'b0;  addr_rom[ 2711]='h00001558;  wr_data_rom[ 2711]='h00000000;
    rd_cycle[ 2712] = 1'b1;  wr_cycle[ 2712] = 1'b0;  addr_rom[ 2712]='h000008cc;  wr_data_rom[ 2712]='h00000000;
    rd_cycle[ 2713] = 1'b1;  wr_cycle[ 2713] = 1'b0;  addr_rom[ 2713]='h000002c8;  wr_data_rom[ 2713]='h00000000;
    rd_cycle[ 2714] = 1'b1;  wr_cycle[ 2714] = 1'b0;  addr_rom[ 2714]='h00001000;  wr_data_rom[ 2714]='h00000000;
    rd_cycle[ 2715] = 1'b0;  wr_cycle[ 2715] = 1'b1;  addr_rom[ 2715]='h00000280;  wr_data_rom[ 2715]='h00001abb;
    rd_cycle[ 2716] = 1'b1;  wr_cycle[ 2716] = 1'b0;  addr_rom[ 2716]='h0000195c;  wr_data_rom[ 2716]='h00000000;
    rd_cycle[ 2717] = 1'b1;  wr_cycle[ 2717] = 1'b0;  addr_rom[ 2717]='h000006e0;  wr_data_rom[ 2717]='h00000000;
    rd_cycle[ 2718] = 1'b0;  wr_cycle[ 2718] = 1'b1;  addr_rom[ 2718]='h000009d8;  wr_data_rom[ 2718]='h00000bac;
    rd_cycle[ 2719] = 1'b0;  wr_cycle[ 2719] = 1'b1;  addr_rom[ 2719]='h00000410;  wr_data_rom[ 2719]='h00001e8f;
    rd_cycle[ 2720] = 1'b1;  wr_cycle[ 2720] = 1'b0;  addr_rom[ 2720]='h00000e18;  wr_data_rom[ 2720]='h00000000;
    rd_cycle[ 2721] = 1'b0;  wr_cycle[ 2721] = 1'b1;  addr_rom[ 2721]='h00001c24;  wr_data_rom[ 2721]='h000018b4;
    rd_cycle[ 2722] = 1'b0;  wr_cycle[ 2722] = 1'b1;  addr_rom[ 2722]='h00001a44;  wr_data_rom[ 2722]='h000004c6;
    rd_cycle[ 2723] = 1'b0;  wr_cycle[ 2723] = 1'b1;  addr_rom[ 2723]='h00001d80;  wr_data_rom[ 2723]='h0000106e;
    rd_cycle[ 2724] = 1'b1;  wr_cycle[ 2724] = 1'b0;  addr_rom[ 2724]='h00001434;  wr_data_rom[ 2724]='h00000000;
    rd_cycle[ 2725] = 1'b0;  wr_cycle[ 2725] = 1'b1;  addr_rom[ 2725]='h00001328;  wr_data_rom[ 2725]='h00000d02;
    rd_cycle[ 2726] = 1'b1;  wr_cycle[ 2726] = 1'b0;  addr_rom[ 2726]='h000004c0;  wr_data_rom[ 2726]='h00000000;
    rd_cycle[ 2727] = 1'b0;  wr_cycle[ 2727] = 1'b1;  addr_rom[ 2727]='h000003a8;  wr_data_rom[ 2727]='h00001810;
    rd_cycle[ 2728] = 1'b1;  wr_cycle[ 2728] = 1'b0;  addr_rom[ 2728]='h00001c98;  wr_data_rom[ 2728]='h00000000;
    rd_cycle[ 2729] = 1'b1;  wr_cycle[ 2729] = 1'b0;  addr_rom[ 2729]='h00001814;  wr_data_rom[ 2729]='h00000000;
    rd_cycle[ 2730] = 1'b1;  wr_cycle[ 2730] = 1'b0;  addr_rom[ 2730]='h00000304;  wr_data_rom[ 2730]='h00000000;
    rd_cycle[ 2731] = 1'b0;  wr_cycle[ 2731] = 1'b1;  addr_rom[ 2731]='h00001e54;  wr_data_rom[ 2731]='h00000123;
    rd_cycle[ 2732] = 1'b1;  wr_cycle[ 2732] = 1'b0;  addr_rom[ 2732]='h00001cc4;  wr_data_rom[ 2732]='h00000000;
    rd_cycle[ 2733] = 1'b1;  wr_cycle[ 2733] = 1'b0;  addr_rom[ 2733]='h0000054c;  wr_data_rom[ 2733]='h00000000;
    rd_cycle[ 2734] = 1'b1;  wr_cycle[ 2734] = 1'b0;  addr_rom[ 2734]='h00001694;  wr_data_rom[ 2734]='h00000000;
    rd_cycle[ 2735] = 1'b0;  wr_cycle[ 2735] = 1'b1;  addr_rom[ 2735]='h00001394;  wr_data_rom[ 2735]='h00001bd9;
    rd_cycle[ 2736] = 1'b1;  wr_cycle[ 2736] = 1'b0;  addr_rom[ 2736]='h000011d0;  wr_data_rom[ 2736]='h00000000;
    rd_cycle[ 2737] = 1'b1;  wr_cycle[ 2737] = 1'b0;  addr_rom[ 2737]='h00001258;  wr_data_rom[ 2737]='h00000000;
    rd_cycle[ 2738] = 1'b0;  wr_cycle[ 2738] = 1'b1;  addr_rom[ 2738]='h00001314;  wr_data_rom[ 2738]='h00001ea6;
    rd_cycle[ 2739] = 1'b0;  wr_cycle[ 2739] = 1'b1;  addr_rom[ 2739]='h000006e0;  wr_data_rom[ 2739]='h00001166;
    rd_cycle[ 2740] = 1'b0;  wr_cycle[ 2740] = 1'b1;  addr_rom[ 2740]='h0000058c;  wr_data_rom[ 2740]='h00001f0e;
    rd_cycle[ 2741] = 1'b0;  wr_cycle[ 2741] = 1'b1;  addr_rom[ 2741]='h000012f4;  wr_data_rom[ 2741]='h00001963;
    rd_cycle[ 2742] = 1'b1;  wr_cycle[ 2742] = 1'b0;  addr_rom[ 2742]='h0000084c;  wr_data_rom[ 2742]='h00000000;
    rd_cycle[ 2743] = 1'b0;  wr_cycle[ 2743] = 1'b1;  addr_rom[ 2743]='h000007cc;  wr_data_rom[ 2743]='h00001395;
    rd_cycle[ 2744] = 1'b1;  wr_cycle[ 2744] = 1'b0;  addr_rom[ 2744]='h00001620;  wr_data_rom[ 2744]='h00000000;
    rd_cycle[ 2745] = 1'b1;  wr_cycle[ 2745] = 1'b0;  addr_rom[ 2745]='h00001154;  wr_data_rom[ 2745]='h00000000;
    rd_cycle[ 2746] = 1'b0;  wr_cycle[ 2746] = 1'b1;  addr_rom[ 2746]='h00000dbc;  wr_data_rom[ 2746]='h0000021a;
    rd_cycle[ 2747] = 1'b1;  wr_cycle[ 2747] = 1'b0;  addr_rom[ 2747]='h00001e14;  wr_data_rom[ 2747]='h00000000;
    rd_cycle[ 2748] = 1'b0;  wr_cycle[ 2748] = 1'b1;  addr_rom[ 2748]='h0000111c;  wr_data_rom[ 2748]='h000019f4;
    rd_cycle[ 2749] = 1'b0;  wr_cycle[ 2749] = 1'b1;  addr_rom[ 2749]='h000005b4;  wr_data_rom[ 2749]='h00001587;
    rd_cycle[ 2750] = 1'b1;  wr_cycle[ 2750] = 1'b0;  addr_rom[ 2750]='h00000ab4;  wr_data_rom[ 2750]='h00000000;
    rd_cycle[ 2751] = 1'b1;  wr_cycle[ 2751] = 1'b0;  addr_rom[ 2751]='h00000c44;  wr_data_rom[ 2751]='h00000000;
    rd_cycle[ 2752] = 1'b0;  wr_cycle[ 2752] = 1'b1;  addr_rom[ 2752]='h000003cc;  wr_data_rom[ 2752]='h0000173d;
    rd_cycle[ 2753] = 1'b0;  wr_cycle[ 2753] = 1'b1;  addr_rom[ 2753]='h00001e94;  wr_data_rom[ 2753]='h00001642;
    rd_cycle[ 2754] = 1'b0;  wr_cycle[ 2754] = 1'b1;  addr_rom[ 2754]='h0000100c;  wr_data_rom[ 2754]='h00000baf;
    rd_cycle[ 2755] = 1'b1;  wr_cycle[ 2755] = 1'b0;  addr_rom[ 2755]='h00000848;  wr_data_rom[ 2755]='h00000000;
    rd_cycle[ 2756] = 1'b0;  wr_cycle[ 2756] = 1'b1;  addr_rom[ 2756]='h00000d54;  wr_data_rom[ 2756]='h00000c25;
    rd_cycle[ 2757] = 1'b1;  wr_cycle[ 2757] = 1'b0;  addr_rom[ 2757]='h000013bc;  wr_data_rom[ 2757]='h00000000;
    rd_cycle[ 2758] = 1'b1;  wr_cycle[ 2758] = 1'b0;  addr_rom[ 2758]='h000014cc;  wr_data_rom[ 2758]='h00000000;
    rd_cycle[ 2759] = 1'b1;  wr_cycle[ 2759] = 1'b0;  addr_rom[ 2759]='h00001594;  wr_data_rom[ 2759]='h00000000;
    rd_cycle[ 2760] = 1'b1;  wr_cycle[ 2760] = 1'b0;  addr_rom[ 2760]='h00000594;  wr_data_rom[ 2760]='h00000000;
    rd_cycle[ 2761] = 1'b0;  wr_cycle[ 2761] = 1'b1;  addr_rom[ 2761]='h00001afc;  wr_data_rom[ 2761]='h000016f7;
    rd_cycle[ 2762] = 1'b0;  wr_cycle[ 2762] = 1'b1;  addr_rom[ 2762]='h00000400;  wr_data_rom[ 2762]='h00000541;
    rd_cycle[ 2763] = 1'b1;  wr_cycle[ 2763] = 1'b0;  addr_rom[ 2763]='h00000790;  wr_data_rom[ 2763]='h00000000;
    rd_cycle[ 2764] = 1'b0;  wr_cycle[ 2764] = 1'b1;  addr_rom[ 2764]='h000001d0;  wr_data_rom[ 2764]='h00001dcc;
    rd_cycle[ 2765] = 1'b1;  wr_cycle[ 2765] = 1'b0;  addr_rom[ 2765]='h0000088c;  wr_data_rom[ 2765]='h00000000;
    rd_cycle[ 2766] = 1'b0;  wr_cycle[ 2766] = 1'b1;  addr_rom[ 2766]='h00001a5c;  wr_data_rom[ 2766]='h00000341;
    rd_cycle[ 2767] = 1'b0;  wr_cycle[ 2767] = 1'b1;  addr_rom[ 2767]='h00000d3c;  wr_data_rom[ 2767]='h00001ce0;
    rd_cycle[ 2768] = 1'b1;  wr_cycle[ 2768] = 1'b0;  addr_rom[ 2768]='h000014e8;  wr_data_rom[ 2768]='h00000000;
    rd_cycle[ 2769] = 1'b0;  wr_cycle[ 2769] = 1'b1;  addr_rom[ 2769]='h00001d94;  wr_data_rom[ 2769]='h00001f11;
    rd_cycle[ 2770] = 1'b0;  wr_cycle[ 2770] = 1'b1;  addr_rom[ 2770]='h00001530;  wr_data_rom[ 2770]='h00001b03;
    rd_cycle[ 2771] = 1'b1;  wr_cycle[ 2771] = 1'b0;  addr_rom[ 2771]='h0000149c;  wr_data_rom[ 2771]='h00000000;
    rd_cycle[ 2772] = 1'b0;  wr_cycle[ 2772] = 1'b1;  addr_rom[ 2772]='h00000fa4;  wr_data_rom[ 2772]='h000003d6;
    rd_cycle[ 2773] = 1'b1;  wr_cycle[ 2773] = 1'b0;  addr_rom[ 2773]='h00001e88;  wr_data_rom[ 2773]='h00000000;
    rd_cycle[ 2774] = 1'b0;  wr_cycle[ 2774] = 1'b1;  addr_rom[ 2774]='h00000078;  wr_data_rom[ 2774]='h0000036a;
    rd_cycle[ 2775] = 1'b0;  wr_cycle[ 2775] = 1'b1;  addr_rom[ 2775]='h000016fc;  wr_data_rom[ 2775]='h00001098;
    rd_cycle[ 2776] = 1'b0;  wr_cycle[ 2776] = 1'b1;  addr_rom[ 2776]='h0000079c;  wr_data_rom[ 2776]='h00000d06;
    rd_cycle[ 2777] = 1'b1;  wr_cycle[ 2777] = 1'b0;  addr_rom[ 2777]='h0000066c;  wr_data_rom[ 2777]='h00000000;
    rd_cycle[ 2778] = 1'b1;  wr_cycle[ 2778] = 1'b0;  addr_rom[ 2778]='h000015cc;  wr_data_rom[ 2778]='h00000000;
    rd_cycle[ 2779] = 1'b1;  wr_cycle[ 2779] = 1'b0;  addr_rom[ 2779]='h0000143c;  wr_data_rom[ 2779]='h00000000;
    rd_cycle[ 2780] = 1'b0;  wr_cycle[ 2780] = 1'b1;  addr_rom[ 2780]='h00000974;  wr_data_rom[ 2780]='h00000dc9;
    rd_cycle[ 2781] = 1'b0;  wr_cycle[ 2781] = 1'b1;  addr_rom[ 2781]='h00000780;  wr_data_rom[ 2781]='h00000d39;
    rd_cycle[ 2782] = 1'b1;  wr_cycle[ 2782] = 1'b0;  addr_rom[ 2782]='h00000bbc;  wr_data_rom[ 2782]='h00000000;
    rd_cycle[ 2783] = 1'b0;  wr_cycle[ 2783] = 1'b1;  addr_rom[ 2783]='h00000fd8;  wr_data_rom[ 2783]='h00000619;
    rd_cycle[ 2784] = 1'b1;  wr_cycle[ 2784] = 1'b0;  addr_rom[ 2784]='h0000145c;  wr_data_rom[ 2784]='h00000000;
    rd_cycle[ 2785] = 1'b0;  wr_cycle[ 2785] = 1'b1;  addr_rom[ 2785]='h00001a20;  wr_data_rom[ 2785]='h00000b64;
    rd_cycle[ 2786] = 1'b1;  wr_cycle[ 2786] = 1'b0;  addr_rom[ 2786]='h00000dbc;  wr_data_rom[ 2786]='h00000000;
    rd_cycle[ 2787] = 1'b0;  wr_cycle[ 2787] = 1'b1;  addr_rom[ 2787]='h00001874;  wr_data_rom[ 2787]='h00000349;
    rd_cycle[ 2788] = 1'b1;  wr_cycle[ 2788] = 1'b0;  addr_rom[ 2788]='h0000190c;  wr_data_rom[ 2788]='h00000000;
    rd_cycle[ 2789] = 1'b0;  wr_cycle[ 2789] = 1'b1;  addr_rom[ 2789]='h00000b00;  wr_data_rom[ 2789]='h0000158e;
    rd_cycle[ 2790] = 1'b0;  wr_cycle[ 2790] = 1'b1;  addr_rom[ 2790]='h000014b0;  wr_data_rom[ 2790]='h000009fe;
    rd_cycle[ 2791] = 1'b0;  wr_cycle[ 2791] = 1'b1;  addr_rom[ 2791]='h0000044c;  wr_data_rom[ 2791]='h0000058f;
    rd_cycle[ 2792] = 1'b1;  wr_cycle[ 2792] = 1'b0;  addr_rom[ 2792]='h00001198;  wr_data_rom[ 2792]='h00000000;
    rd_cycle[ 2793] = 1'b1;  wr_cycle[ 2793] = 1'b0;  addr_rom[ 2793]='h00000ebc;  wr_data_rom[ 2793]='h00000000;
    rd_cycle[ 2794] = 1'b0;  wr_cycle[ 2794] = 1'b1;  addr_rom[ 2794]='h00001398;  wr_data_rom[ 2794]='h000010db;
    rd_cycle[ 2795] = 1'b0;  wr_cycle[ 2795] = 1'b1;  addr_rom[ 2795]='h000019c4;  wr_data_rom[ 2795]='h00000181;
    rd_cycle[ 2796] = 1'b1;  wr_cycle[ 2796] = 1'b0;  addr_rom[ 2796]='h00000068;  wr_data_rom[ 2796]='h00000000;
    rd_cycle[ 2797] = 1'b0;  wr_cycle[ 2797] = 1'b1;  addr_rom[ 2797]='h000018d8;  wr_data_rom[ 2797]='h0000160b;
    rd_cycle[ 2798] = 1'b1;  wr_cycle[ 2798] = 1'b0;  addr_rom[ 2798]='h00000544;  wr_data_rom[ 2798]='h00000000;
    rd_cycle[ 2799] = 1'b1;  wr_cycle[ 2799] = 1'b0;  addr_rom[ 2799]='h000004d8;  wr_data_rom[ 2799]='h00000000;
    rd_cycle[ 2800] = 1'b0;  wr_cycle[ 2800] = 1'b1;  addr_rom[ 2800]='h00001464;  wr_data_rom[ 2800]='h00001d89;
    rd_cycle[ 2801] = 1'b1;  wr_cycle[ 2801] = 1'b0;  addr_rom[ 2801]='h00001ab4;  wr_data_rom[ 2801]='h00000000;
    rd_cycle[ 2802] = 1'b0;  wr_cycle[ 2802] = 1'b1;  addr_rom[ 2802]='h0000041c;  wr_data_rom[ 2802]='h000019ce;
    rd_cycle[ 2803] = 1'b1;  wr_cycle[ 2803] = 1'b0;  addr_rom[ 2803]='h00001010;  wr_data_rom[ 2803]='h00000000;
    rd_cycle[ 2804] = 1'b1;  wr_cycle[ 2804] = 1'b0;  addr_rom[ 2804]='h00000188;  wr_data_rom[ 2804]='h00000000;
    rd_cycle[ 2805] = 1'b0;  wr_cycle[ 2805] = 1'b1;  addr_rom[ 2805]='h00001108;  wr_data_rom[ 2805]='h000008ae;
    rd_cycle[ 2806] = 1'b0;  wr_cycle[ 2806] = 1'b1;  addr_rom[ 2806]='h00000258;  wr_data_rom[ 2806]='h0000169e;
    rd_cycle[ 2807] = 1'b1;  wr_cycle[ 2807] = 1'b0;  addr_rom[ 2807]='h000015e0;  wr_data_rom[ 2807]='h00000000;
    rd_cycle[ 2808] = 1'b1;  wr_cycle[ 2808] = 1'b0;  addr_rom[ 2808]='h000017e0;  wr_data_rom[ 2808]='h00000000;
    rd_cycle[ 2809] = 1'b0;  wr_cycle[ 2809] = 1'b1;  addr_rom[ 2809]='h000013b8;  wr_data_rom[ 2809]='h00000ad4;
    rd_cycle[ 2810] = 1'b1;  wr_cycle[ 2810] = 1'b0;  addr_rom[ 2810]='h0000067c;  wr_data_rom[ 2810]='h00000000;
    rd_cycle[ 2811] = 1'b0;  wr_cycle[ 2811] = 1'b1;  addr_rom[ 2811]='h00001e7c;  wr_data_rom[ 2811]='h00000edd;
    rd_cycle[ 2812] = 1'b0;  wr_cycle[ 2812] = 1'b1;  addr_rom[ 2812]='h00001780;  wr_data_rom[ 2812]='h000010f7;
    rd_cycle[ 2813] = 1'b0;  wr_cycle[ 2813] = 1'b1;  addr_rom[ 2813]='h000014b8;  wr_data_rom[ 2813]='h00001a49;
    rd_cycle[ 2814] = 1'b1;  wr_cycle[ 2814] = 1'b0;  addr_rom[ 2814]='h000002f8;  wr_data_rom[ 2814]='h00000000;
    rd_cycle[ 2815] = 1'b0;  wr_cycle[ 2815] = 1'b1;  addr_rom[ 2815]='h00001130;  wr_data_rom[ 2815]='h000001df;
    rd_cycle[ 2816] = 1'b0;  wr_cycle[ 2816] = 1'b1;  addr_rom[ 2816]='h0000072c;  wr_data_rom[ 2816]='h00001c05;
    rd_cycle[ 2817] = 1'b1;  wr_cycle[ 2817] = 1'b0;  addr_rom[ 2817]='h00001254;  wr_data_rom[ 2817]='h00000000;
    rd_cycle[ 2818] = 1'b1;  wr_cycle[ 2818] = 1'b0;  addr_rom[ 2818]='h00000f04;  wr_data_rom[ 2818]='h00000000;
    rd_cycle[ 2819] = 1'b0;  wr_cycle[ 2819] = 1'b1;  addr_rom[ 2819]='h00001ef8;  wr_data_rom[ 2819]='h000005d3;
    rd_cycle[ 2820] = 1'b1;  wr_cycle[ 2820] = 1'b0;  addr_rom[ 2820]='h00000e64;  wr_data_rom[ 2820]='h00000000;
    rd_cycle[ 2821] = 1'b0;  wr_cycle[ 2821] = 1'b1;  addr_rom[ 2821]='h0000073c;  wr_data_rom[ 2821]='h00001361;
    rd_cycle[ 2822] = 1'b0;  wr_cycle[ 2822] = 1'b1;  addr_rom[ 2822]='h00001cc4;  wr_data_rom[ 2822]='h0000147d;
    rd_cycle[ 2823] = 1'b0;  wr_cycle[ 2823] = 1'b1;  addr_rom[ 2823]='h000012a4;  wr_data_rom[ 2823]='h00000af4;
    rd_cycle[ 2824] = 1'b1;  wr_cycle[ 2824] = 1'b0;  addr_rom[ 2824]='h00000d58;  wr_data_rom[ 2824]='h00000000;
    rd_cycle[ 2825] = 1'b1;  wr_cycle[ 2825] = 1'b0;  addr_rom[ 2825]='h000011b0;  wr_data_rom[ 2825]='h00000000;
    rd_cycle[ 2826] = 1'b1;  wr_cycle[ 2826] = 1'b0;  addr_rom[ 2826]='h00000078;  wr_data_rom[ 2826]='h00000000;
    rd_cycle[ 2827] = 1'b1;  wr_cycle[ 2827] = 1'b0;  addr_rom[ 2827]='h00001cbc;  wr_data_rom[ 2827]='h00000000;
    rd_cycle[ 2828] = 1'b0;  wr_cycle[ 2828] = 1'b1;  addr_rom[ 2828]='h00001bb8;  wr_data_rom[ 2828]='h000002a7;
    rd_cycle[ 2829] = 1'b1;  wr_cycle[ 2829] = 1'b0;  addr_rom[ 2829]='h00001d08;  wr_data_rom[ 2829]='h00000000;
    rd_cycle[ 2830] = 1'b0;  wr_cycle[ 2830] = 1'b1;  addr_rom[ 2830]='h00000840;  wr_data_rom[ 2830]='h0000127c;
    rd_cycle[ 2831] = 1'b1;  wr_cycle[ 2831] = 1'b0;  addr_rom[ 2831]='h00001aa8;  wr_data_rom[ 2831]='h00000000;
    rd_cycle[ 2832] = 1'b1;  wr_cycle[ 2832] = 1'b0;  addr_rom[ 2832]='h00001194;  wr_data_rom[ 2832]='h00000000;
    rd_cycle[ 2833] = 1'b1;  wr_cycle[ 2833] = 1'b0;  addr_rom[ 2833]='h00000004;  wr_data_rom[ 2833]='h00000000;
    rd_cycle[ 2834] = 1'b1;  wr_cycle[ 2834] = 1'b0;  addr_rom[ 2834]='h00001eb4;  wr_data_rom[ 2834]='h00000000;
    rd_cycle[ 2835] = 1'b1;  wr_cycle[ 2835] = 1'b0;  addr_rom[ 2835]='h000008bc;  wr_data_rom[ 2835]='h00000000;
    rd_cycle[ 2836] = 1'b1;  wr_cycle[ 2836] = 1'b0;  addr_rom[ 2836]='h00001040;  wr_data_rom[ 2836]='h00000000;
    rd_cycle[ 2837] = 1'b0;  wr_cycle[ 2837] = 1'b1;  addr_rom[ 2837]='h00001a50;  wr_data_rom[ 2837]='h00000e16;
    rd_cycle[ 2838] = 1'b0;  wr_cycle[ 2838] = 1'b1;  addr_rom[ 2838]='h000007ac;  wr_data_rom[ 2838]='h00001ace;
    rd_cycle[ 2839] = 1'b1;  wr_cycle[ 2839] = 1'b0;  addr_rom[ 2839]='h000008a0;  wr_data_rom[ 2839]='h00000000;
    rd_cycle[ 2840] = 1'b1;  wr_cycle[ 2840] = 1'b0;  addr_rom[ 2840]='h00001664;  wr_data_rom[ 2840]='h00000000;
    rd_cycle[ 2841] = 1'b0;  wr_cycle[ 2841] = 1'b1;  addr_rom[ 2841]='h00000d48;  wr_data_rom[ 2841]='h00001b87;
    rd_cycle[ 2842] = 1'b0;  wr_cycle[ 2842] = 1'b1;  addr_rom[ 2842]='h00001d44;  wr_data_rom[ 2842]='h00000e43;
    rd_cycle[ 2843] = 1'b0;  wr_cycle[ 2843] = 1'b1;  addr_rom[ 2843]='h00001278;  wr_data_rom[ 2843]='h00000bd8;
    rd_cycle[ 2844] = 1'b0;  wr_cycle[ 2844] = 1'b1;  addr_rom[ 2844]='h000010b8;  wr_data_rom[ 2844]='h00001aa4;
    rd_cycle[ 2845] = 1'b1;  wr_cycle[ 2845] = 1'b0;  addr_rom[ 2845]='h00000138;  wr_data_rom[ 2845]='h00000000;
    rd_cycle[ 2846] = 1'b0;  wr_cycle[ 2846] = 1'b1;  addr_rom[ 2846]='h00000310;  wr_data_rom[ 2846]='h0000019b;
    rd_cycle[ 2847] = 1'b0;  wr_cycle[ 2847] = 1'b1;  addr_rom[ 2847]='h00000f10;  wr_data_rom[ 2847]='h00000a8d;
    rd_cycle[ 2848] = 1'b0;  wr_cycle[ 2848] = 1'b1;  addr_rom[ 2848]='h00000b68;  wr_data_rom[ 2848]='h000008dc;
    rd_cycle[ 2849] = 1'b0;  wr_cycle[ 2849] = 1'b1;  addr_rom[ 2849]='h00000c7c;  wr_data_rom[ 2849]='h00001a92;
    rd_cycle[ 2850] = 1'b0;  wr_cycle[ 2850] = 1'b1;  addr_rom[ 2850]='h00000f18;  wr_data_rom[ 2850]='h0000085e;
    rd_cycle[ 2851] = 1'b0;  wr_cycle[ 2851] = 1'b1;  addr_rom[ 2851]='h000012d0;  wr_data_rom[ 2851]='h00001e5c;
    rd_cycle[ 2852] = 1'b1;  wr_cycle[ 2852] = 1'b0;  addr_rom[ 2852]='h00001bd4;  wr_data_rom[ 2852]='h00000000;
    rd_cycle[ 2853] = 1'b1;  wr_cycle[ 2853] = 1'b0;  addr_rom[ 2853]='h00000318;  wr_data_rom[ 2853]='h00000000;
    rd_cycle[ 2854] = 1'b1;  wr_cycle[ 2854] = 1'b0;  addr_rom[ 2854]='h00000458;  wr_data_rom[ 2854]='h00000000;
    rd_cycle[ 2855] = 1'b0;  wr_cycle[ 2855] = 1'b1;  addr_rom[ 2855]='h00001828;  wr_data_rom[ 2855]='h00000b21;
    rd_cycle[ 2856] = 1'b0;  wr_cycle[ 2856] = 1'b1;  addr_rom[ 2856]='h000003ac;  wr_data_rom[ 2856]='h000015f7;
    rd_cycle[ 2857] = 1'b0;  wr_cycle[ 2857] = 1'b1;  addr_rom[ 2857]='h000015e0;  wr_data_rom[ 2857]='h00001596;
    rd_cycle[ 2858] = 1'b0;  wr_cycle[ 2858] = 1'b1;  addr_rom[ 2858]='h00000a48;  wr_data_rom[ 2858]='h0000013e;
    rd_cycle[ 2859] = 1'b1;  wr_cycle[ 2859] = 1'b0;  addr_rom[ 2859]='h000016b8;  wr_data_rom[ 2859]='h00000000;
    rd_cycle[ 2860] = 1'b0;  wr_cycle[ 2860] = 1'b1;  addr_rom[ 2860]='h000013c8;  wr_data_rom[ 2860]='h00000095;
    rd_cycle[ 2861] = 1'b0;  wr_cycle[ 2861] = 1'b1;  addr_rom[ 2861]='h00001864;  wr_data_rom[ 2861]='h0000191c;
    rd_cycle[ 2862] = 1'b1;  wr_cycle[ 2862] = 1'b0;  addr_rom[ 2862]='h00000da4;  wr_data_rom[ 2862]='h00000000;
    rd_cycle[ 2863] = 1'b0;  wr_cycle[ 2863] = 1'b1;  addr_rom[ 2863]='h000012cc;  wr_data_rom[ 2863]='h00000259;
    rd_cycle[ 2864] = 1'b1;  wr_cycle[ 2864] = 1'b0;  addr_rom[ 2864]='h00000904;  wr_data_rom[ 2864]='h00000000;
    rd_cycle[ 2865] = 1'b0;  wr_cycle[ 2865] = 1'b1;  addr_rom[ 2865]='h00000d28;  wr_data_rom[ 2865]='h00000508;
    rd_cycle[ 2866] = 1'b1;  wr_cycle[ 2866] = 1'b0;  addr_rom[ 2866]='h00001e20;  wr_data_rom[ 2866]='h00000000;
    rd_cycle[ 2867] = 1'b1;  wr_cycle[ 2867] = 1'b0;  addr_rom[ 2867]='h00001090;  wr_data_rom[ 2867]='h00000000;
    rd_cycle[ 2868] = 1'b0;  wr_cycle[ 2868] = 1'b1;  addr_rom[ 2868]='h00000318;  wr_data_rom[ 2868]='h00001e9f;
    rd_cycle[ 2869] = 1'b1;  wr_cycle[ 2869] = 1'b0;  addr_rom[ 2869]='h000002f4;  wr_data_rom[ 2869]='h00000000;
    rd_cycle[ 2870] = 1'b1;  wr_cycle[ 2870] = 1'b0;  addr_rom[ 2870]='h00000920;  wr_data_rom[ 2870]='h00000000;
    rd_cycle[ 2871] = 1'b0;  wr_cycle[ 2871] = 1'b1;  addr_rom[ 2871]='h000003cc;  wr_data_rom[ 2871]='h00000b9c;
    rd_cycle[ 2872] = 1'b0;  wr_cycle[ 2872] = 1'b1;  addr_rom[ 2872]='h00000b80;  wr_data_rom[ 2872]='h000000ff;
    rd_cycle[ 2873] = 1'b1;  wr_cycle[ 2873] = 1'b0;  addr_rom[ 2873]='h00000adc;  wr_data_rom[ 2873]='h00000000;
    rd_cycle[ 2874] = 1'b0;  wr_cycle[ 2874] = 1'b1;  addr_rom[ 2874]='h00001eb8;  wr_data_rom[ 2874]='h00000844;
    rd_cycle[ 2875] = 1'b1;  wr_cycle[ 2875] = 1'b0;  addr_rom[ 2875]='h00000a20;  wr_data_rom[ 2875]='h00000000;
    rd_cycle[ 2876] = 1'b0;  wr_cycle[ 2876] = 1'b1;  addr_rom[ 2876]='h00001d90;  wr_data_rom[ 2876]='h0000083d;
    rd_cycle[ 2877] = 1'b1;  wr_cycle[ 2877] = 1'b0;  addr_rom[ 2877]='h00000f78;  wr_data_rom[ 2877]='h00000000;
    rd_cycle[ 2878] = 1'b1;  wr_cycle[ 2878] = 1'b0;  addr_rom[ 2878]='h00001b6c;  wr_data_rom[ 2878]='h00000000;
    rd_cycle[ 2879] = 1'b0;  wr_cycle[ 2879] = 1'b1;  addr_rom[ 2879]='h00000158;  wr_data_rom[ 2879]='h00000f08;
    rd_cycle[ 2880] = 1'b1;  wr_cycle[ 2880] = 1'b0;  addr_rom[ 2880]='h000010c4;  wr_data_rom[ 2880]='h00000000;
    rd_cycle[ 2881] = 1'b1;  wr_cycle[ 2881] = 1'b0;  addr_rom[ 2881]='h00001b7c;  wr_data_rom[ 2881]='h00000000;
    rd_cycle[ 2882] = 1'b0;  wr_cycle[ 2882] = 1'b1;  addr_rom[ 2882]='h00001f34;  wr_data_rom[ 2882]='h0000171a;
    rd_cycle[ 2883] = 1'b0;  wr_cycle[ 2883] = 1'b1;  addr_rom[ 2883]='h00000f20;  wr_data_rom[ 2883]='h00001d90;
    rd_cycle[ 2884] = 1'b1;  wr_cycle[ 2884] = 1'b0;  addr_rom[ 2884]='h00001080;  wr_data_rom[ 2884]='h00000000;
    rd_cycle[ 2885] = 1'b0;  wr_cycle[ 2885] = 1'b1;  addr_rom[ 2885]='h000000d0;  wr_data_rom[ 2885]='h00001180;
    rd_cycle[ 2886] = 1'b0;  wr_cycle[ 2886] = 1'b1;  addr_rom[ 2886]='h0000056c;  wr_data_rom[ 2886]='h00000db7;
    rd_cycle[ 2887] = 1'b0;  wr_cycle[ 2887] = 1'b1;  addr_rom[ 2887]='h00000e30;  wr_data_rom[ 2887]='h00001322;
    rd_cycle[ 2888] = 1'b1;  wr_cycle[ 2888] = 1'b0;  addr_rom[ 2888]='h000016c8;  wr_data_rom[ 2888]='h00000000;
    rd_cycle[ 2889] = 1'b0;  wr_cycle[ 2889] = 1'b1;  addr_rom[ 2889]='h00000a30;  wr_data_rom[ 2889]='h000018c7;
    rd_cycle[ 2890] = 1'b1;  wr_cycle[ 2890] = 1'b0;  addr_rom[ 2890]='h00000c74;  wr_data_rom[ 2890]='h00000000;
    rd_cycle[ 2891] = 1'b1;  wr_cycle[ 2891] = 1'b0;  addr_rom[ 2891]='h00000050;  wr_data_rom[ 2891]='h00000000;
    rd_cycle[ 2892] = 1'b1;  wr_cycle[ 2892] = 1'b0;  addr_rom[ 2892]='h00001864;  wr_data_rom[ 2892]='h00000000;
    rd_cycle[ 2893] = 1'b1;  wr_cycle[ 2893] = 1'b0;  addr_rom[ 2893]='h00001390;  wr_data_rom[ 2893]='h00000000;
    rd_cycle[ 2894] = 1'b0;  wr_cycle[ 2894] = 1'b1;  addr_rom[ 2894]='h000001a4;  wr_data_rom[ 2894]='h000018e4;
    rd_cycle[ 2895] = 1'b0;  wr_cycle[ 2895] = 1'b1;  addr_rom[ 2895]='h00000254;  wr_data_rom[ 2895]='h00000378;
    rd_cycle[ 2896] = 1'b1;  wr_cycle[ 2896] = 1'b0;  addr_rom[ 2896]='h00001370;  wr_data_rom[ 2896]='h00000000;
    rd_cycle[ 2897] = 1'b0;  wr_cycle[ 2897] = 1'b1;  addr_rom[ 2897]='h00001d38;  wr_data_rom[ 2897]='h00000f16;
    rd_cycle[ 2898] = 1'b0;  wr_cycle[ 2898] = 1'b1;  addr_rom[ 2898]='h00000ca8;  wr_data_rom[ 2898]='h00000f07;
    rd_cycle[ 2899] = 1'b0;  wr_cycle[ 2899] = 1'b1;  addr_rom[ 2899]='h000003f8;  wr_data_rom[ 2899]='h00000c0a;
    rd_cycle[ 2900] = 1'b0;  wr_cycle[ 2900] = 1'b1;  addr_rom[ 2900]='h00001748;  wr_data_rom[ 2900]='h00001acc;
    rd_cycle[ 2901] = 1'b0;  wr_cycle[ 2901] = 1'b1;  addr_rom[ 2901]='h00000fcc;  wr_data_rom[ 2901]='h000006a5;
    rd_cycle[ 2902] = 1'b0;  wr_cycle[ 2902] = 1'b1;  addr_rom[ 2902]='h00000a64;  wr_data_rom[ 2902]='h00000ba2;
    rd_cycle[ 2903] = 1'b1;  wr_cycle[ 2903] = 1'b0;  addr_rom[ 2903]='h00000cc0;  wr_data_rom[ 2903]='h00000000;
    rd_cycle[ 2904] = 1'b1;  wr_cycle[ 2904] = 1'b0;  addr_rom[ 2904]='h00001b18;  wr_data_rom[ 2904]='h00000000;
    rd_cycle[ 2905] = 1'b0;  wr_cycle[ 2905] = 1'b1;  addr_rom[ 2905]='h000014ac;  wr_data_rom[ 2905]='h0000179c;
    rd_cycle[ 2906] = 1'b0;  wr_cycle[ 2906] = 1'b1;  addr_rom[ 2906]='h0000073c;  wr_data_rom[ 2906]='h000002ad;
    rd_cycle[ 2907] = 1'b1;  wr_cycle[ 2907] = 1'b0;  addr_rom[ 2907]='h00001138;  wr_data_rom[ 2907]='h00000000;
    rd_cycle[ 2908] = 1'b0;  wr_cycle[ 2908] = 1'b1;  addr_rom[ 2908]='h00000e1c;  wr_data_rom[ 2908]='h0000170c;
    rd_cycle[ 2909] = 1'b0;  wr_cycle[ 2909] = 1'b1;  addr_rom[ 2909]='h00001f3c;  wr_data_rom[ 2909]='h00001427;
    rd_cycle[ 2910] = 1'b0;  wr_cycle[ 2910] = 1'b1;  addr_rom[ 2910]='h000007f0;  wr_data_rom[ 2910]='h00000133;
    rd_cycle[ 2911] = 1'b1;  wr_cycle[ 2911] = 1'b0;  addr_rom[ 2911]='h000015b8;  wr_data_rom[ 2911]='h00000000;
    rd_cycle[ 2912] = 1'b1;  wr_cycle[ 2912] = 1'b0;  addr_rom[ 2912]='h0000089c;  wr_data_rom[ 2912]='h00000000;
    rd_cycle[ 2913] = 1'b0;  wr_cycle[ 2913] = 1'b1;  addr_rom[ 2913]='h00001de0;  wr_data_rom[ 2913]='h0000148b;
    rd_cycle[ 2914] = 1'b0;  wr_cycle[ 2914] = 1'b1;  addr_rom[ 2914]='h00000bd8;  wr_data_rom[ 2914]='h00000d3d;
    rd_cycle[ 2915] = 1'b0;  wr_cycle[ 2915] = 1'b1;  addr_rom[ 2915]='h00001f38;  wr_data_rom[ 2915]='h0000054e;
    rd_cycle[ 2916] = 1'b1;  wr_cycle[ 2916] = 1'b0;  addr_rom[ 2916]='h00000538;  wr_data_rom[ 2916]='h00000000;
    rd_cycle[ 2917] = 1'b0;  wr_cycle[ 2917] = 1'b1;  addr_rom[ 2917]='h00001e44;  wr_data_rom[ 2917]='h00000d78;
    rd_cycle[ 2918] = 1'b1;  wr_cycle[ 2918] = 1'b0;  addr_rom[ 2918]='h00001aa4;  wr_data_rom[ 2918]='h00000000;
    rd_cycle[ 2919] = 1'b1;  wr_cycle[ 2919] = 1'b0;  addr_rom[ 2919]='h00000bb8;  wr_data_rom[ 2919]='h00000000;
    rd_cycle[ 2920] = 1'b0;  wr_cycle[ 2920] = 1'b1;  addr_rom[ 2920]='h000018ac;  wr_data_rom[ 2920]='h00001b99;
    rd_cycle[ 2921] = 1'b0;  wr_cycle[ 2921] = 1'b1;  addr_rom[ 2921]='h00001618;  wr_data_rom[ 2921]='h0000107e;
    rd_cycle[ 2922] = 1'b1;  wr_cycle[ 2922] = 1'b0;  addr_rom[ 2922]='h00001db4;  wr_data_rom[ 2922]='h00000000;
    rd_cycle[ 2923] = 1'b0;  wr_cycle[ 2923] = 1'b1;  addr_rom[ 2923]='h00000ab0;  wr_data_rom[ 2923]='h0000110c;
    rd_cycle[ 2924] = 1'b0;  wr_cycle[ 2924] = 1'b1;  addr_rom[ 2924]='h000004fc;  wr_data_rom[ 2924]='h00000797;
    rd_cycle[ 2925] = 1'b1;  wr_cycle[ 2925] = 1'b0;  addr_rom[ 2925]='h00000ea0;  wr_data_rom[ 2925]='h00000000;
    rd_cycle[ 2926] = 1'b0;  wr_cycle[ 2926] = 1'b1;  addr_rom[ 2926]='h00000b40;  wr_data_rom[ 2926]='h000011e0;
    rd_cycle[ 2927] = 1'b1;  wr_cycle[ 2927] = 1'b0;  addr_rom[ 2927]='h00001b44;  wr_data_rom[ 2927]='h00000000;
    rd_cycle[ 2928] = 1'b0;  wr_cycle[ 2928] = 1'b1;  addr_rom[ 2928]='h000007c0;  wr_data_rom[ 2928]='h000003a5;
    rd_cycle[ 2929] = 1'b0;  wr_cycle[ 2929] = 1'b1;  addr_rom[ 2929]='h0000084c;  wr_data_rom[ 2929]='h000002aa;
    rd_cycle[ 2930] = 1'b1;  wr_cycle[ 2930] = 1'b0;  addr_rom[ 2930]='h000019a4;  wr_data_rom[ 2930]='h00000000;
    rd_cycle[ 2931] = 1'b1;  wr_cycle[ 2931] = 1'b0;  addr_rom[ 2931]='h00000a60;  wr_data_rom[ 2931]='h00000000;
    rd_cycle[ 2932] = 1'b0;  wr_cycle[ 2932] = 1'b1;  addr_rom[ 2932]='h00000e0c;  wr_data_rom[ 2932]='h00000462;
    rd_cycle[ 2933] = 1'b1;  wr_cycle[ 2933] = 1'b0;  addr_rom[ 2933]='h00001834;  wr_data_rom[ 2933]='h00000000;
    rd_cycle[ 2934] = 1'b0;  wr_cycle[ 2934] = 1'b1;  addr_rom[ 2934]='h00001470;  wr_data_rom[ 2934]='h00000f97;
    rd_cycle[ 2935] = 1'b1;  wr_cycle[ 2935] = 1'b0;  addr_rom[ 2935]='h00001be0;  wr_data_rom[ 2935]='h00000000;
    rd_cycle[ 2936] = 1'b1;  wr_cycle[ 2936] = 1'b0;  addr_rom[ 2936]='h00001b38;  wr_data_rom[ 2936]='h00000000;
    rd_cycle[ 2937] = 1'b1;  wr_cycle[ 2937] = 1'b0;  addr_rom[ 2937]='h000018a4;  wr_data_rom[ 2937]='h00000000;
    rd_cycle[ 2938] = 1'b1;  wr_cycle[ 2938] = 1'b0;  addr_rom[ 2938]='h00000e40;  wr_data_rom[ 2938]='h00000000;
    rd_cycle[ 2939] = 1'b0;  wr_cycle[ 2939] = 1'b1;  addr_rom[ 2939]='h0000053c;  wr_data_rom[ 2939]='h000007da;
    rd_cycle[ 2940] = 1'b0;  wr_cycle[ 2940] = 1'b1;  addr_rom[ 2940]='h0000070c;  wr_data_rom[ 2940]='h00000eed;
    rd_cycle[ 2941] = 1'b0;  wr_cycle[ 2941] = 1'b1;  addr_rom[ 2941]='h0000133c;  wr_data_rom[ 2941]='h00000c28;
    rd_cycle[ 2942] = 1'b1;  wr_cycle[ 2942] = 1'b0;  addr_rom[ 2942]='h000001ec;  wr_data_rom[ 2942]='h00000000;
    rd_cycle[ 2943] = 1'b0;  wr_cycle[ 2943] = 1'b1;  addr_rom[ 2943]='h0000189c;  wr_data_rom[ 2943]='h00001531;
    rd_cycle[ 2944] = 1'b1;  wr_cycle[ 2944] = 1'b0;  addr_rom[ 2944]='h000013e0;  wr_data_rom[ 2944]='h00000000;
    rd_cycle[ 2945] = 1'b0;  wr_cycle[ 2945] = 1'b1;  addr_rom[ 2945]='h00000808;  wr_data_rom[ 2945]='h0000021b;
    rd_cycle[ 2946] = 1'b1;  wr_cycle[ 2946] = 1'b0;  addr_rom[ 2946]='h0000085c;  wr_data_rom[ 2946]='h00000000;
    rd_cycle[ 2947] = 1'b1;  wr_cycle[ 2947] = 1'b0;  addr_rom[ 2947]='h00000e88;  wr_data_rom[ 2947]='h00000000;
    rd_cycle[ 2948] = 1'b1;  wr_cycle[ 2948] = 1'b0;  addr_rom[ 2948]='h00000e94;  wr_data_rom[ 2948]='h00000000;
    rd_cycle[ 2949] = 1'b0;  wr_cycle[ 2949] = 1'b1;  addr_rom[ 2949]='h000012c8;  wr_data_rom[ 2949]='h00000abf;
    rd_cycle[ 2950] = 1'b1;  wr_cycle[ 2950] = 1'b0;  addr_rom[ 2950]='h000004ac;  wr_data_rom[ 2950]='h00000000;
    rd_cycle[ 2951] = 1'b0;  wr_cycle[ 2951] = 1'b1;  addr_rom[ 2951]='h00001194;  wr_data_rom[ 2951]='h000018a1;
    rd_cycle[ 2952] = 1'b1;  wr_cycle[ 2952] = 1'b0;  addr_rom[ 2952]='h00001c78;  wr_data_rom[ 2952]='h00000000;
    rd_cycle[ 2953] = 1'b1;  wr_cycle[ 2953] = 1'b0;  addr_rom[ 2953]='h00000464;  wr_data_rom[ 2953]='h00000000;
    rd_cycle[ 2954] = 1'b0;  wr_cycle[ 2954] = 1'b1;  addr_rom[ 2954]='h00000ec8;  wr_data_rom[ 2954]='h00001437;
    rd_cycle[ 2955] = 1'b0;  wr_cycle[ 2955] = 1'b1;  addr_rom[ 2955]='h000010dc;  wr_data_rom[ 2955]='h000008ca;
    rd_cycle[ 2956] = 1'b0;  wr_cycle[ 2956] = 1'b1;  addr_rom[ 2956]='h0000179c;  wr_data_rom[ 2956]='h00001e00;
    rd_cycle[ 2957] = 1'b1;  wr_cycle[ 2957] = 1'b0;  addr_rom[ 2957]='h00000e30;  wr_data_rom[ 2957]='h00000000;
    rd_cycle[ 2958] = 1'b1;  wr_cycle[ 2958] = 1'b0;  addr_rom[ 2958]='h00000370;  wr_data_rom[ 2958]='h00000000;
    rd_cycle[ 2959] = 1'b1;  wr_cycle[ 2959] = 1'b0;  addr_rom[ 2959]='h00001708;  wr_data_rom[ 2959]='h00000000;
    rd_cycle[ 2960] = 1'b0;  wr_cycle[ 2960] = 1'b1;  addr_rom[ 2960]='h0000009c;  wr_data_rom[ 2960]='h000016fa;
    rd_cycle[ 2961] = 1'b0;  wr_cycle[ 2961] = 1'b1;  addr_rom[ 2961]='h00001cb8;  wr_data_rom[ 2961]='h00001965;
    rd_cycle[ 2962] = 1'b0;  wr_cycle[ 2962] = 1'b1;  addr_rom[ 2962]='h00001034;  wr_data_rom[ 2962]='h00001aab;
    rd_cycle[ 2963] = 1'b1;  wr_cycle[ 2963] = 1'b0;  addr_rom[ 2963]='h00000bc4;  wr_data_rom[ 2963]='h00000000;
    rd_cycle[ 2964] = 1'b0;  wr_cycle[ 2964] = 1'b1;  addr_rom[ 2964]='h00001b14;  wr_data_rom[ 2964]='h00001333;
    rd_cycle[ 2965] = 1'b0;  wr_cycle[ 2965] = 1'b1;  addr_rom[ 2965]='h00000a58;  wr_data_rom[ 2965]='h00000c3b;
    rd_cycle[ 2966] = 1'b1;  wr_cycle[ 2966] = 1'b0;  addr_rom[ 2966]='h000010c0;  wr_data_rom[ 2966]='h00000000;
    rd_cycle[ 2967] = 1'b0;  wr_cycle[ 2967] = 1'b1;  addr_rom[ 2967]='h000002cc;  wr_data_rom[ 2967]='h00000885;
    rd_cycle[ 2968] = 1'b0;  wr_cycle[ 2968] = 1'b1;  addr_rom[ 2968]='h000005d0;  wr_data_rom[ 2968]='h0000146e;
    rd_cycle[ 2969] = 1'b1;  wr_cycle[ 2969] = 1'b0;  addr_rom[ 2969]='h0000096c;  wr_data_rom[ 2969]='h00000000;
    rd_cycle[ 2970] = 1'b1;  wr_cycle[ 2970] = 1'b0;  addr_rom[ 2970]='h00000b80;  wr_data_rom[ 2970]='h00000000;
    rd_cycle[ 2971] = 1'b0;  wr_cycle[ 2971] = 1'b1;  addr_rom[ 2971]='h00001f2c;  wr_data_rom[ 2971]='h00001148;
    rd_cycle[ 2972] = 1'b1;  wr_cycle[ 2972] = 1'b0;  addr_rom[ 2972]='h00001d98;  wr_data_rom[ 2972]='h00000000;
    rd_cycle[ 2973] = 1'b0;  wr_cycle[ 2973] = 1'b1;  addr_rom[ 2973]='h000019a8;  wr_data_rom[ 2973]='h00000f43;
    rd_cycle[ 2974] = 1'b1;  wr_cycle[ 2974] = 1'b0;  addr_rom[ 2974]='h000004bc;  wr_data_rom[ 2974]='h00000000;
    rd_cycle[ 2975] = 1'b1;  wr_cycle[ 2975] = 1'b0;  addr_rom[ 2975]='h00000f2c;  wr_data_rom[ 2975]='h00000000;
    rd_cycle[ 2976] = 1'b0;  wr_cycle[ 2976] = 1'b1;  addr_rom[ 2976]='h000018e4;  wr_data_rom[ 2976]='h0000100e;
    rd_cycle[ 2977] = 1'b0;  wr_cycle[ 2977] = 1'b1;  addr_rom[ 2977]='h00001cb0;  wr_data_rom[ 2977]='h00001329;
    rd_cycle[ 2978] = 1'b1;  wr_cycle[ 2978] = 1'b0;  addr_rom[ 2978]='h00001190;  wr_data_rom[ 2978]='h00000000;
    rd_cycle[ 2979] = 1'b1;  wr_cycle[ 2979] = 1'b0;  addr_rom[ 2979]='h00001574;  wr_data_rom[ 2979]='h00000000;
    rd_cycle[ 2980] = 1'b0;  wr_cycle[ 2980] = 1'b1;  addr_rom[ 2980]='h00000650;  wr_data_rom[ 2980]='h000000d2;
    rd_cycle[ 2981] = 1'b0;  wr_cycle[ 2981] = 1'b1;  addr_rom[ 2981]='h00000e20;  wr_data_rom[ 2981]='h000010f1;
    rd_cycle[ 2982] = 1'b1;  wr_cycle[ 2982] = 1'b0;  addr_rom[ 2982]='h00001494;  wr_data_rom[ 2982]='h00000000;
    rd_cycle[ 2983] = 1'b1;  wr_cycle[ 2983] = 1'b0;  addr_rom[ 2983]='h00001da0;  wr_data_rom[ 2983]='h00000000;
    rd_cycle[ 2984] = 1'b1;  wr_cycle[ 2984] = 1'b0;  addr_rom[ 2984]='h000007c4;  wr_data_rom[ 2984]='h00000000;
    rd_cycle[ 2985] = 1'b1;  wr_cycle[ 2985] = 1'b0;  addr_rom[ 2985]='h00001cd8;  wr_data_rom[ 2985]='h00000000;
    rd_cycle[ 2986] = 1'b1;  wr_cycle[ 2986] = 1'b0;  addr_rom[ 2986]='h00001954;  wr_data_rom[ 2986]='h00000000;
    rd_cycle[ 2987] = 1'b0;  wr_cycle[ 2987] = 1'b1;  addr_rom[ 2987]='h00000604;  wr_data_rom[ 2987]='h0000194a;
    rd_cycle[ 2988] = 1'b1;  wr_cycle[ 2988] = 1'b0;  addr_rom[ 2988]='h000015ac;  wr_data_rom[ 2988]='h00000000;
    rd_cycle[ 2989] = 1'b0;  wr_cycle[ 2989] = 1'b1;  addr_rom[ 2989]='h00001484;  wr_data_rom[ 2989]='h00000237;
    rd_cycle[ 2990] = 1'b1;  wr_cycle[ 2990] = 1'b0;  addr_rom[ 2990]='h000008d4;  wr_data_rom[ 2990]='h00000000;
    rd_cycle[ 2991] = 1'b1;  wr_cycle[ 2991] = 1'b0;  addr_rom[ 2991]='h00001d44;  wr_data_rom[ 2991]='h00000000;
    rd_cycle[ 2992] = 1'b0;  wr_cycle[ 2992] = 1'b1;  addr_rom[ 2992]='h00001778;  wr_data_rom[ 2992]='h00000a59;
    rd_cycle[ 2993] = 1'b0;  wr_cycle[ 2993] = 1'b1;  addr_rom[ 2993]='h000012c0;  wr_data_rom[ 2993]='h00000853;
    rd_cycle[ 2994] = 1'b1;  wr_cycle[ 2994] = 1'b0;  addr_rom[ 2994]='h00000328;  wr_data_rom[ 2994]='h00000000;
    rd_cycle[ 2995] = 1'b0;  wr_cycle[ 2995] = 1'b1;  addr_rom[ 2995]='h00000d4c;  wr_data_rom[ 2995]='h000015bd;
    rd_cycle[ 2996] = 1'b1;  wr_cycle[ 2996] = 1'b0;  addr_rom[ 2996]='h00001c50;  wr_data_rom[ 2996]='h00000000;
    rd_cycle[ 2997] = 1'b1;  wr_cycle[ 2997] = 1'b0;  addr_rom[ 2997]='h00001794;  wr_data_rom[ 2997]='h00000000;
    rd_cycle[ 2998] = 1'b0;  wr_cycle[ 2998] = 1'b1;  addr_rom[ 2998]='h00001350;  wr_data_rom[ 2998]='h00001d76;
    rd_cycle[ 2999] = 1'b0;  wr_cycle[ 2999] = 1'b1;  addr_rom[ 2999]='h00001040;  wr_data_rom[ 2999]='h0000126f;
    rd_cycle[ 3000] = 1'b0;  wr_cycle[ 3000] = 1'b1;  addr_rom[ 3000]='h00000ca8;  wr_data_rom[ 3000]='h00001577;
    rd_cycle[ 3001] = 1'b1;  wr_cycle[ 3001] = 1'b0;  addr_rom[ 3001]='h00001e4c;  wr_data_rom[ 3001]='h00000000;
    rd_cycle[ 3002] = 1'b0;  wr_cycle[ 3002] = 1'b1;  addr_rom[ 3002]='h000007d8;  wr_data_rom[ 3002]='h00000f34;
    rd_cycle[ 3003] = 1'b0;  wr_cycle[ 3003] = 1'b1;  addr_rom[ 3003]='h00001298;  wr_data_rom[ 3003]='h00001537;
    rd_cycle[ 3004] = 1'b0;  wr_cycle[ 3004] = 1'b1;  addr_rom[ 3004]='h00001d18;  wr_data_rom[ 3004]='h000011ca;
    rd_cycle[ 3005] = 1'b0;  wr_cycle[ 3005] = 1'b1;  addr_rom[ 3005]='h00001454;  wr_data_rom[ 3005]='h00001abc;
    rd_cycle[ 3006] = 1'b1;  wr_cycle[ 3006] = 1'b0;  addr_rom[ 3006]='h00000a44;  wr_data_rom[ 3006]='h00000000;
    rd_cycle[ 3007] = 1'b1;  wr_cycle[ 3007] = 1'b0;  addr_rom[ 3007]='h0000172c;  wr_data_rom[ 3007]='h00000000;
    rd_cycle[ 3008] = 1'b0;  wr_cycle[ 3008] = 1'b1;  addr_rom[ 3008]='h0000009c;  wr_data_rom[ 3008]='h0000076a;
    rd_cycle[ 3009] = 1'b0;  wr_cycle[ 3009] = 1'b1;  addr_rom[ 3009]='h00000188;  wr_data_rom[ 3009]='h00001978;
    rd_cycle[ 3010] = 1'b0;  wr_cycle[ 3010] = 1'b1;  addr_rom[ 3010]='h00001cd4;  wr_data_rom[ 3010]='h00001356;
    rd_cycle[ 3011] = 1'b1;  wr_cycle[ 3011] = 1'b0;  addr_rom[ 3011]='h00000fa8;  wr_data_rom[ 3011]='h00000000;
    rd_cycle[ 3012] = 1'b1;  wr_cycle[ 3012] = 1'b0;  addr_rom[ 3012]='h000010bc;  wr_data_rom[ 3012]='h00000000;
    rd_cycle[ 3013] = 1'b0;  wr_cycle[ 3013] = 1'b1;  addr_rom[ 3013]='h000014b4;  wr_data_rom[ 3013]='h000012b2;
    rd_cycle[ 3014] = 1'b1;  wr_cycle[ 3014] = 1'b0;  addr_rom[ 3014]='h00001a18;  wr_data_rom[ 3014]='h00000000;
    rd_cycle[ 3015] = 1'b0;  wr_cycle[ 3015] = 1'b1;  addr_rom[ 3015]='h000008c4;  wr_data_rom[ 3015]='h00000ce3;
    rd_cycle[ 3016] = 1'b1;  wr_cycle[ 3016] = 1'b0;  addr_rom[ 3016]='h00000b60;  wr_data_rom[ 3016]='h00000000;
    rd_cycle[ 3017] = 1'b0;  wr_cycle[ 3017] = 1'b1;  addr_rom[ 3017]='h00001444;  wr_data_rom[ 3017]='h000014cb;
    rd_cycle[ 3018] = 1'b1;  wr_cycle[ 3018] = 1'b0;  addr_rom[ 3018]='h00001558;  wr_data_rom[ 3018]='h00000000;
    rd_cycle[ 3019] = 1'b0;  wr_cycle[ 3019] = 1'b1;  addr_rom[ 3019]='h000009ec;  wr_data_rom[ 3019]='h00001e4a;
    rd_cycle[ 3020] = 1'b1;  wr_cycle[ 3020] = 1'b0;  addr_rom[ 3020]='h00001040;  wr_data_rom[ 3020]='h00000000;
    rd_cycle[ 3021] = 1'b0;  wr_cycle[ 3021] = 1'b1;  addr_rom[ 3021]='h0000136c;  wr_data_rom[ 3021]='h00000c83;
    rd_cycle[ 3022] = 1'b1;  wr_cycle[ 3022] = 1'b0;  addr_rom[ 3022]='h00001dfc;  wr_data_rom[ 3022]='h00000000;
    rd_cycle[ 3023] = 1'b0;  wr_cycle[ 3023] = 1'b1;  addr_rom[ 3023]='h00000978;  wr_data_rom[ 3023]='h00001ba0;
    rd_cycle[ 3024] = 1'b1;  wr_cycle[ 3024] = 1'b0;  addr_rom[ 3024]='h00001b0c;  wr_data_rom[ 3024]='h00000000;
    rd_cycle[ 3025] = 1'b1;  wr_cycle[ 3025] = 1'b0;  addr_rom[ 3025]='h00001500;  wr_data_rom[ 3025]='h00000000;
    rd_cycle[ 3026] = 1'b1;  wr_cycle[ 3026] = 1'b0;  addr_rom[ 3026]='h00000ee8;  wr_data_rom[ 3026]='h00000000;
    rd_cycle[ 3027] = 1'b0;  wr_cycle[ 3027] = 1'b1;  addr_rom[ 3027]='h00001c48;  wr_data_rom[ 3027]='h0000104a;
    rd_cycle[ 3028] = 1'b0;  wr_cycle[ 3028] = 1'b1;  addr_rom[ 3028]='h000013c8;  wr_data_rom[ 3028]='h00000295;
    rd_cycle[ 3029] = 1'b0;  wr_cycle[ 3029] = 1'b1;  addr_rom[ 3029]='h00000224;  wr_data_rom[ 3029]='h00000e52;
    rd_cycle[ 3030] = 1'b1;  wr_cycle[ 3030] = 1'b0;  addr_rom[ 3030]='h00001ce8;  wr_data_rom[ 3030]='h00000000;
    rd_cycle[ 3031] = 1'b0;  wr_cycle[ 3031] = 1'b1;  addr_rom[ 3031]='h00001f28;  wr_data_rom[ 3031]='h000013f9;
    rd_cycle[ 3032] = 1'b0;  wr_cycle[ 3032] = 1'b1;  addr_rom[ 3032]='h00001d60;  wr_data_rom[ 3032]='h00001f13;
    rd_cycle[ 3033] = 1'b1;  wr_cycle[ 3033] = 1'b0;  addr_rom[ 3033]='h000007b0;  wr_data_rom[ 3033]='h00000000;
    rd_cycle[ 3034] = 1'b1;  wr_cycle[ 3034] = 1'b0;  addr_rom[ 3034]='h0000153c;  wr_data_rom[ 3034]='h00000000;
    rd_cycle[ 3035] = 1'b0;  wr_cycle[ 3035] = 1'b1;  addr_rom[ 3035]='h000014b8;  wr_data_rom[ 3035]='h00001177;
    rd_cycle[ 3036] = 1'b1;  wr_cycle[ 3036] = 1'b0;  addr_rom[ 3036]='h00001e40;  wr_data_rom[ 3036]='h00000000;
    rd_cycle[ 3037] = 1'b0;  wr_cycle[ 3037] = 1'b1;  addr_rom[ 3037]='h00001e14;  wr_data_rom[ 3037]='h000000d2;
    rd_cycle[ 3038] = 1'b1;  wr_cycle[ 3038] = 1'b0;  addr_rom[ 3038]='h0000021c;  wr_data_rom[ 3038]='h00000000;
    rd_cycle[ 3039] = 1'b1;  wr_cycle[ 3039] = 1'b0;  addr_rom[ 3039]='h000001d0;  wr_data_rom[ 3039]='h00000000;
    rd_cycle[ 3040] = 1'b0;  wr_cycle[ 3040] = 1'b1;  addr_rom[ 3040]='h00001074;  wr_data_rom[ 3040]='h00001ce6;
    rd_cycle[ 3041] = 1'b0;  wr_cycle[ 3041] = 1'b1;  addr_rom[ 3041]='h00000d7c;  wr_data_rom[ 3041]='h00000ebb;
    rd_cycle[ 3042] = 1'b1;  wr_cycle[ 3042] = 1'b0;  addr_rom[ 3042]='h000019b4;  wr_data_rom[ 3042]='h00000000;
    rd_cycle[ 3043] = 1'b0;  wr_cycle[ 3043] = 1'b1;  addr_rom[ 3043]='h00001ef0;  wr_data_rom[ 3043]='h00001c2c;
    rd_cycle[ 3044] = 1'b0;  wr_cycle[ 3044] = 1'b1;  addr_rom[ 3044]='h00000830;  wr_data_rom[ 3044]='h0000035c;
    rd_cycle[ 3045] = 1'b0;  wr_cycle[ 3045] = 1'b1;  addr_rom[ 3045]='h00000edc;  wr_data_rom[ 3045]='h0000109b;
    rd_cycle[ 3046] = 1'b1;  wr_cycle[ 3046] = 1'b0;  addr_rom[ 3046]='h0000183c;  wr_data_rom[ 3046]='h00000000;
    rd_cycle[ 3047] = 1'b1;  wr_cycle[ 3047] = 1'b0;  addr_rom[ 3047]='h00001610;  wr_data_rom[ 3047]='h00000000;
    rd_cycle[ 3048] = 1'b1;  wr_cycle[ 3048] = 1'b0;  addr_rom[ 3048]='h00000a68;  wr_data_rom[ 3048]='h00000000;
    rd_cycle[ 3049] = 1'b0;  wr_cycle[ 3049] = 1'b1;  addr_rom[ 3049]='h00000004;  wr_data_rom[ 3049]='h000011e3;
    rd_cycle[ 3050] = 1'b0;  wr_cycle[ 3050] = 1'b1;  addr_rom[ 3050]='h000001f8;  wr_data_rom[ 3050]='h000008c7;
    rd_cycle[ 3051] = 1'b1;  wr_cycle[ 3051] = 1'b0;  addr_rom[ 3051]='h00001614;  wr_data_rom[ 3051]='h00000000;
    rd_cycle[ 3052] = 1'b1;  wr_cycle[ 3052] = 1'b0;  addr_rom[ 3052]='h000018b0;  wr_data_rom[ 3052]='h00000000;
    rd_cycle[ 3053] = 1'b1;  wr_cycle[ 3053] = 1'b0;  addr_rom[ 3053]='h00000478;  wr_data_rom[ 3053]='h00000000;
    rd_cycle[ 3054] = 1'b1;  wr_cycle[ 3054] = 1'b0;  addr_rom[ 3054]='h00001334;  wr_data_rom[ 3054]='h00000000;
    rd_cycle[ 3055] = 1'b0;  wr_cycle[ 3055] = 1'b1;  addr_rom[ 3055]='h000015a0;  wr_data_rom[ 3055]='h00001206;
    rd_cycle[ 3056] = 1'b0;  wr_cycle[ 3056] = 1'b1;  addr_rom[ 3056]='h00000c60;  wr_data_rom[ 3056]='h00000f20;
    rd_cycle[ 3057] = 1'b0;  wr_cycle[ 3057] = 1'b1;  addr_rom[ 3057]='h00000700;  wr_data_rom[ 3057]='h00000ec0;
    rd_cycle[ 3058] = 1'b1;  wr_cycle[ 3058] = 1'b0;  addr_rom[ 3058]='h000004f8;  wr_data_rom[ 3058]='h00000000;
    rd_cycle[ 3059] = 1'b0;  wr_cycle[ 3059] = 1'b1;  addr_rom[ 3059]='h00001478;  wr_data_rom[ 3059]='h0000125a;
    rd_cycle[ 3060] = 1'b1;  wr_cycle[ 3060] = 1'b0;  addr_rom[ 3060]='h000006d8;  wr_data_rom[ 3060]='h00000000;
    rd_cycle[ 3061] = 1'b0;  wr_cycle[ 3061] = 1'b1;  addr_rom[ 3061]='h00000be8;  wr_data_rom[ 3061]='h00001828;
    rd_cycle[ 3062] = 1'b1;  wr_cycle[ 3062] = 1'b0;  addr_rom[ 3062]='h00001894;  wr_data_rom[ 3062]='h00000000;
    rd_cycle[ 3063] = 1'b0;  wr_cycle[ 3063] = 1'b1;  addr_rom[ 3063]='h00001ba4;  wr_data_rom[ 3063]='h00001457;
    rd_cycle[ 3064] = 1'b0;  wr_cycle[ 3064] = 1'b1;  addr_rom[ 3064]='h00001588;  wr_data_rom[ 3064]='h00001ba3;
    rd_cycle[ 3065] = 1'b1;  wr_cycle[ 3065] = 1'b0;  addr_rom[ 3065]='h00001d30;  wr_data_rom[ 3065]='h00000000;
    rd_cycle[ 3066] = 1'b1;  wr_cycle[ 3066] = 1'b0;  addr_rom[ 3066]='h000018d8;  wr_data_rom[ 3066]='h00000000;
    rd_cycle[ 3067] = 1'b0;  wr_cycle[ 3067] = 1'b1;  addr_rom[ 3067]='h00000b24;  wr_data_rom[ 3067]='h000001b2;
    rd_cycle[ 3068] = 1'b1;  wr_cycle[ 3068] = 1'b0;  addr_rom[ 3068]='h0000001c;  wr_data_rom[ 3068]='h00000000;
    rd_cycle[ 3069] = 1'b0;  wr_cycle[ 3069] = 1'b1;  addr_rom[ 3069]='h00000864;  wr_data_rom[ 3069]='h00001cb9;
    rd_cycle[ 3070] = 1'b0;  wr_cycle[ 3070] = 1'b1;  addr_rom[ 3070]='h00000964;  wr_data_rom[ 3070]='h000009b9;
    rd_cycle[ 3071] = 1'b1;  wr_cycle[ 3071] = 1'b0;  addr_rom[ 3071]='h000006f4;  wr_data_rom[ 3071]='h00000000;
    rd_cycle[ 3072] = 1'b1;  wr_cycle[ 3072] = 1'b0;  addr_rom[ 3072]='h00001a98;  wr_data_rom[ 3072]='h00000000;
    rd_cycle[ 3073] = 1'b1;  wr_cycle[ 3073] = 1'b0;  addr_rom[ 3073]='h00000724;  wr_data_rom[ 3073]='h00000000;
    rd_cycle[ 3074] = 1'b0;  wr_cycle[ 3074] = 1'b1;  addr_rom[ 3074]='h00001bd0;  wr_data_rom[ 3074]='h00001c40;
    rd_cycle[ 3075] = 1'b1;  wr_cycle[ 3075] = 1'b0;  addr_rom[ 3075]='h00001a10;  wr_data_rom[ 3075]='h00000000;
    rd_cycle[ 3076] = 1'b0;  wr_cycle[ 3076] = 1'b1;  addr_rom[ 3076]='h000013c8;  wr_data_rom[ 3076]='h00001083;
    rd_cycle[ 3077] = 1'b1;  wr_cycle[ 3077] = 1'b0;  addr_rom[ 3077]='h0000081c;  wr_data_rom[ 3077]='h00000000;
    rd_cycle[ 3078] = 1'b1;  wr_cycle[ 3078] = 1'b0;  addr_rom[ 3078]='h00001958;  wr_data_rom[ 3078]='h00000000;
    rd_cycle[ 3079] = 1'b0;  wr_cycle[ 3079] = 1'b1;  addr_rom[ 3079]='h00000934;  wr_data_rom[ 3079]='h00000d2f;
    rd_cycle[ 3080] = 1'b1;  wr_cycle[ 3080] = 1'b0;  addr_rom[ 3080]='h000010fc;  wr_data_rom[ 3080]='h00000000;
    rd_cycle[ 3081] = 1'b1;  wr_cycle[ 3081] = 1'b0;  addr_rom[ 3081]='h000005d8;  wr_data_rom[ 3081]='h00000000;
    rd_cycle[ 3082] = 1'b1;  wr_cycle[ 3082] = 1'b0;  addr_rom[ 3082]='h00000900;  wr_data_rom[ 3082]='h00000000;
    rd_cycle[ 3083] = 1'b0;  wr_cycle[ 3083] = 1'b1;  addr_rom[ 3083]='h00001090;  wr_data_rom[ 3083]='h00001595;
    rd_cycle[ 3084] = 1'b0;  wr_cycle[ 3084] = 1'b1;  addr_rom[ 3084]='h00000288;  wr_data_rom[ 3084]='h00001879;
    rd_cycle[ 3085] = 1'b0;  wr_cycle[ 3085] = 1'b1;  addr_rom[ 3085]='h00000810;  wr_data_rom[ 3085]='h000004cc;
    rd_cycle[ 3086] = 1'b1;  wr_cycle[ 3086] = 1'b0;  addr_rom[ 3086]='h000007ec;  wr_data_rom[ 3086]='h00000000;
    rd_cycle[ 3087] = 1'b1;  wr_cycle[ 3087] = 1'b0;  addr_rom[ 3087]='h000018cc;  wr_data_rom[ 3087]='h00000000;
    rd_cycle[ 3088] = 1'b0;  wr_cycle[ 3088] = 1'b1;  addr_rom[ 3088]='h00000e34;  wr_data_rom[ 3088]='h000014b2;
    rd_cycle[ 3089] = 1'b1;  wr_cycle[ 3089] = 1'b0;  addr_rom[ 3089]='h00000e24;  wr_data_rom[ 3089]='h00000000;
    rd_cycle[ 3090] = 1'b0;  wr_cycle[ 3090] = 1'b1;  addr_rom[ 3090]='h00001d3c;  wr_data_rom[ 3090]='h000007ba;
    rd_cycle[ 3091] = 1'b0;  wr_cycle[ 3091] = 1'b1;  addr_rom[ 3091]='h0000034c;  wr_data_rom[ 3091]='h00000000;
    rd_cycle[ 3092] = 1'b1;  wr_cycle[ 3092] = 1'b0;  addr_rom[ 3092]='h00001ad4;  wr_data_rom[ 3092]='h00000000;
    rd_cycle[ 3093] = 1'b1;  wr_cycle[ 3093] = 1'b0;  addr_rom[ 3093]='h00001210;  wr_data_rom[ 3093]='h00000000;
    rd_cycle[ 3094] = 1'b0;  wr_cycle[ 3094] = 1'b1;  addr_rom[ 3094]='h00001e1c;  wr_data_rom[ 3094]='h00000ee3;
    rd_cycle[ 3095] = 1'b1;  wr_cycle[ 3095] = 1'b0;  addr_rom[ 3095]='h00000e3c;  wr_data_rom[ 3095]='h00000000;
    rd_cycle[ 3096] = 1'b1;  wr_cycle[ 3096] = 1'b0;  addr_rom[ 3096]='h00000fb0;  wr_data_rom[ 3096]='h00000000;
    rd_cycle[ 3097] = 1'b1;  wr_cycle[ 3097] = 1'b0;  addr_rom[ 3097]='h0000112c;  wr_data_rom[ 3097]='h00000000;
    rd_cycle[ 3098] = 1'b0;  wr_cycle[ 3098] = 1'b1;  addr_rom[ 3098]='h00000388;  wr_data_rom[ 3098]='h00001b68;
    rd_cycle[ 3099] = 1'b1;  wr_cycle[ 3099] = 1'b0;  addr_rom[ 3099]='h0000012c;  wr_data_rom[ 3099]='h00000000;
    rd_cycle[ 3100] = 1'b0;  wr_cycle[ 3100] = 1'b1;  addr_rom[ 3100]='h00001c98;  wr_data_rom[ 3100]='h00001516;
    rd_cycle[ 3101] = 1'b1;  wr_cycle[ 3101] = 1'b0;  addr_rom[ 3101]='h0000186c;  wr_data_rom[ 3101]='h00000000;
    rd_cycle[ 3102] = 1'b0;  wr_cycle[ 3102] = 1'b1;  addr_rom[ 3102]='h0000187c;  wr_data_rom[ 3102]='h00000e1a;
    rd_cycle[ 3103] = 1'b0;  wr_cycle[ 3103] = 1'b1;  addr_rom[ 3103]='h00001d0c;  wr_data_rom[ 3103]='h00001028;
    rd_cycle[ 3104] = 1'b1;  wr_cycle[ 3104] = 1'b0;  addr_rom[ 3104]='h00000e78;  wr_data_rom[ 3104]='h00000000;
    rd_cycle[ 3105] = 1'b0;  wr_cycle[ 3105] = 1'b1;  addr_rom[ 3105]='h00001294;  wr_data_rom[ 3105]='h00000fbc;
    rd_cycle[ 3106] = 1'b1;  wr_cycle[ 3106] = 1'b0;  addr_rom[ 3106]='h000009f8;  wr_data_rom[ 3106]='h00000000;
    rd_cycle[ 3107] = 1'b1;  wr_cycle[ 3107] = 1'b0;  addr_rom[ 3107]='h000005a0;  wr_data_rom[ 3107]='h00000000;
    rd_cycle[ 3108] = 1'b0;  wr_cycle[ 3108] = 1'b1;  addr_rom[ 3108]='h000006dc;  wr_data_rom[ 3108]='h00000dfc;
    rd_cycle[ 3109] = 1'b1;  wr_cycle[ 3109] = 1'b0;  addr_rom[ 3109]='h00001394;  wr_data_rom[ 3109]='h00000000;
    rd_cycle[ 3110] = 1'b0;  wr_cycle[ 3110] = 1'b1;  addr_rom[ 3110]='h000010b0;  wr_data_rom[ 3110]='h0000017f;
    rd_cycle[ 3111] = 1'b0;  wr_cycle[ 3111] = 1'b1;  addr_rom[ 3111]='h00000dac;  wr_data_rom[ 3111]='h00000182;
    rd_cycle[ 3112] = 1'b1;  wr_cycle[ 3112] = 1'b0;  addr_rom[ 3112]='h000009fc;  wr_data_rom[ 3112]='h00000000;
    rd_cycle[ 3113] = 1'b1;  wr_cycle[ 3113] = 1'b0;  addr_rom[ 3113]='h00001728;  wr_data_rom[ 3113]='h00000000;
    rd_cycle[ 3114] = 1'b0;  wr_cycle[ 3114] = 1'b1;  addr_rom[ 3114]='h00000ae4;  wr_data_rom[ 3114]='h00001751;
    rd_cycle[ 3115] = 1'b1;  wr_cycle[ 3115] = 1'b0;  addr_rom[ 3115]='h0000196c;  wr_data_rom[ 3115]='h00000000;
    rd_cycle[ 3116] = 1'b0;  wr_cycle[ 3116] = 1'b1;  addr_rom[ 3116]='h0000107c;  wr_data_rom[ 3116]='h00001748;
    rd_cycle[ 3117] = 1'b1;  wr_cycle[ 3117] = 1'b0;  addr_rom[ 3117]='h000010fc;  wr_data_rom[ 3117]='h00000000;
    rd_cycle[ 3118] = 1'b0;  wr_cycle[ 3118] = 1'b1;  addr_rom[ 3118]='h00000300;  wr_data_rom[ 3118]='h000007a0;
    rd_cycle[ 3119] = 1'b1;  wr_cycle[ 3119] = 1'b0;  addr_rom[ 3119]='h00001220;  wr_data_rom[ 3119]='h00000000;
    rd_cycle[ 3120] = 1'b0;  wr_cycle[ 3120] = 1'b1;  addr_rom[ 3120]='h00000e00;  wr_data_rom[ 3120]='h0000181a;
    rd_cycle[ 3121] = 1'b1;  wr_cycle[ 3121] = 1'b0;  addr_rom[ 3121]='h00000128;  wr_data_rom[ 3121]='h00000000;
    rd_cycle[ 3122] = 1'b0;  wr_cycle[ 3122] = 1'b1;  addr_rom[ 3122]='h000005d8;  wr_data_rom[ 3122]='h000011f3;
    rd_cycle[ 3123] = 1'b1;  wr_cycle[ 3123] = 1'b0;  addr_rom[ 3123]='h000004c8;  wr_data_rom[ 3123]='h00000000;
    rd_cycle[ 3124] = 1'b1;  wr_cycle[ 3124] = 1'b0;  addr_rom[ 3124]='h000000ec;  wr_data_rom[ 3124]='h00000000;
    rd_cycle[ 3125] = 1'b0;  wr_cycle[ 3125] = 1'b1;  addr_rom[ 3125]='h00000c20;  wr_data_rom[ 3125]='h0000121c;
    rd_cycle[ 3126] = 1'b0;  wr_cycle[ 3126] = 1'b1;  addr_rom[ 3126]='h00001de8;  wr_data_rom[ 3126]='h000002d4;
    rd_cycle[ 3127] = 1'b1;  wr_cycle[ 3127] = 1'b0;  addr_rom[ 3127]='h00001338;  wr_data_rom[ 3127]='h00000000;
    rd_cycle[ 3128] = 1'b0;  wr_cycle[ 3128] = 1'b1;  addr_rom[ 3128]='h000017d0;  wr_data_rom[ 3128]='h0000116a;
    rd_cycle[ 3129] = 1'b0;  wr_cycle[ 3129] = 1'b1;  addr_rom[ 3129]='h000006ec;  wr_data_rom[ 3129]='h0000096e;
    rd_cycle[ 3130] = 1'b0;  wr_cycle[ 3130] = 1'b1;  addr_rom[ 3130]='h000001c0;  wr_data_rom[ 3130]='h0000191d;
    rd_cycle[ 3131] = 1'b1;  wr_cycle[ 3131] = 1'b0;  addr_rom[ 3131]='h0000166c;  wr_data_rom[ 3131]='h00000000;
    rd_cycle[ 3132] = 1'b1;  wr_cycle[ 3132] = 1'b0;  addr_rom[ 3132]='h000016d0;  wr_data_rom[ 3132]='h00000000;
    rd_cycle[ 3133] = 1'b0;  wr_cycle[ 3133] = 1'b1;  addr_rom[ 3133]='h00000134;  wr_data_rom[ 3133]='h000018eb;
    rd_cycle[ 3134] = 1'b0;  wr_cycle[ 3134] = 1'b1;  addr_rom[ 3134]='h00000e68;  wr_data_rom[ 3134]='h0000174b;
    rd_cycle[ 3135] = 1'b1;  wr_cycle[ 3135] = 1'b0;  addr_rom[ 3135]='h00000e88;  wr_data_rom[ 3135]='h00000000;
    rd_cycle[ 3136] = 1'b1;  wr_cycle[ 3136] = 1'b0;  addr_rom[ 3136]='h000016e4;  wr_data_rom[ 3136]='h00000000;
    rd_cycle[ 3137] = 1'b0;  wr_cycle[ 3137] = 1'b1;  addr_rom[ 3137]='h000010d0;  wr_data_rom[ 3137]='h00001e6e;
    rd_cycle[ 3138] = 1'b1;  wr_cycle[ 3138] = 1'b0;  addr_rom[ 3138]='h0000198c;  wr_data_rom[ 3138]='h00000000;
    rd_cycle[ 3139] = 1'b0;  wr_cycle[ 3139] = 1'b1;  addr_rom[ 3139]='h000015a8;  wr_data_rom[ 3139]='h00000de4;
    rd_cycle[ 3140] = 1'b1;  wr_cycle[ 3140] = 1'b0;  addr_rom[ 3140]='h00001640;  wr_data_rom[ 3140]='h00000000;
    rd_cycle[ 3141] = 1'b1;  wr_cycle[ 3141] = 1'b0;  addr_rom[ 3141]='h00001008;  wr_data_rom[ 3141]='h00000000;
    rd_cycle[ 3142] = 1'b0;  wr_cycle[ 3142] = 1'b1;  addr_rom[ 3142]='h000001c0;  wr_data_rom[ 3142]='h00000080;
    rd_cycle[ 3143] = 1'b0;  wr_cycle[ 3143] = 1'b1;  addr_rom[ 3143]='h0000127c;  wr_data_rom[ 3143]='h00001e8c;
    rd_cycle[ 3144] = 1'b0;  wr_cycle[ 3144] = 1'b1;  addr_rom[ 3144]='h00001d2c;  wr_data_rom[ 3144]='h00001a54;
    rd_cycle[ 3145] = 1'b0;  wr_cycle[ 3145] = 1'b1;  addr_rom[ 3145]='h0000048c;  wr_data_rom[ 3145]='h00001345;
    rd_cycle[ 3146] = 1'b0;  wr_cycle[ 3146] = 1'b1;  addr_rom[ 3146]='h000001c0;  wr_data_rom[ 3146]='h00000c0a;
    rd_cycle[ 3147] = 1'b1;  wr_cycle[ 3147] = 1'b0;  addr_rom[ 3147]='h00001dac;  wr_data_rom[ 3147]='h00000000;
    rd_cycle[ 3148] = 1'b1;  wr_cycle[ 3148] = 1'b0;  addr_rom[ 3148]='h00000740;  wr_data_rom[ 3148]='h00000000;
    rd_cycle[ 3149] = 1'b0;  wr_cycle[ 3149] = 1'b1;  addr_rom[ 3149]='h00000fd8;  wr_data_rom[ 3149]='h0000006d;
    rd_cycle[ 3150] = 1'b0;  wr_cycle[ 3150] = 1'b1;  addr_rom[ 3150]='h000016e0;  wr_data_rom[ 3150]='h00000648;
    rd_cycle[ 3151] = 1'b1;  wr_cycle[ 3151] = 1'b0;  addr_rom[ 3151]='h00000824;  wr_data_rom[ 3151]='h00000000;
    rd_cycle[ 3152] = 1'b0;  wr_cycle[ 3152] = 1'b1;  addr_rom[ 3152]='h00001744;  wr_data_rom[ 3152]='h00000f43;
    rd_cycle[ 3153] = 1'b0;  wr_cycle[ 3153] = 1'b1;  addr_rom[ 3153]='h000012b4;  wr_data_rom[ 3153]='h00001e20;
    rd_cycle[ 3154] = 1'b1;  wr_cycle[ 3154] = 1'b0;  addr_rom[ 3154]='h0000144c;  wr_data_rom[ 3154]='h00000000;
    rd_cycle[ 3155] = 1'b1;  wr_cycle[ 3155] = 1'b0;  addr_rom[ 3155]='h00000aa4;  wr_data_rom[ 3155]='h00000000;
    rd_cycle[ 3156] = 1'b1;  wr_cycle[ 3156] = 1'b0;  addr_rom[ 3156]='h0000017c;  wr_data_rom[ 3156]='h00000000;
    rd_cycle[ 3157] = 1'b1;  wr_cycle[ 3157] = 1'b0;  addr_rom[ 3157]='h00001dec;  wr_data_rom[ 3157]='h00000000;
    rd_cycle[ 3158] = 1'b1;  wr_cycle[ 3158] = 1'b0;  addr_rom[ 3158]='h00001bd8;  wr_data_rom[ 3158]='h00000000;
    rd_cycle[ 3159] = 1'b0;  wr_cycle[ 3159] = 1'b1;  addr_rom[ 3159]='h00001c60;  wr_data_rom[ 3159]='h00000670;
    rd_cycle[ 3160] = 1'b0;  wr_cycle[ 3160] = 1'b1;  addr_rom[ 3160]='h00000d38;  wr_data_rom[ 3160]='h00000b7f;
    rd_cycle[ 3161] = 1'b0;  wr_cycle[ 3161] = 1'b1;  addr_rom[ 3161]='h00001a84;  wr_data_rom[ 3161]='h00000987;
    rd_cycle[ 3162] = 1'b1;  wr_cycle[ 3162] = 1'b0;  addr_rom[ 3162]='h00001838;  wr_data_rom[ 3162]='h00000000;
    rd_cycle[ 3163] = 1'b1;  wr_cycle[ 3163] = 1'b0;  addr_rom[ 3163]='h000008d0;  wr_data_rom[ 3163]='h00000000;
    rd_cycle[ 3164] = 1'b0;  wr_cycle[ 3164] = 1'b1;  addr_rom[ 3164]='h000008c8;  wr_data_rom[ 3164]='h00000815;
    rd_cycle[ 3165] = 1'b0;  wr_cycle[ 3165] = 1'b1;  addr_rom[ 3165]='h0000099c;  wr_data_rom[ 3165]='h00001c96;
    rd_cycle[ 3166] = 1'b1;  wr_cycle[ 3166] = 1'b0;  addr_rom[ 3166]='h000009cc;  wr_data_rom[ 3166]='h00000000;
    rd_cycle[ 3167] = 1'b0;  wr_cycle[ 3167] = 1'b1;  addr_rom[ 3167]='h00001190;  wr_data_rom[ 3167]='h000013e3;
    rd_cycle[ 3168] = 1'b0;  wr_cycle[ 3168] = 1'b1;  addr_rom[ 3168]='h00001178;  wr_data_rom[ 3168]='h0000151f;
    rd_cycle[ 3169] = 1'b1;  wr_cycle[ 3169] = 1'b0;  addr_rom[ 3169]='h00001b7c;  wr_data_rom[ 3169]='h00000000;
    rd_cycle[ 3170] = 1'b0;  wr_cycle[ 3170] = 1'b1;  addr_rom[ 3170]='h00001184;  wr_data_rom[ 3170]='h00001635;
    rd_cycle[ 3171] = 1'b1;  wr_cycle[ 3171] = 1'b0;  addr_rom[ 3171]='h0000082c;  wr_data_rom[ 3171]='h00000000;
    rd_cycle[ 3172] = 1'b0;  wr_cycle[ 3172] = 1'b1;  addr_rom[ 3172]='h00000a6c;  wr_data_rom[ 3172]='h00001833;
    rd_cycle[ 3173] = 1'b1;  wr_cycle[ 3173] = 1'b0;  addr_rom[ 3173]='h000000d0;  wr_data_rom[ 3173]='h00000000;
    rd_cycle[ 3174] = 1'b1;  wr_cycle[ 3174] = 1'b0;  addr_rom[ 3174]='h00000454;  wr_data_rom[ 3174]='h00000000;
    rd_cycle[ 3175] = 1'b1;  wr_cycle[ 3175] = 1'b0;  addr_rom[ 3175]='h0000006c;  wr_data_rom[ 3175]='h00000000;
    rd_cycle[ 3176] = 1'b1;  wr_cycle[ 3176] = 1'b0;  addr_rom[ 3176]='h00001394;  wr_data_rom[ 3176]='h00000000;
    rd_cycle[ 3177] = 1'b0;  wr_cycle[ 3177] = 1'b1;  addr_rom[ 3177]='h000012b8;  wr_data_rom[ 3177]='h00001aac;
    rd_cycle[ 3178] = 1'b1;  wr_cycle[ 3178] = 1'b0;  addr_rom[ 3178]='h00000ef8;  wr_data_rom[ 3178]='h00000000;
    rd_cycle[ 3179] = 1'b1;  wr_cycle[ 3179] = 1'b0;  addr_rom[ 3179]='h00001ddc;  wr_data_rom[ 3179]='h00000000;
    rd_cycle[ 3180] = 1'b0;  wr_cycle[ 3180] = 1'b1;  addr_rom[ 3180]='h00001618;  wr_data_rom[ 3180]='h00000f3c;
    rd_cycle[ 3181] = 1'b0;  wr_cycle[ 3181] = 1'b1;  addr_rom[ 3181]='h0000089c;  wr_data_rom[ 3181]='h0000112c;
    rd_cycle[ 3182] = 1'b0;  wr_cycle[ 3182] = 1'b1;  addr_rom[ 3182]='h00001e74;  wr_data_rom[ 3182]='h00001de5;
    rd_cycle[ 3183] = 1'b0;  wr_cycle[ 3183] = 1'b1;  addr_rom[ 3183]='h000002a8;  wr_data_rom[ 3183]='h00001dfd;
    rd_cycle[ 3184] = 1'b1;  wr_cycle[ 3184] = 1'b0;  addr_rom[ 3184]='h00001bfc;  wr_data_rom[ 3184]='h00000000;
    rd_cycle[ 3185] = 1'b1;  wr_cycle[ 3185] = 1'b0;  addr_rom[ 3185]='h00001904;  wr_data_rom[ 3185]='h00000000;
    rd_cycle[ 3186] = 1'b0;  wr_cycle[ 3186] = 1'b1;  addr_rom[ 3186]='h000010ac;  wr_data_rom[ 3186]='h000018a5;
    rd_cycle[ 3187] = 1'b0;  wr_cycle[ 3187] = 1'b1;  addr_rom[ 3187]='h00000048;  wr_data_rom[ 3187]='h0000011e;
    rd_cycle[ 3188] = 1'b0;  wr_cycle[ 3188] = 1'b1;  addr_rom[ 3188]='h00001a10;  wr_data_rom[ 3188]='h00000606;
    rd_cycle[ 3189] = 1'b1;  wr_cycle[ 3189] = 1'b0;  addr_rom[ 3189]='h00001af4;  wr_data_rom[ 3189]='h00000000;
    rd_cycle[ 3190] = 1'b1;  wr_cycle[ 3190] = 1'b0;  addr_rom[ 3190]='h000009d8;  wr_data_rom[ 3190]='h00000000;
    rd_cycle[ 3191] = 1'b1;  wr_cycle[ 3191] = 1'b0;  addr_rom[ 3191]='h0000066c;  wr_data_rom[ 3191]='h00000000;
    rd_cycle[ 3192] = 1'b1;  wr_cycle[ 3192] = 1'b0;  addr_rom[ 3192]='h00001afc;  wr_data_rom[ 3192]='h00000000;
    rd_cycle[ 3193] = 1'b0;  wr_cycle[ 3193] = 1'b1;  addr_rom[ 3193]='h00000fe0;  wr_data_rom[ 3193]='h00000fd5;
    rd_cycle[ 3194] = 1'b0;  wr_cycle[ 3194] = 1'b1;  addr_rom[ 3194]='h00000d00;  wr_data_rom[ 3194]='h00001de4;
    rd_cycle[ 3195] = 1'b0;  wr_cycle[ 3195] = 1'b1;  addr_rom[ 3195]='h00001630;  wr_data_rom[ 3195]='h00001025;
    rd_cycle[ 3196] = 1'b0;  wr_cycle[ 3196] = 1'b1;  addr_rom[ 3196]='h000007a8;  wr_data_rom[ 3196]='h00000934;
    rd_cycle[ 3197] = 1'b0;  wr_cycle[ 3197] = 1'b1;  addr_rom[ 3197]='h00001678;  wr_data_rom[ 3197]='h00001c88;
    rd_cycle[ 3198] = 1'b0;  wr_cycle[ 3198] = 1'b1;  addr_rom[ 3198]='h000005d8;  wr_data_rom[ 3198]='h000019e1;
    rd_cycle[ 3199] = 1'b0;  wr_cycle[ 3199] = 1'b1;  addr_rom[ 3199]='h00000b14;  wr_data_rom[ 3199]='h00000ceb;
    rd_cycle[ 3200] = 1'b0;  wr_cycle[ 3200] = 1'b1;  addr_rom[ 3200]='h00001c78;  wr_data_rom[ 3200]='h00000728;
    rd_cycle[ 3201] = 1'b0;  wr_cycle[ 3201] = 1'b1;  addr_rom[ 3201]='h00001584;  wr_data_rom[ 3201]='h000004fb;
    rd_cycle[ 3202] = 1'b1;  wr_cycle[ 3202] = 1'b0;  addr_rom[ 3202]='h000013a0;  wr_data_rom[ 3202]='h00000000;
    rd_cycle[ 3203] = 1'b0;  wr_cycle[ 3203] = 1'b1;  addr_rom[ 3203]='h000017f8;  wr_data_rom[ 3203]='h000015f8;
    rd_cycle[ 3204] = 1'b1;  wr_cycle[ 3204] = 1'b0;  addr_rom[ 3204]='h000016dc;  wr_data_rom[ 3204]='h00000000;
    rd_cycle[ 3205] = 1'b1;  wr_cycle[ 3205] = 1'b0;  addr_rom[ 3205]='h00000944;  wr_data_rom[ 3205]='h00000000;
    rd_cycle[ 3206] = 1'b0;  wr_cycle[ 3206] = 1'b1;  addr_rom[ 3206]='h00000aa8;  wr_data_rom[ 3206]='h000014cc;
    rd_cycle[ 3207] = 1'b0;  wr_cycle[ 3207] = 1'b1;  addr_rom[ 3207]='h00001e7c;  wr_data_rom[ 3207]='h00001285;
    rd_cycle[ 3208] = 1'b1;  wr_cycle[ 3208] = 1'b0;  addr_rom[ 3208]='h000006ac;  wr_data_rom[ 3208]='h00000000;
    rd_cycle[ 3209] = 1'b1;  wr_cycle[ 3209] = 1'b0;  addr_rom[ 3209]='h0000025c;  wr_data_rom[ 3209]='h00000000;
    rd_cycle[ 3210] = 1'b0;  wr_cycle[ 3210] = 1'b1;  addr_rom[ 3210]='h00001360;  wr_data_rom[ 3210]='h00001155;
    rd_cycle[ 3211] = 1'b1;  wr_cycle[ 3211] = 1'b0;  addr_rom[ 3211]='h00000e44;  wr_data_rom[ 3211]='h00000000;
    rd_cycle[ 3212] = 1'b1;  wr_cycle[ 3212] = 1'b0;  addr_rom[ 3212]='h00000db4;  wr_data_rom[ 3212]='h00000000;
    rd_cycle[ 3213] = 1'b1;  wr_cycle[ 3213] = 1'b0;  addr_rom[ 3213]='h00000e24;  wr_data_rom[ 3213]='h00000000;
    rd_cycle[ 3214] = 1'b1;  wr_cycle[ 3214] = 1'b0;  addr_rom[ 3214]='h0000149c;  wr_data_rom[ 3214]='h00000000;
    rd_cycle[ 3215] = 1'b0;  wr_cycle[ 3215] = 1'b1;  addr_rom[ 3215]='h0000198c;  wr_data_rom[ 3215]='h00001ad6;
    rd_cycle[ 3216] = 1'b1;  wr_cycle[ 3216] = 1'b0;  addr_rom[ 3216]='h000014e0;  wr_data_rom[ 3216]='h00000000;
    rd_cycle[ 3217] = 1'b0;  wr_cycle[ 3217] = 1'b1;  addr_rom[ 3217]='h00000700;  wr_data_rom[ 3217]='h00000d8a;
    rd_cycle[ 3218] = 1'b1;  wr_cycle[ 3218] = 1'b0;  addr_rom[ 3218]='h0000092c;  wr_data_rom[ 3218]='h00000000;
    rd_cycle[ 3219] = 1'b0;  wr_cycle[ 3219] = 1'b1;  addr_rom[ 3219]='h00000370;  wr_data_rom[ 3219]='h000008e6;
    rd_cycle[ 3220] = 1'b0;  wr_cycle[ 3220] = 1'b1;  addr_rom[ 3220]='h00001744;  wr_data_rom[ 3220]='h00001219;
    rd_cycle[ 3221] = 1'b0;  wr_cycle[ 3221] = 1'b1;  addr_rom[ 3221]='h0000083c;  wr_data_rom[ 3221]='h00000890;
    rd_cycle[ 3222] = 1'b0;  wr_cycle[ 3222] = 1'b1;  addr_rom[ 3222]='h0000111c;  wr_data_rom[ 3222]='h00000612;
    rd_cycle[ 3223] = 1'b1;  wr_cycle[ 3223] = 1'b0;  addr_rom[ 3223]='h00001aec;  wr_data_rom[ 3223]='h00000000;
    rd_cycle[ 3224] = 1'b1;  wr_cycle[ 3224] = 1'b0;  addr_rom[ 3224]='h00001c84;  wr_data_rom[ 3224]='h00000000;
    rd_cycle[ 3225] = 1'b0;  wr_cycle[ 3225] = 1'b1;  addr_rom[ 3225]='h000001bc;  wr_data_rom[ 3225]='h00000fee;
    rd_cycle[ 3226] = 1'b0;  wr_cycle[ 3226] = 1'b1;  addr_rom[ 3226]='h00000474;  wr_data_rom[ 3226]='h0000159e;
    rd_cycle[ 3227] = 1'b1;  wr_cycle[ 3227] = 1'b0;  addr_rom[ 3227]='h000002a8;  wr_data_rom[ 3227]='h00000000;
    rd_cycle[ 3228] = 1'b1;  wr_cycle[ 3228] = 1'b0;  addr_rom[ 3228]='h00000a68;  wr_data_rom[ 3228]='h00000000;
    rd_cycle[ 3229] = 1'b0;  wr_cycle[ 3229] = 1'b1;  addr_rom[ 3229]='h00000220;  wr_data_rom[ 3229]='h00000dfa;
    rd_cycle[ 3230] = 1'b1;  wr_cycle[ 3230] = 1'b0;  addr_rom[ 3230]='h00000748;  wr_data_rom[ 3230]='h00000000;
    rd_cycle[ 3231] = 1'b0;  wr_cycle[ 3231] = 1'b1;  addr_rom[ 3231]='h0000038c;  wr_data_rom[ 3231]='h0000021f;
    rd_cycle[ 3232] = 1'b0;  wr_cycle[ 3232] = 1'b1;  addr_rom[ 3232]='h000018b4;  wr_data_rom[ 3232]='h0000135a;
    rd_cycle[ 3233] = 1'b0;  wr_cycle[ 3233] = 1'b1;  addr_rom[ 3233]='h00000284;  wr_data_rom[ 3233]='h00001252;
    rd_cycle[ 3234] = 1'b0;  wr_cycle[ 3234] = 1'b1;  addr_rom[ 3234]='h00000e44;  wr_data_rom[ 3234]='h000006c0;
    rd_cycle[ 3235] = 1'b0;  wr_cycle[ 3235] = 1'b1;  addr_rom[ 3235]='h00000858;  wr_data_rom[ 3235]='h000006de;
    rd_cycle[ 3236] = 1'b1;  wr_cycle[ 3236] = 1'b0;  addr_rom[ 3236]='h00001e64;  wr_data_rom[ 3236]='h00000000;
    rd_cycle[ 3237] = 1'b0;  wr_cycle[ 3237] = 1'b1;  addr_rom[ 3237]='h00001bd0;  wr_data_rom[ 3237]='h00000fb9;
    rd_cycle[ 3238] = 1'b0;  wr_cycle[ 3238] = 1'b1;  addr_rom[ 3238]='h0000084c;  wr_data_rom[ 3238]='h0000188f;
    rd_cycle[ 3239] = 1'b0;  wr_cycle[ 3239] = 1'b1;  addr_rom[ 3239]='h000018f4;  wr_data_rom[ 3239]='h0000140e;
    rd_cycle[ 3240] = 1'b0;  wr_cycle[ 3240] = 1'b1;  addr_rom[ 3240]='h00001e5c;  wr_data_rom[ 3240]='h00001a9d;
    rd_cycle[ 3241] = 1'b1;  wr_cycle[ 3241] = 1'b0;  addr_rom[ 3241]='h000011f8;  wr_data_rom[ 3241]='h00000000;
    rd_cycle[ 3242] = 1'b0;  wr_cycle[ 3242] = 1'b1;  addr_rom[ 3242]='h00001e88;  wr_data_rom[ 3242]='h00000442;
    rd_cycle[ 3243] = 1'b1;  wr_cycle[ 3243] = 1'b0;  addr_rom[ 3243]='h000007bc;  wr_data_rom[ 3243]='h00000000;
    rd_cycle[ 3244] = 1'b0;  wr_cycle[ 3244] = 1'b1;  addr_rom[ 3244]='h00001bdc;  wr_data_rom[ 3244]='h000013f3;
    rd_cycle[ 3245] = 1'b0;  wr_cycle[ 3245] = 1'b1;  addr_rom[ 3245]='h00000038;  wr_data_rom[ 3245]='h00000e73;
    rd_cycle[ 3246] = 1'b1;  wr_cycle[ 3246] = 1'b0;  addr_rom[ 3246]='h00001bd4;  wr_data_rom[ 3246]='h00000000;
    rd_cycle[ 3247] = 1'b0;  wr_cycle[ 3247] = 1'b1;  addr_rom[ 3247]='h00000198;  wr_data_rom[ 3247]='h00001232;
    rd_cycle[ 3248] = 1'b1;  wr_cycle[ 3248] = 1'b0;  addr_rom[ 3248]='h00000a44;  wr_data_rom[ 3248]='h00000000;
    rd_cycle[ 3249] = 1'b1;  wr_cycle[ 3249] = 1'b0;  addr_rom[ 3249]='h00001de0;  wr_data_rom[ 3249]='h00000000;
    rd_cycle[ 3250] = 1'b0;  wr_cycle[ 3250] = 1'b1;  addr_rom[ 3250]='h00000320;  wr_data_rom[ 3250]='h000008b6;
    rd_cycle[ 3251] = 1'b0;  wr_cycle[ 3251] = 1'b1;  addr_rom[ 3251]='h00000378;  wr_data_rom[ 3251]='h0000187f;
    rd_cycle[ 3252] = 1'b1;  wr_cycle[ 3252] = 1'b0;  addr_rom[ 3252]='h00001a80;  wr_data_rom[ 3252]='h00000000;
    rd_cycle[ 3253] = 1'b1;  wr_cycle[ 3253] = 1'b0;  addr_rom[ 3253]='h0000057c;  wr_data_rom[ 3253]='h00000000;
    rd_cycle[ 3254] = 1'b0;  wr_cycle[ 3254] = 1'b1;  addr_rom[ 3254]='h00000c90;  wr_data_rom[ 3254]='h0000001e;
    rd_cycle[ 3255] = 1'b1;  wr_cycle[ 3255] = 1'b0;  addr_rom[ 3255]='h0000150c;  wr_data_rom[ 3255]='h00000000;
    rd_cycle[ 3256] = 1'b0;  wr_cycle[ 3256] = 1'b1;  addr_rom[ 3256]='h00000400;  wr_data_rom[ 3256]='h0000105a;
    rd_cycle[ 3257] = 1'b0;  wr_cycle[ 3257] = 1'b1;  addr_rom[ 3257]='h00001204;  wr_data_rom[ 3257]='h000000fa;
    rd_cycle[ 3258] = 1'b0;  wr_cycle[ 3258] = 1'b1;  addr_rom[ 3258]='h000016f8;  wr_data_rom[ 3258]='h00000345;
    rd_cycle[ 3259] = 1'b0;  wr_cycle[ 3259] = 1'b1;  addr_rom[ 3259]='h000000dc;  wr_data_rom[ 3259]='h0000014e;
    rd_cycle[ 3260] = 1'b0;  wr_cycle[ 3260] = 1'b1;  addr_rom[ 3260]='h00001a04;  wr_data_rom[ 3260]='h0000007a;
    rd_cycle[ 3261] = 1'b1;  wr_cycle[ 3261] = 1'b0;  addr_rom[ 3261]='h000004e0;  wr_data_rom[ 3261]='h00000000;
    rd_cycle[ 3262] = 1'b1;  wr_cycle[ 3262] = 1'b0;  addr_rom[ 3262]='h00001cec;  wr_data_rom[ 3262]='h00000000;
    rd_cycle[ 3263] = 1'b1;  wr_cycle[ 3263] = 1'b0;  addr_rom[ 3263]='h00000914;  wr_data_rom[ 3263]='h00000000;
    rd_cycle[ 3264] = 1'b0;  wr_cycle[ 3264] = 1'b1;  addr_rom[ 3264]='h0000172c;  wr_data_rom[ 3264]='h00001b0e;
    rd_cycle[ 3265] = 1'b0;  wr_cycle[ 3265] = 1'b1;  addr_rom[ 3265]='h000005b4;  wr_data_rom[ 3265]='h00001b4d;
    rd_cycle[ 3266] = 1'b1;  wr_cycle[ 3266] = 1'b0;  addr_rom[ 3266]='h00000a38;  wr_data_rom[ 3266]='h00000000;
    rd_cycle[ 3267] = 1'b0;  wr_cycle[ 3267] = 1'b1;  addr_rom[ 3267]='h00000b08;  wr_data_rom[ 3267]='h00001e5c;
    rd_cycle[ 3268] = 1'b1;  wr_cycle[ 3268] = 1'b0;  addr_rom[ 3268]='h00001ca4;  wr_data_rom[ 3268]='h00000000;
    rd_cycle[ 3269] = 1'b0;  wr_cycle[ 3269] = 1'b1;  addr_rom[ 3269]='h00001460;  wr_data_rom[ 3269]='h00000f02;
    rd_cycle[ 3270] = 1'b1;  wr_cycle[ 3270] = 1'b0;  addr_rom[ 3270]='h00000444;  wr_data_rom[ 3270]='h00000000;
    rd_cycle[ 3271] = 1'b1;  wr_cycle[ 3271] = 1'b0;  addr_rom[ 3271]='h00001a0c;  wr_data_rom[ 3271]='h00000000;
    rd_cycle[ 3272] = 1'b1;  wr_cycle[ 3272] = 1'b0;  addr_rom[ 3272]='h00000898;  wr_data_rom[ 3272]='h00000000;
    rd_cycle[ 3273] = 1'b0;  wr_cycle[ 3273] = 1'b1;  addr_rom[ 3273]='h000008c4;  wr_data_rom[ 3273]='h00000f30;
    rd_cycle[ 3274] = 1'b0;  wr_cycle[ 3274] = 1'b1;  addr_rom[ 3274]='h0000057c;  wr_data_rom[ 3274]='h00000b52;
    rd_cycle[ 3275] = 1'b0;  wr_cycle[ 3275] = 1'b1;  addr_rom[ 3275]='h000004c0;  wr_data_rom[ 3275]='h00000deb;
    rd_cycle[ 3276] = 1'b1;  wr_cycle[ 3276] = 1'b0;  addr_rom[ 3276]='h00001a3c;  wr_data_rom[ 3276]='h00000000;
    rd_cycle[ 3277] = 1'b0;  wr_cycle[ 3277] = 1'b1;  addr_rom[ 3277]='h00001a24;  wr_data_rom[ 3277]='h00001816;
    rd_cycle[ 3278] = 1'b0;  wr_cycle[ 3278] = 1'b1;  addr_rom[ 3278]='h0000083c;  wr_data_rom[ 3278]='h000004c5;
    rd_cycle[ 3279] = 1'b0;  wr_cycle[ 3279] = 1'b1;  addr_rom[ 3279]='h00000df8;  wr_data_rom[ 3279]='h00001399;
    rd_cycle[ 3280] = 1'b0;  wr_cycle[ 3280] = 1'b1;  addr_rom[ 3280]='h00000a6c;  wr_data_rom[ 3280]='h00001d32;
    rd_cycle[ 3281] = 1'b0;  wr_cycle[ 3281] = 1'b1;  addr_rom[ 3281]='h00000858;  wr_data_rom[ 3281]='h000013fa;
    rd_cycle[ 3282] = 1'b1;  wr_cycle[ 3282] = 1'b0;  addr_rom[ 3282]='h000012f4;  wr_data_rom[ 3282]='h00000000;
    rd_cycle[ 3283] = 1'b0;  wr_cycle[ 3283] = 1'b1;  addr_rom[ 3283]='h00001ea8;  wr_data_rom[ 3283]='h00000600;
    rd_cycle[ 3284] = 1'b1;  wr_cycle[ 3284] = 1'b0;  addr_rom[ 3284]='h00000770;  wr_data_rom[ 3284]='h00000000;
    rd_cycle[ 3285] = 1'b0;  wr_cycle[ 3285] = 1'b1;  addr_rom[ 3285]='h00000c2c;  wr_data_rom[ 3285]='h00001e05;
    rd_cycle[ 3286] = 1'b0;  wr_cycle[ 3286] = 1'b1;  addr_rom[ 3286]='h00000fdc;  wr_data_rom[ 3286]='h00001261;
    rd_cycle[ 3287] = 1'b1;  wr_cycle[ 3287] = 1'b0;  addr_rom[ 3287]='h00001e0c;  wr_data_rom[ 3287]='h00000000;
    rd_cycle[ 3288] = 1'b1;  wr_cycle[ 3288] = 1'b0;  addr_rom[ 3288]='h00000d34;  wr_data_rom[ 3288]='h00000000;
    rd_cycle[ 3289] = 1'b0;  wr_cycle[ 3289] = 1'b1;  addr_rom[ 3289]='h00001470;  wr_data_rom[ 3289]='h00001c93;
    rd_cycle[ 3290] = 1'b0;  wr_cycle[ 3290] = 1'b1;  addr_rom[ 3290]='h000012e0;  wr_data_rom[ 3290]='h0000031f;
    rd_cycle[ 3291] = 1'b1;  wr_cycle[ 3291] = 1'b0;  addr_rom[ 3291]='h00001f28;  wr_data_rom[ 3291]='h00000000;
    rd_cycle[ 3292] = 1'b0;  wr_cycle[ 3292] = 1'b1;  addr_rom[ 3292]='h0000102c;  wr_data_rom[ 3292]='h00001c05;
    rd_cycle[ 3293] = 1'b0;  wr_cycle[ 3293] = 1'b1;  addr_rom[ 3293]='h00001adc;  wr_data_rom[ 3293]='h00001e22;
    rd_cycle[ 3294] = 1'b0;  wr_cycle[ 3294] = 1'b1;  addr_rom[ 3294]='h00001864;  wr_data_rom[ 3294]='h00000916;
    rd_cycle[ 3295] = 1'b0;  wr_cycle[ 3295] = 1'b1;  addr_rom[ 3295]='h000001b4;  wr_data_rom[ 3295]='h00000629;
    rd_cycle[ 3296] = 1'b1;  wr_cycle[ 3296] = 1'b0;  addr_rom[ 3296]='h0000142c;  wr_data_rom[ 3296]='h00000000;
    rd_cycle[ 3297] = 1'b1;  wr_cycle[ 3297] = 1'b0;  addr_rom[ 3297]='h00001b3c;  wr_data_rom[ 3297]='h00000000;
    rd_cycle[ 3298] = 1'b0;  wr_cycle[ 3298] = 1'b1;  addr_rom[ 3298]='h00000ad8;  wr_data_rom[ 3298]='h00001df0;
    rd_cycle[ 3299] = 1'b0;  wr_cycle[ 3299] = 1'b1;  addr_rom[ 3299]='h00001e30;  wr_data_rom[ 3299]='h00001d2e;
    rd_cycle[ 3300] = 1'b1;  wr_cycle[ 3300] = 1'b0;  addr_rom[ 3300]='h00000e44;  wr_data_rom[ 3300]='h00000000;
    rd_cycle[ 3301] = 1'b0;  wr_cycle[ 3301] = 1'b1;  addr_rom[ 3301]='h00001704;  wr_data_rom[ 3301]='h00000749;
    rd_cycle[ 3302] = 1'b0;  wr_cycle[ 3302] = 1'b1;  addr_rom[ 3302]='h00000370;  wr_data_rom[ 3302]='h00000cb6;
    rd_cycle[ 3303] = 1'b0;  wr_cycle[ 3303] = 1'b1;  addr_rom[ 3303]='h000015bc;  wr_data_rom[ 3303]='h000009f8;
    rd_cycle[ 3304] = 1'b0;  wr_cycle[ 3304] = 1'b1;  addr_rom[ 3304]='h00001430;  wr_data_rom[ 3304]='h00001d38;
    rd_cycle[ 3305] = 1'b0;  wr_cycle[ 3305] = 1'b1;  addr_rom[ 3305]='h0000176c;  wr_data_rom[ 3305]='h000006d6;
    rd_cycle[ 3306] = 1'b0;  wr_cycle[ 3306] = 1'b1;  addr_rom[ 3306]='h0000171c;  wr_data_rom[ 3306]='h00001130;
    rd_cycle[ 3307] = 1'b1;  wr_cycle[ 3307] = 1'b0;  addr_rom[ 3307]='h00000f80;  wr_data_rom[ 3307]='h00000000;
    rd_cycle[ 3308] = 1'b1;  wr_cycle[ 3308] = 1'b0;  addr_rom[ 3308]='h000007fc;  wr_data_rom[ 3308]='h00000000;
    rd_cycle[ 3309] = 1'b0;  wr_cycle[ 3309] = 1'b1;  addr_rom[ 3309]='h00001c58;  wr_data_rom[ 3309]='h000010d2;
    rd_cycle[ 3310] = 1'b1;  wr_cycle[ 3310] = 1'b0;  addr_rom[ 3310]='h00000734;  wr_data_rom[ 3310]='h00000000;
    rd_cycle[ 3311] = 1'b1;  wr_cycle[ 3311] = 1'b0;  addr_rom[ 3311]='h00001ca8;  wr_data_rom[ 3311]='h00000000;
    rd_cycle[ 3312] = 1'b0;  wr_cycle[ 3312] = 1'b1;  addr_rom[ 3312]='h00001be4;  wr_data_rom[ 3312]='h0000190d;
    rd_cycle[ 3313] = 1'b1;  wr_cycle[ 3313] = 1'b0;  addr_rom[ 3313]='h00001b1c;  wr_data_rom[ 3313]='h00000000;
    rd_cycle[ 3314] = 1'b0;  wr_cycle[ 3314] = 1'b1;  addr_rom[ 3314]='h00000334;  wr_data_rom[ 3314]='h000009d0;
    rd_cycle[ 3315] = 1'b1;  wr_cycle[ 3315] = 1'b0;  addr_rom[ 3315]='h00000ea0;  wr_data_rom[ 3315]='h00000000;
    rd_cycle[ 3316] = 1'b0;  wr_cycle[ 3316] = 1'b1;  addr_rom[ 3316]='h00000efc;  wr_data_rom[ 3316]='h000014eb;
    rd_cycle[ 3317] = 1'b0;  wr_cycle[ 3317] = 1'b1;  addr_rom[ 3317]='h00001400;  wr_data_rom[ 3317]='h00000e89;
    rd_cycle[ 3318] = 1'b1;  wr_cycle[ 3318] = 1'b0;  addr_rom[ 3318]='h000000b4;  wr_data_rom[ 3318]='h00000000;
    rd_cycle[ 3319] = 1'b1;  wr_cycle[ 3319] = 1'b0;  addr_rom[ 3319]='h00000c14;  wr_data_rom[ 3319]='h00000000;
    rd_cycle[ 3320] = 1'b0;  wr_cycle[ 3320] = 1'b1;  addr_rom[ 3320]='h000002c0;  wr_data_rom[ 3320]='h00001e54;
    rd_cycle[ 3321] = 1'b0;  wr_cycle[ 3321] = 1'b1;  addr_rom[ 3321]='h00000894;  wr_data_rom[ 3321]='h00001017;
    rd_cycle[ 3322] = 1'b1;  wr_cycle[ 3322] = 1'b0;  addr_rom[ 3322]='h00000288;  wr_data_rom[ 3322]='h00000000;
    rd_cycle[ 3323] = 1'b0;  wr_cycle[ 3323] = 1'b1;  addr_rom[ 3323]='h000002c8;  wr_data_rom[ 3323]='h00000dfe;
    rd_cycle[ 3324] = 1'b1;  wr_cycle[ 3324] = 1'b0;  addr_rom[ 3324]='h00000290;  wr_data_rom[ 3324]='h00000000;
    rd_cycle[ 3325] = 1'b0;  wr_cycle[ 3325] = 1'b1;  addr_rom[ 3325]='h00001474;  wr_data_rom[ 3325]='h000005d7;
    rd_cycle[ 3326] = 1'b1;  wr_cycle[ 3326] = 1'b0;  addr_rom[ 3326]='h000000c4;  wr_data_rom[ 3326]='h00000000;
    rd_cycle[ 3327] = 1'b0;  wr_cycle[ 3327] = 1'b1;  addr_rom[ 3327]='h00001bdc;  wr_data_rom[ 3327]='h00000c15;
    rd_cycle[ 3328] = 1'b1;  wr_cycle[ 3328] = 1'b0;  addr_rom[ 3328]='h000004b0;  wr_data_rom[ 3328]='h00000000;
    rd_cycle[ 3329] = 1'b0;  wr_cycle[ 3329] = 1'b1;  addr_rom[ 3329]='h000008e4;  wr_data_rom[ 3329]='h00001414;
    rd_cycle[ 3330] = 1'b0;  wr_cycle[ 3330] = 1'b1;  addr_rom[ 3330]='h0000172c;  wr_data_rom[ 3330]='h000017c5;
    rd_cycle[ 3331] = 1'b0;  wr_cycle[ 3331] = 1'b1;  addr_rom[ 3331]='h00001de8;  wr_data_rom[ 3331]='h00000083;
    rd_cycle[ 3332] = 1'b0;  wr_cycle[ 3332] = 1'b1;  addr_rom[ 3332]='h0000133c;  wr_data_rom[ 3332]='h00001a01;
    rd_cycle[ 3333] = 1'b1;  wr_cycle[ 3333] = 1'b0;  addr_rom[ 3333]='h000012dc;  wr_data_rom[ 3333]='h00000000;
    rd_cycle[ 3334] = 1'b0;  wr_cycle[ 3334] = 1'b1;  addr_rom[ 3334]='h0000183c;  wr_data_rom[ 3334]='h0000075f;
    rd_cycle[ 3335] = 1'b0;  wr_cycle[ 3335] = 1'b1;  addr_rom[ 3335]='h00001160;  wr_data_rom[ 3335]='h00000a39;
    rd_cycle[ 3336] = 1'b1;  wr_cycle[ 3336] = 1'b0;  addr_rom[ 3336]='h00001d24;  wr_data_rom[ 3336]='h00000000;
    rd_cycle[ 3337] = 1'b1;  wr_cycle[ 3337] = 1'b0;  addr_rom[ 3337]='h00001bec;  wr_data_rom[ 3337]='h00000000;
    rd_cycle[ 3338] = 1'b0;  wr_cycle[ 3338] = 1'b1;  addr_rom[ 3338]='h0000089c;  wr_data_rom[ 3338]='h00001e8d;
    rd_cycle[ 3339] = 1'b1;  wr_cycle[ 3339] = 1'b0;  addr_rom[ 3339]='h000012f8;  wr_data_rom[ 3339]='h00000000;
    rd_cycle[ 3340] = 1'b1;  wr_cycle[ 3340] = 1'b0;  addr_rom[ 3340]='h00001418;  wr_data_rom[ 3340]='h00000000;
    rd_cycle[ 3341] = 1'b1;  wr_cycle[ 3341] = 1'b0;  addr_rom[ 3341]='h00001b5c;  wr_data_rom[ 3341]='h00000000;
    rd_cycle[ 3342] = 1'b1;  wr_cycle[ 3342] = 1'b0;  addr_rom[ 3342]='h00001e6c;  wr_data_rom[ 3342]='h00000000;
    rd_cycle[ 3343] = 1'b1;  wr_cycle[ 3343] = 1'b0;  addr_rom[ 3343]='h0000123c;  wr_data_rom[ 3343]='h00000000;
    rd_cycle[ 3344] = 1'b1;  wr_cycle[ 3344] = 1'b0;  addr_rom[ 3344]='h00000408;  wr_data_rom[ 3344]='h00000000;
    rd_cycle[ 3345] = 1'b1;  wr_cycle[ 3345] = 1'b0;  addr_rom[ 3345]='h000015c4;  wr_data_rom[ 3345]='h00000000;
    rd_cycle[ 3346] = 1'b1;  wr_cycle[ 3346] = 1'b0;  addr_rom[ 3346]='h000001e0;  wr_data_rom[ 3346]='h00000000;
    rd_cycle[ 3347] = 1'b0;  wr_cycle[ 3347] = 1'b1;  addr_rom[ 3347]='h00000160;  wr_data_rom[ 3347]='h000006ae;
    rd_cycle[ 3348] = 1'b1;  wr_cycle[ 3348] = 1'b0;  addr_rom[ 3348]='h00000284;  wr_data_rom[ 3348]='h00000000;
    rd_cycle[ 3349] = 1'b1;  wr_cycle[ 3349] = 1'b0;  addr_rom[ 3349]='h000004a0;  wr_data_rom[ 3349]='h00000000;
    rd_cycle[ 3350] = 1'b0;  wr_cycle[ 3350] = 1'b1;  addr_rom[ 3350]='h00001608;  wr_data_rom[ 3350]='h00000e50;
    rd_cycle[ 3351] = 1'b1;  wr_cycle[ 3351] = 1'b0;  addr_rom[ 3351]='h00000a6c;  wr_data_rom[ 3351]='h00000000;
    rd_cycle[ 3352] = 1'b0;  wr_cycle[ 3352] = 1'b1;  addr_rom[ 3352]='h00001920;  wr_data_rom[ 3352]='h00000fa2;
    rd_cycle[ 3353] = 1'b1;  wr_cycle[ 3353] = 1'b0;  addr_rom[ 3353]='h00001f14;  wr_data_rom[ 3353]='h00000000;
    rd_cycle[ 3354] = 1'b1;  wr_cycle[ 3354] = 1'b0;  addr_rom[ 3354]='h000010b8;  wr_data_rom[ 3354]='h00000000;
    rd_cycle[ 3355] = 1'b0;  wr_cycle[ 3355] = 1'b1;  addr_rom[ 3355]='h000013d4;  wr_data_rom[ 3355]='h000001c8;
    rd_cycle[ 3356] = 1'b1;  wr_cycle[ 3356] = 1'b0;  addr_rom[ 3356]='h00000244;  wr_data_rom[ 3356]='h00000000;
    rd_cycle[ 3357] = 1'b1;  wr_cycle[ 3357] = 1'b0;  addr_rom[ 3357]='h00001e60;  wr_data_rom[ 3357]='h00000000;
    rd_cycle[ 3358] = 1'b0;  wr_cycle[ 3358] = 1'b1;  addr_rom[ 3358]='h00001a00;  wr_data_rom[ 3358]='h00001878;
    rd_cycle[ 3359] = 1'b0;  wr_cycle[ 3359] = 1'b1;  addr_rom[ 3359]='h00001440;  wr_data_rom[ 3359]='h00001a4d;
    rd_cycle[ 3360] = 1'b1;  wr_cycle[ 3360] = 1'b0;  addr_rom[ 3360]='h000017fc;  wr_data_rom[ 3360]='h00000000;
    rd_cycle[ 3361] = 1'b0;  wr_cycle[ 3361] = 1'b1;  addr_rom[ 3361]='h0000030c;  wr_data_rom[ 3361]='h00000d6c;
    rd_cycle[ 3362] = 1'b0;  wr_cycle[ 3362] = 1'b1;  addr_rom[ 3362]='h00000298;  wr_data_rom[ 3362]='h00000325;
    rd_cycle[ 3363] = 1'b0;  wr_cycle[ 3363] = 1'b1;  addr_rom[ 3363]='h00000bb4;  wr_data_rom[ 3363]='h0000040d;
    rd_cycle[ 3364] = 1'b1;  wr_cycle[ 3364] = 1'b0;  addr_rom[ 3364]='h00000964;  wr_data_rom[ 3364]='h00000000;
    rd_cycle[ 3365] = 1'b1;  wr_cycle[ 3365] = 1'b0;  addr_rom[ 3365]='h00001ab4;  wr_data_rom[ 3365]='h00000000;
    rd_cycle[ 3366] = 1'b0;  wr_cycle[ 3366] = 1'b1;  addr_rom[ 3366]='h000001e8;  wr_data_rom[ 3366]='h00000137;
    rd_cycle[ 3367] = 1'b1;  wr_cycle[ 3367] = 1'b0;  addr_rom[ 3367]='h000014b4;  wr_data_rom[ 3367]='h00000000;
    rd_cycle[ 3368] = 1'b1;  wr_cycle[ 3368] = 1'b0;  addr_rom[ 3368]='h00001e3c;  wr_data_rom[ 3368]='h00000000;
    rd_cycle[ 3369] = 1'b0;  wr_cycle[ 3369] = 1'b1;  addr_rom[ 3369]='h000009ac;  wr_data_rom[ 3369]='h00001bf8;
    rd_cycle[ 3370] = 1'b0;  wr_cycle[ 3370] = 1'b1;  addr_rom[ 3370]='h00001a1c;  wr_data_rom[ 3370]='h00001044;
    rd_cycle[ 3371] = 1'b1;  wr_cycle[ 3371] = 1'b0;  addr_rom[ 3371]='h00000d5c;  wr_data_rom[ 3371]='h00000000;
    rd_cycle[ 3372] = 1'b0;  wr_cycle[ 3372] = 1'b1;  addr_rom[ 3372]='h000002a0;  wr_data_rom[ 3372]='h00000272;
    rd_cycle[ 3373] = 1'b0;  wr_cycle[ 3373] = 1'b1;  addr_rom[ 3373]='h00000494;  wr_data_rom[ 3373]='h00001132;
    rd_cycle[ 3374] = 1'b0;  wr_cycle[ 3374] = 1'b1;  addr_rom[ 3374]='h00000f54;  wr_data_rom[ 3374]='h000007aa;
    rd_cycle[ 3375] = 1'b0;  wr_cycle[ 3375] = 1'b1;  addr_rom[ 3375]='h00000964;  wr_data_rom[ 3375]='h00000379;
    rd_cycle[ 3376] = 1'b1;  wr_cycle[ 3376] = 1'b0;  addr_rom[ 3376]='h00001a68;  wr_data_rom[ 3376]='h00000000;
    rd_cycle[ 3377] = 1'b0;  wr_cycle[ 3377] = 1'b1;  addr_rom[ 3377]='h00001758;  wr_data_rom[ 3377]='h000011ae;
    rd_cycle[ 3378] = 1'b0;  wr_cycle[ 3378] = 1'b1;  addr_rom[ 3378]='h00001250;  wr_data_rom[ 3378]='h00000388;
    rd_cycle[ 3379] = 1'b0;  wr_cycle[ 3379] = 1'b1;  addr_rom[ 3379]='h0000127c;  wr_data_rom[ 3379]='h000001f6;
    rd_cycle[ 3380] = 1'b0;  wr_cycle[ 3380] = 1'b1;  addr_rom[ 3380]='h00000598;  wr_data_rom[ 3380]='h000009c9;
    rd_cycle[ 3381] = 1'b0;  wr_cycle[ 3381] = 1'b1;  addr_rom[ 3381]='h00001aa4;  wr_data_rom[ 3381]='h00001a41;
    rd_cycle[ 3382] = 1'b0;  wr_cycle[ 3382] = 1'b1;  addr_rom[ 3382]='h00001864;  wr_data_rom[ 3382]='h0000162f;
    rd_cycle[ 3383] = 1'b1;  wr_cycle[ 3383] = 1'b0;  addr_rom[ 3383]='h00000cf0;  wr_data_rom[ 3383]='h00000000;
    rd_cycle[ 3384] = 1'b0;  wr_cycle[ 3384] = 1'b1;  addr_rom[ 3384]='h00000480;  wr_data_rom[ 3384]='h0000172a;
    rd_cycle[ 3385] = 1'b1;  wr_cycle[ 3385] = 1'b0;  addr_rom[ 3385]='h000005c4;  wr_data_rom[ 3385]='h00000000;
    rd_cycle[ 3386] = 1'b0;  wr_cycle[ 3386] = 1'b1;  addr_rom[ 3386]='h00001d68;  wr_data_rom[ 3386]='h00001900;
    rd_cycle[ 3387] = 1'b1;  wr_cycle[ 3387] = 1'b0;  addr_rom[ 3387]='h000006ec;  wr_data_rom[ 3387]='h00000000;
    rd_cycle[ 3388] = 1'b0;  wr_cycle[ 3388] = 1'b1;  addr_rom[ 3388]='h00001cc4;  wr_data_rom[ 3388]='h0000049f;
    rd_cycle[ 3389] = 1'b1;  wr_cycle[ 3389] = 1'b0;  addr_rom[ 3389]='h000008cc;  wr_data_rom[ 3389]='h00000000;
    rd_cycle[ 3390] = 1'b1;  wr_cycle[ 3390] = 1'b0;  addr_rom[ 3390]='h000018fc;  wr_data_rom[ 3390]='h00000000;
    rd_cycle[ 3391] = 1'b1;  wr_cycle[ 3391] = 1'b0;  addr_rom[ 3391]='h00001694;  wr_data_rom[ 3391]='h00000000;
    rd_cycle[ 3392] = 1'b1;  wr_cycle[ 3392] = 1'b0;  addr_rom[ 3392]='h00000bd8;  wr_data_rom[ 3392]='h00000000;
    rd_cycle[ 3393] = 1'b1;  wr_cycle[ 3393] = 1'b0;  addr_rom[ 3393]='h00001e78;  wr_data_rom[ 3393]='h00000000;
    rd_cycle[ 3394] = 1'b1;  wr_cycle[ 3394] = 1'b0;  addr_rom[ 3394]='h00000b7c;  wr_data_rom[ 3394]='h00000000;
    rd_cycle[ 3395] = 1'b0;  wr_cycle[ 3395] = 1'b1;  addr_rom[ 3395]='h00000068;  wr_data_rom[ 3395]='h000011ae;
    rd_cycle[ 3396] = 1'b1;  wr_cycle[ 3396] = 1'b0;  addr_rom[ 3396]='h00000d00;  wr_data_rom[ 3396]='h00000000;
    rd_cycle[ 3397] = 1'b0;  wr_cycle[ 3397] = 1'b1;  addr_rom[ 3397]='h00000450;  wr_data_rom[ 3397]='h00001370;
    rd_cycle[ 3398] = 1'b1;  wr_cycle[ 3398] = 1'b0;  addr_rom[ 3398]='h00000954;  wr_data_rom[ 3398]='h00000000;
    rd_cycle[ 3399] = 1'b0;  wr_cycle[ 3399] = 1'b1;  addr_rom[ 3399]='h00000528;  wr_data_rom[ 3399]='h00001970;
    rd_cycle[ 3400] = 1'b0;  wr_cycle[ 3400] = 1'b1;  addr_rom[ 3400]='h00000874;  wr_data_rom[ 3400]='h00000c3c;
    rd_cycle[ 3401] = 1'b1;  wr_cycle[ 3401] = 1'b0;  addr_rom[ 3401]='h00000760;  wr_data_rom[ 3401]='h00000000;
    rd_cycle[ 3402] = 1'b1;  wr_cycle[ 3402] = 1'b0;  addr_rom[ 3402]='h00000f5c;  wr_data_rom[ 3402]='h00000000;
    rd_cycle[ 3403] = 1'b0;  wr_cycle[ 3403] = 1'b1;  addr_rom[ 3403]='h000009b8;  wr_data_rom[ 3403]='h000009fe;
    rd_cycle[ 3404] = 1'b0;  wr_cycle[ 3404] = 1'b1;  addr_rom[ 3404]='h00000250;  wr_data_rom[ 3404]='h00000548;
    rd_cycle[ 3405] = 1'b0;  wr_cycle[ 3405] = 1'b1;  addr_rom[ 3405]='h000005cc;  wr_data_rom[ 3405]='h00000f53;
    rd_cycle[ 3406] = 1'b1;  wr_cycle[ 3406] = 1'b0;  addr_rom[ 3406]='h000016fc;  wr_data_rom[ 3406]='h00000000;
    rd_cycle[ 3407] = 1'b1;  wr_cycle[ 3407] = 1'b0;  addr_rom[ 3407]='h000007e8;  wr_data_rom[ 3407]='h00000000;
    rd_cycle[ 3408] = 1'b0;  wr_cycle[ 3408] = 1'b1;  addr_rom[ 3408]='h0000117c;  wr_data_rom[ 3408]='h0000095b;
    rd_cycle[ 3409] = 1'b0;  wr_cycle[ 3409] = 1'b1;  addr_rom[ 3409]='h00000f58;  wr_data_rom[ 3409]='h0000045b;
    rd_cycle[ 3410] = 1'b1;  wr_cycle[ 3410] = 1'b0;  addr_rom[ 3410]='h00001150;  wr_data_rom[ 3410]='h00000000;
    rd_cycle[ 3411] = 1'b0;  wr_cycle[ 3411] = 1'b1;  addr_rom[ 3411]='h00001b6c;  wr_data_rom[ 3411]='h00001350;
    rd_cycle[ 3412] = 1'b0;  wr_cycle[ 3412] = 1'b1;  addr_rom[ 3412]='h0000145c;  wr_data_rom[ 3412]='h0000082b;
    rd_cycle[ 3413] = 1'b1;  wr_cycle[ 3413] = 1'b0;  addr_rom[ 3413]='h00000f20;  wr_data_rom[ 3413]='h00000000;
    rd_cycle[ 3414] = 1'b0;  wr_cycle[ 3414] = 1'b1;  addr_rom[ 3414]='h0000107c;  wr_data_rom[ 3414]='h00000668;
    rd_cycle[ 3415] = 1'b0;  wr_cycle[ 3415] = 1'b1;  addr_rom[ 3415]='h00001928;  wr_data_rom[ 3415]='h00001557;
    rd_cycle[ 3416] = 1'b1;  wr_cycle[ 3416] = 1'b0;  addr_rom[ 3416]='h00000888;  wr_data_rom[ 3416]='h00000000;
    rd_cycle[ 3417] = 1'b1;  wr_cycle[ 3417] = 1'b0;  addr_rom[ 3417]='h00001990;  wr_data_rom[ 3417]='h00000000;
    rd_cycle[ 3418] = 1'b0;  wr_cycle[ 3418] = 1'b1;  addr_rom[ 3418]='h00001af8;  wr_data_rom[ 3418]='h000000fe;
    rd_cycle[ 3419] = 1'b1;  wr_cycle[ 3419] = 1'b0;  addr_rom[ 3419]='h0000155c;  wr_data_rom[ 3419]='h00000000;
    rd_cycle[ 3420] = 1'b1;  wr_cycle[ 3420] = 1'b0;  addr_rom[ 3420]='h00000228;  wr_data_rom[ 3420]='h00000000;
    rd_cycle[ 3421] = 1'b1;  wr_cycle[ 3421] = 1'b0;  addr_rom[ 3421]='h00000590;  wr_data_rom[ 3421]='h00000000;
    rd_cycle[ 3422] = 1'b1;  wr_cycle[ 3422] = 1'b0;  addr_rom[ 3422]='h0000129c;  wr_data_rom[ 3422]='h00000000;
    rd_cycle[ 3423] = 1'b1;  wr_cycle[ 3423] = 1'b0;  addr_rom[ 3423]='h00000a28;  wr_data_rom[ 3423]='h00000000;
    rd_cycle[ 3424] = 1'b1;  wr_cycle[ 3424] = 1'b0;  addr_rom[ 3424]='h000008cc;  wr_data_rom[ 3424]='h00000000;
    rd_cycle[ 3425] = 1'b0;  wr_cycle[ 3425] = 1'b1;  addr_rom[ 3425]='h0000026c;  wr_data_rom[ 3425]='h00000d92;
    rd_cycle[ 3426] = 1'b0;  wr_cycle[ 3426] = 1'b1;  addr_rom[ 3426]='h00000158;  wr_data_rom[ 3426]='h00000315;
    rd_cycle[ 3427] = 1'b0;  wr_cycle[ 3427] = 1'b1;  addr_rom[ 3427]='h0000095c;  wr_data_rom[ 3427]='h00001a4d;
    rd_cycle[ 3428] = 1'b0;  wr_cycle[ 3428] = 1'b1;  addr_rom[ 3428]='h00001538;  wr_data_rom[ 3428]='h00000dab;
    rd_cycle[ 3429] = 1'b1;  wr_cycle[ 3429] = 1'b0;  addr_rom[ 3429]='h00001e00;  wr_data_rom[ 3429]='h00000000;
    rd_cycle[ 3430] = 1'b0;  wr_cycle[ 3430] = 1'b1;  addr_rom[ 3430]='h00001348;  wr_data_rom[ 3430]='h00001127;
    rd_cycle[ 3431] = 1'b0;  wr_cycle[ 3431] = 1'b1;  addr_rom[ 3431]='h00001024;  wr_data_rom[ 3431]='h00001df6;
    rd_cycle[ 3432] = 1'b1;  wr_cycle[ 3432] = 1'b0;  addr_rom[ 3432]='h00000b40;  wr_data_rom[ 3432]='h00000000;
    rd_cycle[ 3433] = 1'b0;  wr_cycle[ 3433] = 1'b1;  addr_rom[ 3433]='h00000450;  wr_data_rom[ 3433]='h00001af1;
    rd_cycle[ 3434] = 1'b1;  wr_cycle[ 3434] = 1'b0;  addr_rom[ 3434]='h00000700;  wr_data_rom[ 3434]='h00000000;
    rd_cycle[ 3435] = 1'b0;  wr_cycle[ 3435] = 1'b1;  addr_rom[ 3435]='h000006d8;  wr_data_rom[ 3435]='h0000008b;
    rd_cycle[ 3436] = 1'b0;  wr_cycle[ 3436] = 1'b1;  addr_rom[ 3436]='h000015cc;  wr_data_rom[ 3436]='h0000030d;
    rd_cycle[ 3437] = 1'b1;  wr_cycle[ 3437] = 1'b0;  addr_rom[ 3437]='h000019c4;  wr_data_rom[ 3437]='h00000000;
    rd_cycle[ 3438] = 1'b0;  wr_cycle[ 3438] = 1'b1;  addr_rom[ 3438]='h00001b58;  wr_data_rom[ 3438]='h00000cbc;
    rd_cycle[ 3439] = 1'b0;  wr_cycle[ 3439] = 1'b1;  addr_rom[ 3439]='h00001b44;  wr_data_rom[ 3439]='h0000012e;
    rd_cycle[ 3440] = 1'b0;  wr_cycle[ 3440] = 1'b1;  addr_rom[ 3440]='h000014b8;  wr_data_rom[ 3440]='h00001d88;
    rd_cycle[ 3441] = 1'b0;  wr_cycle[ 3441] = 1'b1;  addr_rom[ 3441]='h000015cc;  wr_data_rom[ 3441]='h0000022b;
    rd_cycle[ 3442] = 1'b0;  wr_cycle[ 3442] = 1'b1;  addr_rom[ 3442]='h00000dc8;  wr_data_rom[ 3442]='h0000044a;
    rd_cycle[ 3443] = 1'b0;  wr_cycle[ 3443] = 1'b1;  addr_rom[ 3443]='h00000950;  wr_data_rom[ 3443]='h000002ee;
    rd_cycle[ 3444] = 1'b1;  wr_cycle[ 3444] = 1'b0;  addr_rom[ 3444]='h000001f8;  wr_data_rom[ 3444]='h00000000;
    rd_cycle[ 3445] = 1'b0;  wr_cycle[ 3445] = 1'b1;  addr_rom[ 3445]='h00001960;  wr_data_rom[ 3445]='h0000001c;
    rd_cycle[ 3446] = 1'b0;  wr_cycle[ 3446] = 1'b1;  addr_rom[ 3446]='h0000074c;  wr_data_rom[ 3446]='h00001dd4;
    rd_cycle[ 3447] = 1'b1;  wr_cycle[ 3447] = 1'b0;  addr_rom[ 3447]='h00000a4c;  wr_data_rom[ 3447]='h00000000;
    rd_cycle[ 3448] = 1'b1;  wr_cycle[ 3448] = 1'b0;  addr_rom[ 3448]='h000005f4;  wr_data_rom[ 3448]='h00000000;
    rd_cycle[ 3449] = 1'b0;  wr_cycle[ 3449] = 1'b1;  addr_rom[ 3449]='h000006f4;  wr_data_rom[ 3449]='h0000148d;
    rd_cycle[ 3450] = 1'b0;  wr_cycle[ 3450] = 1'b1;  addr_rom[ 3450]='h0000019c;  wr_data_rom[ 3450]='h00000370;
    rd_cycle[ 3451] = 1'b1;  wr_cycle[ 3451] = 1'b0;  addr_rom[ 3451]='h00000db0;  wr_data_rom[ 3451]='h00000000;
    rd_cycle[ 3452] = 1'b0;  wr_cycle[ 3452] = 1'b1;  addr_rom[ 3452]='h00001798;  wr_data_rom[ 3452]='h000011e3;
    rd_cycle[ 3453] = 1'b0;  wr_cycle[ 3453] = 1'b1;  addr_rom[ 3453]='h000018a8;  wr_data_rom[ 3453]='h0000091f;
    rd_cycle[ 3454] = 1'b1;  wr_cycle[ 3454] = 1'b0;  addr_rom[ 3454]='h00000cb8;  wr_data_rom[ 3454]='h00000000;
    rd_cycle[ 3455] = 1'b1;  wr_cycle[ 3455] = 1'b0;  addr_rom[ 3455]='h00001b68;  wr_data_rom[ 3455]='h00000000;
    rd_cycle[ 3456] = 1'b1;  wr_cycle[ 3456] = 1'b0;  addr_rom[ 3456]='h00001954;  wr_data_rom[ 3456]='h00000000;
    rd_cycle[ 3457] = 1'b1;  wr_cycle[ 3457] = 1'b0;  addr_rom[ 3457]='h000004b8;  wr_data_rom[ 3457]='h00000000;
    rd_cycle[ 3458] = 1'b1;  wr_cycle[ 3458] = 1'b0;  addr_rom[ 3458]='h00000144;  wr_data_rom[ 3458]='h00000000;
    rd_cycle[ 3459] = 1'b0;  wr_cycle[ 3459] = 1'b1;  addr_rom[ 3459]='h000019b0;  wr_data_rom[ 3459]='h0000169e;
    rd_cycle[ 3460] = 1'b0;  wr_cycle[ 3460] = 1'b1;  addr_rom[ 3460]='h00001544;  wr_data_rom[ 3460]='h00001893;
    rd_cycle[ 3461] = 1'b0;  wr_cycle[ 3461] = 1'b1;  addr_rom[ 3461]='h000003ec;  wr_data_rom[ 3461]='h000001b4;
    rd_cycle[ 3462] = 1'b0;  wr_cycle[ 3462] = 1'b1;  addr_rom[ 3462]='h00000cdc;  wr_data_rom[ 3462]='h000017cf;
    rd_cycle[ 3463] = 1'b0;  wr_cycle[ 3463] = 1'b1;  addr_rom[ 3463]='h00000d7c;  wr_data_rom[ 3463]='h00000a6c;
    rd_cycle[ 3464] = 1'b1;  wr_cycle[ 3464] = 1'b0;  addr_rom[ 3464]='h000006d8;  wr_data_rom[ 3464]='h00000000;
    rd_cycle[ 3465] = 1'b1;  wr_cycle[ 3465] = 1'b0;  addr_rom[ 3465]='h00000514;  wr_data_rom[ 3465]='h00000000;
    rd_cycle[ 3466] = 1'b1;  wr_cycle[ 3466] = 1'b0;  addr_rom[ 3466]='h00001f2c;  wr_data_rom[ 3466]='h00000000;
    rd_cycle[ 3467] = 1'b1;  wr_cycle[ 3467] = 1'b0;  addr_rom[ 3467]='h000012fc;  wr_data_rom[ 3467]='h00000000;
    rd_cycle[ 3468] = 1'b0;  wr_cycle[ 3468] = 1'b1;  addr_rom[ 3468]='h00001774;  wr_data_rom[ 3468]='h00000f36;
    rd_cycle[ 3469] = 1'b0;  wr_cycle[ 3469] = 1'b1;  addr_rom[ 3469]='h000008ac;  wr_data_rom[ 3469]='h000000ef;
    rd_cycle[ 3470] = 1'b1;  wr_cycle[ 3470] = 1'b0;  addr_rom[ 3470]='h00001624;  wr_data_rom[ 3470]='h00000000;
    rd_cycle[ 3471] = 1'b0;  wr_cycle[ 3471] = 1'b1;  addr_rom[ 3471]='h00000ea0;  wr_data_rom[ 3471]='h000013e0;
    rd_cycle[ 3472] = 1'b0;  wr_cycle[ 3472] = 1'b1;  addr_rom[ 3472]='h00000bf4;  wr_data_rom[ 3472]='h00001e10;
    rd_cycle[ 3473] = 1'b1;  wr_cycle[ 3473] = 1'b0;  addr_rom[ 3473]='h0000158c;  wr_data_rom[ 3473]='h00000000;
    rd_cycle[ 3474] = 1'b0;  wr_cycle[ 3474] = 1'b1;  addr_rom[ 3474]='h0000031c;  wr_data_rom[ 3474]='h00000cd0;
    rd_cycle[ 3475] = 1'b1;  wr_cycle[ 3475] = 1'b0;  addr_rom[ 3475]='h00001160;  wr_data_rom[ 3475]='h00000000;
    rd_cycle[ 3476] = 1'b1;  wr_cycle[ 3476] = 1'b0;  addr_rom[ 3476]='h00001630;  wr_data_rom[ 3476]='h00000000;
    rd_cycle[ 3477] = 1'b0;  wr_cycle[ 3477] = 1'b1;  addr_rom[ 3477]='h00000740;  wr_data_rom[ 3477]='h000001a2;
    rd_cycle[ 3478] = 1'b1;  wr_cycle[ 3478] = 1'b0;  addr_rom[ 3478]='h00000850;  wr_data_rom[ 3478]='h00000000;
    rd_cycle[ 3479] = 1'b0;  wr_cycle[ 3479] = 1'b1;  addr_rom[ 3479]='h00001f24;  wr_data_rom[ 3479]='h00001c74;
    rd_cycle[ 3480] = 1'b0;  wr_cycle[ 3480] = 1'b1;  addr_rom[ 3480]='h00001368;  wr_data_rom[ 3480]='h000011e2;
    rd_cycle[ 3481] = 1'b1;  wr_cycle[ 3481] = 1'b0;  addr_rom[ 3481]='h000016bc;  wr_data_rom[ 3481]='h00000000;
    rd_cycle[ 3482] = 1'b1;  wr_cycle[ 3482] = 1'b0;  addr_rom[ 3482]='h0000100c;  wr_data_rom[ 3482]='h00000000;
    rd_cycle[ 3483] = 1'b0;  wr_cycle[ 3483] = 1'b1;  addr_rom[ 3483]='h000008b0;  wr_data_rom[ 3483]='h00000189;
    rd_cycle[ 3484] = 1'b0;  wr_cycle[ 3484] = 1'b1;  addr_rom[ 3484]='h00001374;  wr_data_rom[ 3484]='h000014e3;
    rd_cycle[ 3485] = 1'b1;  wr_cycle[ 3485] = 1'b0;  addr_rom[ 3485]='h00000108;  wr_data_rom[ 3485]='h00000000;
    rd_cycle[ 3486] = 1'b1;  wr_cycle[ 3486] = 1'b0;  addr_rom[ 3486]='h00000664;  wr_data_rom[ 3486]='h00000000;
    rd_cycle[ 3487] = 1'b1;  wr_cycle[ 3487] = 1'b0;  addr_rom[ 3487]='h00001b6c;  wr_data_rom[ 3487]='h00000000;
    rd_cycle[ 3488] = 1'b1;  wr_cycle[ 3488] = 1'b0;  addr_rom[ 3488]='h00000604;  wr_data_rom[ 3488]='h00000000;
    rd_cycle[ 3489] = 1'b1;  wr_cycle[ 3489] = 1'b0;  addr_rom[ 3489]='h00000f94;  wr_data_rom[ 3489]='h00000000;
    rd_cycle[ 3490] = 1'b1;  wr_cycle[ 3490] = 1'b0;  addr_rom[ 3490]='h0000104c;  wr_data_rom[ 3490]='h00000000;
    rd_cycle[ 3491] = 1'b0;  wr_cycle[ 3491] = 1'b1;  addr_rom[ 3491]='h00000eb0;  wr_data_rom[ 3491]='h000000d3;
    rd_cycle[ 3492] = 1'b0;  wr_cycle[ 3492] = 1'b1;  addr_rom[ 3492]='h00000f94;  wr_data_rom[ 3492]='h00000da8;
    rd_cycle[ 3493] = 1'b0;  wr_cycle[ 3493] = 1'b1;  addr_rom[ 3493]='h00000f34;  wr_data_rom[ 3493]='h000010a5;
    rd_cycle[ 3494] = 1'b1;  wr_cycle[ 3494] = 1'b0;  addr_rom[ 3494]='h000009f0;  wr_data_rom[ 3494]='h00000000;
    rd_cycle[ 3495] = 1'b1;  wr_cycle[ 3495] = 1'b0;  addr_rom[ 3495]='h000006dc;  wr_data_rom[ 3495]='h00000000;
    rd_cycle[ 3496] = 1'b1;  wr_cycle[ 3496] = 1'b0;  addr_rom[ 3496]='h00001888;  wr_data_rom[ 3496]='h00000000;
    rd_cycle[ 3497] = 1'b0;  wr_cycle[ 3497] = 1'b1;  addr_rom[ 3497]='h00001c74;  wr_data_rom[ 3497]='h00000429;
    rd_cycle[ 3498] = 1'b1;  wr_cycle[ 3498] = 1'b0;  addr_rom[ 3498]='h00000948;  wr_data_rom[ 3498]='h00000000;
    rd_cycle[ 3499] = 1'b0;  wr_cycle[ 3499] = 1'b1;  addr_rom[ 3499]='h000013dc;  wr_data_rom[ 3499]='h00000e2e;
    rd_cycle[ 3500] = 1'b0;  wr_cycle[ 3500] = 1'b1;  addr_rom[ 3500]='h00001048;  wr_data_rom[ 3500]='h0000140c;
    rd_cycle[ 3501] = 1'b0;  wr_cycle[ 3501] = 1'b1;  addr_rom[ 3501]='h000015c0;  wr_data_rom[ 3501]='h000006bd;
    rd_cycle[ 3502] = 1'b0;  wr_cycle[ 3502] = 1'b1;  addr_rom[ 3502]='h00001310;  wr_data_rom[ 3502]='h0000016b;
    rd_cycle[ 3503] = 1'b0;  wr_cycle[ 3503] = 1'b1;  addr_rom[ 3503]='h00001e68;  wr_data_rom[ 3503]='h000008cd;
    rd_cycle[ 3504] = 1'b1;  wr_cycle[ 3504] = 1'b0;  addr_rom[ 3504]='h0000033c;  wr_data_rom[ 3504]='h00000000;
    rd_cycle[ 3505] = 1'b1;  wr_cycle[ 3505] = 1'b0;  addr_rom[ 3505]='h000008b8;  wr_data_rom[ 3505]='h00000000;
    rd_cycle[ 3506] = 1'b1;  wr_cycle[ 3506] = 1'b0;  addr_rom[ 3506]='h00000978;  wr_data_rom[ 3506]='h00000000;
    rd_cycle[ 3507] = 1'b0;  wr_cycle[ 3507] = 1'b1;  addr_rom[ 3507]='h00001954;  wr_data_rom[ 3507]='h00001283;
    rd_cycle[ 3508] = 1'b0;  wr_cycle[ 3508] = 1'b1;  addr_rom[ 3508]='h00001b0c;  wr_data_rom[ 3508]='h0000168c;
    rd_cycle[ 3509] = 1'b1;  wr_cycle[ 3509] = 1'b0;  addr_rom[ 3509]='h000011d8;  wr_data_rom[ 3509]='h00000000;
    rd_cycle[ 3510] = 1'b1;  wr_cycle[ 3510] = 1'b0;  addr_rom[ 3510]='h00000690;  wr_data_rom[ 3510]='h00000000;
    rd_cycle[ 3511] = 1'b0;  wr_cycle[ 3511] = 1'b1;  addr_rom[ 3511]='h00000fac;  wr_data_rom[ 3511]='h00000298;
    rd_cycle[ 3512] = 1'b0;  wr_cycle[ 3512] = 1'b1;  addr_rom[ 3512]='h00001230;  wr_data_rom[ 3512]='h00000042;
    rd_cycle[ 3513] = 1'b1;  wr_cycle[ 3513] = 1'b0;  addr_rom[ 3513]='h00000e90;  wr_data_rom[ 3513]='h00000000;
    rd_cycle[ 3514] = 1'b1;  wr_cycle[ 3514] = 1'b0;  addr_rom[ 3514]='h00000e8c;  wr_data_rom[ 3514]='h00000000;
    rd_cycle[ 3515] = 1'b1;  wr_cycle[ 3515] = 1'b0;  addr_rom[ 3515]='h00000518;  wr_data_rom[ 3515]='h00000000;
    rd_cycle[ 3516] = 1'b0;  wr_cycle[ 3516] = 1'b1;  addr_rom[ 3516]='h0000068c;  wr_data_rom[ 3516]='h0000101f;
    rd_cycle[ 3517] = 1'b0;  wr_cycle[ 3517] = 1'b1;  addr_rom[ 3517]='h00000b2c;  wr_data_rom[ 3517]='h0000174e;
    rd_cycle[ 3518] = 1'b1;  wr_cycle[ 3518] = 1'b0;  addr_rom[ 3518]='h0000135c;  wr_data_rom[ 3518]='h00000000;
    rd_cycle[ 3519] = 1'b0;  wr_cycle[ 3519] = 1'b1;  addr_rom[ 3519]='h0000050c;  wr_data_rom[ 3519]='h00000c4a;
    rd_cycle[ 3520] = 1'b0;  wr_cycle[ 3520] = 1'b1;  addr_rom[ 3520]='h00000f40;  wr_data_rom[ 3520]='h000009b4;
    rd_cycle[ 3521] = 1'b0;  wr_cycle[ 3521] = 1'b1;  addr_rom[ 3521]='h000019c4;  wr_data_rom[ 3521]='h00001840;
    rd_cycle[ 3522] = 1'b0;  wr_cycle[ 3522] = 1'b1;  addr_rom[ 3522]='h00001910;  wr_data_rom[ 3522]='h00001d54;
    rd_cycle[ 3523] = 1'b1;  wr_cycle[ 3523] = 1'b0;  addr_rom[ 3523]='h00000024;  wr_data_rom[ 3523]='h00000000;
    rd_cycle[ 3524] = 1'b1;  wr_cycle[ 3524] = 1'b0;  addr_rom[ 3524]='h00000e50;  wr_data_rom[ 3524]='h00000000;
    rd_cycle[ 3525] = 1'b0;  wr_cycle[ 3525] = 1'b1;  addr_rom[ 3525]='h00000e20;  wr_data_rom[ 3525]='h00000ed5;
    rd_cycle[ 3526] = 1'b1;  wr_cycle[ 3526] = 1'b0;  addr_rom[ 3526]='h00000d78;  wr_data_rom[ 3526]='h00000000;
    rd_cycle[ 3527] = 1'b0;  wr_cycle[ 3527] = 1'b1;  addr_rom[ 3527]='h000009b8;  wr_data_rom[ 3527]='h00001866;
    rd_cycle[ 3528] = 1'b0;  wr_cycle[ 3528] = 1'b1;  addr_rom[ 3528]='h00001b8c;  wr_data_rom[ 3528]='h000008ad;
    rd_cycle[ 3529] = 1'b0;  wr_cycle[ 3529] = 1'b1;  addr_rom[ 3529]='h000011c4;  wr_data_rom[ 3529]='h00001383;
    rd_cycle[ 3530] = 1'b1;  wr_cycle[ 3530] = 1'b0;  addr_rom[ 3530]='h00001568;  wr_data_rom[ 3530]='h00000000;
    rd_cycle[ 3531] = 1'b0;  wr_cycle[ 3531] = 1'b1;  addr_rom[ 3531]='h00000e38;  wr_data_rom[ 3531]='h000004c1;
    rd_cycle[ 3532] = 1'b1;  wr_cycle[ 3532] = 1'b0;  addr_rom[ 3532]='h00001498;  wr_data_rom[ 3532]='h00000000;
    rd_cycle[ 3533] = 1'b0;  wr_cycle[ 3533] = 1'b1;  addr_rom[ 3533]='h000016e8;  wr_data_rom[ 3533]='h000007b7;
    rd_cycle[ 3534] = 1'b0;  wr_cycle[ 3534] = 1'b1;  addr_rom[ 3534]='h0000120c;  wr_data_rom[ 3534]='h00000791;
    rd_cycle[ 3535] = 1'b0;  wr_cycle[ 3535] = 1'b1;  addr_rom[ 3535]='h00001870;  wr_data_rom[ 3535]='h00000ece;
    rd_cycle[ 3536] = 1'b0;  wr_cycle[ 3536] = 1'b1;  addr_rom[ 3536]='h00001c34;  wr_data_rom[ 3536]='h00000053;
    rd_cycle[ 3537] = 1'b1;  wr_cycle[ 3537] = 1'b0;  addr_rom[ 3537]='h00000e0c;  wr_data_rom[ 3537]='h00000000;
    rd_cycle[ 3538] = 1'b0;  wr_cycle[ 3538] = 1'b1;  addr_rom[ 3538]='h00001d18;  wr_data_rom[ 3538]='h00000052;
    rd_cycle[ 3539] = 1'b1;  wr_cycle[ 3539] = 1'b0;  addr_rom[ 3539]='h00000d8c;  wr_data_rom[ 3539]='h00000000;
    rd_cycle[ 3540] = 1'b0;  wr_cycle[ 3540] = 1'b1;  addr_rom[ 3540]='h00001320;  wr_data_rom[ 3540]='h00000fc1;
    rd_cycle[ 3541] = 1'b1;  wr_cycle[ 3541] = 1'b0;  addr_rom[ 3541]='h00000dd0;  wr_data_rom[ 3541]='h00000000;
    rd_cycle[ 3542] = 1'b1;  wr_cycle[ 3542] = 1'b0;  addr_rom[ 3542]='h000009e4;  wr_data_rom[ 3542]='h00000000;
    rd_cycle[ 3543] = 1'b0;  wr_cycle[ 3543] = 1'b1;  addr_rom[ 3543]='h00000528;  wr_data_rom[ 3543]='h00001a33;
    rd_cycle[ 3544] = 1'b0;  wr_cycle[ 3544] = 1'b1;  addr_rom[ 3544]='h00000ff8;  wr_data_rom[ 3544]='h00000209;
    rd_cycle[ 3545] = 1'b0;  wr_cycle[ 3545] = 1'b1;  addr_rom[ 3545]='h00001470;  wr_data_rom[ 3545]='h00001a01;
    rd_cycle[ 3546] = 1'b0;  wr_cycle[ 3546] = 1'b1;  addr_rom[ 3546]='h000000c0;  wr_data_rom[ 3546]='h00000eb7;
    rd_cycle[ 3547] = 1'b1;  wr_cycle[ 3547] = 1'b0;  addr_rom[ 3547]='h00000e78;  wr_data_rom[ 3547]='h00000000;
    rd_cycle[ 3548] = 1'b0;  wr_cycle[ 3548] = 1'b1;  addr_rom[ 3548]='h00001cd4;  wr_data_rom[ 3548]='h00001064;
    rd_cycle[ 3549] = 1'b0;  wr_cycle[ 3549] = 1'b1;  addr_rom[ 3549]='h00000400;  wr_data_rom[ 3549]='h00001ccb;
    rd_cycle[ 3550] = 1'b1;  wr_cycle[ 3550] = 1'b0;  addr_rom[ 3550]='h00001944;  wr_data_rom[ 3550]='h00000000;
    rd_cycle[ 3551] = 1'b1;  wr_cycle[ 3551] = 1'b0;  addr_rom[ 3551]='h00001bc0;  wr_data_rom[ 3551]='h00000000;
    rd_cycle[ 3552] = 1'b0;  wr_cycle[ 3552] = 1'b1;  addr_rom[ 3552]='h0000008c;  wr_data_rom[ 3552]='h00001c6e;
    rd_cycle[ 3553] = 1'b0;  wr_cycle[ 3553] = 1'b1;  addr_rom[ 3553]='h00000890;  wr_data_rom[ 3553]='h0000110d;
    rd_cycle[ 3554] = 1'b0;  wr_cycle[ 3554] = 1'b1;  addr_rom[ 3554]='h0000045c;  wr_data_rom[ 3554]='h00000fb6;
    rd_cycle[ 3555] = 1'b1;  wr_cycle[ 3555] = 1'b0;  addr_rom[ 3555]='h00001430;  wr_data_rom[ 3555]='h00000000;
    rd_cycle[ 3556] = 1'b0;  wr_cycle[ 3556] = 1'b1;  addr_rom[ 3556]='h00000ad0;  wr_data_rom[ 3556]='h00001c8f;
    rd_cycle[ 3557] = 1'b1;  wr_cycle[ 3557] = 1'b0;  addr_rom[ 3557]='h000008e0;  wr_data_rom[ 3557]='h00000000;
    rd_cycle[ 3558] = 1'b1;  wr_cycle[ 3558] = 1'b0;  addr_rom[ 3558]='h000004e8;  wr_data_rom[ 3558]='h00000000;
    rd_cycle[ 3559] = 1'b1;  wr_cycle[ 3559] = 1'b0;  addr_rom[ 3559]='h00000b04;  wr_data_rom[ 3559]='h00000000;
    rd_cycle[ 3560] = 1'b0;  wr_cycle[ 3560] = 1'b1;  addr_rom[ 3560]='h00000b1c;  wr_data_rom[ 3560]='h00000def;
    rd_cycle[ 3561] = 1'b0;  wr_cycle[ 3561] = 1'b1;  addr_rom[ 3561]='h00000a38;  wr_data_rom[ 3561]='h000007b3;
    rd_cycle[ 3562] = 1'b0;  wr_cycle[ 3562] = 1'b1;  addr_rom[ 3562]='h000002ec;  wr_data_rom[ 3562]='h00001350;
    rd_cycle[ 3563] = 1'b0;  wr_cycle[ 3563] = 1'b1;  addr_rom[ 3563]='h00000f60;  wr_data_rom[ 3563]='h00000370;
    rd_cycle[ 3564] = 1'b1;  wr_cycle[ 3564] = 1'b0;  addr_rom[ 3564]='h000000e8;  wr_data_rom[ 3564]='h00000000;
    rd_cycle[ 3565] = 1'b1;  wr_cycle[ 3565] = 1'b0;  addr_rom[ 3565]='h00001724;  wr_data_rom[ 3565]='h00000000;
    rd_cycle[ 3566] = 1'b1;  wr_cycle[ 3566] = 1'b0;  addr_rom[ 3566]='h00001e6c;  wr_data_rom[ 3566]='h00000000;
    rd_cycle[ 3567] = 1'b0;  wr_cycle[ 3567] = 1'b1;  addr_rom[ 3567]='h00001dc8;  wr_data_rom[ 3567]='h00001a72;
    rd_cycle[ 3568] = 1'b1;  wr_cycle[ 3568] = 1'b0;  addr_rom[ 3568]='h00000b6c;  wr_data_rom[ 3568]='h00000000;
    rd_cycle[ 3569] = 1'b1;  wr_cycle[ 3569] = 1'b0;  addr_rom[ 3569]='h00001190;  wr_data_rom[ 3569]='h00000000;
    rd_cycle[ 3570] = 1'b1;  wr_cycle[ 3570] = 1'b0;  addr_rom[ 3570]='h0000081c;  wr_data_rom[ 3570]='h00000000;
    rd_cycle[ 3571] = 1'b1;  wr_cycle[ 3571] = 1'b0;  addr_rom[ 3571]='h000018d4;  wr_data_rom[ 3571]='h00000000;
    rd_cycle[ 3572] = 1'b1;  wr_cycle[ 3572] = 1'b0;  addr_rom[ 3572]='h00000d10;  wr_data_rom[ 3572]='h00000000;
    rd_cycle[ 3573] = 1'b1;  wr_cycle[ 3573] = 1'b0;  addr_rom[ 3573]='h000009f0;  wr_data_rom[ 3573]='h00000000;
    rd_cycle[ 3574] = 1'b0;  wr_cycle[ 3574] = 1'b1;  addr_rom[ 3574]='h00001304;  wr_data_rom[ 3574]='h0000157a;
    rd_cycle[ 3575] = 1'b1;  wr_cycle[ 3575] = 1'b0;  addr_rom[ 3575]='h0000144c;  wr_data_rom[ 3575]='h00000000;
    rd_cycle[ 3576] = 1'b0;  wr_cycle[ 3576] = 1'b1;  addr_rom[ 3576]='h00000c68;  wr_data_rom[ 3576]='h00000038;
    rd_cycle[ 3577] = 1'b1;  wr_cycle[ 3577] = 1'b0;  addr_rom[ 3577]='h000011a8;  wr_data_rom[ 3577]='h00000000;
    rd_cycle[ 3578] = 1'b1;  wr_cycle[ 3578] = 1'b0;  addr_rom[ 3578]='h00000310;  wr_data_rom[ 3578]='h00000000;
    rd_cycle[ 3579] = 1'b1;  wr_cycle[ 3579] = 1'b0;  addr_rom[ 3579]='h00001a5c;  wr_data_rom[ 3579]='h00000000;
    rd_cycle[ 3580] = 1'b0;  wr_cycle[ 3580] = 1'b1;  addr_rom[ 3580]='h0000187c;  wr_data_rom[ 3580]='h00001d33;
    rd_cycle[ 3581] = 1'b1;  wr_cycle[ 3581] = 1'b0;  addr_rom[ 3581]='h000012d8;  wr_data_rom[ 3581]='h00000000;
    rd_cycle[ 3582] = 1'b1;  wr_cycle[ 3582] = 1'b0;  addr_rom[ 3582]='h00001b4c;  wr_data_rom[ 3582]='h00000000;
    rd_cycle[ 3583] = 1'b1;  wr_cycle[ 3583] = 1'b0;  addr_rom[ 3583]='h00001b70;  wr_data_rom[ 3583]='h00000000;
    rd_cycle[ 3584] = 1'b1;  wr_cycle[ 3584] = 1'b0;  addr_rom[ 3584]='h0000191c;  wr_data_rom[ 3584]='h00000000;
    rd_cycle[ 3585] = 1'b0;  wr_cycle[ 3585] = 1'b1;  addr_rom[ 3585]='h000011d4;  wr_data_rom[ 3585]='h0000184a;
    rd_cycle[ 3586] = 1'b0;  wr_cycle[ 3586] = 1'b1;  addr_rom[ 3586]='h000017e8;  wr_data_rom[ 3586]='h00000aa9;
    rd_cycle[ 3587] = 1'b1;  wr_cycle[ 3587] = 1'b0;  addr_rom[ 3587]='h00000360;  wr_data_rom[ 3587]='h00000000;
    rd_cycle[ 3588] = 1'b1;  wr_cycle[ 3588] = 1'b0;  addr_rom[ 3588]='h00001eb0;  wr_data_rom[ 3588]='h00000000;
    rd_cycle[ 3589] = 1'b0;  wr_cycle[ 3589] = 1'b1;  addr_rom[ 3589]='h00000ce8;  wr_data_rom[ 3589]='h0000170d;
    rd_cycle[ 3590] = 1'b0;  wr_cycle[ 3590] = 1'b1;  addr_rom[ 3590]='h00001454;  wr_data_rom[ 3590]='h00001588;
    rd_cycle[ 3591] = 1'b0;  wr_cycle[ 3591] = 1'b1;  addr_rom[ 3591]='h00001138;  wr_data_rom[ 3591]='h00000b15;
    rd_cycle[ 3592] = 1'b1;  wr_cycle[ 3592] = 1'b0;  addr_rom[ 3592]='h00000cf0;  wr_data_rom[ 3592]='h00000000;
    rd_cycle[ 3593] = 1'b0;  wr_cycle[ 3593] = 1'b1;  addr_rom[ 3593]='h00001a30;  wr_data_rom[ 3593]='h00000fe7;
    rd_cycle[ 3594] = 1'b1;  wr_cycle[ 3594] = 1'b0;  addr_rom[ 3594]='h00000978;  wr_data_rom[ 3594]='h00000000;
    rd_cycle[ 3595] = 1'b0;  wr_cycle[ 3595] = 1'b1;  addr_rom[ 3595]='h00000dc4;  wr_data_rom[ 3595]='h000017f6;
    rd_cycle[ 3596] = 1'b0;  wr_cycle[ 3596] = 1'b1;  addr_rom[ 3596]='h0000101c;  wr_data_rom[ 3596]='h00000b1c;
    rd_cycle[ 3597] = 1'b0;  wr_cycle[ 3597] = 1'b1;  addr_rom[ 3597]='h00000de0;  wr_data_rom[ 3597]='h000012b5;
    rd_cycle[ 3598] = 1'b1;  wr_cycle[ 3598] = 1'b0;  addr_rom[ 3598]='h000004dc;  wr_data_rom[ 3598]='h00000000;
    rd_cycle[ 3599] = 1'b1;  wr_cycle[ 3599] = 1'b0;  addr_rom[ 3599]='h000008ac;  wr_data_rom[ 3599]='h00000000;
    rd_cycle[ 3600] = 1'b0;  wr_cycle[ 3600] = 1'b1;  addr_rom[ 3600]='h00000f40;  wr_data_rom[ 3600]='h00001d03;
    rd_cycle[ 3601] = 1'b1;  wr_cycle[ 3601] = 1'b0;  addr_rom[ 3601]='h00000994;  wr_data_rom[ 3601]='h00000000;
    rd_cycle[ 3602] = 1'b0;  wr_cycle[ 3602] = 1'b1;  addr_rom[ 3602]='h0000191c;  wr_data_rom[ 3602]='h00000ed0;
    rd_cycle[ 3603] = 1'b0;  wr_cycle[ 3603] = 1'b1;  addr_rom[ 3603]='h0000088c;  wr_data_rom[ 3603]='h00001d9a;
    rd_cycle[ 3604] = 1'b0;  wr_cycle[ 3604] = 1'b1;  addr_rom[ 3604]='h00000ff4;  wr_data_rom[ 3604]='h00000f4f;
    rd_cycle[ 3605] = 1'b0;  wr_cycle[ 3605] = 1'b1;  addr_rom[ 3605]='h000010a0;  wr_data_rom[ 3605]='h000001fa;
    rd_cycle[ 3606] = 1'b1;  wr_cycle[ 3606] = 1'b0;  addr_rom[ 3606]='h00001520;  wr_data_rom[ 3606]='h00000000;
    rd_cycle[ 3607] = 1'b1;  wr_cycle[ 3607] = 1'b0;  addr_rom[ 3607]='h00000698;  wr_data_rom[ 3607]='h00000000;
    rd_cycle[ 3608] = 1'b0;  wr_cycle[ 3608] = 1'b1;  addr_rom[ 3608]='h00001934;  wr_data_rom[ 3608]='h00001ece;
    rd_cycle[ 3609] = 1'b0;  wr_cycle[ 3609] = 1'b1;  addr_rom[ 3609]='h00001ef4;  wr_data_rom[ 3609]='h00001c34;
    rd_cycle[ 3610] = 1'b1;  wr_cycle[ 3610] = 1'b0;  addr_rom[ 3610]='h00000acc;  wr_data_rom[ 3610]='h00000000;
    rd_cycle[ 3611] = 1'b0;  wr_cycle[ 3611] = 1'b1;  addr_rom[ 3611]='h00000ee4;  wr_data_rom[ 3611]='h000009b6;
    rd_cycle[ 3612] = 1'b0;  wr_cycle[ 3612] = 1'b1;  addr_rom[ 3612]='h00001bb4;  wr_data_rom[ 3612]='h000011ca;
    rd_cycle[ 3613] = 1'b0;  wr_cycle[ 3613] = 1'b1;  addr_rom[ 3613]='h000008f8;  wr_data_rom[ 3613]='h000011d8;
    rd_cycle[ 3614] = 1'b1;  wr_cycle[ 3614] = 1'b0;  addr_rom[ 3614]='h0000153c;  wr_data_rom[ 3614]='h00000000;
    rd_cycle[ 3615] = 1'b1;  wr_cycle[ 3615] = 1'b0;  addr_rom[ 3615]='h0000024c;  wr_data_rom[ 3615]='h00000000;
    rd_cycle[ 3616] = 1'b1;  wr_cycle[ 3616] = 1'b0;  addr_rom[ 3616]='h00000330;  wr_data_rom[ 3616]='h00000000;
    rd_cycle[ 3617] = 1'b1;  wr_cycle[ 3617] = 1'b0;  addr_rom[ 3617]='h000004dc;  wr_data_rom[ 3617]='h00000000;
    rd_cycle[ 3618] = 1'b1;  wr_cycle[ 3618] = 1'b0;  addr_rom[ 3618]='h00000628;  wr_data_rom[ 3618]='h00000000;
    rd_cycle[ 3619] = 1'b1;  wr_cycle[ 3619] = 1'b0;  addr_rom[ 3619]='h000000ec;  wr_data_rom[ 3619]='h00000000;
    rd_cycle[ 3620] = 1'b0;  wr_cycle[ 3620] = 1'b1;  addr_rom[ 3620]='h00001a0c;  wr_data_rom[ 3620]='h0000130a;
    rd_cycle[ 3621] = 1'b1;  wr_cycle[ 3621] = 1'b0;  addr_rom[ 3621]='h00000014;  wr_data_rom[ 3621]='h00000000;
    rd_cycle[ 3622] = 1'b1;  wr_cycle[ 3622] = 1'b0;  addr_rom[ 3622]='h0000130c;  wr_data_rom[ 3622]='h00000000;
    rd_cycle[ 3623] = 1'b1;  wr_cycle[ 3623] = 1'b0;  addr_rom[ 3623]='h00000be8;  wr_data_rom[ 3623]='h00000000;
    rd_cycle[ 3624] = 1'b1;  wr_cycle[ 3624] = 1'b0;  addr_rom[ 3624]='h00000bc4;  wr_data_rom[ 3624]='h00000000;
    rd_cycle[ 3625] = 1'b1;  wr_cycle[ 3625] = 1'b0;  addr_rom[ 3625]='h000003dc;  wr_data_rom[ 3625]='h00000000;
    rd_cycle[ 3626] = 1'b1;  wr_cycle[ 3626] = 1'b0;  addr_rom[ 3626]='h00000f6c;  wr_data_rom[ 3626]='h00000000;
    rd_cycle[ 3627] = 1'b1;  wr_cycle[ 3627] = 1'b0;  addr_rom[ 3627]='h00001b14;  wr_data_rom[ 3627]='h00000000;
    rd_cycle[ 3628] = 1'b1;  wr_cycle[ 3628] = 1'b0;  addr_rom[ 3628]='h00000e78;  wr_data_rom[ 3628]='h00000000;
    rd_cycle[ 3629] = 1'b0;  wr_cycle[ 3629] = 1'b1;  addr_rom[ 3629]='h0000158c;  wr_data_rom[ 3629]='h000012aa;
    rd_cycle[ 3630] = 1'b0;  wr_cycle[ 3630] = 1'b1;  addr_rom[ 3630]='h0000188c;  wr_data_rom[ 3630]='h0000092c;
    rd_cycle[ 3631] = 1'b0;  wr_cycle[ 3631] = 1'b1;  addr_rom[ 3631]='h00000be0;  wr_data_rom[ 3631]='h000007a5;
    rd_cycle[ 3632] = 1'b0;  wr_cycle[ 3632] = 1'b1;  addr_rom[ 3632]='h00001230;  wr_data_rom[ 3632]='h00000589;
    rd_cycle[ 3633] = 1'b1;  wr_cycle[ 3633] = 1'b0;  addr_rom[ 3633]='h00001258;  wr_data_rom[ 3633]='h00000000;
    rd_cycle[ 3634] = 1'b0;  wr_cycle[ 3634] = 1'b1;  addr_rom[ 3634]='h00001598;  wr_data_rom[ 3634]='h000018e5;
    rd_cycle[ 3635] = 1'b0;  wr_cycle[ 3635] = 1'b1;  addr_rom[ 3635]='h0000102c;  wr_data_rom[ 3635]='h00001267;
    rd_cycle[ 3636] = 1'b0;  wr_cycle[ 3636] = 1'b1;  addr_rom[ 3636]='h00001e0c;  wr_data_rom[ 3636]='h0000062e;
    rd_cycle[ 3637] = 1'b1;  wr_cycle[ 3637] = 1'b0;  addr_rom[ 3637]='h0000133c;  wr_data_rom[ 3637]='h00000000;
    rd_cycle[ 3638] = 1'b1;  wr_cycle[ 3638] = 1'b0;  addr_rom[ 3638]='h0000034c;  wr_data_rom[ 3638]='h00000000;
    rd_cycle[ 3639] = 1'b0;  wr_cycle[ 3639] = 1'b1;  addr_rom[ 3639]='h00000818;  wr_data_rom[ 3639]='h000019be;
    rd_cycle[ 3640] = 1'b1;  wr_cycle[ 3640] = 1'b0;  addr_rom[ 3640]='h0000029c;  wr_data_rom[ 3640]='h00000000;
    rd_cycle[ 3641] = 1'b1;  wr_cycle[ 3641] = 1'b0;  addr_rom[ 3641]='h000008e0;  wr_data_rom[ 3641]='h00000000;
    rd_cycle[ 3642] = 1'b1;  wr_cycle[ 3642] = 1'b0;  addr_rom[ 3642]='h000012f8;  wr_data_rom[ 3642]='h00000000;
    rd_cycle[ 3643] = 1'b0;  wr_cycle[ 3643] = 1'b1;  addr_rom[ 3643]='h00000664;  wr_data_rom[ 3643]='h000018be;
    rd_cycle[ 3644] = 1'b1;  wr_cycle[ 3644] = 1'b0;  addr_rom[ 3644]='h000001b8;  wr_data_rom[ 3644]='h00000000;
    rd_cycle[ 3645] = 1'b1;  wr_cycle[ 3645] = 1'b0;  addr_rom[ 3645]='h00001460;  wr_data_rom[ 3645]='h00000000;
    rd_cycle[ 3646] = 1'b1;  wr_cycle[ 3646] = 1'b0;  addr_rom[ 3646]='h000019f4;  wr_data_rom[ 3646]='h00000000;
    rd_cycle[ 3647] = 1'b0;  wr_cycle[ 3647] = 1'b1;  addr_rom[ 3647]='h00000c14;  wr_data_rom[ 3647]='h00000332;
    rd_cycle[ 3648] = 1'b1;  wr_cycle[ 3648] = 1'b0;  addr_rom[ 3648]='h00000050;  wr_data_rom[ 3648]='h00000000;
    rd_cycle[ 3649] = 1'b0;  wr_cycle[ 3649] = 1'b1;  addr_rom[ 3649]='h00001194;  wr_data_rom[ 3649]='h000019f8;
    rd_cycle[ 3650] = 1'b0;  wr_cycle[ 3650] = 1'b1;  addr_rom[ 3650]='h000000ec;  wr_data_rom[ 3650]='h00000f2a;
    rd_cycle[ 3651] = 1'b0;  wr_cycle[ 3651] = 1'b1;  addr_rom[ 3651]='h00000ce8;  wr_data_rom[ 3651]='h00000220;
    rd_cycle[ 3652] = 1'b0;  wr_cycle[ 3652] = 1'b1;  addr_rom[ 3652]='h00001410;  wr_data_rom[ 3652]='h00001de4;
    rd_cycle[ 3653] = 1'b1;  wr_cycle[ 3653] = 1'b0;  addr_rom[ 3653]='h0000060c;  wr_data_rom[ 3653]='h00000000;
    rd_cycle[ 3654] = 1'b1;  wr_cycle[ 3654] = 1'b0;  addr_rom[ 3654]='h0000107c;  wr_data_rom[ 3654]='h00000000;
    rd_cycle[ 3655] = 1'b0;  wr_cycle[ 3655] = 1'b1;  addr_rom[ 3655]='h00001650;  wr_data_rom[ 3655]='h00000638;
    rd_cycle[ 3656] = 1'b0;  wr_cycle[ 3656] = 1'b1;  addr_rom[ 3656]='h000017e4;  wr_data_rom[ 3656]='h00000a69;
    rd_cycle[ 3657] = 1'b1;  wr_cycle[ 3657] = 1'b0;  addr_rom[ 3657]='h00001eac;  wr_data_rom[ 3657]='h00000000;
    rd_cycle[ 3658] = 1'b0;  wr_cycle[ 3658] = 1'b1;  addr_rom[ 3658]='h0000098c;  wr_data_rom[ 3658]='h00001d17;
    rd_cycle[ 3659] = 1'b0;  wr_cycle[ 3659] = 1'b1;  addr_rom[ 3659]='h00001ed0;  wr_data_rom[ 3659]='h00000851;
    rd_cycle[ 3660] = 1'b1;  wr_cycle[ 3660] = 1'b0;  addr_rom[ 3660]='h000009c8;  wr_data_rom[ 3660]='h00000000;
    rd_cycle[ 3661] = 1'b0;  wr_cycle[ 3661] = 1'b1;  addr_rom[ 3661]='h00001bf8;  wr_data_rom[ 3661]='h00000dc7;
    rd_cycle[ 3662] = 1'b0;  wr_cycle[ 3662] = 1'b1;  addr_rom[ 3662]='h00000bfc;  wr_data_rom[ 3662]='h00000940;
    rd_cycle[ 3663] = 1'b1;  wr_cycle[ 3663] = 1'b0;  addr_rom[ 3663]='h00000858;  wr_data_rom[ 3663]='h00000000;
    rd_cycle[ 3664] = 1'b1;  wr_cycle[ 3664] = 1'b0;  addr_rom[ 3664]='h00001080;  wr_data_rom[ 3664]='h00000000;
    rd_cycle[ 3665] = 1'b1;  wr_cycle[ 3665] = 1'b0;  addr_rom[ 3665]='h000015fc;  wr_data_rom[ 3665]='h00000000;
    rd_cycle[ 3666] = 1'b0;  wr_cycle[ 3666] = 1'b1;  addr_rom[ 3666]='h000018d0;  wr_data_rom[ 3666]='h00001db8;
    rd_cycle[ 3667] = 1'b1;  wr_cycle[ 3667] = 1'b0;  addr_rom[ 3667]='h00001428;  wr_data_rom[ 3667]='h00000000;
    rd_cycle[ 3668] = 1'b0;  wr_cycle[ 3668] = 1'b1;  addr_rom[ 3668]='h00001418;  wr_data_rom[ 3668]='h00001ea9;
    rd_cycle[ 3669] = 1'b1;  wr_cycle[ 3669] = 1'b0;  addr_rom[ 3669]='h00001b38;  wr_data_rom[ 3669]='h00000000;
    rd_cycle[ 3670] = 1'b1;  wr_cycle[ 3670] = 1'b0;  addr_rom[ 3670]='h00001970;  wr_data_rom[ 3670]='h00000000;
    rd_cycle[ 3671] = 1'b0;  wr_cycle[ 3671] = 1'b1;  addr_rom[ 3671]='h00000288;  wr_data_rom[ 3671]='h00000175;
    rd_cycle[ 3672] = 1'b1;  wr_cycle[ 3672] = 1'b0;  addr_rom[ 3672]='h00000488;  wr_data_rom[ 3672]='h00000000;
    rd_cycle[ 3673] = 1'b0;  wr_cycle[ 3673] = 1'b1;  addr_rom[ 3673]='h000017fc;  wr_data_rom[ 3673]='h00001e51;
    rd_cycle[ 3674] = 1'b1;  wr_cycle[ 3674] = 1'b0;  addr_rom[ 3674]='h00000588;  wr_data_rom[ 3674]='h00000000;
    rd_cycle[ 3675] = 1'b1;  wr_cycle[ 3675] = 1'b0;  addr_rom[ 3675]='h000006a0;  wr_data_rom[ 3675]='h00000000;
    rd_cycle[ 3676] = 1'b0;  wr_cycle[ 3676] = 1'b1;  addr_rom[ 3676]='h000014e4;  wr_data_rom[ 3676]='h00001d83;
    rd_cycle[ 3677] = 1'b1;  wr_cycle[ 3677] = 1'b0;  addr_rom[ 3677]='h00001e08;  wr_data_rom[ 3677]='h00000000;
    rd_cycle[ 3678] = 1'b0;  wr_cycle[ 3678] = 1'b1;  addr_rom[ 3678]='h00000eb8;  wr_data_rom[ 3678]='h0000108c;
    rd_cycle[ 3679] = 1'b1;  wr_cycle[ 3679] = 1'b0;  addr_rom[ 3679]='h00001920;  wr_data_rom[ 3679]='h00000000;
    rd_cycle[ 3680] = 1'b1;  wr_cycle[ 3680] = 1'b0;  addr_rom[ 3680]='h000010dc;  wr_data_rom[ 3680]='h00000000;
    rd_cycle[ 3681] = 1'b0;  wr_cycle[ 3681] = 1'b1;  addr_rom[ 3681]='h000014f8;  wr_data_rom[ 3681]='h00000b12;
    rd_cycle[ 3682] = 1'b1;  wr_cycle[ 3682] = 1'b0;  addr_rom[ 3682]='h000002c0;  wr_data_rom[ 3682]='h00000000;
    rd_cycle[ 3683] = 1'b0;  wr_cycle[ 3683] = 1'b1;  addr_rom[ 3683]='h000008e0;  wr_data_rom[ 3683]='h000004c0;
    rd_cycle[ 3684] = 1'b0;  wr_cycle[ 3684] = 1'b1;  addr_rom[ 3684]='h000001c0;  wr_data_rom[ 3684]='h00001d7a;
    rd_cycle[ 3685] = 1'b0;  wr_cycle[ 3685] = 1'b1;  addr_rom[ 3685]='h0000160c;  wr_data_rom[ 3685]='h00001153;
    rd_cycle[ 3686] = 1'b0;  wr_cycle[ 3686] = 1'b1;  addr_rom[ 3686]='h00001e1c;  wr_data_rom[ 3686]='h000004cb;
    rd_cycle[ 3687] = 1'b1;  wr_cycle[ 3687] = 1'b0;  addr_rom[ 3687]='h00001e30;  wr_data_rom[ 3687]='h00000000;
    rd_cycle[ 3688] = 1'b1;  wr_cycle[ 3688] = 1'b0;  addr_rom[ 3688]='h00000068;  wr_data_rom[ 3688]='h00000000;
    rd_cycle[ 3689] = 1'b1;  wr_cycle[ 3689] = 1'b0;  addr_rom[ 3689]='h00000cc4;  wr_data_rom[ 3689]='h00000000;
    rd_cycle[ 3690] = 1'b1;  wr_cycle[ 3690] = 1'b0;  addr_rom[ 3690]='h00001ca0;  wr_data_rom[ 3690]='h00000000;
    rd_cycle[ 3691] = 1'b0;  wr_cycle[ 3691] = 1'b1;  addr_rom[ 3691]='h00001aec;  wr_data_rom[ 3691]='h00000abb;
    rd_cycle[ 3692] = 1'b0;  wr_cycle[ 3692] = 1'b1;  addr_rom[ 3692]='h000008dc;  wr_data_rom[ 3692]='h0000083a;
    rd_cycle[ 3693] = 1'b1;  wr_cycle[ 3693] = 1'b0;  addr_rom[ 3693]='h00001d8c;  wr_data_rom[ 3693]='h00000000;
    rd_cycle[ 3694] = 1'b0;  wr_cycle[ 3694] = 1'b1;  addr_rom[ 3694]='h000019e8;  wr_data_rom[ 3694]='h000004a7;
    rd_cycle[ 3695] = 1'b0;  wr_cycle[ 3695] = 1'b1;  addr_rom[ 3695]='h000014a0;  wr_data_rom[ 3695]='h000014e7;
    rd_cycle[ 3696] = 1'b1;  wr_cycle[ 3696] = 1'b0;  addr_rom[ 3696]='h00000844;  wr_data_rom[ 3696]='h00000000;
    rd_cycle[ 3697] = 1'b0;  wr_cycle[ 3697] = 1'b1;  addr_rom[ 3697]='h000013fc;  wr_data_rom[ 3697]='h0000115b;
    rd_cycle[ 3698] = 1'b1;  wr_cycle[ 3698] = 1'b0;  addr_rom[ 3698]='h00001c64;  wr_data_rom[ 3698]='h00000000;
    rd_cycle[ 3699] = 1'b0;  wr_cycle[ 3699] = 1'b1;  addr_rom[ 3699]='h00001d60;  wr_data_rom[ 3699]='h00000620;
    rd_cycle[ 3700] = 1'b0;  wr_cycle[ 3700] = 1'b1;  addr_rom[ 3700]='h00000e28;  wr_data_rom[ 3700]='h000012b5;
    rd_cycle[ 3701] = 1'b0;  wr_cycle[ 3701] = 1'b1;  addr_rom[ 3701]='h000008d8;  wr_data_rom[ 3701]='h00000724;
    rd_cycle[ 3702] = 1'b1;  wr_cycle[ 3702] = 1'b0;  addr_rom[ 3702]='h000015b4;  wr_data_rom[ 3702]='h00000000;
    rd_cycle[ 3703] = 1'b0;  wr_cycle[ 3703] = 1'b1;  addr_rom[ 3703]='h00000acc;  wr_data_rom[ 3703]='h0000019a;
    rd_cycle[ 3704] = 1'b0;  wr_cycle[ 3704] = 1'b1;  addr_rom[ 3704]='h00000ad8;  wr_data_rom[ 3704]='h00001c84;
    rd_cycle[ 3705] = 1'b0;  wr_cycle[ 3705] = 1'b1;  addr_rom[ 3705]='h000003cc;  wr_data_rom[ 3705]='h0000051d;
    rd_cycle[ 3706] = 1'b0;  wr_cycle[ 3706] = 1'b1;  addr_rom[ 3706]='h00001174;  wr_data_rom[ 3706]='h00001cef;
    rd_cycle[ 3707] = 1'b0;  wr_cycle[ 3707] = 1'b1;  addr_rom[ 3707]='h00001c90;  wr_data_rom[ 3707]='h000010ca;
    rd_cycle[ 3708] = 1'b0;  wr_cycle[ 3708] = 1'b1;  addr_rom[ 3708]='h00001520;  wr_data_rom[ 3708]='h00001605;
    rd_cycle[ 3709] = 1'b0;  wr_cycle[ 3709] = 1'b1;  addr_rom[ 3709]='h0000019c;  wr_data_rom[ 3709]='h000009df;
    rd_cycle[ 3710] = 1'b0;  wr_cycle[ 3710] = 1'b1;  addr_rom[ 3710]='h0000160c;  wr_data_rom[ 3710]='h00000339;
    rd_cycle[ 3711] = 1'b0;  wr_cycle[ 3711] = 1'b1;  addr_rom[ 3711]='h00000a70;  wr_data_rom[ 3711]='h000015ce;
    rd_cycle[ 3712] = 1'b0;  wr_cycle[ 3712] = 1'b1;  addr_rom[ 3712]='h000003c0;  wr_data_rom[ 3712]='h00001b29;
    rd_cycle[ 3713] = 1'b0;  wr_cycle[ 3713] = 1'b1;  addr_rom[ 3713]='h00001950;  wr_data_rom[ 3713]='h000006f5;
    rd_cycle[ 3714] = 1'b1;  wr_cycle[ 3714] = 1'b0;  addr_rom[ 3714]='h000015d4;  wr_data_rom[ 3714]='h00000000;
    rd_cycle[ 3715] = 1'b0;  wr_cycle[ 3715] = 1'b1;  addr_rom[ 3715]='h00000890;  wr_data_rom[ 3715]='h000019ff;
    rd_cycle[ 3716] = 1'b0;  wr_cycle[ 3716] = 1'b1;  addr_rom[ 3716]='h00001478;  wr_data_rom[ 3716]='h000002d7;
    rd_cycle[ 3717] = 1'b1;  wr_cycle[ 3717] = 1'b0;  addr_rom[ 3717]='h00001410;  wr_data_rom[ 3717]='h00000000;
    rd_cycle[ 3718] = 1'b1;  wr_cycle[ 3718] = 1'b0;  addr_rom[ 3718]='h000006ac;  wr_data_rom[ 3718]='h00000000;
    rd_cycle[ 3719] = 1'b1;  wr_cycle[ 3719] = 1'b0;  addr_rom[ 3719]='h00001a14;  wr_data_rom[ 3719]='h00000000;
    rd_cycle[ 3720] = 1'b0;  wr_cycle[ 3720] = 1'b1;  addr_rom[ 3720]='h00000280;  wr_data_rom[ 3720]='h0000004f;
    rd_cycle[ 3721] = 1'b0;  wr_cycle[ 3721] = 1'b1;  addr_rom[ 3721]='h00000fb0;  wr_data_rom[ 3721]='h00001ee4;
    rd_cycle[ 3722] = 1'b0;  wr_cycle[ 3722] = 1'b1;  addr_rom[ 3722]='h00000a38;  wr_data_rom[ 3722]='h0000108e;
    rd_cycle[ 3723] = 1'b0;  wr_cycle[ 3723] = 1'b1;  addr_rom[ 3723]='h000002bc;  wr_data_rom[ 3723]='h000003f3;
    rd_cycle[ 3724] = 1'b0;  wr_cycle[ 3724] = 1'b1;  addr_rom[ 3724]='h00000ba0;  wr_data_rom[ 3724]='h0000068f;
    rd_cycle[ 3725] = 1'b1;  wr_cycle[ 3725] = 1'b0;  addr_rom[ 3725]='h00001dfc;  wr_data_rom[ 3725]='h00000000;
    rd_cycle[ 3726] = 1'b1;  wr_cycle[ 3726] = 1'b0;  addr_rom[ 3726]='h00001d78;  wr_data_rom[ 3726]='h00000000;
    rd_cycle[ 3727] = 1'b1;  wr_cycle[ 3727] = 1'b0;  addr_rom[ 3727]='h000007b4;  wr_data_rom[ 3727]='h00000000;
    rd_cycle[ 3728] = 1'b0;  wr_cycle[ 3728] = 1'b1;  addr_rom[ 3728]='h000008ec;  wr_data_rom[ 3728]='h0000164f;
    rd_cycle[ 3729] = 1'b1;  wr_cycle[ 3729] = 1'b0;  addr_rom[ 3729]='h00000648;  wr_data_rom[ 3729]='h00000000;
    rd_cycle[ 3730] = 1'b0;  wr_cycle[ 3730] = 1'b1;  addr_rom[ 3730]='h00000344;  wr_data_rom[ 3730]='h00001e0f;
    rd_cycle[ 3731] = 1'b0;  wr_cycle[ 3731] = 1'b1;  addr_rom[ 3731]='h00001c1c;  wr_data_rom[ 3731]='h00001e06;
    rd_cycle[ 3732] = 1'b1;  wr_cycle[ 3732] = 1'b0;  addr_rom[ 3732]='h000006a4;  wr_data_rom[ 3732]='h00000000;
    rd_cycle[ 3733] = 1'b0;  wr_cycle[ 3733] = 1'b1;  addr_rom[ 3733]='h000015c4;  wr_data_rom[ 3733]='h00000646;
    rd_cycle[ 3734] = 1'b1;  wr_cycle[ 3734] = 1'b0;  addr_rom[ 3734]='h00001b54;  wr_data_rom[ 3734]='h00000000;
    rd_cycle[ 3735] = 1'b1;  wr_cycle[ 3735] = 1'b0;  addr_rom[ 3735]='h000013dc;  wr_data_rom[ 3735]='h00000000;
    rd_cycle[ 3736] = 1'b0;  wr_cycle[ 3736] = 1'b1;  addr_rom[ 3736]='h0000095c;  wr_data_rom[ 3736]='h000014d9;
    rd_cycle[ 3737] = 1'b0;  wr_cycle[ 3737] = 1'b1;  addr_rom[ 3737]='h00000294;  wr_data_rom[ 3737]='h00000405;
    rd_cycle[ 3738] = 1'b0;  wr_cycle[ 3738] = 1'b1;  addr_rom[ 3738]='h0000038c;  wr_data_rom[ 3738]='h00000379;
    rd_cycle[ 3739] = 1'b1;  wr_cycle[ 3739] = 1'b0;  addr_rom[ 3739]='h00001dfc;  wr_data_rom[ 3739]='h00000000;
    rd_cycle[ 3740] = 1'b0;  wr_cycle[ 3740] = 1'b1;  addr_rom[ 3740]='h00000798;  wr_data_rom[ 3740]='h00001d5d;
    rd_cycle[ 3741] = 1'b0;  wr_cycle[ 3741] = 1'b1;  addr_rom[ 3741]='h00001ddc;  wr_data_rom[ 3741]='h000011ac;
    rd_cycle[ 3742] = 1'b1;  wr_cycle[ 3742] = 1'b0;  addr_rom[ 3742]='h0000029c;  wr_data_rom[ 3742]='h00000000;
    rd_cycle[ 3743] = 1'b1;  wr_cycle[ 3743] = 1'b0;  addr_rom[ 3743]='h000004e4;  wr_data_rom[ 3743]='h00000000;
    rd_cycle[ 3744] = 1'b1;  wr_cycle[ 3744] = 1'b0;  addr_rom[ 3744]='h00000d38;  wr_data_rom[ 3744]='h00000000;
    rd_cycle[ 3745] = 1'b0;  wr_cycle[ 3745] = 1'b1;  addr_rom[ 3745]='h00000ea4;  wr_data_rom[ 3745]='h00001391;
    rd_cycle[ 3746] = 1'b1;  wr_cycle[ 3746] = 1'b0;  addr_rom[ 3746]='h00000c34;  wr_data_rom[ 3746]='h00000000;
    rd_cycle[ 3747] = 1'b1;  wr_cycle[ 3747] = 1'b0;  addr_rom[ 3747]='h00000164;  wr_data_rom[ 3747]='h00000000;
    rd_cycle[ 3748] = 1'b1;  wr_cycle[ 3748] = 1'b0;  addr_rom[ 3748]='h000017b0;  wr_data_rom[ 3748]='h00000000;
    rd_cycle[ 3749] = 1'b1;  wr_cycle[ 3749] = 1'b0;  addr_rom[ 3749]='h00000d04;  wr_data_rom[ 3749]='h00000000;
    rd_cycle[ 3750] = 1'b0;  wr_cycle[ 3750] = 1'b1;  addr_rom[ 3750]='h00000174;  wr_data_rom[ 3750]='h00000600;
    rd_cycle[ 3751] = 1'b1;  wr_cycle[ 3751] = 1'b0;  addr_rom[ 3751]='h00001a3c;  wr_data_rom[ 3751]='h00000000;
    rd_cycle[ 3752] = 1'b1;  wr_cycle[ 3752] = 1'b0;  addr_rom[ 3752]='h000001a8;  wr_data_rom[ 3752]='h00000000;
    rd_cycle[ 3753] = 1'b1;  wr_cycle[ 3753] = 1'b0;  addr_rom[ 3753]='h00000308;  wr_data_rom[ 3753]='h00000000;
    rd_cycle[ 3754] = 1'b0;  wr_cycle[ 3754] = 1'b1;  addr_rom[ 3754]='h00000e14;  wr_data_rom[ 3754]='h000007f5;
    rd_cycle[ 3755] = 1'b1;  wr_cycle[ 3755] = 1'b0;  addr_rom[ 3755]='h00001738;  wr_data_rom[ 3755]='h00000000;
    rd_cycle[ 3756] = 1'b1;  wr_cycle[ 3756] = 1'b0;  addr_rom[ 3756]='h000011f8;  wr_data_rom[ 3756]='h00000000;
    rd_cycle[ 3757] = 1'b0;  wr_cycle[ 3757] = 1'b1;  addr_rom[ 3757]='h000009f0;  wr_data_rom[ 3757]='h000015b6;
    rd_cycle[ 3758] = 1'b0;  wr_cycle[ 3758] = 1'b1;  addr_rom[ 3758]='h0000143c;  wr_data_rom[ 3758]='h000019d0;
    rd_cycle[ 3759] = 1'b0;  wr_cycle[ 3759] = 1'b1;  addr_rom[ 3759]='h00001718;  wr_data_rom[ 3759]='h0000154e;
    rd_cycle[ 3760] = 1'b0;  wr_cycle[ 3760] = 1'b1;  addr_rom[ 3760]='h000011dc;  wr_data_rom[ 3760]='h00000e02;
    rd_cycle[ 3761] = 1'b1;  wr_cycle[ 3761] = 1'b0;  addr_rom[ 3761]='h0000058c;  wr_data_rom[ 3761]='h00000000;
    rd_cycle[ 3762] = 1'b1;  wr_cycle[ 3762] = 1'b0;  addr_rom[ 3762]='h00001de8;  wr_data_rom[ 3762]='h00000000;
    rd_cycle[ 3763] = 1'b0;  wr_cycle[ 3763] = 1'b1;  addr_rom[ 3763]='h00001dac;  wr_data_rom[ 3763]='h00001823;
    rd_cycle[ 3764] = 1'b0;  wr_cycle[ 3764] = 1'b1;  addr_rom[ 3764]='h000016f8;  wr_data_rom[ 3764]='h00000276;
    rd_cycle[ 3765] = 1'b0;  wr_cycle[ 3765] = 1'b1;  addr_rom[ 3765]='h00001330;  wr_data_rom[ 3765]='h00000152;
    rd_cycle[ 3766] = 1'b0;  wr_cycle[ 3766] = 1'b1;  addr_rom[ 3766]='h000010ec;  wr_data_rom[ 3766]='h00000de4;
    rd_cycle[ 3767] = 1'b0;  wr_cycle[ 3767] = 1'b1;  addr_rom[ 3767]='h00001c5c;  wr_data_rom[ 3767]='h00000ec7;
    rd_cycle[ 3768] = 1'b1;  wr_cycle[ 3768] = 1'b0;  addr_rom[ 3768]='h0000117c;  wr_data_rom[ 3768]='h00000000;
    rd_cycle[ 3769] = 1'b0;  wr_cycle[ 3769] = 1'b1;  addr_rom[ 3769]='h00001708;  wr_data_rom[ 3769]='h00000fdd;
    rd_cycle[ 3770] = 1'b0;  wr_cycle[ 3770] = 1'b1;  addr_rom[ 3770]='h00001f34;  wr_data_rom[ 3770]='h0000017d;
    rd_cycle[ 3771] = 1'b0;  wr_cycle[ 3771] = 1'b1;  addr_rom[ 3771]='h00001954;  wr_data_rom[ 3771]='h0000085f;
    rd_cycle[ 3772] = 1'b0;  wr_cycle[ 3772] = 1'b1;  addr_rom[ 3772]='h000018a4;  wr_data_rom[ 3772]='h00000e08;
    rd_cycle[ 3773] = 1'b0;  wr_cycle[ 3773] = 1'b1;  addr_rom[ 3773]='h00000c38;  wr_data_rom[ 3773]='h00000fec;
    rd_cycle[ 3774] = 1'b1;  wr_cycle[ 3774] = 1'b0;  addr_rom[ 3774]='h000014b4;  wr_data_rom[ 3774]='h00000000;
    rd_cycle[ 3775] = 1'b0;  wr_cycle[ 3775] = 1'b1;  addr_rom[ 3775]='h000015fc;  wr_data_rom[ 3775]='h00001d2e;
    rd_cycle[ 3776] = 1'b1;  wr_cycle[ 3776] = 1'b0;  addr_rom[ 3776]='h00000450;  wr_data_rom[ 3776]='h00000000;
    rd_cycle[ 3777] = 1'b1;  wr_cycle[ 3777] = 1'b0;  addr_rom[ 3777]='h0000062c;  wr_data_rom[ 3777]='h00000000;
    rd_cycle[ 3778] = 1'b1;  wr_cycle[ 3778] = 1'b0;  addr_rom[ 3778]='h000009f8;  wr_data_rom[ 3778]='h00000000;
    rd_cycle[ 3779] = 1'b0;  wr_cycle[ 3779] = 1'b1;  addr_rom[ 3779]='h00000fd8;  wr_data_rom[ 3779]='h00000c31;
    rd_cycle[ 3780] = 1'b1;  wr_cycle[ 3780] = 1'b0;  addr_rom[ 3780]='h00001434;  wr_data_rom[ 3780]='h00000000;
    rd_cycle[ 3781] = 1'b0;  wr_cycle[ 3781] = 1'b1;  addr_rom[ 3781]='h0000015c;  wr_data_rom[ 3781]='h00001447;
    rd_cycle[ 3782] = 1'b1;  wr_cycle[ 3782] = 1'b0;  addr_rom[ 3782]='h00000f24;  wr_data_rom[ 3782]='h00000000;
    rd_cycle[ 3783] = 1'b1;  wr_cycle[ 3783] = 1'b0;  addr_rom[ 3783]='h000004c0;  wr_data_rom[ 3783]='h00000000;
    rd_cycle[ 3784] = 1'b0;  wr_cycle[ 3784] = 1'b1;  addr_rom[ 3784]='h00001a3c;  wr_data_rom[ 3784]='h000004a5;
    rd_cycle[ 3785] = 1'b1;  wr_cycle[ 3785] = 1'b0;  addr_rom[ 3785]='h00000350;  wr_data_rom[ 3785]='h00000000;
    rd_cycle[ 3786] = 1'b0;  wr_cycle[ 3786] = 1'b1;  addr_rom[ 3786]='h00000988;  wr_data_rom[ 3786]='h00001d77;
    rd_cycle[ 3787] = 1'b0;  wr_cycle[ 3787] = 1'b1;  addr_rom[ 3787]='h000010f0;  wr_data_rom[ 3787]='h00001007;
    rd_cycle[ 3788] = 1'b1;  wr_cycle[ 3788] = 1'b0;  addr_rom[ 3788]='h00000ce8;  wr_data_rom[ 3788]='h00000000;
    rd_cycle[ 3789] = 1'b0;  wr_cycle[ 3789] = 1'b1;  addr_rom[ 3789]='h00001708;  wr_data_rom[ 3789]='h00001a6c;
    rd_cycle[ 3790] = 1'b1;  wr_cycle[ 3790] = 1'b0;  addr_rom[ 3790]='h00000438;  wr_data_rom[ 3790]='h00000000;
    rd_cycle[ 3791] = 1'b1;  wr_cycle[ 3791] = 1'b0;  addr_rom[ 3791]='h00000878;  wr_data_rom[ 3791]='h00000000;
    rd_cycle[ 3792] = 1'b0;  wr_cycle[ 3792] = 1'b1;  addr_rom[ 3792]='h000016b4;  wr_data_rom[ 3792]='h0000020c;
    rd_cycle[ 3793] = 1'b1;  wr_cycle[ 3793] = 1'b0;  addr_rom[ 3793]='h00000544;  wr_data_rom[ 3793]='h00000000;
    rd_cycle[ 3794] = 1'b1;  wr_cycle[ 3794] = 1'b0;  addr_rom[ 3794]='h00001a58;  wr_data_rom[ 3794]='h00000000;
    rd_cycle[ 3795] = 1'b0;  wr_cycle[ 3795] = 1'b1;  addr_rom[ 3795]='h00000e38;  wr_data_rom[ 3795]='h00000b64;
    rd_cycle[ 3796] = 1'b1;  wr_cycle[ 3796] = 1'b0;  addr_rom[ 3796]='h000005d8;  wr_data_rom[ 3796]='h00000000;
    rd_cycle[ 3797] = 1'b1;  wr_cycle[ 3797] = 1'b0;  addr_rom[ 3797]='h000017a4;  wr_data_rom[ 3797]='h00000000;
    rd_cycle[ 3798] = 1'b0;  wr_cycle[ 3798] = 1'b1;  addr_rom[ 3798]='h0000196c;  wr_data_rom[ 3798]='h000011dd;
    rd_cycle[ 3799] = 1'b0;  wr_cycle[ 3799] = 1'b1;  addr_rom[ 3799]='h0000130c;  wr_data_rom[ 3799]='h0000115f;
    rd_cycle[ 3800] = 1'b0;  wr_cycle[ 3800] = 1'b1;  addr_rom[ 3800]='h000011f0;  wr_data_rom[ 3800]='h00001cd2;
    rd_cycle[ 3801] = 1'b0;  wr_cycle[ 3801] = 1'b1;  addr_rom[ 3801]='h000019fc;  wr_data_rom[ 3801]='h00001e36;
    rd_cycle[ 3802] = 1'b0;  wr_cycle[ 3802] = 1'b1;  addr_rom[ 3802]='h00001dec;  wr_data_rom[ 3802]='h00000975;
    rd_cycle[ 3803] = 1'b0;  wr_cycle[ 3803] = 1'b1;  addr_rom[ 3803]='h0000131c;  wr_data_rom[ 3803]='h00001df2;
    rd_cycle[ 3804] = 1'b0;  wr_cycle[ 3804] = 1'b1;  addr_rom[ 3804]='h000008cc;  wr_data_rom[ 3804]='h00000b4c;
    rd_cycle[ 3805] = 1'b1;  wr_cycle[ 3805] = 1'b0;  addr_rom[ 3805]='h00001704;  wr_data_rom[ 3805]='h00000000;
    rd_cycle[ 3806] = 1'b1;  wr_cycle[ 3806] = 1'b0;  addr_rom[ 3806]='h00000254;  wr_data_rom[ 3806]='h00000000;
    rd_cycle[ 3807] = 1'b0;  wr_cycle[ 3807] = 1'b1;  addr_rom[ 3807]='h00000928;  wr_data_rom[ 3807]='h00001c48;
    rd_cycle[ 3808] = 1'b0;  wr_cycle[ 3808] = 1'b1;  addr_rom[ 3808]='h000013bc;  wr_data_rom[ 3808]='h00000b7d;
    rd_cycle[ 3809] = 1'b0;  wr_cycle[ 3809] = 1'b1;  addr_rom[ 3809]='h00001af4;  wr_data_rom[ 3809]='h00001102;
    rd_cycle[ 3810] = 1'b0;  wr_cycle[ 3810] = 1'b1;  addr_rom[ 3810]='h000007e0;  wr_data_rom[ 3810]='h0000156b;
    rd_cycle[ 3811] = 1'b1;  wr_cycle[ 3811] = 1'b0;  addr_rom[ 3811]='h000015f8;  wr_data_rom[ 3811]='h00000000;
    rd_cycle[ 3812] = 1'b1;  wr_cycle[ 3812] = 1'b0;  addr_rom[ 3812]='h00001934;  wr_data_rom[ 3812]='h00000000;
    rd_cycle[ 3813] = 1'b0;  wr_cycle[ 3813] = 1'b1;  addr_rom[ 3813]='h00001938;  wr_data_rom[ 3813]='h0000107f;
    rd_cycle[ 3814] = 1'b0;  wr_cycle[ 3814] = 1'b1;  addr_rom[ 3814]='h000018a4;  wr_data_rom[ 3814]='h000006b2;
    rd_cycle[ 3815] = 1'b0;  wr_cycle[ 3815] = 1'b1;  addr_rom[ 3815]='h00000718;  wr_data_rom[ 3815]='h000013cf;
    rd_cycle[ 3816] = 1'b1;  wr_cycle[ 3816] = 1'b0;  addr_rom[ 3816]='h0000196c;  wr_data_rom[ 3816]='h00000000;
    rd_cycle[ 3817] = 1'b1;  wr_cycle[ 3817] = 1'b0;  addr_rom[ 3817]='h00000d3c;  wr_data_rom[ 3817]='h00000000;
    rd_cycle[ 3818] = 1'b1;  wr_cycle[ 3818] = 1'b0;  addr_rom[ 3818]='h000018a0;  wr_data_rom[ 3818]='h00000000;
    rd_cycle[ 3819] = 1'b0;  wr_cycle[ 3819] = 1'b1;  addr_rom[ 3819]='h0000017c;  wr_data_rom[ 3819]='h00001881;
    rd_cycle[ 3820] = 1'b1;  wr_cycle[ 3820] = 1'b0;  addr_rom[ 3820]='h00001b74;  wr_data_rom[ 3820]='h00000000;
    rd_cycle[ 3821] = 1'b0;  wr_cycle[ 3821] = 1'b1;  addr_rom[ 3821]='h00000a74;  wr_data_rom[ 3821]='h00000b7f;
    rd_cycle[ 3822] = 1'b1;  wr_cycle[ 3822] = 1'b0;  addr_rom[ 3822]='h00000424;  wr_data_rom[ 3822]='h00000000;
    rd_cycle[ 3823] = 1'b1;  wr_cycle[ 3823] = 1'b0;  addr_rom[ 3823]='h00000844;  wr_data_rom[ 3823]='h00000000;
    rd_cycle[ 3824] = 1'b0;  wr_cycle[ 3824] = 1'b1;  addr_rom[ 3824]='h000005fc;  wr_data_rom[ 3824]='h0000178c;
    rd_cycle[ 3825] = 1'b0;  wr_cycle[ 3825] = 1'b1;  addr_rom[ 3825]='h00001da0;  wr_data_rom[ 3825]='h0000179b;
    rd_cycle[ 3826] = 1'b0;  wr_cycle[ 3826] = 1'b1;  addr_rom[ 3826]='h00001d5c;  wr_data_rom[ 3826]='h00000b53;
    rd_cycle[ 3827] = 1'b1;  wr_cycle[ 3827] = 1'b0;  addr_rom[ 3827]='h00000e9c;  wr_data_rom[ 3827]='h00000000;
    rd_cycle[ 3828] = 1'b0;  wr_cycle[ 3828] = 1'b1;  addr_rom[ 3828]='h00000724;  wr_data_rom[ 3828]='h00000d15;
    rd_cycle[ 3829] = 1'b1;  wr_cycle[ 3829] = 1'b0;  addr_rom[ 3829]='h000010c0;  wr_data_rom[ 3829]='h00000000;
    rd_cycle[ 3830] = 1'b1;  wr_cycle[ 3830] = 1'b0;  addr_rom[ 3830]='h00000a18;  wr_data_rom[ 3830]='h00000000;
    rd_cycle[ 3831] = 1'b0;  wr_cycle[ 3831] = 1'b1;  addr_rom[ 3831]='h00000ce0;  wr_data_rom[ 3831]='h00000883;
    rd_cycle[ 3832] = 1'b0;  wr_cycle[ 3832] = 1'b1;  addr_rom[ 3832]='h0000082c;  wr_data_rom[ 3832]='h00000ef4;
    rd_cycle[ 3833] = 1'b1;  wr_cycle[ 3833] = 1'b0;  addr_rom[ 3833]='h000001b8;  wr_data_rom[ 3833]='h00000000;
    rd_cycle[ 3834] = 1'b1;  wr_cycle[ 3834] = 1'b0;  addr_rom[ 3834]='h00000248;  wr_data_rom[ 3834]='h00000000;
    rd_cycle[ 3835] = 1'b0;  wr_cycle[ 3835] = 1'b1;  addr_rom[ 3835]='h00000ab4;  wr_data_rom[ 3835]='h000016c2;
    rd_cycle[ 3836] = 1'b0;  wr_cycle[ 3836] = 1'b1;  addr_rom[ 3836]='h000010dc;  wr_data_rom[ 3836]='h0000100c;
    rd_cycle[ 3837] = 1'b1;  wr_cycle[ 3837] = 1'b0;  addr_rom[ 3837]='h00001b2c;  wr_data_rom[ 3837]='h00000000;
    rd_cycle[ 3838] = 1'b0;  wr_cycle[ 3838] = 1'b1;  addr_rom[ 3838]='h00000890;  wr_data_rom[ 3838]='h00001e81;
    rd_cycle[ 3839] = 1'b0;  wr_cycle[ 3839] = 1'b1;  addr_rom[ 3839]='h00001d80;  wr_data_rom[ 3839]='h00000584;
    rd_cycle[ 3840] = 1'b0;  wr_cycle[ 3840] = 1'b1;  addr_rom[ 3840]='h00001728;  wr_data_rom[ 3840]='h00001270;
    rd_cycle[ 3841] = 1'b1;  wr_cycle[ 3841] = 1'b0;  addr_rom[ 3841]='h00001960;  wr_data_rom[ 3841]='h00000000;
    rd_cycle[ 3842] = 1'b0;  wr_cycle[ 3842] = 1'b1;  addr_rom[ 3842]='h000015dc;  wr_data_rom[ 3842]='h00001cad;
    rd_cycle[ 3843] = 1'b1;  wr_cycle[ 3843] = 1'b0;  addr_rom[ 3843]='h00001c14;  wr_data_rom[ 3843]='h00000000;
    rd_cycle[ 3844] = 1'b1;  wr_cycle[ 3844] = 1'b0;  addr_rom[ 3844]='h00001018;  wr_data_rom[ 3844]='h00000000;
    rd_cycle[ 3845] = 1'b1;  wr_cycle[ 3845] = 1'b0;  addr_rom[ 3845]='h0000076c;  wr_data_rom[ 3845]='h00000000;
    rd_cycle[ 3846] = 1'b0;  wr_cycle[ 3846] = 1'b1;  addr_rom[ 3846]='h00000ef0;  wr_data_rom[ 3846]='h00001204;
    rd_cycle[ 3847] = 1'b0;  wr_cycle[ 3847] = 1'b1;  addr_rom[ 3847]='h00000ac8;  wr_data_rom[ 3847]='h0000195f;
    rd_cycle[ 3848] = 1'b1;  wr_cycle[ 3848] = 1'b0;  addr_rom[ 3848]='h000006b0;  wr_data_rom[ 3848]='h00000000;
    rd_cycle[ 3849] = 1'b0;  wr_cycle[ 3849] = 1'b1;  addr_rom[ 3849]='h00001284;  wr_data_rom[ 3849]='h000015e1;
    rd_cycle[ 3850] = 1'b1;  wr_cycle[ 3850] = 1'b0;  addr_rom[ 3850]='h00001230;  wr_data_rom[ 3850]='h00000000;
    rd_cycle[ 3851] = 1'b0;  wr_cycle[ 3851] = 1'b1;  addr_rom[ 3851]='h00000e40;  wr_data_rom[ 3851]='h000007fa;
    rd_cycle[ 3852] = 1'b0;  wr_cycle[ 3852] = 1'b1;  addr_rom[ 3852]='h00000c8c;  wr_data_rom[ 3852]='h0000071b;
    rd_cycle[ 3853] = 1'b1;  wr_cycle[ 3853] = 1'b0;  addr_rom[ 3853]='h00001a78;  wr_data_rom[ 3853]='h00000000;
    rd_cycle[ 3854] = 1'b0;  wr_cycle[ 3854] = 1'b1;  addr_rom[ 3854]='h0000021c;  wr_data_rom[ 3854]='h000017cd;
    rd_cycle[ 3855] = 1'b0;  wr_cycle[ 3855] = 1'b1;  addr_rom[ 3855]='h00000168;  wr_data_rom[ 3855]='h00000618;
    rd_cycle[ 3856] = 1'b0;  wr_cycle[ 3856] = 1'b1;  addr_rom[ 3856]='h00001820;  wr_data_rom[ 3856]='h0000143f;
    rd_cycle[ 3857] = 1'b1;  wr_cycle[ 3857] = 1'b0;  addr_rom[ 3857]='h000014d4;  wr_data_rom[ 3857]='h00000000;
    rd_cycle[ 3858] = 1'b1;  wr_cycle[ 3858] = 1'b0;  addr_rom[ 3858]='h00000fc8;  wr_data_rom[ 3858]='h00000000;
    rd_cycle[ 3859] = 1'b1;  wr_cycle[ 3859] = 1'b0;  addr_rom[ 3859]='h00001da4;  wr_data_rom[ 3859]='h00000000;
    rd_cycle[ 3860] = 1'b0;  wr_cycle[ 3860] = 1'b1;  addr_rom[ 3860]='h0000141c;  wr_data_rom[ 3860]='h00000012;
    rd_cycle[ 3861] = 1'b1;  wr_cycle[ 3861] = 1'b0;  addr_rom[ 3861]='h00001e70;  wr_data_rom[ 3861]='h00000000;
    rd_cycle[ 3862] = 1'b1;  wr_cycle[ 3862] = 1'b0;  addr_rom[ 3862]='h00000e7c;  wr_data_rom[ 3862]='h00000000;
    rd_cycle[ 3863] = 1'b1;  wr_cycle[ 3863] = 1'b0;  addr_rom[ 3863]='h00001ea8;  wr_data_rom[ 3863]='h00000000;
    rd_cycle[ 3864] = 1'b1;  wr_cycle[ 3864] = 1'b0;  addr_rom[ 3864]='h000013d4;  wr_data_rom[ 3864]='h00000000;
    rd_cycle[ 3865] = 1'b0;  wr_cycle[ 3865] = 1'b1;  addr_rom[ 3865]='h00001edc;  wr_data_rom[ 3865]='h00001bbf;
    rd_cycle[ 3866] = 1'b0;  wr_cycle[ 3866] = 1'b1;  addr_rom[ 3866]='h00000c60;  wr_data_rom[ 3866]='h000018d6;
    rd_cycle[ 3867] = 1'b0;  wr_cycle[ 3867] = 1'b1;  addr_rom[ 3867]='h000013b8;  wr_data_rom[ 3867]='h00000e81;
    rd_cycle[ 3868] = 1'b1;  wr_cycle[ 3868] = 1'b0;  addr_rom[ 3868]='h0000160c;  wr_data_rom[ 3868]='h00000000;
    rd_cycle[ 3869] = 1'b0;  wr_cycle[ 3869] = 1'b1;  addr_rom[ 3869]='h00001e94;  wr_data_rom[ 3869]='h000015f8;
    rd_cycle[ 3870] = 1'b0;  wr_cycle[ 3870] = 1'b1;  addr_rom[ 3870]='h00000448;  wr_data_rom[ 3870]='h00000dff;
    rd_cycle[ 3871] = 1'b0;  wr_cycle[ 3871] = 1'b1;  addr_rom[ 3871]='h000010f0;  wr_data_rom[ 3871]='h000013af;
    rd_cycle[ 3872] = 1'b0;  wr_cycle[ 3872] = 1'b1;  addr_rom[ 3872]='h00000d10;  wr_data_rom[ 3872]='h00001b3c;
    rd_cycle[ 3873] = 1'b0;  wr_cycle[ 3873] = 1'b1;  addr_rom[ 3873]='h00001794;  wr_data_rom[ 3873]='h00000d1a;
    rd_cycle[ 3874] = 1'b0;  wr_cycle[ 3874] = 1'b1;  addr_rom[ 3874]='h00000090;  wr_data_rom[ 3874]='h00000e19;
    rd_cycle[ 3875] = 1'b1;  wr_cycle[ 3875] = 1'b0;  addr_rom[ 3875]='h00000d88;  wr_data_rom[ 3875]='h00000000;
    rd_cycle[ 3876] = 1'b0;  wr_cycle[ 3876] = 1'b1;  addr_rom[ 3876]='h000017c0;  wr_data_rom[ 3876]='h00000c2b;
    rd_cycle[ 3877] = 1'b0;  wr_cycle[ 3877] = 1'b1;  addr_rom[ 3877]='h000019e4;  wr_data_rom[ 3877]='h0000008f;
    rd_cycle[ 3878] = 1'b1;  wr_cycle[ 3878] = 1'b0;  addr_rom[ 3878]='h00000788;  wr_data_rom[ 3878]='h00000000;
    rd_cycle[ 3879] = 1'b1;  wr_cycle[ 3879] = 1'b0;  addr_rom[ 3879]='h0000061c;  wr_data_rom[ 3879]='h00000000;
    rd_cycle[ 3880] = 1'b0;  wr_cycle[ 3880] = 1'b1;  addr_rom[ 3880]='h00000f6c;  wr_data_rom[ 3880]='h000007ab;
    rd_cycle[ 3881] = 1'b1;  wr_cycle[ 3881] = 1'b0;  addr_rom[ 3881]='h00001280;  wr_data_rom[ 3881]='h00000000;
    rd_cycle[ 3882] = 1'b1;  wr_cycle[ 3882] = 1'b0;  addr_rom[ 3882]='h00001b40;  wr_data_rom[ 3882]='h00000000;
    rd_cycle[ 3883] = 1'b1;  wr_cycle[ 3883] = 1'b0;  addr_rom[ 3883]='h00000240;  wr_data_rom[ 3883]='h00000000;
    rd_cycle[ 3884] = 1'b1;  wr_cycle[ 3884] = 1'b0;  addr_rom[ 3884]='h00000e18;  wr_data_rom[ 3884]='h00000000;
    rd_cycle[ 3885] = 1'b0;  wr_cycle[ 3885] = 1'b1;  addr_rom[ 3885]='h00000764;  wr_data_rom[ 3885]='h00001f3b;
    rd_cycle[ 3886] = 1'b1;  wr_cycle[ 3886] = 1'b0;  addr_rom[ 3886]='h00000af8;  wr_data_rom[ 3886]='h00000000;
    rd_cycle[ 3887] = 1'b0;  wr_cycle[ 3887] = 1'b1;  addr_rom[ 3887]='h000004fc;  wr_data_rom[ 3887]='h0000039b;
    rd_cycle[ 3888] = 1'b0;  wr_cycle[ 3888] = 1'b1;  addr_rom[ 3888]='h000000fc;  wr_data_rom[ 3888]='h00001a37;
    rd_cycle[ 3889] = 1'b1;  wr_cycle[ 3889] = 1'b0;  addr_rom[ 3889]='h00001350;  wr_data_rom[ 3889]='h00000000;
    rd_cycle[ 3890] = 1'b1;  wr_cycle[ 3890] = 1'b0;  addr_rom[ 3890]='h00000dd4;  wr_data_rom[ 3890]='h00000000;
    rd_cycle[ 3891] = 1'b0;  wr_cycle[ 3891] = 1'b1;  addr_rom[ 3891]='h000008c0;  wr_data_rom[ 3891]='h000009e7;
    rd_cycle[ 3892] = 1'b0;  wr_cycle[ 3892] = 1'b1;  addr_rom[ 3892]='h00001914;  wr_data_rom[ 3892]='h00000050;
    rd_cycle[ 3893] = 1'b1;  wr_cycle[ 3893] = 1'b0;  addr_rom[ 3893]='h00000d90;  wr_data_rom[ 3893]='h00000000;
    rd_cycle[ 3894] = 1'b1;  wr_cycle[ 3894] = 1'b0;  addr_rom[ 3894]='h00001114;  wr_data_rom[ 3894]='h00000000;
    rd_cycle[ 3895] = 1'b1;  wr_cycle[ 3895] = 1'b0;  addr_rom[ 3895]='h00000d88;  wr_data_rom[ 3895]='h00000000;
    rd_cycle[ 3896] = 1'b0;  wr_cycle[ 3896] = 1'b1;  addr_rom[ 3896]='h0000122c;  wr_data_rom[ 3896]='h00000be6;
    rd_cycle[ 3897] = 1'b0;  wr_cycle[ 3897] = 1'b1;  addr_rom[ 3897]='h00001210;  wr_data_rom[ 3897]='h00001b1d;
    rd_cycle[ 3898] = 1'b1;  wr_cycle[ 3898] = 1'b0;  addr_rom[ 3898]='h00001b20;  wr_data_rom[ 3898]='h00000000;
    rd_cycle[ 3899] = 1'b1;  wr_cycle[ 3899] = 1'b0;  addr_rom[ 3899]='h00000d20;  wr_data_rom[ 3899]='h00000000;
    rd_cycle[ 3900] = 1'b0;  wr_cycle[ 3900] = 1'b1;  addr_rom[ 3900]='h00001adc;  wr_data_rom[ 3900]='h00001878;
    rd_cycle[ 3901] = 1'b0;  wr_cycle[ 3901] = 1'b1;  addr_rom[ 3901]='h00000380;  wr_data_rom[ 3901]='h00000ca4;
    rd_cycle[ 3902] = 1'b0;  wr_cycle[ 3902] = 1'b1;  addr_rom[ 3902]='h00000708;  wr_data_rom[ 3902]='h00000b7c;
    rd_cycle[ 3903] = 1'b1;  wr_cycle[ 3903] = 1'b0;  addr_rom[ 3903]='h00001ca4;  wr_data_rom[ 3903]='h00000000;
    rd_cycle[ 3904] = 1'b0;  wr_cycle[ 3904] = 1'b1;  addr_rom[ 3904]='h000012d8;  wr_data_rom[ 3904]='h000014e0;
    rd_cycle[ 3905] = 1'b1;  wr_cycle[ 3905] = 1'b0;  addr_rom[ 3905]='h00001840;  wr_data_rom[ 3905]='h00000000;
    rd_cycle[ 3906] = 1'b0;  wr_cycle[ 3906] = 1'b1;  addr_rom[ 3906]='h000002a4;  wr_data_rom[ 3906]='h00000c34;
    rd_cycle[ 3907] = 1'b0;  wr_cycle[ 3907] = 1'b1;  addr_rom[ 3907]='h00000c98;  wr_data_rom[ 3907]='h000016e8;
    rd_cycle[ 3908] = 1'b0;  wr_cycle[ 3908] = 1'b1;  addr_rom[ 3908]='h00001b00;  wr_data_rom[ 3908]='h00000257;
    rd_cycle[ 3909] = 1'b0;  wr_cycle[ 3909] = 1'b1;  addr_rom[ 3909]='h00001984;  wr_data_rom[ 3909]='h000017a1;
    rd_cycle[ 3910] = 1'b1;  wr_cycle[ 3910] = 1'b0;  addr_rom[ 3910]='h00000f50;  wr_data_rom[ 3910]='h00000000;
    rd_cycle[ 3911] = 1'b0;  wr_cycle[ 3911] = 1'b1;  addr_rom[ 3911]='h00000580;  wr_data_rom[ 3911]='h0000093d;
    rd_cycle[ 3912] = 1'b1;  wr_cycle[ 3912] = 1'b0;  addr_rom[ 3912]='h00000854;  wr_data_rom[ 3912]='h00000000;
    rd_cycle[ 3913] = 1'b1;  wr_cycle[ 3913] = 1'b0;  addr_rom[ 3913]='h000011f0;  wr_data_rom[ 3913]='h00000000;
    rd_cycle[ 3914] = 1'b1;  wr_cycle[ 3914] = 1'b0;  addr_rom[ 3914]='h00000d74;  wr_data_rom[ 3914]='h00000000;
    rd_cycle[ 3915] = 1'b1;  wr_cycle[ 3915] = 1'b0;  addr_rom[ 3915]='h000011fc;  wr_data_rom[ 3915]='h00000000;
    rd_cycle[ 3916] = 1'b0;  wr_cycle[ 3916] = 1'b1;  addr_rom[ 3916]='h00000c90;  wr_data_rom[ 3916]='h0000045c;
    rd_cycle[ 3917] = 1'b0;  wr_cycle[ 3917] = 1'b1;  addr_rom[ 3917]='h0000069c;  wr_data_rom[ 3917]='h00000fae;
    rd_cycle[ 3918] = 1'b0;  wr_cycle[ 3918] = 1'b1;  addr_rom[ 3918]='h00001f08;  wr_data_rom[ 3918]='h000008b5;
    rd_cycle[ 3919] = 1'b0;  wr_cycle[ 3919] = 1'b1;  addr_rom[ 3919]='h00000800;  wr_data_rom[ 3919]='h00000dc4;
    rd_cycle[ 3920] = 1'b1;  wr_cycle[ 3920] = 1'b0;  addr_rom[ 3920]='h000008a0;  wr_data_rom[ 3920]='h00000000;
    rd_cycle[ 3921] = 1'b1;  wr_cycle[ 3921] = 1'b0;  addr_rom[ 3921]='h00000d9c;  wr_data_rom[ 3921]='h00000000;
    rd_cycle[ 3922] = 1'b0;  wr_cycle[ 3922] = 1'b1;  addr_rom[ 3922]='h0000181c;  wr_data_rom[ 3922]='h00001d2a;
    rd_cycle[ 3923] = 1'b0;  wr_cycle[ 3923] = 1'b1;  addr_rom[ 3923]='h00001488;  wr_data_rom[ 3923]='h00001a34;
    rd_cycle[ 3924] = 1'b0;  wr_cycle[ 3924] = 1'b1;  addr_rom[ 3924]='h00001ce4;  wr_data_rom[ 3924]='h00000807;
    rd_cycle[ 3925] = 1'b1;  wr_cycle[ 3925] = 1'b0;  addr_rom[ 3925]='h0000096c;  wr_data_rom[ 3925]='h00000000;
    rd_cycle[ 3926] = 1'b0;  wr_cycle[ 3926] = 1'b1;  addr_rom[ 3926]='h00000900;  wr_data_rom[ 3926]='h00000165;
    rd_cycle[ 3927] = 1'b1;  wr_cycle[ 3927] = 1'b0;  addr_rom[ 3927]='h00000ed8;  wr_data_rom[ 3927]='h00000000;
    rd_cycle[ 3928] = 1'b0;  wr_cycle[ 3928] = 1'b1;  addr_rom[ 3928]='h0000058c;  wr_data_rom[ 3928]='h00000cc4;
    rd_cycle[ 3929] = 1'b1;  wr_cycle[ 3929] = 1'b0;  addr_rom[ 3929]='h000009a4;  wr_data_rom[ 3929]='h00000000;
    rd_cycle[ 3930] = 1'b0;  wr_cycle[ 3930] = 1'b1;  addr_rom[ 3930]='h000009f0;  wr_data_rom[ 3930]='h00000ca5;
    rd_cycle[ 3931] = 1'b1;  wr_cycle[ 3931] = 1'b0;  addr_rom[ 3931]='h000009f4;  wr_data_rom[ 3931]='h00000000;
    rd_cycle[ 3932] = 1'b0;  wr_cycle[ 3932] = 1'b1;  addr_rom[ 3932]='h0000019c;  wr_data_rom[ 3932]='h00001220;
    rd_cycle[ 3933] = 1'b1;  wr_cycle[ 3933] = 1'b0;  addr_rom[ 3933]='h000018f4;  wr_data_rom[ 3933]='h00000000;
    rd_cycle[ 3934] = 1'b1;  wr_cycle[ 3934] = 1'b0;  addr_rom[ 3934]='h00001cbc;  wr_data_rom[ 3934]='h00000000;
    rd_cycle[ 3935] = 1'b0;  wr_cycle[ 3935] = 1'b1;  addr_rom[ 3935]='h000019e4;  wr_data_rom[ 3935]='h00000434;
    rd_cycle[ 3936] = 1'b0;  wr_cycle[ 3936] = 1'b1;  addr_rom[ 3936]='h00001894;  wr_data_rom[ 3936]='h00000b65;
    rd_cycle[ 3937] = 1'b1;  wr_cycle[ 3937] = 1'b0;  addr_rom[ 3937]='h00000ee0;  wr_data_rom[ 3937]='h00000000;
    rd_cycle[ 3938] = 1'b1;  wr_cycle[ 3938] = 1'b0;  addr_rom[ 3938]='h00000f38;  wr_data_rom[ 3938]='h00000000;
    rd_cycle[ 3939] = 1'b0;  wr_cycle[ 3939] = 1'b1;  addr_rom[ 3939]='h00001a54;  wr_data_rom[ 3939]='h000012a1;
    rd_cycle[ 3940] = 1'b0;  wr_cycle[ 3940] = 1'b1;  addr_rom[ 3940]='h000013d4;  wr_data_rom[ 3940]='h00001e94;
    rd_cycle[ 3941] = 1'b1;  wr_cycle[ 3941] = 1'b0;  addr_rom[ 3941]='h000003a4;  wr_data_rom[ 3941]='h00000000;
    rd_cycle[ 3942] = 1'b0;  wr_cycle[ 3942] = 1'b1;  addr_rom[ 3942]='h00000338;  wr_data_rom[ 3942]='h00000654;
    rd_cycle[ 3943] = 1'b1;  wr_cycle[ 3943] = 1'b0;  addr_rom[ 3943]='h000019cc;  wr_data_rom[ 3943]='h00000000;
    rd_cycle[ 3944] = 1'b1;  wr_cycle[ 3944] = 1'b0;  addr_rom[ 3944]='h00000eec;  wr_data_rom[ 3944]='h00000000;
    rd_cycle[ 3945] = 1'b1;  wr_cycle[ 3945] = 1'b0;  addr_rom[ 3945]='h00001444;  wr_data_rom[ 3945]='h00000000;
    rd_cycle[ 3946] = 1'b1;  wr_cycle[ 3946] = 1'b0;  addr_rom[ 3946]='h00000c18;  wr_data_rom[ 3946]='h00000000;
    rd_cycle[ 3947] = 1'b1;  wr_cycle[ 3947] = 1'b0;  addr_rom[ 3947]='h00001ea8;  wr_data_rom[ 3947]='h00000000;
    rd_cycle[ 3948] = 1'b1;  wr_cycle[ 3948] = 1'b0;  addr_rom[ 3948]='h000001d0;  wr_data_rom[ 3948]='h00000000;
    rd_cycle[ 3949] = 1'b1;  wr_cycle[ 3949] = 1'b0;  addr_rom[ 3949]='h000010ec;  wr_data_rom[ 3949]='h00000000;
    rd_cycle[ 3950] = 1'b0;  wr_cycle[ 3950] = 1'b1;  addr_rom[ 3950]='h00001120;  wr_data_rom[ 3950]='h000018c7;
    rd_cycle[ 3951] = 1'b1;  wr_cycle[ 3951] = 1'b0;  addr_rom[ 3951]='h000006cc;  wr_data_rom[ 3951]='h00000000;
    rd_cycle[ 3952] = 1'b1;  wr_cycle[ 3952] = 1'b0;  addr_rom[ 3952]='h00000410;  wr_data_rom[ 3952]='h00000000;
    rd_cycle[ 3953] = 1'b1;  wr_cycle[ 3953] = 1'b0;  addr_rom[ 3953]='h00001b7c;  wr_data_rom[ 3953]='h00000000;
    rd_cycle[ 3954] = 1'b1;  wr_cycle[ 3954] = 1'b0;  addr_rom[ 3954]='h00001378;  wr_data_rom[ 3954]='h00000000;
    rd_cycle[ 3955] = 1'b0;  wr_cycle[ 3955] = 1'b1;  addr_rom[ 3955]='h00000b04;  wr_data_rom[ 3955]='h00000983;
    rd_cycle[ 3956] = 1'b0;  wr_cycle[ 3956] = 1'b1;  addr_rom[ 3956]='h00000aa0;  wr_data_rom[ 3956]='h00001c4d;
    rd_cycle[ 3957] = 1'b1;  wr_cycle[ 3957] = 1'b0;  addr_rom[ 3957]='h00001b98;  wr_data_rom[ 3957]='h00000000;
    rd_cycle[ 3958] = 1'b0;  wr_cycle[ 3958] = 1'b1;  addr_rom[ 3958]='h00000d68;  wr_data_rom[ 3958]='h000012ef;
    rd_cycle[ 3959] = 1'b0;  wr_cycle[ 3959] = 1'b1;  addr_rom[ 3959]='h00000350;  wr_data_rom[ 3959]='h00001296;
    rd_cycle[ 3960] = 1'b0;  wr_cycle[ 3960] = 1'b1;  addr_rom[ 3960]='h000016dc;  wr_data_rom[ 3960]='h000003a6;
    rd_cycle[ 3961] = 1'b0;  wr_cycle[ 3961] = 1'b1;  addr_rom[ 3961]='h00001294;  wr_data_rom[ 3961]='h0000059a;
    rd_cycle[ 3962] = 1'b1;  wr_cycle[ 3962] = 1'b0;  addr_rom[ 3962]='h000002e8;  wr_data_rom[ 3962]='h00000000;
    rd_cycle[ 3963] = 1'b1;  wr_cycle[ 3963] = 1'b0;  addr_rom[ 3963]='h00000a4c;  wr_data_rom[ 3963]='h00000000;
    rd_cycle[ 3964] = 1'b1;  wr_cycle[ 3964] = 1'b0;  addr_rom[ 3964]='h00000360;  wr_data_rom[ 3964]='h00000000;
    rd_cycle[ 3965] = 1'b1;  wr_cycle[ 3965] = 1'b0;  addr_rom[ 3965]='h00000b3c;  wr_data_rom[ 3965]='h00000000;
    rd_cycle[ 3966] = 1'b1;  wr_cycle[ 3966] = 1'b0;  addr_rom[ 3966]='h00000b14;  wr_data_rom[ 3966]='h00000000;
    rd_cycle[ 3967] = 1'b1;  wr_cycle[ 3967] = 1'b0;  addr_rom[ 3967]='h00000d80;  wr_data_rom[ 3967]='h00000000;
    rd_cycle[ 3968] = 1'b0;  wr_cycle[ 3968] = 1'b1;  addr_rom[ 3968]='h00000c7c;  wr_data_rom[ 3968]='h00000ac0;
    rd_cycle[ 3969] = 1'b0;  wr_cycle[ 3969] = 1'b1;  addr_rom[ 3969]='h0000154c;  wr_data_rom[ 3969]='h000008aa;
    rd_cycle[ 3970] = 1'b1;  wr_cycle[ 3970] = 1'b0;  addr_rom[ 3970]='h00001554;  wr_data_rom[ 3970]='h00000000;
    rd_cycle[ 3971] = 1'b0;  wr_cycle[ 3971] = 1'b1;  addr_rom[ 3971]='h000003f8;  wr_data_rom[ 3971]='h000007f9;
    rd_cycle[ 3972] = 1'b0;  wr_cycle[ 3972] = 1'b1;  addr_rom[ 3972]='h000016d0;  wr_data_rom[ 3972]='h000007ed;
    rd_cycle[ 3973] = 1'b1;  wr_cycle[ 3973] = 1'b0;  addr_rom[ 3973]='h000008dc;  wr_data_rom[ 3973]='h00000000;
    rd_cycle[ 3974] = 1'b1;  wr_cycle[ 3974] = 1'b0;  addr_rom[ 3974]='h0000111c;  wr_data_rom[ 3974]='h00000000;
    rd_cycle[ 3975] = 1'b0;  wr_cycle[ 3975] = 1'b1;  addr_rom[ 3975]='h00000a30;  wr_data_rom[ 3975]='h0000143d;
    rd_cycle[ 3976] = 1'b0;  wr_cycle[ 3976] = 1'b1;  addr_rom[ 3976]='h00001ad8;  wr_data_rom[ 3976]='h00000889;
    rd_cycle[ 3977] = 1'b1;  wr_cycle[ 3977] = 1'b0;  addr_rom[ 3977]='h00000db4;  wr_data_rom[ 3977]='h00000000;
    rd_cycle[ 3978] = 1'b0;  wr_cycle[ 3978] = 1'b1;  addr_rom[ 3978]='h000008d4;  wr_data_rom[ 3978]='h000014fe;
    rd_cycle[ 3979] = 1'b0;  wr_cycle[ 3979] = 1'b1;  addr_rom[ 3979]='h0000059c;  wr_data_rom[ 3979]='h00001741;
    rd_cycle[ 3980] = 1'b0;  wr_cycle[ 3980] = 1'b1;  addr_rom[ 3980]='h00001304;  wr_data_rom[ 3980]='h0000021b;
    rd_cycle[ 3981] = 1'b0;  wr_cycle[ 3981] = 1'b1;  addr_rom[ 3981]='h00000b0c;  wr_data_rom[ 3981]='h00000dd6;
    rd_cycle[ 3982] = 1'b1;  wr_cycle[ 3982] = 1'b0;  addr_rom[ 3982]='h0000146c;  wr_data_rom[ 3982]='h00000000;
    rd_cycle[ 3983] = 1'b1;  wr_cycle[ 3983] = 1'b0;  addr_rom[ 3983]='h0000158c;  wr_data_rom[ 3983]='h00000000;
    rd_cycle[ 3984] = 1'b1;  wr_cycle[ 3984] = 1'b0;  addr_rom[ 3984]='h000014e8;  wr_data_rom[ 3984]='h00000000;
    rd_cycle[ 3985] = 1'b1;  wr_cycle[ 3985] = 1'b0;  addr_rom[ 3985]='h00000a24;  wr_data_rom[ 3985]='h00000000;
    rd_cycle[ 3986] = 1'b0;  wr_cycle[ 3986] = 1'b1;  addr_rom[ 3986]='h000017c0;  wr_data_rom[ 3986]='h00000250;
    rd_cycle[ 3987] = 1'b0;  wr_cycle[ 3987] = 1'b1;  addr_rom[ 3987]='h00001484;  wr_data_rom[ 3987]='h00001afc;
    rd_cycle[ 3988] = 1'b0;  wr_cycle[ 3988] = 1'b1;  addr_rom[ 3988]='h00001c8c;  wr_data_rom[ 3988]='h00000a69;
    rd_cycle[ 3989] = 1'b0;  wr_cycle[ 3989] = 1'b1;  addr_rom[ 3989]='h00001aa0;  wr_data_rom[ 3989]='h00001aab;
    rd_cycle[ 3990] = 1'b1;  wr_cycle[ 3990] = 1'b0;  addr_rom[ 3990]='h00001a18;  wr_data_rom[ 3990]='h00000000;
    rd_cycle[ 3991] = 1'b1;  wr_cycle[ 3991] = 1'b0;  addr_rom[ 3991]='h000014b4;  wr_data_rom[ 3991]='h00000000;
    rd_cycle[ 3992] = 1'b0;  wr_cycle[ 3992] = 1'b1;  addr_rom[ 3992]='h00001b14;  wr_data_rom[ 3992]='h00001717;
    rd_cycle[ 3993] = 1'b1;  wr_cycle[ 3993] = 1'b0;  addr_rom[ 3993]='h0000176c;  wr_data_rom[ 3993]='h00000000;
    rd_cycle[ 3994] = 1'b1;  wr_cycle[ 3994] = 1'b0;  addr_rom[ 3994]='h00001eb0;  wr_data_rom[ 3994]='h00000000;
    rd_cycle[ 3995] = 1'b0;  wr_cycle[ 3995] = 1'b1;  addr_rom[ 3995]='h000011f8;  wr_data_rom[ 3995]='h000019e8;
    rd_cycle[ 3996] = 1'b1;  wr_cycle[ 3996] = 1'b0;  addr_rom[ 3996]='h000007fc;  wr_data_rom[ 3996]='h00000000;
    rd_cycle[ 3997] = 1'b1;  wr_cycle[ 3997] = 1'b0;  addr_rom[ 3997]='h00000dcc;  wr_data_rom[ 3997]='h00000000;
    rd_cycle[ 3998] = 1'b0;  wr_cycle[ 3998] = 1'b1;  addr_rom[ 3998]='h000003b4;  wr_data_rom[ 3998]='h000011bb;
    rd_cycle[ 3999] = 1'b0;  wr_cycle[ 3999] = 1'b1;  addr_rom[ 3999]='h00001174;  wr_data_rom[ 3999]='h00000db6;
    rd_cycle[ 4000] = 1'b1;  wr_cycle[ 4000] = 1'b0;  addr_rom[ 4000]='h000017ac;  wr_data_rom[ 4000]='h00000000;
    rd_cycle[ 4001] = 1'b0;  wr_cycle[ 4001] = 1'b1;  addr_rom[ 4001]='h00000b64;  wr_data_rom[ 4001]='h0000012b;
    rd_cycle[ 4002] = 1'b1;  wr_cycle[ 4002] = 1'b0;  addr_rom[ 4002]='h00001a1c;  wr_data_rom[ 4002]='h00000000;
    rd_cycle[ 4003] = 1'b1;  wr_cycle[ 4003] = 1'b0;  addr_rom[ 4003]='h00000d4c;  wr_data_rom[ 4003]='h00000000;
    rd_cycle[ 4004] = 1'b1;  wr_cycle[ 4004] = 1'b0;  addr_rom[ 4004]='h00001844;  wr_data_rom[ 4004]='h00000000;
    rd_cycle[ 4005] = 1'b1;  wr_cycle[ 4005] = 1'b0;  addr_rom[ 4005]='h00000b18;  wr_data_rom[ 4005]='h00000000;
    rd_cycle[ 4006] = 1'b0;  wr_cycle[ 4006] = 1'b1;  addr_rom[ 4006]='h00001628;  wr_data_rom[ 4006]='h00001d3d;
    rd_cycle[ 4007] = 1'b0;  wr_cycle[ 4007] = 1'b1;  addr_rom[ 4007]='h0000174c;  wr_data_rom[ 4007]='h00001562;
    rd_cycle[ 4008] = 1'b0;  wr_cycle[ 4008] = 1'b1;  addr_rom[ 4008]='h000017fc;  wr_data_rom[ 4008]='h00000626;
    rd_cycle[ 4009] = 1'b1;  wr_cycle[ 4009] = 1'b0;  addr_rom[ 4009]='h00001be8;  wr_data_rom[ 4009]='h00000000;
    rd_cycle[ 4010] = 1'b0;  wr_cycle[ 4010] = 1'b1;  addr_rom[ 4010]='h000000d0;  wr_data_rom[ 4010]='h00000cf0;
    rd_cycle[ 4011] = 1'b0;  wr_cycle[ 4011] = 1'b1;  addr_rom[ 4011]='h000013dc;  wr_data_rom[ 4011]='h0000152f;
    rd_cycle[ 4012] = 1'b0;  wr_cycle[ 4012] = 1'b1;  addr_rom[ 4012]='h000015f4;  wr_data_rom[ 4012]='h00001e06;
    rd_cycle[ 4013] = 1'b0;  wr_cycle[ 4013] = 1'b1;  addr_rom[ 4013]='h00001eec;  wr_data_rom[ 4013]='h00001bf4;
    rd_cycle[ 4014] = 1'b0;  wr_cycle[ 4014] = 1'b1;  addr_rom[ 4014]='h00000afc;  wr_data_rom[ 4014]='h00000a9d;
    rd_cycle[ 4015] = 1'b1;  wr_cycle[ 4015] = 1'b0;  addr_rom[ 4015]='h00001624;  wr_data_rom[ 4015]='h00000000;
    rd_cycle[ 4016] = 1'b0;  wr_cycle[ 4016] = 1'b1;  addr_rom[ 4016]='h000019dc;  wr_data_rom[ 4016]='h000011a6;
    rd_cycle[ 4017] = 1'b0;  wr_cycle[ 4017] = 1'b1;  addr_rom[ 4017]='h0000097c;  wr_data_rom[ 4017]='h00001c13;
    rd_cycle[ 4018] = 1'b1;  wr_cycle[ 4018] = 1'b0;  addr_rom[ 4018]='h00000118;  wr_data_rom[ 4018]='h00000000;
    rd_cycle[ 4019] = 1'b0;  wr_cycle[ 4019] = 1'b1;  addr_rom[ 4019]='h00001cac;  wr_data_rom[ 4019]='h0000049d;
    rd_cycle[ 4020] = 1'b0;  wr_cycle[ 4020] = 1'b1;  addr_rom[ 4020]='h00000010;  wr_data_rom[ 4020]='h00000c86;
    rd_cycle[ 4021] = 1'b1;  wr_cycle[ 4021] = 1'b0;  addr_rom[ 4021]='h00001818;  wr_data_rom[ 4021]='h00000000;
    rd_cycle[ 4022] = 1'b1;  wr_cycle[ 4022] = 1'b0;  addr_rom[ 4022]='h000009b0;  wr_data_rom[ 4022]='h00000000;
    rd_cycle[ 4023] = 1'b1;  wr_cycle[ 4023] = 1'b0;  addr_rom[ 4023]='h00001ca0;  wr_data_rom[ 4023]='h00000000;
    rd_cycle[ 4024] = 1'b0;  wr_cycle[ 4024] = 1'b1;  addr_rom[ 4024]='h000019ac;  wr_data_rom[ 4024]='h000000cb;
    rd_cycle[ 4025] = 1'b0;  wr_cycle[ 4025] = 1'b1;  addr_rom[ 4025]='h00001418;  wr_data_rom[ 4025]='h00000e51;
    rd_cycle[ 4026] = 1'b1;  wr_cycle[ 4026] = 1'b0;  addr_rom[ 4026]='h00000314;  wr_data_rom[ 4026]='h00000000;
    rd_cycle[ 4027] = 1'b0;  wr_cycle[ 4027] = 1'b1;  addr_rom[ 4027]='h00000044;  wr_data_rom[ 4027]='h0000152e;
    rd_cycle[ 4028] = 1'b0;  wr_cycle[ 4028] = 1'b1;  addr_rom[ 4028]='h00000a5c;  wr_data_rom[ 4028]='h00000875;
    rd_cycle[ 4029] = 1'b0;  wr_cycle[ 4029] = 1'b1;  addr_rom[ 4029]='h000003c4;  wr_data_rom[ 4029]='h0000046c;
    rd_cycle[ 4030] = 1'b1;  wr_cycle[ 4030] = 1'b0;  addr_rom[ 4030]='h00000528;  wr_data_rom[ 4030]='h00000000;
    rd_cycle[ 4031] = 1'b0;  wr_cycle[ 4031] = 1'b1;  addr_rom[ 4031]='h000014cc;  wr_data_rom[ 4031]='h00001c64;
    rd_cycle[ 4032] = 1'b0;  wr_cycle[ 4032] = 1'b1;  addr_rom[ 4032]='h000013e8;  wr_data_rom[ 4032]='h00000b9b;
    rd_cycle[ 4033] = 1'b0;  wr_cycle[ 4033] = 1'b1;  addr_rom[ 4033]='h00000bdc;  wr_data_rom[ 4033]='h0000145d;
    rd_cycle[ 4034] = 1'b0;  wr_cycle[ 4034] = 1'b1;  addr_rom[ 4034]='h00000918;  wr_data_rom[ 4034]='h00001c9c;
    rd_cycle[ 4035] = 1'b0;  wr_cycle[ 4035] = 1'b1;  addr_rom[ 4035]='h00000328;  wr_data_rom[ 4035]='h00001b52;
    rd_cycle[ 4036] = 1'b0;  wr_cycle[ 4036] = 1'b1;  addr_rom[ 4036]='h000014a0;  wr_data_rom[ 4036]='h0000111e;
    rd_cycle[ 4037] = 1'b0;  wr_cycle[ 4037] = 1'b1;  addr_rom[ 4037]='h0000049c;  wr_data_rom[ 4037]='h00001239;
    rd_cycle[ 4038] = 1'b1;  wr_cycle[ 4038] = 1'b0;  addr_rom[ 4038]='h00000390;  wr_data_rom[ 4038]='h00000000;
    rd_cycle[ 4039] = 1'b0;  wr_cycle[ 4039] = 1'b1;  addr_rom[ 4039]='h00001ab4;  wr_data_rom[ 4039]='h0000007c;
    rd_cycle[ 4040] = 1'b1;  wr_cycle[ 4040] = 1'b0;  addr_rom[ 4040]='h0000032c;  wr_data_rom[ 4040]='h00000000;
    rd_cycle[ 4041] = 1'b1;  wr_cycle[ 4041] = 1'b0;  addr_rom[ 4041]='h00001254;  wr_data_rom[ 4041]='h00000000;
    rd_cycle[ 4042] = 1'b1;  wr_cycle[ 4042] = 1'b0;  addr_rom[ 4042]='h000019a8;  wr_data_rom[ 4042]='h00000000;
    rd_cycle[ 4043] = 1'b0;  wr_cycle[ 4043] = 1'b1;  addr_rom[ 4043]='h000002ac;  wr_data_rom[ 4043]='h00000240;
    rd_cycle[ 4044] = 1'b0;  wr_cycle[ 4044] = 1'b1;  addr_rom[ 4044]='h000005c8;  wr_data_rom[ 4044]='h000010ff;
    rd_cycle[ 4045] = 1'b0;  wr_cycle[ 4045] = 1'b1;  addr_rom[ 4045]='h00001038;  wr_data_rom[ 4045]='h00001d11;
    rd_cycle[ 4046] = 1'b1;  wr_cycle[ 4046] = 1'b0;  addr_rom[ 4046]='h00000d68;  wr_data_rom[ 4046]='h00000000;
    rd_cycle[ 4047] = 1'b0;  wr_cycle[ 4047] = 1'b1;  addr_rom[ 4047]='h00000840;  wr_data_rom[ 4047]='h00000415;
    rd_cycle[ 4048] = 1'b0;  wr_cycle[ 4048] = 1'b1;  addr_rom[ 4048]='h00001524;  wr_data_rom[ 4048]='h000019be;
    rd_cycle[ 4049] = 1'b1;  wr_cycle[ 4049] = 1'b0;  addr_rom[ 4049]='h00000b10;  wr_data_rom[ 4049]='h00000000;
    rd_cycle[ 4050] = 1'b1;  wr_cycle[ 4050] = 1'b0;  addr_rom[ 4050]='h00001e94;  wr_data_rom[ 4050]='h00000000;
    rd_cycle[ 4051] = 1'b1;  wr_cycle[ 4051] = 1'b0;  addr_rom[ 4051]='h00001d10;  wr_data_rom[ 4051]='h00000000;
    rd_cycle[ 4052] = 1'b1;  wr_cycle[ 4052] = 1'b0;  addr_rom[ 4052]='h00001eb0;  wr_data_rom[ 4052]='h00000000;
    rd_cycle[ 4053] = 1'b1;  wr_cycle[ 4053] = 1'b0;  addr_rom[ 4053]='h00001aac;  wr_data_rom[ 4053]='h00000000;
    rd_cycle[ 4054] = 1'b1;  wr_cycle[ 4054] = 1'b0;  addr_rom[ 4054]='h00001ef0;  wr_data_rom[ 4054]='h00000000;
    rd_cycle[ 4055] = 1'b0;  wr_cycle[ 4055] = 1'b1;  addr_rom[ 4055]='h000018fc;  wr_data_rom[ 4055]='h00000b6d;
    rd_cycle[ 4056] = 1'b1;  wr_cycle[ 4056] = 1'b0;  addr_rom[ 4056]='h0000035c;  wr_data_rom[ 4056]='h00000000;
    rd_cycle[ 4057] = 1'b1;  wr_cycle[ 4057] = 1'b0;  addr_rom[ 4057]='h00000ec4;  wr_data_rom[ 4057]='h00000000;
    rd_cycle[ 4058] = 1'b0;  wr_cycle[ 4058] = 1'b1;  addr_rom[ 4058]='h00001ea4;  wr_data_rom[ 4058]='h00001ad0;
    rd_cycle[ 4059] = 1'b1;  wr_cycle[ 4059] = 1'b0;  addr_rom[ 4059]='h00000b60;  wr_data_rom[ 4059]='h00000000;
    rd_cycle[ 4060] = 1'b1;  wr_cycle[ 4060] = 1'b0;  addr_rom[ 4060]='h00001110;  wr_data_rom[ 4060]='h00000000;
    rd_cycle[ 4061] = 1'b0;  wr_cycle[ 4061] = 1'b1;  addr_rom[ 4061]='h000008a8;  wr_data_rom[ 4061]='h000016cc;
    rd_cycle[ 4062] = 1'b0;  wr_cycle[ 4062] = 1'b1;  addr_rom[ 4062]='h000006c8;  wr_data_rom[ 4062]='h00000266;
    rd_cycle[ 4063] = 1'b1;  wr_cycle[ 4063] = 1'b0;  addr_rom[ 4063]='h00000e18;  wr_data_rom[ 4063]='h00000000;
    rd_cycle[ 4064] = 1'b1;  wr_cycle[ 4064] = 1'b0;  addr_rom[ 4064]='h00001514;  wr_data_rom[ 4064]='h00000000;
    rd_cycle[ 4065] = 1'b1;  wr_cycle[ 4065] = 1'b0;  addr_rom[ 4065]='h00000358;  wr_data_rom[ 4065]='h00000000;
    rd_cycle[ 4066] = 1'b0;  wr_cycle[ 4066] = 1'b1;  addr_rom[ 4066]='h000019dc;  wr_data_rom[ 4066]='h00000ea6;
    rd_cycle[ 4067] = 1'b0;  wr_cycle[ 4067] = 1'b1;  addr_rom[ 4067]='h0000121c;  wr_data_rom[ 4067]='h00000b23;
    rd_cycle[ 4068] = 1'b0;  wr_cycle[ 4068] = 1'b1;  addr_rom[ 4068]='h00000304;  wr_data_rom[ 4068]='h00001c02;
    rd_cycle[ 4069] = 1'b0;  wr_cycle[ 4069] = 1'b1;  addr_rom[ 4069]='h00000b84;  wr_data_rom[ 4069]='h00000781;
    rd_cycle[ 4070] = 1'b1;  wr_cycle[ 4070] = 1'b0;  addr_rom[ 4070]='h00000a00;  wr_data_rom[ 4070]='h00000000;
    rd_cycle[ 4071] = 1'b0;  wr_cycle[ 4071] = 1'b1;  addr_rom[ 4071]='h00001f14;  wr_data_rom[ 4071]='h00000c45;
    rd_cycle[ 4072] = 1'b1;  wr_cycle[ 4072] = 1'b0;  addr_rom[ 4072]='h00001014;  wr_data_rom[ 4072]='h00000000;
    rd_cycle[ 4073] = 1'b1;  wr_cycle[ 4073] = 1'b0;  addr_rom[ 4073]='h000001ec;  wr_data_rom[ 4073]='h00000000;
    rd_cycle[ 4074] = 1'b0;  wr_cycle[ 4074] = 1'b1;  addr_rom[ 4074]='h000014c8;  wr_data_rom[ 4074]='h0000042c;
    rd_cycle[ 4075] = 1'b1;  wr_cycle[ 4075] = 1'b0;  addr_rom[ 4075]='h000000e0;  wr_data_rom[ 4075]='h00000000;
    rd_cycle[ 4076] = 1'b1;  wr_cycle[ 4076] = 1'b0;  addr_rom[ 4076]='h00001ea4;  wr_data_rom[ 4076]='h00000000;
    rd_cycle[ 4077] = 1'b0;  wr_cycle[ 4077] = 1'b1;  addr_rom[ 4077]='h000001cc;  wr_data_rom[ 4077]='h00000411;
    rd_cycle[ 4078] = 1'b0;  wr_cycle[ 4078] = 1'b1;  addr_rom[ 4078]='h00001aa8;  wr_data_rom[ 4078]='h00000651;
    rd_cycle[ 4079] = 1'b0;  wr_cycle[ 4079] = 1'b1;  addr_rom[ 4079]='h00001184;  wr_data_rom[ 4079]='h00000116;
    rd_cycle[ 4080] = 1'b1;  wr_cycle[ 4080] = 1'b0;  addr_rom[ 4080]='h00001630;  wr_data_rom[ 4080]='h00000000;
    rd_cycle[ 4081] = 1'b1;  wr_cycle[ 4081] = 1'b0;  addr_rom[ 4081]='h00001348;  wr_data_rom[ 4081]='h00000000;
    rd_cycle[ 4082] = 1'b1;  wr_cycle[ 4082] = 1'b0;  addr_rom[ 4082]='h00001b80;  wr_data_rom[ 4082]='h00000000;
    rd_cycle[ 4083] = 1'b1;  wr_cycle[ 4083] = 1'b0;  addr_rom[ 4083]='h00001018;  wr_data_rom[ 4083]='h00000000;
    rd_cycle[ 4084] = 1'b1;  wr_cycle[ 4084] = 1'b0;  addr_rom[ 4084]='h000002c4;  wr_data_rom[ 4084]='h00000000;
    rd_cycle[ 4085] = 1'b1;  wr_cycle[ 4085] = 1'b0;  addr_rom[ 4085]='h00000ad4;  wr_data_rom[ 4085]='h00000000;
    rd_cycle[ 4086] = 1'b0;  wr_cycle[ 4086] = 1'b1;  addr_rom[ 4086]='h000016f8;  wr_data_rom[ 4086]='h0000051b;
    rd_cycle[ 4087] = 1'b0;  wr_cycle[ 4087] = 1'b1;  addr_rom[ 4087]='h00001764;  wr_data_rom[ 4087]='h000000c2;
    rd_cycle[ 4088] = 1'b0;  wr_cycle[ 4088] = 1'b1;  addr_rom[ 4088]='h00000fb0;  wr_data_rom[ 4088]='h00000857;
    rd_cycle[ 4089] = 1'b0;  wr_cycle[ 4089] = 1'b1;  addr_rom[ 4089]='h00000728;  wr_data_rom[ 4089]='h00001bf3;
    rd_cycle[ 4090] = 1'b1;  wr_cycle[ 4090] = 1'b0;  addr_rom[ 4090]='h0000060c;  wr_data_rom[ 4090]='h00000000;
    rd_cycle[ 4091] = 1'b0;  wr_cycle[ 4091] = 1'b1;  addr_rom[ 4091]='h00001a24;  wr_data_rom[ 4091]='h00000c2e;
    rd_cycle[ 4092] = 1'b1;  wr_cycle[ 4092] = 1'b0;  addr_rom[ 4092]='h000007b0;  wr_data_rom[ 4092]='h00000000;
    rd_cycle[ 4093] = 1'b1;  wr_cycle[ 4093] = 1'b0;  addr_rom[ 4093]='h000007c8;  wr_data_rom[ 4093]='h00000000;
    rd_cycle[ 4094] = 1'b0;  wr_cycle[ 4094] = 1'b1;  addr_rom[ 4094]='h000018d4;  wr_data_rom[ 4094]='h00001d2d;
    rd_cycle[ 4095] = 1'b1;  wr_cycle[ 4095] = 1'b0;  addr_rom[ 4095]='h00000264;  wr_data_rom[ 4095]='h00000000;
    rd_cycle[ 4096] = 1'b1;  wr_cycle[ 4096] = 1'b0;  addr_rom[ 4096]='h00001570;  wr_data_rom[ 4096]='h00000000;
    rd_cycle[ 4097] = 1'b1;  wr_cycle[ 4097] = 1'b0;  addr_rom[ 4097]='h00001560;  wr_data_rom[ 4097]='h00000000;
    rd_cycle[ 4098] = 1'b0;  wr_cycle[ 4098] = 1'b1;  addr_rom[ 4098]='h00000378;  wr_data_rom[ 4098]='h00001aa0;
    rd_cycle[ 4099] = 1'b1;  wr_cycle[ 4099] = 1'b0;  addr_rom[ 4099]='h00001a98;  wr_data_rom[ 4099]='h00000000;
    rd_cycle[ 4100] = 1'b1;  wr_cycle[ 4100] = 1'b0;  addr_rom[ 4100]='h000014e0;  wr_data_rom[ 4100]='h00000000;
    rd_cycle[ 4101] = 1'b1;  wr_cycle[ 4101] = 1'b0;  addr_rom[ 4101]='h000005b8;  wr_data_rom[ 4101]='h00000000;
    rd_cycle[ 4102] = 1'b0;  wr_cycle[ 4102] = 1'b1;  addr_rom[ 4102]='h00001124;  wr_data_rom[ 4102]='h00000021;
    rd_cycle[ 4103] = 1'b0;  wr_cycle[ 4103] = 1'b1;  addr_rom[ 4103]='h00000808;  wr_data_rom[ 4103]='h000012a4;
    rd_cycle[ 4104] = 1'b1;  wr_cycle[ 4104] = 1'b0;  addr_rom[ 4104]='h00000ba0;  wr_data_rom[ 4104]='h00000000;
    rd_cycle[ 4105] = 1'b1;  wr_cycle[ 4105] = 1'b0;  addr_rom[ 4105]='h0000107c;  wr_data_rom[ 4105]='h00000000;
    rd_cycle[ 4106] = 1'b1;  wr_cycle[ 4106] = 1'b0;  addr_rom[ 4106]='h000019d0;  wr_data_rom[ 4106]='h00000000;
    rd_cycle[ 4107] = 1'b1;  wr_cycle[ 4107] = 1'b0;  addr_rom[ 4107]='h00001584;  wr_data_rom[ 4107]='h00000000;
    rd_cycle[ 4108] = 1'b1;  wr_cycle[ 4108] = 1'b0;  addr_rom[ 4108]='h000016b8;  wr_data_rom[ 4108]='h00000000;
    rd_cycle[ 4109] = 1'b1;  wr_cycle[ 4109] = 1'b0;  addr_rom[ 4109]='h000016ac;  wr_data_rom[ 4109]='h00000000;
    rd_cycle[ 4110] = 1'b0;  wr_cycle[ 4110] = 1'b1;  addr_rom[ 4110]='h00000b28;  wr_data_rom[ 4110]='h0000064f;
    rd_cycle[ 4111] = 1'b0;  wr_cycle[ 4111] = 1'b1;  addr_rom[ 4111]='h00001c7c;  wr_data_rom[ 4111]='h000016fa;
    rd_cycle[ 4112] = 1'b1;  wr_cycle[ 4112] = 1'b0;  addr_rom[ 4112]='h00000334;  wr_data_rom[ 4112]='h00000000;
    rd_cycle[ 4113] = 1'b0;  wr_cycle[ 4113] = 1'b1;  addr_rom[ 4113]='h000011d4;  wr_data_rom[ 4113]='h0000110b;
    rd_cycle[ 4114] = 1'b0;  wr_cycle[ 4114] = 1'b1;  addr_rom[ 4114]='h00000ce0;  wr_data_rom[ 4114]='h00001c37;
    rd_cycle[ 4115] = 1'b1;  wr_cycle[ 4115] = 1'b0;  addr_rom[ 4115]='h00000440;  wr_data_rom[ 4115]='h00000000;
    rd_cycle[ 4116] = 1'b0;  wr_cycle[ 4116] = 1'b1;  addr_rom[ 4116]='h00001848;  wr_data_rom[ 4116]='h00000e4f;
    rd_cycle[ 4117] = 1'b1;  wr_cycle[ 4117] = 1'b0;  addr_rom[ 4117]='h00000914;  wr_data_rom[ 4117]='h00000000;
    rd_cycle[ 4118] = 1'b1;  wr_cycle[ 4118] = 1'b0;  addr_rom[ 4118]='h00001018;  wr_data_rom[ 4118]='h00000000;
    rd_cycle[ 4119] = 1'b0;  wr_cycle[ 4119] = 1'b1;  addr_rom[ 4119]='h0000083c;  wr_data_rom[ 4119]='h00000cdb;
    rd_cycle[ 4120] = 1'b0;  wr_cycle[ 4120] = 1'b1;  addr_rom[ 4120]='h00001e80;  wr_data_rom[ 4120]='h0000117c;
    rd_cycle[ 4121] = 1'b0;  wr_cycle[ 4121] = 1'b1;  addr_rom[ 4121]='h00001db4;  wr_data_rom[ 4121]='h00001126;
    rd_cycle[ 4122] = 1'b1;  wr_cycle[ 4122] = 1'b0;  addr_rom[ 4122]='h000005c0;  wr_data_rom[ 4122]='h00000000;
    rd_cycle[ 4123] = 1'b1;  wr_cycle[ 4123] = 1'b0;  addr_rom[ 4123]='h00000060;  wr_data_rom[ 4123]='h00000000;
    rd_cycle[ 4124] = 1'b1;  wr_cycle[ 4124] = 1'b0;  addr_rom[ 4124]='h000011b4;  wr_data_rom[ 4124]='h00000000;
    rd_cycle[ 4125] = 1'b0;  wr_cycle[ 4125] = 1'b1;  addr_rom[ 4125]='h00001c4c;  wr_data_rom[ 4125]='h00001b7d;
    rd_cycle[ 4126] = 1'b1;  wr_cycle[ 4126] = 1'b0;  addr_rom[ 4126]='h00000eac;  wr_data_rom[ 4126]='h00000000;
    rd_cycle[ 4127] = 1'b0;  wr_cycle[ 4127] = 1'b1;  addr_rom[ 4127]='h00001e3c;  wr_data_rom[ 4127]='h00001227;
    rd_cycle[ 4128] = 1'b0;  wr_cycle[ 4128] = 1'b1;  addr_rom[ 4128]='h00000aa0;  wr_data_rom[ 4128]='h00000090;
    rd_cycle[ 4129] = 1'b1;  wr_cycle[ 4129] = 1'b0;  addr_rom[ 4129]='h000006b8;  wr_data_rom[ 4129]='h00000000;
    rd_cycle[ 4130] = 1'b1;  wr_cycle[ 4130] = 1'b0;  addr_rom[ 4130]='h00001a70;  wr_data_rom[ 4130]='h00000000;
    rd_cycle[ 4131] = 1'b0;  wr_cycle[ 4131] = 1'b1;  addr_rom[ 4131]='h00000a40;  wr_data_rom[ 4131]='h000001a9;
    rd_cycle[ 4132] = 1'b1;  wr_cycle[ 4132] = 1'b0;  addr_rom[ 4132]='h00001c9c;  wr_data_rom[ 4132]='h00000000;
    rd_cycle[ 4133] = 1'b0;  wr_cycle[ 4133] = 1'b1;  addr_rom[ 4133]='h0000093c;  wr_data_rom[ 4133]='h000005ab;
    rd_cycle[ 4134] = 1'b1;  wr_cycle[ 4134] = 1'b0;  addr_rom[ 4134]='h00000938;  wr_data_rom[ 4134]='h00000000;
    rd_cycle[ 4135] = 1'b1;  wr_cycle[ 4135] = 1'b0;  addr_rom[ 4135]='h00001ba4;  wr_data_rom[ 4135]='h00000000;
    rd_cycle[ 4136] = 1'b0;  wr_cycle[ 4136] = 1'b1;  addr_rom[ 4136]='h000017fc;  wr_data_rom[ 4136]='h00001adf;
    rd_cycle[ 4137] = 1'b1;  wr_cycle[ 4137] = 1'b0;  addr_rom[ 4137]='h00001a68;  wr_data_rom[ 4137]='h00000000;
    rd_cycle[ 4138] = 1'b0;  wr_cycle[ 4138] = 1'b1;  addr_rom[ 4138]='h0000111c;  wr_data_rom[ 4138]='h000016ce;
    rd_cycle[ 4139] = 1'b0;  wr_cycle[ 4139] = 1'b1;  addr_rom[ 4139]='h0000027c;  wr_data_rom[ 4139]='h00001098;
    rd_cycle[ 4140] = 1'b0;  wr_cycle[ 4140] = 1'b1;  addr_rom[ 4140]='h000011fc;  wr_data_rom[ 4140]='h00001068;
    rd_cycle[ 4141] = 1'b1;  wr_cycle[ 4141] = 1'b0;  addr_rom[ 4141]='h00001dec;  wr_data_rom[ 4141]='h00000000;
    rd_cycle[ 4142] = 1'b0;  wr_cycle[ 4142] = 1'b1;  addr_rom[ 4142]='h00000f54;  wr_data_rom[ 4142]='h0000072d;
    rd_cycle[ 4143] = 1'b1;  wr_cycle[ 4143] = 1'b0;  addr_rom[ 4143]='h0000114c;  wr_data_rom[ 4143]='h00000000;
    rd_cycle[ 4144] = 1'b0;  wr_cycle[ 4144] = 1'b1;  addr_rom[ 4144]='h00000844;  wr_data_rom[ 4144]='h0000134c;
    rd_cycle[ 4145] = 1'b1;  wr_cycle[ 4145] = 1'b0;  addr_rom[ 4145]='h00000cc0;  wr_data_rom[ 4145]='h00000000;
    rd_cycle[ 4146] = 1'b0;  wr_cycle[ 4146] = 1'b1;  addr_rom[ 4146]='h00000440;  wr_data_rom[ 4146]='h00001502;
    rd_cycle[ 4147] = 1'b0;  wr_cycle[ 4147] = 1'b1;  addr_rom[ 4147]='h000016d0;  wr_data_rom[ 4147]='h00001a1a;
    rd_cycle[ 4148] = 1'b1;  wr_cycle[ 4148] = 1'b0;  addr_rom[ 4148]='h000008dc;  wr_data_rom[ 4148]='h00000000;
    rd_cycle[ 4149] = 1'b1;  wr_cycle[ 4149] = 1'b0;  addr_rom[ 4149]='h00001910;  wr_data_rom[ 4149]='h00000000;
    rd_cycle[ 4150] = 1'b0;  wr_cycle[ 4150] = 1'b1;  addr_rom[ 4150]='h00000328;  wr_data_rom[ 4150]='h00001423;
    rd_cycle[ 4151] = 1'b1;  wr_cycle[ 4151] = 1'b0;  addr_rom[ 4151]='h000014f8;  wr_data_rom[ 4151]='h00000000;
    rd_cycle[ 4152] = 1'b0;  wr_cycle[ 4152] = 1'b1;  addr_rom[ 4152]='h00001ce4;  wr_data_rom[ 4152]='h00001c31;
    rd_cycle[ 4153] = 1'b1;  wr_cycle[ 4153] = 1'b0;  addr_rom[ 4153]='h000006d8;  wr_data_rom[ 4153]='h00000000;
    rd_cycle[ 4154] = 1'b1;  wr_cycle[ 4154] = 1'b0;  addr_rom[ 4154]='h00001334;  wr_data_rom[ 4154]='h00000000;
    rd_cycle[ 4155] = 1'b1;  wr_cycle[ 4155] = 1'b0;  addr_rom[ 4155]='h0000045c;  wr_data_rom[ 4155]='h00000000;
    rd_cycle[ 4156] = 1'b0;  wr_cycle[ 4156] = 1'b1;  addr_rom[ 4156]='h00001560;  wr_data_rom[ 4156]='h000002ed;
    rd_cycle[ 4157] = 1'b0;  wr_cycle[ 4157] = 1'b1;  addr_rom[ 4157]='h00000b5c;  wr_data_rom[ 4157]='h0000141d;
    rd_cycle[ 4158] = 1'b0;  wr_cycle[ 4158] = 1'b1;  addr_rom[ 4158]='h00001ed4;  wr_data_rom[ 4158]='h0000154f;
    rd_cycle[ 4159] = 1'b0;  wr_cycle[ 4159] = 1'b1;  addr_rom[ 4159]='h00001258;  wr_data_rom[ 4159]='h00000905;
    rd_cycle[ 4160] = 1'b1;  wr_cycle[ 4160] = 1'b0;  addr_rom[ 4160]='h00000ff8;  wr_data_rom[ 4160]='h00000000;
    rd_cycle[ 4161] = 1'b0;  wr_cycle[ 4161] = 1'b1;  addr_rom[ 4161]='h00000fe8;  wr_data_rom[ 4161]='h000013b6;
    rd_cycle[ 4162] = 1'b0;  wr_cycle[ 4162] = 1'b1;  addr_rom[ 4162]='h00001bc4;  wr_data_rom[ 4162]='h0000169c;
    rd_cycle[ 4163] = 1'b1;  wr_cycle[ 4163] = 1'b0;  addr_rom[ 4163]='h000017dc;  wr_data_rom[ 4163]='h00000000;
    rd_cycle[ 4164] = 1'b0;  wr_cycle[ 4164] = 1'b1;  addr_rom[ 4164]='h000019b4;  wr_data_rom[ 4164]='h000007f2;
    rd_cycle[ 4165] = 1'b0;  wr_cycle[ 4165] = 1'b1;  addr_rom[ 4165]='h00000374;  wr_data_rom[ 4165]='h00001117;
    rd_cycle[ 4166] = 1'b1;  wr_cycle[ 4166] = 1'b0;  addr_rom[ 4166]='h00000e00;  wr_data_rom[ 4166]='h00000000;
    rd_cycle[ 4167] = 1'b1;  wr_cycle[ 4167] = 1'b0;  addr_rom[ 4167]='h000003f8;  wr_data_rom[ 4167]='h00000000;
    rd_cycle[ 4168] = 1'b0;  wr_cycle[ 4168] = 1'b1;  addr_rom[ 4168]='h00000f40;  wr_data_rom[ 4168]='h00001254;
    rd_cycle[ 4169] = 1'b0;  wr_cycle[ 4169] = 1'b1;  addr_rom[ 4169]='h000005b4;  wr_data_rom[ 4169]='h00001488;
    rd_cycle[ 4170] = 1'b0;  wr_cycle[ 4170] = 1'b1;  addr_rom[ 4170]='h00000fc4;  wr_data_rom[ 4170]='h00000179;
    rd_cycle[ 4171] = 1'b1;  wr_cycle[ 4171] = 1'b0;  addr_rom[ 4171]='h00001da8;  wr_data_rom[ 4171]='h00000000;
    rd_cycle[ 4172] = 1'b1;  wr_cycle[ 4172] = 1'b0;  addr_rom[ 4172]='h000013e4;  wr_data_rom[ 4172]='h00000000;
    rd_cycle[ 4173] = 1'b0;  wr_cycle[ 4173] = 1'b1;  addr_rom[ 4173]='h0000085c;  wr_data_rom[ 4173]='h00000376;
    rd_cycle[ 4174] = 1'b1;  wr_cycle[ 4174] = 1'b0;  addr_rom[ 4174]='h00001b10;  wr_data_rom[ 4174]='h00000000;
    rd_cycle[ 4175] = 1'b0;  wr_cycle[ 4175] = 1'b1;  addr_rom[ 4175]='h00001cc8;  wr_data_rom[ 4175]='h000011c0;
    rd_cycle[ 4176] = 1'b1;  wr_cycle[ 4176] = 1'b0;  addr_rom[ 4176]='h0000068c;  wr_data_rom[ 4176]='h00000000;
    rd_cycle[ 4177] = 1'b0;  wr_cycle[ 4177] = 1'b1;  addr_rom[ 4177]='h00000970;  wr_data_rom[ 4177]='h0000144c;
    rd_cycle[ 4178] = 1'b1;  wr_cycle[ 4178] = 1'b0;  addr_rom[ 4178]='h00000fc0;  wr_data_rom[ 4178]='h00000000;
    rd_cycle[ 4179] = 1'b1;  wr_cycle[ 4179] = 1'b0;  addr_rom[ 4179]='h00000d18;  wr_data_rom[ 4179]='h00000000;
    rd_cycle[ 4180] = 1'b0;  wr_cycle[ 4180] = 1'b1;  addr_rom[ 4180]='h000003c8;  wr_data_rom[ 4180]='h00000d23;
    rd_cycle[ 4181] = 1'b1;  wr_cycle[ 4181] = 1'b0;  addr_rom[ 4181]='h000018ac;  wr_data_rom[ 4181]='h00000000;
    rd_cycle[ 4182] = 1'b1;  wr_cycle[ 4182] = 1'b0;  addr_rom[ 4182]='h00001af8;  wr_data_rom[ 4182]='h00000000;
    rd_cycle[ 4183] = 1'b1;  wr_cycle[ 4183] = 1'b0;  addr_rom[ 4183]='h0000129c;  wr_data_rom[ 4183]='h00000000;
    rd_cycle[ 4184] = 1'b1;  wr_cycle[ 4184] = 1'b0;  addr_rom[ 4184]='h00001a74;  wr_data_rom[ 4184]='h00000000;
    rd_cycle[ 4185] = 1'b0;  wr_cycle[ 4185] = 1'b1;  addr_rom[ 4185]='h000012cc;  wr_data_rom[ 4185]='h00001834;
    rd_cycle[ 4186] = 1'b0;  wr_cycle[ 4186] = 1'b1;  addr_rom[ 4186]='h0000077c;  wr_data_rom[ 4186]='h00000eb0;
    rd_cycle[ 4187] = 1'b0;  wr_cycle[ 4187] = 1'b1;  addr_rom[ 4187]='h00001628;  wr_data_rom[ 4187]='h00001ba8;
    rd_cycle[ 4188] = 1'b1;  wr_cycle[ 4188] = 1'b0;  addr_rom[ 4188]='h00001f30;  wr_data_rom[ 4188]='h00000000;
    rd_cycle[ 4189] = 1'b1;  wr_cycle[ 4189] = 1'b0;  addr_rom[ 4189]='h00000b50;  wr_data_rom[ 4189]='h00000000;
    rd_cycle[ 4190] = 1'b1;  wr_cycle[ 4190] = 1'b0;  addr_rom[ 4190]='h0000154c;  wr_data_rom[ 4190]='h00000000;
    rd_cycle[ 4191] = 1'b1;  wr_cycle[ 4191] = 1'b0;  addr_rom[ 4191]='h000007a8;  wr_data_rom[ 4191]='h00000000;
    rd_cycle[ 4192] = 1'b0;  wr_cycle[ 4192] = 1'b1;  addr_rom[ 4192]='h00000528;  wr_data_rom[ 4192]='h000017c3;
    rd_cycle[ 4193] = 1'b0;  wr_cycle[ 4193] = 1'b1;  addr_rom[ 4193]='h00000f7c;  wr_data_rom[ 4193]='h0000011b;
    rd_cycle[ 4194] = 1'b0;  wr_cycle[ 4194] = 1'b1;  addr_rom[ 4194]='h00000178;  wr_data_rom[ 4194]='h000016d9;
    rd_cycle[ 4195] = 1'b0;  wr_cycle[ 4195] = 1'b1;  addr_rom[ 4195]='h00000588;  wr_data_rom[ 4195]='h00000b0f;
    rd_cycle[ 4196] = 1'b0;  wr_cycle[ 4196] = 1'b1;  addr_rom[ 4196]='h00000580;  wr_data_rom[ 4196]='h00001d7b;
    rd_cycle[ 4197] = 1'b1;  wr_cycle[ 4197] = 1'b0;  addr_rom[ 4197]='h000005b8;  wr_data_rom[ 4197]='h00000000;
    rd_cycle[ 4198] = 1'b1;  wr_cycle[ 4198] = 1'b0;  addr_rom[ 4198]='h000004d8;  wr_data_rom[ 4198]='h00000000;
    rd_cycle[ 4199] = 1'b0;  wr_cycle[ 4199] = 1'b1;  addr_rom[ 4199]='h0000076c;  wr_data_rom[ 4199]='h0000197f;
    rd_cycle[ 4200] = 1'b0;  wr_cycle[ 4200] = 1'b1;  addr_rom[ 4200]='h00001194;  wr_data_rom[ 4200]='h000011e4;
    rd_cycle[ 4201] = 1'b0;  wr_cycle[ 4201] = 1'b1;  addr_rom[ 4201]='h00000834;  wr_data_rom[ 4201]='h00000902;
    rd_cycle[ 4202] = 1'b0;  wr_cycle[ 4202] = 1'b1;  addr_rom[ 4202]='h00000374;  wr_data_rom[ 4202]='h00000521;
    rd_cycle[ 4203] = 1'b0;  wr_cycle[ 4203] = 1'b1;  addr_rom[ 4203]='h000000e8;  wr_data_rom[ 4203]='h00000f0d;
    rd_cycle[ 4204] = 1'b1;  wr_cycle[ 4204] = 1'b0;  addr_rom[ 4204]='h00001870;  wr_data_rom[ 4204]='h00000000;
    rd_cycle[ 4205] = 1'b1;  wr_cycle[ 4205] = 1'b0;  addr_rom[ 4205]='h00001398;  wr_data_rom[ 4205]='h00000000;
    rd_cycle[ 4206] = 1'b0;  wr_cycle[ 4206] = 1'b1;  addr_rom[ 4206]='h00001410;  wr_data_rom[ 4206]='h00001d38;
    rd_cycle[ 4207] = 1'b1;  wr_cycle[ 4207] = 1'b0;  addr_rom[ 4207]='h00000d28;  wr_data_rom[ 4207]='h00000000;
    rd_cycle[ 4208] = 1'b0;  wr_cycle[ 4208] = 1'b1;  addr_rom[ 4208]='h00000dcc;  wr_data_rom[ 4208]='h00000b43;
    rd_cycle[ 4209] = 1'b1;  wr_cycle[ 4209] = 1'b0;  addr_rom[ 4209]='h00001848;  wr_data_rom[ 4209]='h00000000;
    rd_cycle[ 4210] = 1'b0;  wr_cycle[ 4210] = 1'b1;  addr_rom[ 4210]='h00001534;  wr_data_rom[ 4210]='h00001732;
    rd_cycle[ 4211] = 1'b0;  wr_cycle[ 4211] = 1'b1;  addr_rom[ 4211]='h0000099c;  wr_data_rom[ 4211]='h00001ea9;
    rd_cycle[ 4212] = 1'b1;  wr_cycle[ 4212] = 1'b0;  addr_rom[ 4212]='h00001ef4;  wr_data_rom[ 4212]='h00000000;
    rd_cycle[ 4213] = 1'b0;  wr_cycle[ 4213] = 1'b1;  addr_rom[ 4213]='h000001e8;  wr_data_rom[ 4213]='h000016f7;
    rd_cycle[ 4214] = 1'b0;  wr_cycle[ 4214] = 1'b1;  addr_rom[ 4214]='h00001810;  wr_data_rom[ 4214]='h000010b6;
    rd_cycle[ 4215] = 1'b0;  wr_cycle[ 4215] = 1'b1;  addr_rom[ 4215]='h00001e6c;  wr_data_rom[ 4215]='h0000008e;
    rd_cycle[ 4216] = 1'b0;  wr_cycle[ 4216] = 1'b1;  addr_rom[ 4216]='h000018e8;  wr_data_rom[ 4216]='h000012a4;
    rd_cycle[ 4217] = 1'b0;  wr_cycle[ 4217] = 1'b1;  addr_rom[ 4217]='h00000ce4;  wr_data_rom[ 4217]='h000007f0;
    rd_cycle[ 4218] = 1'b0;  wr_cycle[ 4218] = 1'b1;  addr_rom[ 4218]='h00000f74;  wr_data_rom[ 4218]='h00000728;
    rd_cycle[ 4219] = 1'b0;  wr_cycle[ 4219] = 1'b1;  addr_rom[ 4219]='h00000198;  wr_data_rom[ 4219]='h00000616;
    rd_cycle[ 4220] = 1'b1;  wr_cycle[ 4220] = 1'b0;  addr_rom[ 4220]='h00001dc0;  wr_data_rom[ 4220]='h00000000;
    rd_cycle[ 4221] = 1'b0;  wr_cycle[ 4221] = 1'b1;  addr_rom[ 4221]='h000015d4;  wr_data_rom[ 4221]='h00000a1c;
    rd_cycle[ 4222] = 1'b1;  wr_cycle[ 4222] = 1'b0;  addr_rom[ 4222]='h000008f0;  wr_data_rom[ 4222]='h00000000;
    rd_cycle[ 4223] = 1'b1;  wr_cycle[ 4223] = 1'b0;  addr_rom[ 4223]='h00000e98;  wr_data_rom[ 4223]='h00000000;
    rd_cycle[ 4224] = 1'b1;  wr_cycle[ 4224] = 1'b0;  addr_rom[ 4224]='h00001f0c;  wr_data_rom[ 4224]='h00000000;
    rd_cycle[ 4225] = 1'b0;  wr_cycle[ 4225] = 1'b1;  addr_rom[ 4225]='h000018a0;  wr_data_rom[ 4225]='h000008e5;
    rd_cycle[ 4226] = 1'b1;  wr_cycle[ 4226] = 1'b0;  addr_rom[ 4226]='h000016d4;  wr_data_rom[ 4226]='h00000000;
    rd_cycle[ 4227] = 1'b1;  wr_cycle[ 4227] = 1'b0;  addr_rom[ 4227]='h00001370;  wr_data_rom[ 4227]='h00000000;
    rd_cycle[ 4228] = 1'b1;  wr_cycle[ 4228] = 1'b0;  addr_rom[ 4228]='h00000844;  wr_data_rom[ 4228]='h00000000;
    rd_cycle[ 4229] = 1'b0;  wr_cycle[ 4229] = 1'b1;  addr_rom[ 4229]='h000003b4;  wr_data_rom[ 4229]='h00001d79;
    rd_cycle[ 4230] = 1'b0;  wr_cycle[ 4230] = 1'b1;  addr_rom[ 4230]='h000010e4;  wr_data_rom[ 4230]='h0000143e;
    rd_cycle[ 4231] = 1'b0;  wr_cycle[ 4231] = 1'b1;  addr_rom[ 4231]='h000011bc;  wr_data_rom[ 4231]='h000002c0;
    rd_cycle[ 4232] = 1'b1;  wr_cycle[ 4232] = 1'b0;  addr_rom[ 4232]='h00000bac;  wr_data_rom[ 4232]='h00000000;
    rd_cycle[ 4233] = 1'b0;  wr_cycle[ 4233] = 1'b1;  addr_rom[ 4233]='h000004b8;  wr_data_rom[ 4233]='h0000070d;
    rd_cycle[ 4234] = 1'b1;  wr_cycle[ 4234] = 1'b0;  addr_rom[ 4234]='h000010c0;  wr_data_rom[ 4234]='h00000000;
    rd_cycle[ 4235] = 1'b0;  wr_cycle[ 4235] = 1'b1;  addr_rom[ 4235]='h00000f90;  wr_data_rom[ 4235]='h000011b8;
    rd_cycle[ 4236] = 1'b1;  wr_cycle[ 4236] = 1'b0;  addr_rom[ 4236]='h00000f84;  wr_data_rom[ 4236]='h00000000;
    rd_cycle[ 4237] = 1'b0;  wr_cycle[ 4237] = 1'b1;  addr_rom[ 4237]='h000001a8;  wr_data_rom[ 4237]='h0000039b;
    rd_cycle[ 4238] = 1'b0;  wr_cycle[ 4238] = 1'b1;  addr_rom[ 4238]='h00000494;  wr_data_rom[ 4238]='h0000075e;
    rd_cycle[ 4239] = 1'b0;  wr_cycle[ 4239] = 1'b1;  addr_rom[ 4239]='h00000ae8;  wr_data_rom[ 4239]='h000009b1;
    rd_cycle[ 4240] = 1'b0;  wr_cycle[ 4240] = 1'b1;  addr_rom[ 4240]='h00001edc;  wr_data_rom[ 4240]='h000003c2;
    rd_cycle[ 4241] = 1'b0;  wr_cycle[ 4241] = 1'b1;  addr_rom[ 4241]='h0000120c;  wr_data_rom[ 4241]='h00001167;
    rd_cycle[ 4242] = 1'b0;  wr_cycle[ 4242] = 1'b1;  addr_rom[ 4242]='h00000674;  wr_data_rom[ 4242]='h00000dae;
    rd_cycle[ 4243] = 1'b1;  wr_cycle[ 4243] = 1'b0;  addr_rom[ 4243]='h000008dc;  wr_data_rom[ 4243]='h00000000;
    rd_cycle[ 4244] = 1'b0;  wr_cycle[ 4244] = 1'b1;  addr_rom[ 4244]='h000000b4;  wr_data_rom[ 4244]='h00001e58;
    rd_cycle[ 4245] = 1'b0;  wr_cycle[ 4245] = 1'b1;  addr_rom[ 4245]='h000005ec;  wr_data_rom[ 4245]='h00000609;
    rd_cycle[ 4246] = 1'b1;  wr_cycle[ 4246] = 1'b0;  addr_rom[ 4246]='h00000a50;  wr_data_rom[ 4246]='h00000000;
    rd_cycle[ 4247] = 1'b1;  wr_cycle[ 4247] = 1'b0;  addr_rom[ 4247]='h00001914;  wr_data_rom[ 4247]='h00000000;
    rd_cycle[ 4248] = 1'b0;  wr_cycle[ 4248] = 1'b1;  addr_rom[ 4248]='h00000dd8;  wr_data_rom[ 4248]='h00001824;
    rd_cycle[ 4249] = 1'b0;  wr_cycle[ 4249] = 1'b1;  addr_rom[ 4249]='h000003ec;  wr_data_rom[ 4249]='h0000006c;
    rd_cycle[ 4250] = 1'b1;  wr_cycle[ 4250] = 1'b0;  addr_rom[ 4250]='h00000dec;  wr_data_rom[ 4250]='h00000000;
    rd_cycle[ 4251] = 1'b0;  wr_cycle[ 4251] = 1'b1;  addr_rom[ 4251]='h00001a54;  wr_data_rom[ 4251]='h000013c6;
    rd_cycle[ 4252] = 1'b1;  wr_cycle[ 4252] = 1'b0;  addr_rom[ 4252]='h00001424;  wr_data_rom[ 4252]='h00000000;
    rd_cycle[ 4253] = 1'b0;  wr_cycle[ 4253] = 1'b1;  addr_rom[ 4253]='h00000f90;  wr_data_rom[ 4253]='h00001d99;
    rd_cycle[ 4254] = 1'b1;  wr_cycle[ 4254] = 1'b0;  addr_rom[ 4254]='h00000124;  wr_data_rom[ 4254]='h00000000;
    rd_cycle[ 4255] = 1'b1;  wr_cycle[ 4255] = 1'b0;  addr_rom[ 4255]='h000009b8;  wr_data_rom[ 4255]='h00000000;
    rd_cycle[ 4256] = 1'b0;  wr_cycle[ 4256] = 1'b1;  addr_rom[ 4256]='h00000874;  wr_data_rom[ 4256]='h00001471;
    rd_cycle[ 4257] = 1'b0;  wr_cycle[ 4257] = 1'b1;  addr_rom[ 4257]='h000000fc;  wr_data_rom[ 4257]='h000005a1;
    rd_cycle[ 4258] = 1'b1;  wr_cycle[ 4258] = 1'b0;  addr_rom[ 4258]='h000007c0;  wr_data_rom[ 4258]='h00000000;
    rd_cycle[ 4259] = 1'b1;  wr_cycle[ 4259] = 1'b0;  addr_rom[ 4259]='h00001e40;  wr_data_rom[ 4259]='h00000000;
    rd_cycle[ 4260] = 1'b0;  wr_cycle[ 4260] = 1'b1;  addr_rom[ 4260]='h000010b4;  wr_data_rom[ 4260]='h00001ac6;
    rd_cycle[ 4261] = 1'b0;  wr_cycle[ 4261] = 1'b1;  addr_rom[ 4261]='h00000f5c;  wr_data_rom[ 4261]='h00000fa1;
    rd_cycle[ 4262] = 1'b0;  wr_cycle[ 4262] = 1'b1;  addr_rom[ 4262]='h00001718;  wr_data_rom[ 4262]='h00001b07;
    rd_cycle[ 4263] = 1'b1;  wr_cycle[ 4263] = 1'b0;  addr_rom[ 4263]='h000016e4;  wr_data_rom[ 4263]='h00000000;
    rd_cycle[ 4264] = 1'b1;  wr_cycle[ 4264] = 1'b0;  addr_rom[ 4264]='h00001c14;  wr_data_rom[ 4264]='h00000000;
    rd_cycle[ 4265] = 1'b0;  wr_cycle[ 4265] = 1'b1;  addr_rom[ 4265]='h0000079c;  wr_data_rom[ 4265]='h000015f3;
    rd_cycle[ 4266] = 1'b0;  wr_cycle[ 4266] = 1'b1;  addr_rom[ 4266]='h0000040c;  wr_data_rom[ 4266]='h0000170f;
    rd_cycle[ 4267] = 1'b1;  wr_cycle[ 4267] = 1'b0;  addr_rom[ 4267]='h00001aa0;  wr_data_rom[ 4267]='h00000000;
    rd_cycle[ 4268] = 1'b1;  wr_cycle[ 4268] = 1'b0;  addr_rom[ 4268]='h00000454;  wr_data_rom[ 4268]='h00000000;
    rd_cycle[ 4269] = 1'b1;  wr_cycle[ 4269] = 1'b0;  addr_rom[ 4269]='h00001ba0;  wr_data_rom[ 4269]='h00000000;
    rd_cycle[ 4270] = 1'b0;  wr_cycle[ 4270] = 1'b1;  addr_rom[ 4270]='h0000113c;  wr_data_rom[ 4270]='h0000104f;
    rd_cycle[ 4271] = 1'b1;  wr_cycle[ 4271] = 1'b0;  addr_rom[ 4271]='h0000129c;  wr_data_rom[ 4271]='h00000000;
    rd_cycle[ 4272] = 1'b0;  wr_cycle[ 4272] = 1'b1;  addr_rom[ 4272]='h00000ef0;  wr_data_rom[ 4272]='h00001f09;
    rd_cycle[ 4273] = 1'b1;  wr_cycle[ 4273] = 1'b0;  addr_rom[ 4273]='h0000141c;  wr_data_rom[ 4273]='h00000000;
    rd_cycle[ 4274] = 1'b0;  wr_cycle[ 4274] = 1'b1;  addr_rom[ 4274]='h00000328;  wr_data_rom[ 4274]='h00000320;
    rd_cycle[ 4275] = 1'b1;  wr_cycle[ 4275] = 1'b0;  addr_rom[ 4275]='h00000e98;  wr_data_rom[ 4275]='h00000000;
    rd_cycle[ 4276] = 1'b0;  wr_cycle[ 4276] = 1'b1;  addr_rom[ 4276]='h00001824;  wr_data_rom[ 4276]='h00001d81;
    rd_cycle[ 4277] = 1'b1;  wr_cycle[ 4277] = 1'b0;  addr_rom[ 4277]='h00001990;  wr_data_rom[ 4277]='h00000000;
    rd_cycle[ 4278] = 1'b1;  wr_cycle[ 4278] = 1'b0;  addr_rom[ 4278]='h00000fe0;  wr_data_rom[ 4278]='h00000000;
    rd_cycle[ 4279] = 1'b0;  wr_cycle[ 4279] = 1'b1;  addr_rom[ 4279]='h000001b8;  wr_data_rom[ 4279]='h00001040;
    rd_cycle[ 4280] = 1'b1;  wr_cycle[ 4280] = 1'b0;  addr_rom[ 4280]='h00000a70;  wr_data_rom[ 4280]='h00000000;
    rd_cycle[ 4281] = 1'b1;  wr_cycle[ 4281] = 1'b0;  addr_rom[ 4281]='h00001b98;  wr_data_rom[ 4281]='h00000000;
    rd_cycle[ 4282] = 1'b1;  wr_cycle[ 4282] = 1'b0;  addr_rom[ 4282]='h00000f84;  wr_data_rom[ 4282]='h00000000;
    rd_cycle[ 4283] = 1'b1;  wr_cycle[ 4283] = 1'b0;  addr_rom[ 4283]='h0000164c;  wr_data_rom[ 4283]='h00000000;
    rd_cycle[ 4284] = 1'b1;  wr_cycle[ 4284] = 1'b0;  addr_rom[ 4284]='h0000044c;  wr_data_rom[ 4284]='h00000000;
    rd_cycle[ 4285] = 1'b0;  wr_cycle[ 4285] = 1'b1;  addr_rom[ 4285]='h00001894;  wr_data_rom[ 4285]='h00000094;
    rd_cycle[ 4286] = 1'b1;  wr_cycle[ 4286] = 1'b0;  addr_rom[ 4286]='h00000dc4;  wr_data_rom[ 4286]='h00000000;
    rd_cycle[ 4287] = 1'b1;  wr_cycle[ 4287] = 1'b0;  addr_rom[ 4287]='h00000714;  wr_data_rom[ 4287]='h00000000;
    rd_cycle[ 4288] = 1'b0;  wr_cycle[ 4288] = 1'b1;  addr_rom[ 4288]='h00000fa4;  wr_data_rom[ 4288]='h000000c9;
    rd_cycle[ 4289] = 1'b0;  wr_cycle[ 4289] = 1'b1;  addr_rom[ 4289]='h00001f1c;  wr_data_rom[ 4289]='h00001384;
    rd_cycle[ 4290] = 1'b0;  wr_cycle[ 4290] = 1'b1;  addr_rom[ 4290]='h0000127c;  wr_data_rom[ 4290]='h00001f23;
    rd_cycle[ 4291] = 1'b0;  wr_cycle[ 4291] = 1'b1;  addr_rom[ 4291]='h0000002c;  wr_data_rom[ 4291]='h0000086f;
    rd_cycle[ 4292] = 1'b1;  wr_cycle[ 4292] = 1'b0;  addr_rom[ 4292]='h0000028c;  wr_data_rom[ 4292]='h00000000;
    rd_cycle[ 4293] = 1'b1;  wr_cycle[ 4293] = 1'b0;  addr_rom[ 4293]='h00001cd4;  wr_data_rom[ 4293]='h00000000;
    rd_cycle[ 4294] = 1'b0;  wr_cycle[ 4294] = 1'b1;  addr_rom[ 4294]='h000019b0;  wr_data_rom[ 4294]='h00001887;
    rd_cycle[ 4295] = 1'b1;  wr_cycle[ 4295] = 1'b0;  addr_rom[ 4295]='h000006c0;  wr_data_rom[ 4295]='h00000000;
    rd_cycle[ 4296] = 1'b1;  wr_cycle[ 4296] = 1'b0;  addr_rom[ 4296]='h00001d4c;  wr_data_rom[ 4296]='h00000000;
    rd_cycle[ 4297] = 1'b0;  wr_cycle[ 4297] = 1'b1;  addr_rom[ 4297]='h00000944;  wr_data_rom[ 4297]='h00000d1c;
    rd_cycle[ 4298] = 1'b0;  wr_cycle[ 4298] = 1'b1;  addr_rom[ 4298]='h00001b28;  wr_data_rom[ 4298]='h00001bcb;
    rd_cycle[ 4299] = 1'b1;  wr_cycle[ 4299] = 1'b0;  addr_rom[ 4299]='h00001b98;  wr_data_rom[ 4299]='h00000000;
    rd_cycle[ 4300] = 1'b1;  wr_cycle[ 4300] = 1'b0;  addr_rom[ 4300]='h00000314;  wr_data_rom[ 4300]='h00000000;
    rd_cycle[ 4301] = 1'b0;  wr_cycle[ 4301] = 1'b1;  addr_rom[ 4301]='h00001a58;  wr_data_rom[ 4301]='h000000c6;
    rd_cycle[ 4302] = 1'b1;  wr_cycle[ 4302] = 1'b0;  addr_rom[ 4302]='h00000d7c;  wr_data_rom[ 4302]='h00000000;
    rd_cycle[ 4303] = 1'b1;  wr_cycle[ 4303] = 1'b0;  addr_rom[ 4303]='h00000dd4;  wr_data_rom[ 4303]='h00000000;
    rd_cycle[ 4304] = 1'b1;  wr_cycle[ 4304] = 1'b0;  addr_rom[ 4304]='h00001ce0;  wr_data_rom[ 4304]='h00000000;
    rd_cycle[ 4305] = 1'b1;  wr_cycle[ 4305] = 1'b0;  addr_rom[ 4305]='h00000d60;  wr_data_rom[ 4305]='h00000000;
    rd_cycle[ 4306] = 1'b1;  wr_cycle[ 4306] = 1'b0;  addr_rom[ 4306]='h000008fc;  wr_data_rom[ 4306]='h00000000;
    rd_cycle[ 4307] = 1'b0;  wr_cycle[ 4307] = 1'b1;  addr_rom[ 4307]='h000005e8;  wr_data_rom[ 4307]='h00000343;
    rd_cycle[ 4308] = 1'b0;  wr_cycle[ 4308] = 1'b1;  addr_rom[ 4308]='h00000f64;  wr_data_rom[ 4308]='h00000815;
    rd_cycle[ 4309] = 1'b0;  wr_cycle[ 4309] = 1'b1;  addr_rom[ 4309]='h00000d0c;  wr_data_rom[ 4309]='h00000197;
    rd_cycle[ 4310] = 1'b1;  wr_cycle[ 4310] = 1'b0;  addr_rom[ 4310]='h00001998;  wr_data_rom[ 4310]='h00000000;
    rd_cycle[ 4311] = 1'b0;  wr_cycle[ 4311] = 1'b1;  addr_rom[ 4311]='h00000cfc;  wr_data_rom[ 4311]='h00001770;
    rd_cycle[ 4312] = 1'b1;  wr_cycle[ 4312] = 1'b0;  addr_rom[ 4312]='h00001014;  wr_data_rom[ 4312]='h00000000;
    rd_cycle[ 4313] = 1'b1;  wr_cycle[ 4313] = 1'b0;  addr_rom[ 4313]='h00000f04;  wr_data_rom[ 4313]='h00000000;
    rd_cycle[ 4314] = 1'b0;  wr_cycle[ 4314] = 1'b1;  addr_rom[ 4314]='h00001290;  wr_data_rom[ 4314]='h00001c70;
    rd_cycle[ 4315] = 1'b0;  wr_cycle[ 4315] = 1'b1;  addr_rom[ 4315]='h000006f4;  wr_data_rom[ 4315]='h0000051c;
    rd_cycle[ 4316] = 1'b1;  wr_cycle[ 4316] = 1'b0;  addr_rom[ 4316]='h00000488;  wr_data_rom[ 4316]='h00000000;
    rd_cycle[ 4317] = 1'b1;  wr_cycle[ 4317] = 1'b0;  addr_rom[ 4317]='h0000165c;  wr_data_rom[ 4317]='h00000000;
    rd_cycle[ 4318] = 1'b1;  wr_cycle[ 4318] = 1'b0;  addr_rom[ 4318]='h00001070;  wr_data_rom[ 4318]='h00000000;
    rd_cycle[ 4319] = 1'b1;  wr_cycle[ 4319] = 1'b0;  addr_rom[ 4319]='h00000e74;  wr_data_rom[ 4319]='h00000000;
    rd_cycle[ 4320] = 1'b1;  wr_cycle[ 4320] = 1'b0;  addr_rom[ 4320]='h0000025c;  wr_data_rom[ 4320]='h00000000;
    rd_cycle[ 4321] = 1'b0;  wr_cycle[ 4321] = 1'b1;  addr_rom[ 4321]='h00000dd4;  wr_data_rom[ 4321]='h000016e8;
    rd_cycle[ 4322] = 1'b1;  wr_cycle[ 4322] = 1'b0;  addr_rom[ 4322]='h0000086c;  wr_data_rom[ 4322]='h00000000;
    rd_cycle[ 4323] = 1'b1;  wr_cycle[ 4323] = 1'b0;  addr_rom[ 4323]='h000010e0;  wr_data_rom[ 4323]='h00000000;
    rd_cycle[ 4324] = 1'b1;  wr_cycle[ 4324] = 1'b0;  addr_rom[ 4324]='h000016e0;  wr_data_rom[ 4324]='h00000000;
    rd_cycle[ 4325] = 1'b1;  wr_cycle[ 4325] = 1'b0;  addr_rom[ 4325]='h00000980;  wr_data_rom[ 4325]='h00000000;
    rd_cycle[ 4326] = 1'b1;  wr_cycle[ 4326] = 1'b0;  addr_rom[ 4326]='h00000f5c;  wr_data_rom[ 4326]='h00000000;
    rd_cycle[ 4327] = 1'b1;  wr_cycle[ 4327] = 1'b0;  addr_rom[ 4327]='h00000f54;  wr_data_rom[ 4327]='h00000000;
    rd_cycle[ 4328] = 1'b0;  wr_cycle[ 4328] = 1'b1;  addr_rom[ 4328]='h00001268;  wr_data_rom[ 4328]='h000015fb;
    rd_cycle[ 4329] = 1'b0;  wr_cycle[ 4329] = 1'b1;  addr_rom[ 4329]='h00000f98;  wr_data_rom[ 4329]='h0000104b;
    rd_cycle[ 4330] = 1'b1;  wr_cycle[ 4330] = 1'b0;  addr_rom[ 4330]='h00000d0c;  wr_data_rom[ 4330]='h00000000;
    rd_cycle[ 4331] = 1'b0;  wr_cycle[ 4331] = 1'b1;  addr_rom[ 4331]='h00001590;  wr_data_rom[ 4331]='h00001b9d;
    rd_cycle[ 4332] = 1'b0;  wr_cycle[ 4332] = 1'b1;  addr_rom[ 4332]='h000002c8;  wr_data_rom[ 4332]='h00000902;
    rd_cycle[ 4333] = 1'b0;  wr_cycle[ 4333] = 1'b1;  addr_rom[ 4333]='h00001d00;  wr_data_rom[ 4333]='h00001a32;
    rd_cycle[ 4334] = 1'b1;  wr_cycle[ 4334] = 1'b0;  addr_rom[ 4334]='h00001d3c;  wr_data_rom[ 4334]='h00000000;
    rd_cycle[ 4335] = 1'b1;  wr_cycle[ 4335] = 1'b0;  addr_rom[ 4335]='h00000a20;  wr_data_rom[ 4335]='h00000000;
    rd_cycle[ 4336] = 1'b1;  wr_cycle[ 4336] = 1'b0;  addr_rom[ 4336]='h00001008;  wr_data_rom[ 4336]='h00000000;
    rd_cycle[ 4337] = 1'b1;  wr_cycle[ 4337] = 1'b0;  addr_rom[ 4337]='h00000a70;  wr_data_rom[ 4337]='h00000000;
    rd_cycle[ 4338] = 1'b1;  wr_cycle[ 4338] = 1'b0;  addr_rom[ 4338]='h000011ec;  wr_data_rom[ 4338]='h00000000;
    rd_cycle[ 4339] = 1'b0;  wr_cycle[ 4339] = 1'b1;  addr_rom[ 4339]='h00000248;  wr_data_rom[ 4339]='h000019e8;
    rd_cycle[ 4340] = 1'b1;  wr_cycle[ 4340] = 1'b0;  addr_rom[ 4340]='h000000fc;  wr_data_rom[ 4340]='h00000000;
    rd_cycle[ 4341] = 1'b1;  wr_cycle[ 4341] = 1'b0;  addr_rom[ 4341]='h000007e4;  wr_data_rom[ 4341]='h00000000;
    rd_cycle[ 4342] = 1'b1;  wr_cycle[ 4342] = 1'b0;  addr_rom[ 4342]='h0000173c;  wr_data_rom[ 4342]='h00000000;
    rd_cycle[ 4343] = 1'b1;  wr_cycle[ 4343] = 1'b0;  addr_rom[ 4343]='h0000125c;  wr_data_rom[ 4343]='h00000000;
    rd_cycle[ 4344] = 1'b0;  wr_cycle[ 4344] = 1'b1;  addr_rom[ 4344]='h00000230;  wr_data_rom[ 4344]='h00000579;
    rd_cycle[ 4345] = 1'b0;  wr_cycle[ 4345] = 1'b1;  addr_rom[ 4345]='h00001c44;  wr_data_rom[ 4345]='h00000da1;
    rd_cycle[ 4346] = 1'b0;  wr_cycle[ 4346] = 1'b1;  addr_rom[ 4346]='h00000cb4;  wr_data_rom[ 4346]='h000016b5;
    rd_cycle[ 4347] = 1'b0;  wr_cycle[ 4347] = 1'b1;  addr_rom[ 4347]='h000003b4;  wr_data_rom[ 4347]='h00001a2d;
    rd_cycle[ 4348] = 1'b1;  wr_cycle[ 4348] = 1'b0;  addr_rom[ 4348]='h000002c0;  wr_data_rom[ 4348]='h00000000;
    rd_cycle[ 4349] = 1'b1;  wr_cycle[ 4349] = 1'b0;  addr_rom[ 4349]='h000008f8;  wr_data_rom[ 4349]='h00000000;
    rd_cycle[ 4350] = 1'b0;  wr_cycle[ 4350] = 1'b1;  addr_rom[ 4350]='h000017b0;  wr_data_rom[ 4350]='h000001ed;
    rd_cycle[ 4351] = 1'b0;  wr_cycle[ 4351] = 1'b1;  addr_rom[ 4351]='h00001834;  wr_data_rom[ 4351]='h0000108d;
    rd_cycle[ 4352] = 1'b0;  wr_cycle[ 4352] = 1'b1;  addr_rom[ 4352]='h00000094;  wr_data_rom[ 4352]='h00000ae5;
    rd_cycle[ 4353] = 1'b0;  wr_cycle[ 4353] = 1'b1;  addr_rom[ 4353]='h00001b70;  wr_data_rom[ 4353]='h000011d7;
    rd_cycle[ 4354] = 1'b0;  wr_cycle[ 4354] = 1'b1;  addr_rom[ 4354]='h00001b08;  wr_data_rom[ 4354]='h000001e7;
    rd_cycle[ 4355] = 1'b1;  wr_cycle[ 4355] = 1'b0;  addr_rom[ 4355]='h00000c5c;  wr_data_rom[ 4355]='h00000000;
    rd_cycle[ 4356] = 1'b1;  wr_cycle[ 4356] = 1'b0;  addr_rom[ 4356]='h00001158;  wr_data_rom[ 4356]='h00000000;
    rd_cycle[ 4357] = 1'b0;  wr_cycle[ 4357] = 1'b1;  addr_rom[ 4357]='h000000e0;  wr_data_rom[ 4357]='h00001bbe;
    rd_cycle[ 4358] = 1'b0;  wr_cycle[ 4358] = 1'b1;  addr_rom[ 4358]='h00000654;  wr_data_rom[ 4358]='h00000865;
    rd_cycle[ 4359] = 1'b0;  wr_cycle[ 4359] = 1'b1;  addr_rom[ 4359]='h00001f1c;  wr_data_rom[ 4359]='h0000067b;
    rd_cycle[ 4360] = 1'b1;  wr_cycle[ 4360] = 1'b0;  addr_rom[ 4360]='h00001564;  wr_data_rom[ 4360]='h00000000;
    rd_cycle[ 4361] = 1'b0;  wr_cycle[ 4361] = 1'b1;  addr_rom[ 4361]='h00001ad4;  wr_data_rom[ 4361]='h00000b72;
    rd_cycle[ 4362] = 1'b1;  wr_cycle[ 4362] = 1'b0;  addr_rom[ 4362]='h00000ba4;  wr_data_rom[ 4362]='h00000000;
    rd_cycle[ 4363] = 1'b1;  wr_cycle[ 4363] = 1'b0;  addr_rom[ 4363]='h00001dd0;  wr_data_rom[ 4363]='h00000000;
    rd_cycle[ 4364] = 1'b1;  wr_cycle[ 4364] = 1'b0;  addr_rom[ 4364]='h00001f20;  wr_data_rom[ 4364]='h00000000;
    rd_cycle[ 4365] = 1'b1;  wr_cycle[ 4365] = 1'b0;  addr_rom[ 4365]='h00000cac;  wr_data_rom[ 4365]='h00000000;
    rd_cycle[ 4366] = 1'b0;  wr_cycle[ 4366] = 1'b1;  addr_rom[ 4366]='h00001690;  wr_data_rom[ 4366]='h00000013;
    rd_cycle[ 4367] = 1'b1;  wr_cycle[ 4367] = 1'b0;  addr_rom[ 4367]='h00001dcc;  wr_data_rom[ 4367]='h00000000;
    rd_cycle[ 4368] = 1'b0;  wr_cycle[ 4368] = 1'b1;  addr_rom[ 4368]='h0000118c;  wr_data_rom[ 4368]='h00000e2a;
    rd_cycle[ 4369] = 1'b1;  wr_cycle[ 4369] = 1'b0;  addr_rom[ 4369]='h00001a70;  wr_data_rom[ 4369]='h00000000;
    rd_cycle[ 4370] = 1'b0;  wr_cycle[ 4370] = 1'b1;  addr_rom[ 4370]='h00000068;  wr_data_rom[ 4370]='h00000665;
    rd_cycle[ 4371] = 1'b0;  wr_cycle[ 4371] = 1'b1;  addr_rom[ 4371]='h00000218;  wr_data_rom[ 4371]='h00000de0;
    rd_cycle[ 4372] = 1'b1;  wr_cycle[ 4372] = 1'b0;  addr_rom[ 4372]='h000016e0;  wr_data_rom[ 4372]='h00000000;
    rd_cycle[ 4373] = 1'b0;  wr_cycle[ 4373] = 1'b1;  addr_rom[ 4373]='h0000083c;  wr_data_rom[ 4373]='h00000661;
    rd_cycle[ 4374] = 1'b0;  wr_cycle[ 4374] = 1'b1;  addr_rom[ 4374]='h0000093c;  wr_data_rom[ 4374]='h0000190f;
    rd_cycle[ 4375] = 1'b1;  wr_cycle[ 4375] = 1'b0;  addr_rom[ 4375]='h00001534;  wr_data_rom[ 4375]='h00000000;
    rd_cycle[ 4376] = 1'b0;  wr_cycle[ 4376] = 1'b1;  addr_rom[ 4376]='h00000e68;  wr_data_rom[ 4376]='h00001013;
    rd_cycle[ 4377] = 1'b0;  wr_cycle[ 4377] = 1'b1;  addr_rom[ 4377]='h000019e8;  wr_data_rom[ 4377]='h0000003f;
    rd_cycle[ 4378] = 1'b1;  wr_cycle[ 4378] = 1'b0;  addr_rom[ 4378]='h00001aac;  wr_data_rom[ 4378]='h00000000;
    rd_cycle[ 4379] = 1'b1;  wr_cycle[ 4379] = 1'b0;  addr_rom[ 4379]='h000000e0;  wr_data_rom[ 4379]='h00000000;
    rd_cycle[ 4380] = 1'b0;  wr_cycle[ 4380] = 1'b1;  addr_rom[ 4380]='h000002d8;  wr_data_rom[ 4380]='h0000022e;
    rd_cycle[ 4381] = 1'b1;  wr_cycle[ 4381] = 1'b0;  addr_rom[ 4381]='h00000608;  wr_data_rom[ 4381]='h00000000;
    rd_cycle[ 4382] = 1'b0;  wr_cycle[ 4382] = 1'b1;  addr_rom[ 4382]='h00001480;  wr_data_rom[ 4382]='h0000158f;
    rd_cycle[ 4383] = 1'b0;  wr_cycle[ 4383] = 1'b1;  addr_rom[ 4383]='h00001974;  wr_data_rom[ 4383]='h000016d1;
    rd_cycle[ 4384] = 1'b1;  wr_cycle[ 4384] = 1'b0;  addr_rom[ 4384]='h00001c20;  wr_data_rom[ 4384]='h00000000;
    rd_cycle[ 4385] = 1'b0;  wr_cycle[ 4385] = 1'b1;  addr_rom[ 4385]='h00000d04;  wr_data_rom[ 4385]='h00000d52;
    rd_cycle[ 4386] = 1'b1;  wr_cycle[ 4386] = 1'b0;  addr_rom[ 4386]='h00001e60;  wr_data_rom[ 4386]='h00000000;
    rd_cycle[ 4387] = 1'b1;  wr_cycle[ 4387] = 1'b0;  addr_rom[ 4387]='h00000354;  wr_data_rom[ 4387]='h00000000;
    rd_cycle[ 4388] = 1'b1;  wr_cycle[ 4388] = 1'b0;  addr_rom[ 4388]='h00001d30;  wr_data_rom[ 4388]='h00000000;
    rd_cycle[ 4389] = 1'b1;  wr_cycle[ 4389] = 1'b0;  addr_rom[ 4389]='h0000041c;  wr_data_rom[ 4389]='h00000000;
    rd_cycle[ 4390] = 1'b1;  wr_cycle[ 4390] = 1'b0;  addr_rom[ 4390]='h000004a0;  wr_data_rom[ 4390]='h00000000;
    rd_cycle[ 4391] = 1'b0;  wr_cycle[ 4391] = 1'b1;  addr_rom[ 4391]='h00001e88;  wr_data_rom[ 4391]='h00000928;
    rd_cycle[ 4392] = 1'b1;  wr_cycle[ 4392] = 1'b0;  addr_rom[ 4392]='h00001988;  wr_data_rom[ 4392]='h00000000;
    rd_cycle[ 4393] = 1'b0;  wr_cycle[ 4393] = 1'b1;  addr_rom[ 4393]='h00000284;  wr_data_rom[ 4393]='h00000ed2;
    rd_cycle[ 4394] = 1'b0;  wr_cycle[ 4394] = 1'b1;  addr_rom[ 4394]='h00000b7c;  wr_data_rom[ 4394]='h00000d34;
    rd_cycle[ 4395] = 1'b0;  wr_cycle[ 4395] = 1'b1;  addr_rom[ 4395]='h00000004;  wr_data_rom[ 4395]='h00000cf0;
    rd_cycle[ 4396] = 1'b0;  wr_cycle[ 4396] = 1'b1;  addr_rom[ 4396]='h00000270;  wr_data_rom[ 4396]='h00001629;
    rd_cycle[ 4397] = 1'b1;  wr_cycle[ 4397] = 1'b0;  addr_rom[ 4397]='h00001938;  wr_data_rom[ 4397]='h00000000;
    rd_cycle[ 4398] = 1'b1;  wr_cycle[ 4398] = 1'b0;  addr_rom[ 4398]='h00001604;  wr_data_rom[ 4398]='h00000000;
    rd_cycle[ 4399] = 1'b1;  wr_cycle[ 4399] = 1'b0;  addr_rom[ 4399]='h00000738;  wr_data_rom[ 4399]='h00000000;
    rd_cycle[ 4400] = 1'b0;  wr_cycle[ 4400] = 1'b1;  addr_rom[ 4400]='h00000b58;  wr_data_rom[ 4400]='h00000b45;
    rd_cycle[ 4401] = 1'b1;  wr_cycle[ 4401] = 1'b0;  addr_rom[ 4401]='h00000f18;  wr_data_rom[ 4401]='h00000000;
    rd_cycle[ 4402] = 1'b1;  wr_cycle[ 4402] = 1'b0;  addr_rom[ 4402]='h00001718;  wr_data_rom[ 4402]='h00000000;
    rd_cycle[ 4403] = 1'b0;  wr_cycle[ 4403] = 1'b1;  addr_rom[ 4403]='h00001e44;  wr_data_rom[ 4403]='h0000047e;
    rd_cycle[ 4404] = 1'b1;  wr_cycle[ 4404] = 1'b0;  addr_rom[ 4404]='h00001b00;  wr_data_rom[ 4404]='h00000000;
    rd_cycle[ 4405] = 1'b1;  wr_cycle[ 4405] = 1'b0;  addr_rom[ 4405]='h00001c14;  wr_data_rom[ 4405]='h00000000;
    rd_cycle[ 4406] = 1'b0;  wr_cycle[ 4406] = 1'b1;  addr_rom[ 4406]='h0000030c;  wr_data_rom[ 4406]='h00001079;
    rd_cycle[ 4407] = 1'b0;  wr_cycle[ 4407] = 1'b1;  addr_rom[ 4407]='h000015f8;  wr_data_rom[ 4407]='h000006fe;
    rd_cycle[ 4408] = 1'b0;  wr_cycle[ 4408] = 1'b1;  addr_rom[ 4408]='h00000658;  wr_data_rom[ 4408]='h00001d2a;
    rd_cycle[ 4409] = 1'b0;  wr_cycle[ 4409] = 1'b1;  addr_rom[ 4409]='h00001500;  wr_data_rom[ 4409]='h00001ca7;
    rd_cycle[ 4410] = 1'b0;  wr_cycle[ 4410] = 1'b1;  addr_rom[ 4410]='h00000768;  wr_data_rom[ 4410]='h00000c5b;
    rd_cycle[ 4411] = 1'b1;  wr_cycle[ 4411] = 1'b0;  addr_rom[ 4411]='h00001368;  wr_data_rom[ 4411]='h00000000;
    rd_cycle[ 4412] = 1'b0;  wr_cycle[ 4412] = 1'b1;  addr_rom[ 4412]='h00000ad8;  wr_data_rom[ 4412]='h00000c4f;
    rd_cycle[ 4413] = 1'b1;  wr_cycle[ 4413] = 1'b0;  addr_rom[ 4413]='h0000017c;  wr_data_rom[ 4413]='h00000000;
    rd_cycle[ 4414] = 1'b0;  wr_cycle[ 4414] = 1'b1;  addr_rom[ 4414]='h0000077c;  wr_data_rom[ 4414]='h00001a48;
    rd_cycle[ 4415] = 1'b1;  wr_cycle[ 4415] = 1'b0;  addr_rom[ 4415]='h00001a98;  wr_data_rom[ 4415]='h00000000;
    rd_cycle[ 4416] = 1'b0;  wr_cycle[ 4416] = 1'b1;  addr_rom[ 4416]='h00000c18;  wr_data_rom[ 4416]='h000001d2;
    rd_cycle[ 4417] = 1'b1;  wr_cycle[ 4417] = 1'b0;  addr_rom[ 4417]='h00000628;  wr_data_rom[ 4417]='h00000000;
    rd_cycle[ 4418] = 1'b0;  wr_cycle[ 4418] = 1'b1;  addr_rom[ 4418]='h00001038;  wr_data_rom[ 4418]='h00001462;
    rd_cycle[ 4419] = 1'b1;  wr_cycle[ 4419] = 1'b0;  addr_rom[ 4419]='h000016d0;  wr_data_rom[ 4419]='h00000000;
    rd_cycle[ 4420] = 1'b1;  wr_cycle[ 4420] = 1'b0;  addr_rom[ 4420]='h00000034;  wr_data_rom[ 4420]='h00000000;
    rd_cycle[ 4421] = 1'b0;  wr_cycle[ 4421] = 1'b1;  addr_rom[ 4421]='h00000c58;  wr_data_rom[ 4421]='h00000c83;
    rd_cycle[ 4422] = 1'b1;  wr_cycle[ 4422] = 1'b0;  addr_rom[ 4422]='h000007fc;  wr_data_rom[ 4422]='h00000000;
    rd_cycle[ 4423] = 1'b0;  wr_cycle[ 4423] = 1'b1;  addr_rom[ 4423]='h00000cf4;  wr_data_rom[ 4423]='h000018c2;
    rd_cycle[ 4424] = 1'b1;  wr_cycle[ 4424] = 1'b0;  addr_rom[ 4424]='h000007b0;  wr_data_rom[ 4424]='h00000000;
    rd_cycle[ 4425] = 1'b1;  wr_cycle[ 4425] = 1'b0;  addr_rom[ 4425]='h00000efc;  wr_data_rom[ 4425]='h00000000;
    rd_cycle[ 4426] = 1'b1;  wr_cycle[ 4426] = 1'b0;  addr_rom[ 4426]='h00000604;  wr_data_rom[ 4426]='h00000000;
    rd_cycle[ 4427] = 1'b0;  wr_cycle[ 4427] = 1'b1;  addr_rom[ 4427]='h00000ea0;  wr_data_rom[ 4427]='h00000946;
    rd_cycle[ 4428] = 1'b1;  wr_cycle[ 4428] = 1'b0;  addr_rom[ 4428]='h00000d9c;  wr_data_rom[ 4428]='h00000000;
    rd_cycle[ 4429] = 1'b1;  wr_cycle[ 4429] = 1'b0;  addr_rom[ 4429]='h000018f0;  wr_data_rom[ 4429]='h00000000;
    rd_cycle[ 4430] = 1'b0;  wr_cycle[ 4430] = 1'b1;  addr_rom[ 4430]='h00000de4;  wr_data_rom[ 4430]='h00001a9a;
    rd_cycle[ 4431] = 1'b1;  wr_cycle[ 4431] = 1'b0;  addr_rom[ 4431]='h00000c5c;  wr_data_rom[ 4431]='h00000000;
    rd_cycle[ 4432] = 1'b1;  wr_cycle[ 4432] = 1'b0;  addr_rom[ 4432]='h0000006c;  wr_data_rom[ 4432]='h00000000;
    rd_cycle[ 4433] = 1'b0;  wr_cycle[ 4433] = 1'b1;  addr_rom[ 4433]='h000010f4;  wr_data_rom[ 4433]='h00001216;
    rd_cycle[ 4434] = 1'b1;  wr_cycle[ 4434] = 1'b0;  addr_rom[ 4434]='h00000370;  wr_data_rom[ 4434]='h00000000;
    rd_cycle[ 4435] = 1'b0;  wr_cycle[ 4435] = 1'b1;  addr_rom[ 4435]='h00000c68;  wr_data_rom[ 4435]='h000007bd;
    rd_cycle[ 4436] = 1'b0;  wr_cycle[ 4436] = 1'b1;  addr_rom[ 4436]='h00001a14;  wr_data_rom[ 4436]='h0000038a;
    rd_cycle[ 4437] = 1'b0;  wr_cycle[ 4437] = 1'b1;  addr_rom[ 4437]='h0000047c;  wr_data_rom[ 4437]='h00001658;
    rd_cycle[ 4438] = 1'b0;  wr_cycle[ 4438] = 1'b1;  addr_rom[ 4438]='h00001e94;  wr_data_rom[ 4438]='h0000155c;
    rd_cycle[ 4439] = 1'b0;  wr_cycle[ 4439] = 1'b1;  addr_rom[ 4439]='h000016d4;  wr_data_rom[ 4439]='h00001b62;
    rd_cycle[ 4440] = 1'b0;  wr_cycle[ 4440] = 1'b1;  addr_rom[ 4440]='h000003ac;  wr_data_rom[ 4440]='h00001200;
    rd_cycle[ 4441] = 1'b1;  wr_cycle[ 4441] = 1'b0;  addr_rom[ 4441]='h00000070;  wr_data_rom[ 4441]='h00000000;
    rd_cycle[ 4442] = 1'b1;  wr_cycle[ 4442] = 1'b0;  addr_rom[ 4442]='h00000b7c;  wr_data_rom[ 4442]='h00000000;
    rd_cycle[ 4443] = 1'b0;  wr_cycle[ 4443] = 1'b1;  addr_rom[ 4443]='h00000b94;  wr_data_rom[ 4443]='h0000163c;
    rd_cycle[ 4444] = 1'b0;  wr_cycle[ 4444] = 1'b1;  addr_rom[ 4444]='h00000238;  wr_data_rom[ 4444]='h0000134c;
    rd_cycle[ 4445] = 1'b0;  wr_cycle[ 4445] = 1'b1;  addr_rom[ 4445]='h00001b90;  wr_data_rom[ 4445]='h00001dd5;
    rd_cycle[ 4446] = 1'b0;  wr_cycle[ 4446] = 1'b1;  addr_rom[ 4446]='h00000af4;  wr_data_rom[ 4446]='h00000f66;
    rd_cycle[ 4447] = 1'b1;  wr_cycle[ 4447] = 1'b0;  addr_rom[ 4447]='h00000508;  wr_data_rom[ 4447]='h00000000;
    rd_cycle[ 4448] = 1'b0;  wr_cycle[ 4448] = 1'b1;  addr_rom[ 4448]='h000018bc;  wr_data_rom[ 4448]='h00000a95;
    rd_cycle[ 4449] = 1'b1;  wr_cycle[ 4449] = 1'b0;  addr_rom[ 4449]='h00000a30;  wr_data_rom[ 4449]='h00000000;
    rd_cycle[ 4450] = 1'b0;  wr_cycle[ 4450] = 1'b1;  addr_rom[ 4450]='h00000b80;  wr_data_rom[ 4450]='h00001dde;
    rd_cycle[ 4451] = 1'b0;  wr_cycle[ 4451] = 1'b1;  addr_rom[ 4451]='h00000490;  wr_data_rom[ 4451]='h00000967;
    rd_cycle[ 4452] = 1'b1;  wr_cycle[ 4452] = 1'b0;  addr_rom[ 4452]='h00001f08;  wr_data_rom[ 4452]='h00000000;
    rd_cycle[ 4453] = 1'b1;  wr_cycle[ 4453] = 1'b0;  addr_rom[ 4453]='h00001000;  wr_data_rom[ 4453]='h00000000;
    rd_cycle[ 4454] = 1'b0;  wr_cycle[ 4454] = 1'b1;  addr_rom[ 4454]='h00000040;  wr_data_rom[ 4454]='h00000c17;
    rd_cycle[ 4455] = 1'b1;  wr_cycle[ 4455] = 1'b0;  addr_rom[ 4455]='h00001274;  wr_data_rom[ 4455]='h00000000;
    rd_cycle[ 4456] = 1'b1;  wr_cycle[ 4456] = 1'b0;  addr_rom[ 4456]='h00000be8;  wr_data_rom[ 4456]='h00000000;
    rd_cycle[ 4457] = 1'b0;  wr_cycle[ 4457] = 1'b1;  addr_rom[ 4457]='h00001170;  wr_data_rom[ 4457]='h000014f0;
    rd_cycle[ 4458] = 1'b1;  wr_cycle[ 4458] = 1'b0;  addr_rom[ 4458]='h00000420;  wr_data_rom[ 4458]='h00000000;
    rd_cycle[ 4459] = 1'b0;  wr_cycle[ 4459] = 1'b1;  addr_rom[ 4459]='h00001330;  wr_data_rom[ 4459]='h000018f8;
    rd_cycle[ 4460] = 1'b0;  wr_cycle[ 4460] = 1'b1;  addr_rom[ 4460]='h00001410;  wr_data_rom[ 4460]='h00000484;
    rd_cycle[ 4461] = 1'b1;  wr_cycle[ 4461] = 1'b0;  addr_rom[ 4461]='h00001980;  wr_data_rom[ 4461]='h00000000;
    rd_cycle[ 4462] = 1'b0;  wr_cycle[ 4462] = 1'b1;  addr_rom[ 4462]='h0000164c;  wr_data_rom[ 4462]='h00001760;
    rd_cycle[ 4463] = 1'b0;  wr_cycle[ 4463] = 1'b1;  addr_rom[ 4463]='h00000088;  wr_data_rom[ 4463]='h00000c2a;
    rd_cycle[ 4464] = 1'b1;  wr_cycle[ 4464] = 1'b0;  addr_rom[ 4464]='h00001d04;  wr_data_rom[ 4464]='h00000000;
    rd_cycle[ 4465] = 1'b0;  wr_cycle[ 4465] = 1'b1;  addr_rom[ 4465]='h00001108;  wr_data_rom[ 4465]='h000001dd;
    rd_cycle[ 4466] = 1'b0;  wr_cycle[ 4466] = 1'b1;  addr_rom[ 4466]='h00000c18;  wr_data_rom[ 4466]='h000001d0;
    rd_cycle[ 4467] = 1'b1;  wr_cycle[ 4467] = 1'b0;  addr_rom[ 4467]='h00000e84;  wr_data_rom[ 4467]='h00000000;
    rd_cycle[ 4468] = 1'b1;  wr_cycle[ 4468] = 1'b0;  addr_rom[ 4468]='h000019b8;  wr_data_rom[ 4468]='h00000000;
    rd_cycle[ 4469] = 1'b1;  wr_cycle[ 4469] = 1'b0;  addr_rom[ 4469]='h00000170;  wr_data_rom[ 4469]='h00000000;
    rd_cycle[ 4470] = 1'b1;  wr_cycle[ 4470] = 1'b0;  addr_rom[ 4470]='h0000064c;  wr_data_rom[ 4470]='h00000000;
    rd_cycle[ 4471] = 1'b0;  wr_cycle[ 4471] = 1'b1;  addr_rom[ 4471]='h00001268;  wr_data_rom[ 4471]='h000004c8;
    rd_cycle[ 4472] = 1'b0;  wr_cycle[ 4472] = 1'b1;  addr_rom[ 4472]='h00000654;  wr_data_rom[ 4472]='h000007af;
    rd_cycle[ 4473] = 1'b0;  wr_cycle[ 4473] = 1'b1;  addr_rom[ 4473]='h000010d4;  wr_data_rom[ 4473]='h00000f74;
    rd_cycle[ 4474] = 1'b0;  wr_cycle[ 4474] = 1'b1;  addr_rom[ 4474]='h000017a4;  wr_data_rom[ 4474]='h00001355;
    rd_cycle[ 4475] = 1'b0;  wr_cycle[ 4475] = 1'b1;  addr_rom[ 4475]='h000004c4;  wr_data_rom[ 4475]='h00000584;
    rd_cycle[ 4476] = 1'b1;  wr_cycle[ 4476] = 1'b0;  addr_rom[ 4476]='h00001ed0;  wr_data_rom[ 4476]='h00000000;
    rd_cycle[ 4477] = 1'b1;  wr_cycle[ 4477] = 1'b0;  addr_rom[ 4477]='h0000082c;  wr_data_rom[ 4477]='h00000000;
    rd_cycle[ 4478] = 1'b0;  wr_cycle[ 4478] = 1'b1;  addr_rom[ 4478]='h00000890;  wr_data_rom[ 4478]='h00001877;
    rd_cycle[ 4479] = 1'b0;  wr_cycle[ 4479] = 1'b1;  addr_rom[ 4479]='h00000340;  wr_data_rom[ 4479]='h00000bc8;
    rd_cycle[ 4480] = 1'b1;  wr_cycle[ 4480] = 1'b0;  addr_rom[ 4480]='h000017ec;  wr_data_rom[ 4480]='h00000000;
    rd_cycle[ 4481] = 1'b0;  wr_cycle[ 4481] = 1'b1;  addr_rom[ 4481]='h00001544;  wr_data_rom[ 4481]='h00001cba;
    rd_cycle[ 4482] = 1'b0;  wr_cycle[ 4482] = 1'b1;  addr_rom[ 4482]='h000009a4;  wr_data_rom[ 4482]='h00000e22;
    rd_cycle[ 4483] = 1'b1;  wr_cycle[ 4483] = 1'b0;  addr_rom[ 4483]='h00001ab8;  wr_data_rom[ 4483]='h00000000;
    rd_cycle[ 4484] = 1'b0;  wr_cycle[ 4484] = 1'b1;  addr_rom[ 4484]='h00001f24;  wr_data_rom[ 4484]='h00000160;
    rd_cycle[ 4485] = 1'b1;  wr_cycle[ 4485] = 1'b0;  addr_rom[ 4485]='h00000574;  wr_data_rom[ 4485]='h00000000;
    rd_cycle[ 4486] = 1'b1;  wr_cycle[ 4486] = 1'b0;  addr_rom[ 4486]='h000010cc;  wr_data_rom[ 4486]='h00000000;
    rd_cycle[ 4487] = 1'b0;  wr_cycle[ 4487] = 1'b1;  addr_rom[ 4487]='h000009bc;  wr_data_rom[ 4487]='h000001be;
    rd_cycle[ 4488] = 1'b0;  wr_cycle[ 4488] = 1'b1;  addr_rom[ 4488]='h000000e0;  wr_data_rom[ 4488]='h00001449;
    rd_cycle[ 4489] = 1'b1;  wr_cycle[ 4489] = 1'b0;  addr_rom[ 4489]='h00000c28;  wr_data_rom[ 4489]='h00000000;
    rd_cycle[ 4490] = 1'b0;  wr_cycle[ 4490] = 1'b1;  addr_rom[ 4490]='h00000ac4;  wr_data_rom[ 4490]='h000007e7;
    rd_cycle[ 4491] = 1'b0;  wr_cycle[ 4491] = 1'b1;  addr_rom[ 4491]='h00001e94;  wr_data_rom[ 4491]='h00000005;
    rd_cycle[ 4492] = 1'b1;  wr_cycle[ 4492] = 1'b0;  addr_rom[ 4492]='h00000554;  wr_data_rom[ 4492]='h00000000;
    rd_cycle[ 4493] = 1'b0;  wr_cycle[ 4493] = 1'b1;  addr_rom[ 4493]='h00000dec;  wr_data_rom[ 4493]='h00000ffd;
    rd_cycle[ 4494] = 1'b0;  wr_cycle[ 4494] = 1'b1;  addr_rom[ 4494]='h00000bb4;  wr_data_rom[ 4494]='h00001165;
    rd_cycle[ 4495] = 1'b1;  wr_cycle[ 4495] = 1'b0;  addr_rom[ 4495]='h00000e9c;  wr_data_rom[ 4495]='h00000000;
    rd_cycle[ 4496] = 1'b0;  wr_cycle[ 4496] = 1'b1;  addr_rom[ 4496]='h00000030;  wr_data_rom[ 4496]='h00001f14;
    rd_cycle[ 4497] = 1'b0;  wr_cycle[ 4497] = 1'b1;  addr_rom[ 4497]='h00001e60;  wr_data_rom[ 4497]='h00001c18;
    rd_cycle[ 4498] = 1'b1;  wr_cycle[ 4498] = 1'b0;  addr_rom[ 4498]='h00001b8c;  wr_data_rom[ 4498]='h00000000;
    rd_cycle[ 4499] = 1'b0;  wr_cycle[ 4499] = 1'b1;  addr_rom[ 4499]='h000005b0;  wr_data_rom[ 4499]='h0000103a;
    rd_cycle[ 4500] = 1'b0;  wr_cycle[ 4500] = 1'b1;  addr_rom[ 4500]='h00001b40;  wr_data_rom[ 4500]='h00000001;
    rd_cycle[ 4501] = 1'b1;  wr_cycle[ 4501] = 1'b0;  addr_rom[ 4501]='h00000024;  wr_data_rom[ 4501]='h00000000;
    rd_cycle[ 4502] = 1'b0;  wr_cycle[ 4502] = 1'b1;  addr_rom[ 4502]='h0000179c;  wr_data_rom[ 4502]='h00001cc5;
    rd_cycle[ 4503] = 1'b0;  wr_cycle[ 4503] = 1'b1;  addr_rom[ 4503]='h000008a4;  wr_data_rom[ 4503]='h000015ac;
    rd_cycle[ 4504] = 1'b1;  wr_cycle[ 4504] = 1'b0;  addr_rom[ 4504]='h00001854;  wr_data_rom[ 4504]='h00000000;
    rd_cycle[ 4505] = 1'b0;  wr_cycle[ 4505] = 1'b1;  addr_rom[ 4505]='h00000b7c;  wr_data_rom[ 4505]='h000012e3;
    rd_cycle[ 4506] = 1'b0;  wr_cycle[ 4506] = 1'b1;  addr_rom[ 4506]='h000014c0;  wr_data_rom[ 4506]='h00000d85;
    rd_cycle[ 4507] = 1'b1;  wr_cycle[ 4507] = 1'b0;  addr_rom[ 4507]='h00000c44;  wr_data_rom[ 4507]='h00000000;
    rd_cycle[ 4508] = 1'b0;  wr_cycle[ 4508] = 1'b1;  addr_rom[ 4508]='h000006c8;  wr_data_rom[ 4508]='h000004df;
    rd_cycle[ 4509] = 1'b1;  wr_cycle[ 4509] = 1'b0;  addr_rom[ 4509]='h00000908;  wr_data_rom[ 4509]='h00000000;
    rd_cycle[ 4510] = 1'b1;  wr_cycle[ 4510] = 1'b0;  addr_rom[ 4510]='h00000bb4;  wr_data_rom[ 4510]='h00000000;
    rd_cycle[ 4511] = 1'b0;  wr_cycle[ 4511] = 1'b1;  addr_rom[ 4511]='h000011e0;  wr_data_rom[ 4511]='h0000050a;
    rd_cycle[ 4512] = 1'b0;  wr_cycle[ 4512] = 1'b1;  addr_rom[ 4512]='h000008e4;  wr_data_rom[ 4512]='h00001905;
    rd_cycle[ 4513] = 1'b0;  wr_cycle[ 4513] = 1'b1;  addr_rom[ 4513]='h00001900;  wr_data_rom[ 4513]='h00000a32;
    rd_cycle[ 4514] = 1'b0;  wr_cycle[ 4514] = 1'b1;  addr_rom[ 4514]='h00001148;  wr_data_rom[ 4514]='h000004d1;
    rd_cycle[ 4515] = 1'b1;  wr_cycle[ 4515] = 1'b0;  addr_rom[ 4515]='h0000016c;  wr_data_rom[ 4515]='h00000000;
    rd_cycle[ 4516] = 1'b0;  wr_cycle[ 4516] = 1'b1;  addr_rom[ 4516]='h00000ccc;  wr_data_rom[ 4516]='h00001e6f;
    rd_cycle[ 4517] = 1'b1;  wr_cycle[ 4517] = 1'b0;  addr_rom[ 4517]='h00001620;  wr_data_rom[ 4517]='h00000000;
    rd_cycle[ 4518] = 1'b0;  wr_cycle[ 4518] = 1'b1;  addr_rom[ 4518]='h00000bc0;  wr_data_rom[ 4518]='h00000846;
    rd_cycle[ 4519] = 1'b1;  wr_cycle[ 4519] = 1'b0;  addr_rom[ 4519]='h00001854;  wr_data_rom[ 4519]='h00000000;
    rd_cycle[ 4520] = 1'b0;  wr_cycle[ 4520] = 1'b1;  addr_rom[ 4520]='h00000408;  wr_data_rom[ 4520]='h00001ccf;
    rd_cycle[ 4521] = 1'b1;  wr_cycle[ 4521] = 1'b0;  addr_rom[ 4521]='h00000ec8;  wr_data_rom[ 4521]='h00000000;
    rd_cycle[ 4522] = 1'b0;  wr_cycle[ 4522] = 1'b1;  addr_rom[ 4522]='h00001938;  wr_data_rom[ 4522]='h00001436;
    rd_cycle[ 4523] = 1'b0;  wr_cycle[ 4523] = 1'b1;  addr_rom[ 4523]='h000015f8;  wr_data_rom[ 4523]='h00001a13;
    rd_cycle[ 4524] = 1'b0;  wr_cycle[ 4524] = 1'b1;  addr_rom[ 4524]='h000004a4;  wr_data_rom[ 4524]='h00000635;
    rd_cycle[ 4525] = 1'b0;  wr_cycle[ 4525] = 1'b1;  addr_rom[ 4525]='h00000744;  wr_data_rom[ 4525]='h000001a7;
    rd_cycle[ 4526] = 1'b0;  wr_cycle[ 4526] = 1'b1;  addr_rom[ 4526]='h000017f0;  wr_data_rom[ 4526]='h00001652;
    rd_cycle[ 4527] = 1'b1;  wr_cycle[ 4527] = 1'b0;  addr_rom[ 4527]='h00001ee0;  wr_data_rom[ 4527]='h00000000;
    rd_cycle[ 4528] = 1'b0;  wr_cycle[ 4528] = 1'b1;  addr_rom[ 4528]='h000006f8;  wr_data_rom[ 4528]='h00001146;
    rd_cycle[ 4529] = 1'b1;  wr_cycle[ 4529] = 1'b0;  addr_rom[ 4529]='h00000788;  wr_data_rom[ 4529]='h00000000;
    rd_cycle[ 4530] = 1'b1;  wr_cycle[ 4530] = 1'b0;  addr_rom[ 4530]='h00001824;  wr_data_rom[ 4530]='h00000000;
    rd_cycle[ 4531] = 1'b0;  wr_cycle[ 4531] = 1'b1;  addr_rom[ 4531]='h00001944;  wr_data_rom[ 4531]='h0000001c;
    rd_cycle[ 4532] = 1'b1;  wr_cycle[ 4532] = 1'b0;  addr_rom[ 4532]='h00000014;  wr_data_rom[ 4532]='h00000000;
    rd_cycle[ 4533] = 1'b0;  wr_cycle[ 4533] = 1'b1;  addr_rom[ 4533]='h00000698;  wr_data_rom[ 4533]='h00000661;
    rd_cycle[ 4534] = 1'b0;  wr_cycle[ 4534] = 1'b1;  addr_rom[ 4534]='h00001af0;  wr_data_rom[ 4534]='h00000df5;
    rd_cycle[ 4535] = 1'b1;  wr_cycle[ 4535] = 1'b0;  addr_rom[ 4535]='h000012bc;  wr_data_rom[ 4535]='h00000000;
    rd_cycle[ 4536] = 1'b0;  wr_cycle[ 4536] = 1'b1;  addr_rom[ 4536]='h00000968;  wr_data_rom[ 4536]='h00001328;
    rd_cycle[ 4537] = 1'b1;  wr_cycle[ 4537] = 1'b0;  addr_rom[ 4537]='h00000798;  wr_data_rom[ 4537]='h00000000;
    rd_cycle[ 4538] = 1'b0;  wr_cycle[ 4538] = 1'b1;  addr_rom[ 4538]='h0000193c;  wr_data_rom[ 4538]='h00001464;
    rd_cycle[ 4539] = 1'b0;  wr_cycle[ 4539] = 1'b1;  addr_rom[ 4539]='h00001138;  wr_data_rom[ 4539]='h00000f6c;
    rd_cycle[ 4540] = 1'b0;  wr_cycle[ 4540] = 1'b1;  addr_rom[ 4540]='h000007bc;  wr_data_rom[ 4540]='h0000080d;
    rd_cycle[ 4541] = 1'b1;  wr_cycle[ 4541] = 1'b0;  addr_rom[ 4541]='h00001c2c;  wr_data_rom[ 4541]='h00000000;
    rd_cycle[ 4542] = 1'b0;  wr_cycle[ 4542] = 1'b1;  addr_rom[ 4542]='h000008dc;  wr_data_rom[ 4542]='h0000150d;
    rd_cycle[ 4543] = 1'b0;  wr_cycle[ 4543] = 1'b1;  addr_rom[ 4543]='h00001cac;  wr_data_rom[ 4543]='h000012a4;
    rd_cycle[ 4544] = 1'b0;  wr_cycle[ 4544] = 1'b1;  addr_rom[ 4544]='h00000da0;  wr_data_rom[ 4544]='h000017fd;
    rd_cycle[ 4545] = 1'b1;  wr_cycle[ 4545] = 1'b0;  addr_rom[ 4545]='h000012f0;  wr_data_rom[ 4545]='h00000000;
    rd_cycle[ 4546] = 1'b1;  wr_cycle[ 4546] = 1'b0;  addr_rom[ 4546]='h00001c20;  wr_data_rom[ 4546]='h00000000;
    rd_cycle[ 4547] = 1'b0;  wr_cycle[ 4547] = 1'b1;  addr_rom[ 4547]='h000016e8;  wr_data_rom[ 4547]='h000007fe;
    rd_cycle[ 4548] = 1'b0;  wr_cycle[ 4548] = 1'b1;  addr_rom[ 4548]='h00001ed8;  wr_data_rom[ 4548]='h00000665;
    rd_cycle[ 4549] = 1'b0;  wr_cycle[ 4549] = 1'b1;  addr_rom[ 4549]='h00000490;  wr_data_rom[ 4549]='h00001285;
    rd_cycle[ 4550] = 1'b1;  wr_cycle[ 4550] = 1'b0;  addr_rom[ 4550]='h00001668;  wr_data_rom[ 4550]='h00000000;
    rd_cycle[ 4551] = 1'b1;  wr_cycle[ 4551] = 1'b0;  addr_rom[ 4551]='h000018c8;  wr_data_rom[ 4551]='h00000000;
    rd_cycle[ 4552] = 1'b0;  wr_cycle[ 4552] = 1'b1;  addr_rom[ 4552]='h00001860;  wr_data_rom[ 4552]='h000002ad;
    rd_cycle[ 4553] = 1'b0;  wr_cycle[ 4553] = 1'b1;  addr_rom[ 4553]='h00001db8;  wr_data_rom[ 4553]='h000002f9;
    rd_cycle[ 4554] = 1'b0;  wr_cycle[ 4554] = 1'b1;  addr_rom[ 4554]='h000015f8;  wr_data_rom[ 4554]='h00000c3c;
    rd_cycle[ 4555] = 1'b1;  wr_cycle[ 4555] = 1'b0;  addr_rom[ 4555]='h00001a50;  wr_data_rom[ 4555]='h00000000;
    rd_cycle[ 4556] = 1'b0;  wr_cycle[ 4556] = 1'b1;  addr_rom[ 4556]='h00000a4c;  wr_data_rom[ 4556]='h0000163a;
    rd_cycle[ 4557] = 1'b0;  wr_cycle[ 4557] = 1'b1;  addr_rom[ 4557]='h000010c4;  wr_data_rom[ 4557]='h0000023f;
    rd_cycle[ 4558] = 1'b0;  wr_cycle[ 4558] = 1'b1;  addr_rom[ 4558]='h000007fc;  wr_data_rom[ 4558]='h00001cab;
    rd_cycle[ 4559] = 1'b0;  wr_cycle[ 4559] = 1'b1;  addr_rom[ 4559]='h00000710;  wr_data_rom[ 4559]='h0000190e;
    rd_cycle[ 4560] = 1'b1;  wr_cycle[ 4560] = 1'b0;  addr_rom[ 4560]='h00000604;  wr_data_rom[ 4560]='h00000000;
    rd_cycle[ 4561] = 1'b1;  wr_cycle[ 4561] = 1'b0;  addr_rom[ 4561]='h00001234;  wr_data_rom[ 4561]='h00000000;
    rd_cycle[ 4562] = 1'b0;  wr_cycle[ 4562] = 1'b1;  addr_rom[ 4562]='h0000172c;  wr_data_rom[ 4562]='h0000179f;
    rd_cycle[ 4563] = 1'b0;  wr_cycle[ 4563] = 1'b1;  addr_rom[ 4563]='h00000b6c;  wr_data_rom[ 4563]='h00001403;
    rd_cycle[ 4564] = 1'b0;  wr_cycle[ 4564] = 1'b1;  addr_rom[ 4564]='h00001ee4;  wr_data_rom[ 4564]='h00001ad8;
    rd_cycle[ 4565] = 1'b1;  wr_cycle[ 4565] = 1'b0;  addr_rom[ 4565]='h00000608;  wr_data_rom[ 4565]='h00000000;
    rd_cycle[ 4566] = 1'b0;  wr_cycle[ 4566] = 1'b1;  addr_rom[ 4566]='h000011bc;  wr_data_rom[ 4566]='h00001d10;
    rd_cycle[ 4567] = 1'b0;  wr_cycle[ 4567] = 1'b1;  addr_rom[ 4567]='h00000ddc;  wr_data_rom[ 4567]='h000000d6;
    rd_cycle[ 4568] = 1'b1;  wr_cycle[ 4568] = 1'b0;  addr_rom[ 4568]='h00001ad8;  wr_data_rom[ 4568]='h00000000;
    rd_cycle[ 4569] = 1'b0;  wr_cycle[ 4569] = 1'b1;  addr_rom[ 4569]='h0000153c;  wr_data_rom[ 4569]='h00000a26;
    rd_cycle[ 4570] = 1'b0;  wr_cycle[ 4570] = 1'b1;  addr_rom[ 4570]='h00001570;  wr_data_rom[ 4570]='h00000b55;
    rd_cycle[ 4571] = 1'b1;  wr_cycle[ 4571] = 1'b0;  addr_rom[ 4571]='h000001a4;  wr_data_rom[ 4571]='h00000000;
    rd_cycle[ 4572] = 1'b0;  wr_cycle[ 4572] = 1'b1;  addr_rom[ 4572]='h000019cc;  wr_data_rom[ 4572]='h000001da;
    rd_cycle[ 4573] = 1'b1;  wr_cycle[ 4573] = 1'b0;  addr_rom[ 4573]='h00001f20;  wr_data_rom[ 4573]='h00000000;
    rd_cycle[ 4574] = 1'b0;  wr_cycle[ 4574] = 1'b1;  addr_rom[ 4574]='h00000e08;  wr_data_rom[ 4574]='h000018f1;
    rd_cycle[ 4575] = 1'b1;  wr_cycle[ 4575] = 1'b0;  addr_rom[ 4575]='h00001b1c;  wr_data_rom[ 4575]='h00000000;
    rd_cycle[ 4576] = 1'b1;  wr_cycle[ 4576] = 1'b0;  addr_rom[ 4576]='h00001d94;  wr_data_rom[ 4576]='h00000000;
    rd_cycle[ 4577] = 1'b0;  wr_cycle[ 4577] = 1'b1;  addr_rom[ 4577]='h0000036c;  wr_data_rom[ 4577]='h00000348;
    rd_cycle[ 4578] = 1'b1;  wr_cycle[ 4578] = 1'b0;  addr_rom[ 4578]='h000000c0;  wr_data_rom[ 4578]='h00000000;
    rd_cycle[ 4579] = 1'b1;  wr_cycle[ 4579] = 1'b0;  addr_rom[ 4579]='h00000ec4;  wr_data_rom[ 4579]='h00000000;
    rd_cycle[ 4580] = 1'b1;  wr_cycle[ 4580] = 1'b0;  addr_rom[ 4580]='h000005ac;  wr_data_rom[ 4580]='h00000000;
    rd_cycle[ 4581] = 1'b0;  wr_cycle[ 4581] = 1'b1;  addr_rom[ 4581]='h000013f8;  wr_data_rom[ 4581]='h00000c69;
    rd_cycle[ 4582] = 1'b1;  wr_cycle[ 4582] = 1'b0;  addr_rom[ 4582]='h00000de4;  wr_data_rom[ 4582]='h00000000;
    rd_cycle[ 4583] = 1'b1;  wr_cycle[ 4583] = 1'b0;  addr_rom[ 4583]='h00001454;  wr_data_rom[ 4583]='h00000000;
    rd_cycle[ 4584] = 1'b1;  wr_cycle[ 4584] = 1'b0;  addr_rom[ 4584]='h0000060c;  wr_data_rom[ 4584]='h00000000;
    rd_cycle[ 4585] = 1'b0;  wr_cycle[ 4585] = 1'b1;  addr_rom[ 4585]='h00001c48;  wr_data_rom[ 4585]='h00001192;
    rd_cycle[ 4586] = 1'b1;  wr_cycle[ 4586] = 1'b0;  addr_rom[ 4586]='h000002ac;  wr_data_rom[ 4586]='h00000000;
    rd_cycle[ 4587] = 1'b0;  wr_cycle[ 4587] = 1'b1;  addr_rom[ 4587]='h000012a8;  wr_data_rom[ 4587]='h000017bc;
    rd_cycle[ 4588] = 1'b1;  wr_cycle[ 4588] = 1'b0;  addr_rom[ 4588]='h0000006c;  wr_data_rom[ 4588]='h00000000;
    rd_cycle[ 4589] = 1'b1;  wr_cycle[ 4589] = 1'b0;  addr_rom[ 4589]='h00001540;  wr_data_rom[ 4589]='h00000000;
    rd_cycle[ 4590] = 1'b1;  wr_cycle[ 4590] = 1'b0;  addr_rom[ 4590]='h0000033c;  wr_data_rom[ 4590]='h00000000;
    rd_cycle[ 4591] = 1'b0;  wr_cycle[ 4591] = 1'b1;  addr_rom[ 4591]='h00000d28;  wr_data_rom[ 4591]='h000000a3;
    rd_cycle[ 4592] = 1'b1;  wr_cycle[ 4592] = 1'b0;  addr_rom[ 4592]='h000011cc;  wr_data_rom[ 4592]='h00000000;
    rd_cycle[ 4593] = 1'b1;  wr_cycle[ 4593] = 1'b0;  addr_rom[ 4593]='h00000874;  wr_data_rom[ 4593]='h00000000;
    rd_cycle[ 4594] = 1'b1;  wr_cycle[ 4594] = 1'b0;  addr_rom[ 4594]='h00001b6c;  wr_data_rom[ 4594]='h00000000;
    rd_cycle[ 4595] = 1'b0;  wr_cycle[ 4595] = 1'b1;  addr_rom[ 4595]='h00001050;  wr_data_rom[ 4595]='h0000128c;
    rd_cycle[ 4596] = 1'b1;  wr_cycle[ 4596] = 1'b0;  addr_rom[ 4596]='h00001614;  wr_data_rom[ 4596]='h00000000;
    rd_cycle[ 4597] = 1'b0;  wr_cycle[ 4597] = 1'b1;  addr_rom[ 4597]='h00001e00;  wr_data_rom[ 4597]='h000000d4;
    rd_cycle[ 4598] = 1'b0;  wr_cycle[ 4598] = 1'b1;  addr_rom[ 4598]='h000010c4;  wr_data_rom[ 4598]='h00001df7;
    rd_cycle[ 4599] = 1'b1;  wr_cycle[ 4599] = 1'b0;  addr_rom[ 4599]='h00001394;  wr_data_rom[ 4599]='h00000000;
    rd_cycle[ 4600] = 1'b1;  wr_cycle[ 4600] = 1'b0;  addr_rom[ 4600]='h00000a5c;  wr_data_rom[ 4600]='h00000000;
    rd_cycle[ 4601] = 1'b0;  wr_cycle[ 4601] = 1'b1;  addr_rom[ 4601]='h000015d4;  wr_data_rom[ 4601]='h0000097e;
    rd_cycle[ 4602] = 1'b1;  wr_cycle[ 4602] = 1'b0;  addr_rom[ 4602]='h000003cc;  wr_data_rom[ 4602]='h00000000;
    rd_cycle[ 4603] = 1'b0;  wr_cycle[ 4603] = 1'b1;  addr_rom[ 4603]='h00000304;  wr_data_rom[ 4603]='h0000096b;
    rd_cycle[ 4604] = 1'b1;  wr_cycle[ 4604] = 1'b0;  addr_rom[ 4604]='h00001798;  wr_data_rom[ 4604]='h00000000;
    rd_cycle[ 4605] = 1'b0;  wr_cycle[ 4605] = 1'b1;  addr_rom[ 4605]='h00001cb0;  wr_data_rom[ 4605]='h00000e04;
    rd_cycle[ 4606] = 1'b1;  wr_cycle[ 4606] = 1'b0;  addr_rom[ 4606]='h000019c4;  wr_data_rom[ 4606]='h00000000;
    rd_cycle[ 4607] = 1'b1;  wr_cycle[ 4607] = 1'b0;  addr_rom[ 4607]='h00000ed0;  wr_data_rom[ 4607]='h00000000;
    rd_cycle[ 4608] = 1'b0;  wr_cycle[ 4608] = 1'b1;  addr_rom[ 4608]='h00001b54;  wr_data_rom[ 4608]='h00000a59;
    rd_cycle[ 4609] = 1'b0;  wr_cycle[ 4609] = 1'b1;  addr_rom[ 4609]='h000019cc;  wr_data_rom[ 4609]='h000002f1;
    rd_cycle[ 4610] = 1'b0;  wr_cycle[ 4610] = 1'b1;  addr_rom[ 4610]='h00000eb4;  wr_data_rom[ 4610]='h0000048e;
    rd_cycle[ 4611] = 1'b1;  wr_cycle[ 4611] = 1'b0;  addr_rom[ 4611]='h00001568;  wr_data_rom[ 4611]='h00000000;
    rd_cycle[ 4612] = 1'b1;  wr_cycle[ 4612] = 1'b0;  addr_rom[ 4612]='h000011b4;  wr_data_rom[ 4612]='h00000000;
    rd_cycle[ 4613] = 1'b0;  wr_cycle[ 4613] = 1'b1;  addr_rom[ 4613]='h00001a04;  wr_data_rom[ 4613]='h000001cd;
    rd_cycle[ 4614] = 1'b1;  wr_cycle[ 4614] = 1'b0;  addr_rom[ 4614]='h00000488;  wr_data_rom[ 4614]='h00000000;
    rd_cycle[ 4615] = 1'b1;  wr_cycle[ 4615] = 1'b0;  addr_rom[ 4615]='h000014c0;  wr_data_rom[ 4615]='h00000000;
    rd_cycle[ 4616] = 1'b1;  wr_cycle[ 4616] = 1'b0;  addr_rom[ 4616]='h00001218;  wr_data_rom[ 4616]='h00000000;
    rd_cycle[ 4617] = 1'b1;  wr_cycle[ 4617] = 1'b0;  addr_rom[ 4617]='h00001014;  wr_data_rom[ 4617]='h00000000;
    rd_cycle[ 4618] = 1'b1;  wr_cycle[ 4618] = 1'b0;  addr_rom[ 4618]='h00000c8c;  wr_data_rom[ 4618]='h00000000;
    rd_cycle[ 4619] = 1'b1;  wr_cycle[ 4619] = 1'b0;  addr_rom[ 4619]='h000007e8;  wr_data_rom[ 4619]='h00000000;
    rd_cycle[ 4620] = 1'b0;  wr_cycle[ 4620] = 1'b1;  addr_rom[ 4620]='h00000164;  wr_data_rom[ 4620]='h000007c2;
    rd_cycle[ 4621] = 1'b1;  wr_cycle[ 4621] = 1'b0;  addr_rom[ 4621]='h000014ec;  wr_data_rom[ 4621]='h00000000;
    rd_cycle[ 4622] = 1'b1;  wr_cycle[ 4622] = 1'b0;  addr_rom[ 4622]='h0000147c;  wr_data_rom[ 4622]='h00000000;
    rd_cycle[ 4623] = 1'b0;  wr_cycle[ 4623] = 1'b1;  addr_rom[ 4623]='h00000a10;  wr_data_rom[ 4623]='h00001526;
    rd_cycle[ 4624] = 1'b0;  wr_cycle[ 4624] = 1'b1;  addr_rom[ 4624]='h0000189c;  wr_data_rom[ 4624]='h00000d44;
    rd_cycle[ 4625] = 1'b1;  wr_cycle[ 4625] = 1'b0;  addr_rom[ 4625]='h000010ac;  wr_data_rom[ 4625]='h00000000;
    rd_cycle[ 4626] = 1'b1;  wr_cycle[ 4626] = 1'b0;  addr_rom[ 4626]='h000011d4;  wr_data_rom[ 4626]='h00000000;
    rd_cycle[ 4627] = 1'b0;  wr_cycle[ 4627] = 1'b1;  addr_rom[ 4627]='h0000129c;  wr_data_rom[ 4627]='h00001bee;
    rd_cycle[ 4628] = 1'b0;  wr_cycle[ 4628] = 1'b1;  addr_rom[ 4628]='h00001550;  wr_data_rom[ 4628]='h0000068c;
    rd_cycle[ 4629] = 1'b0;  wr_cycle[ 4629] = 1'b1;  addr_rom[ 4629]='h00001718;  wr_data_rom[ 4629]='h000004e0;
    rd_cycle[ 4630] = 1'b1;  wr_cycle[ 4630] = 1'b0;  addr_rom[ 4630]='h00001898;  wr_data_rom[ 4630]='h00000000;
    rd_cycle[ 4631] = 1'b0;  wr_cycle[ 4631] = 1'b1;  addr_rom[ 4631]='h0000038c;  wr_data_rom[ 4631]='h000007c1;
    rd_cycle[ 4632] = 1'b0;  wr_cycle[ 4632] = 1'b1;  addr_rom[ 4632]='h000017e0;  wr_data_rom[ 4632]='h000015c5;
    rd_cycle[ 4633] = 1'b0;  wr_cycle[ 4633] = 1'b1;  addr_rom[ 4633]='h00001a74;  wr_data_rom[ 4633]='h00001084;
    rd_cycle[ 4634] = 1'b0;  wr_cycle[ 4634] = 1'b1;  addr_rom[ 4634]='h00000864;  wr_data_rom[ 4634]='h00001b75;
    rd_cycle[ 4635] = 1'b0;  wr_cycle[ 4635] = 1'b1;  addr_rom[ 4635]='h00001bd0;  wr_data_rom[ 4635]='h00001c2a;
    rd_cycle[ 4636] = 1'b1;  wr_cycle[ 4636] = 1'b0;  addr_rom[ 4636]='h00000b50;  wr_data_rom[ 4636]='h00000000;
    rd_cycle[ 4637] = 1'b0;  wr_cycle[ 4637] = 1'b1;  addr_rom[ 4637]='h0000042c;  wr_data_rom[ 4637]='h00000493;
    rd_cycle[ 4638] = 1'b0;  wr_cycle[ 4638] = 1'b1;  addr_rom[ 4638]='h00000be0;  wr_data_rom[ 4638]='h0000142c;
    rd_cycle[ 4639] = 1'b0;  wr_cycle[ 4639] = 1'b1;  addr_rom[ 4639]='h00001b98;  wr_data_rom[ 4639]='h000010d6;
    rd_cycle[ 4640] = 1'b0;  wr_cycle[ 4640] = 1'b1;  addr_rom[ 4640]='h0000147c;  wr_data_rom[ 4640]='h000014cc;
    rd_cycle[ 4641] = 1'b0;  wr_cycle[ 4641] = 1'b1;  addr_rom[ 4641]='h00001acc;  wr_data_rom[ 4641]='h00000209;
    rd_cycle[ 4642] = 1'b0;  wr_cycle[ 4642] = 1'b1;  addr_rom[ 4642]='h00000e74;  wr_data_rom[ 4642]='h0000103b;
    rd_cycle[ 4643] = 1'b1;  wr_cycle[ 4643] = 1'b0;  addr_rom[ 4643]='h000001a4;  wr_data_rom[ 4643]='h00000000;
    rd_cycle[ 4644] = 1'b1;  wr_cycle[ 4644] = 1'b0;  addr_rom[ 4644]='h000011cc;  wr_data_rom[ 4644]='h00000000;
    rd_cycle[ 4645] = 1'b1;  wr_cycle[ 4645] = 1'b0;  addr_rom[ 4645]='h00000c94;  wr_data_rom[ 4645]='h00000000;
    rd_cycle[ 4646] = 1'b0;  wr_cycle[ 4646] = 1'b1;  addr_rom[ 4646]='h00001e64;  wr_data_rom[ 4646]='h00001f2a;
    rd_cycle[ 4647] = 1'b0;  wr_cycle[ 4647] = 1'b1;  addr_rom[ 4647]='h000009fc;  wr_data_rom[ 4647]='h000006d0;
    rd_cycle[ 4648] = 1'b0;  wr_cycle[ 4648] = 1'b1;  addr_rom[ 4648]='h00001ef8;  wr_data_rom[ 4648]='h00000e67;
    rd_cycle[ 4649] = 1'b0;  wr_cycle[ 4649] = 1'b1;  addr_rom[ 4649]='h00001928;  wr_data_rom[ 4649]='h00001349;
    rd_cycle[ 4650] = 1'b0;  wr_cycle[ 4650] = 1'b1;  addr_rom[ 4650]='h00001b28;  wr_data_rom[ 4650]='h00001ec3;
    rd_cycle[ 4651] = 1'b0;  wr_cycle[ 4651] = 1'b1;  addr_rom[ 4651]='h00000c60;  wr_data_rom[ 4651]='h00000c61;
    rd_cycle[ 4652] = 1'b1;  wr_cycle[ 4652] = 1'b0;  addr_rom[ 4652]='h00001bd4;  wr_data_rom[ 4652]='h00000000;
    rd_cycle[ 4653] = 1'b1;  wr_cycle[ 4653] = 1'b0;  addr_rom[ 4653]='h000017d8;  wr_data_rom[ 4653]='h00000000;
    rd_cycle[ 4654] = 1'b1;  wr_cycle[ 4654] = 1'b0;  addr_rom[ 4654]='h00001414;  wr_data_rom[ 4654]='h00000000;
    rd_cycle[ 4655] = 1'b0;  wr_cycle[ 4655] = 1'b1;  addr_rom[ 4655]='h000005b8;  wr_data_rom[ 4655]='h000019ad;
    rd_cycle[ 4656] = 1'b1;  wr_cycle[ 4656] = 1'b0;  addr_rom[ 4656]='h0000176c;  wr_data_rom[ 4656]='h00000000;
    rd_cycle[ 4657] = 1'b1;  wr_cycle[ 4657] = 1'b0;  addr_rom[ 4657]='h00001cf0;  wr_data_rom[ 4657]='h00000000;
    rd_cycle[ 4658] = 1'b1;  wr_cycle[ 4658] = 1'b0;  addr_rom[ 4658]='h00001284;  wr_data_rom[ 4658]='h00000000;
    rd_cycle[ 4659] = 1'b0;  wr_cycle[ 4659] = 1'b1;  addr_rom[ 4659]='h00000f28;  wr_data_rom[ 4659]='h000006e6;
    rd_cycle[ 4660] = 1'b1;  wr_cycle[ 4660] = 1'b0;  addr_rom[ 4660]='h000015f0;  wr_data_rom[ 4660]='h00000000;
    rd_cycle[ 4661] = 1'b0;  wr_cycle[ 4661] = 1'b1;  addr_rom[ 4661]='h00001af4;  wr_data_rom[ 4661]='h000013ed;
    rd_cycle[ 4662] = 1'b1;  wr_cycle[ 4662] = 1'b0;  addr_rom[ 4662]='h00001be0;  wr_data_rom[ 4662]='h00000000;
    rd_cycle[ 4663] = 1'b0;  wr_cycle[ 4663] = 1'b1;  addr_rom[ 4663]='h00000b30;  wr_data_rom[ 4663]='h000015d6;
    rd_cycle[ 4664] = 1'b1;  wr_cycle[ 4664] = 1'b0;  addr_rom[ 4664]='h0000077c;  wr_data_rom[ 4664]='h00000000;
    rd_cycle[ 4665] = 1'b1;  wr_cycle[ 4665] = 1'b0;  addr_rom[ 4665]='h00000fb8;  wr_data_rom[ 4665]='h00000000;
    rd_cycle[ 4666] = 1'b0;  wr_cycle[ 4666] = 1'b1;  addr_rom[ 4666]='h0000001c;  wr_data_rom[ 4666]='h00000f20;
    rd_cycle[ 4667] = 1'b0;  wr_cycle[ 4667] = 1'b1;  addr_rom[ 4667]='h00000874;  wr_data_rom[ 4667]='h00001b85;
    rd_cycle[ 4668] = 1'b0;  wr_cycle[ 4668] = 1'b1;  addr_rom[ 4668]='h000010e0;  wr_data_rom[ 4668]='h0000033f;
    rd_cycle[ 4669] = 1'b0;  wr_cycle[ 4669] = 1'b1;  addr_rom[ 4669]='h00001b14;  wr_data_rom[ 4669]='h000019cb;
    rd_cycle[ 4670] = 1'b1;  wr_cycle[ 4670] = 1'b0;  addr_rom[ 4670]='h000019c0;  wr_data_rom[ 4670]='h00000000;
    rd_cycle[ 4671] = 1'b1;  wr_cycle[ 4671] = 1'b0;  addr_rom[ 4671]='h00000b60;  wr_data_rom[ 4671]='h00000000;
    rd_cycle[ 4672] = 1'b0;  wr_cycle[ 4672] = 1'b1;  addr_rom[ 4672]='h00000a98;  wr_data_rom[ 4672]='h00000755;
    rd_cycle[ 4673] = 1'b1;  wr_cycle[ 4673] = 1'b0;  addr_rom[ 4673]='h00001624;  wr_data_rom[ 4673]='h00000000;
    rd_cycle[ 4674] = 1'b1;  wr_cycle[ 4674] = 1'b0;  addr_rom[ 4674]='h000006f8;  wr_data_rom[ 4674]='h00000000;
    rd_cycle[ 4675] = 1'b0;  wr_cycle[ 4675] = 1'b1;  addr_rom[ 4675]='h00000420;  wr_data_rom[ 4675]='h000011cd;
    rd_cycle[ 4676] = 1'b0;  wr_cycle[ 4676] = 1'b1;  addr_rom[ 4676]='h000005b8;  wr_data_rom[ 4676]='h000003f7;
    rd_cycle[ 4677] = 1'b0;  wr_cycle[ 4677] = 1'b1;  addr_rom[ 4677]='h00000acc;  wr_data_rom[ 4677]='h000006ac;
    rd_cycle[ 4678] = 1'b0;  wr_cycle[ 4678] = 1'b1;  addr_rom[ 4678]='h00000594;  wr_data_rom[ 4678]='h00001783;
    rd_cycle[ 4679] = 1'b0;  wr_cycle[ 4679] = 1'b1;  addr_rom[ 4679]='h000008bc;  wr_data_rom[ 4679]='h00001a9e;
    rd_cycle[ 4680] = 1'b1;  wr_cycle[ 4680] = 1'b0;  addr_rom[ 4680]='h0000174c;  wr_data_rom[ 4680]='h00000000;
    rd_cycle[ 4681] = 1'b0;  wr_cycle[ 4681] = 1'b1;  addr_rom[ 4681]='h00000d50;  wr_data_rom[ 4681]='h00000750;
    rd_cycle[ 4682] = 1'b1;  wr_cycle[ 4682] = 1'b0;  addr_rom[ 4682]='h00000ea0;  wr_data_rom[ 4682]='h00000000;
    rd_cycle[ 4683] = 1'b0;  wr_cycle[ 4683] = 1'b1;  addr_rom[ 4683]='h0000069c;  wr_data_rom[ 4683]='h00001d43;
    rd_cycle[ 4684] = 1'b0;  wr_cycle[ 4684] = 1'b1;  addr_rom[ 4684]='h00001194;  wr_data_rom[ 4684]='h00000b08;
    rd_cycle[ 4685] = 1'b0;  wr_cycle[ 4685] = 1'b1;  addr_rom[ 4685]='h000007cc;  wr_data_rom[ 4685]='h00000846;
    rd_cycle[ 4686] = 1'b0;  wr_cycle[ 4686] = 1'b1;  addr_rom[ 4686]='h000018c8;  wr_data_rom[ 4686]='h000013d3;
    rd_cycle[ 4687] = 1'b0;  wr_cycle[ 4687] = 1'b1;  addr_rom[ 4687]='h000002a0;  wr_data_rom[ 4687]='h00000ac4;
    rd_cycle[ 4688] = 1'b1;  wr_cycle[ 4688] = 1'b0;  addr_rom[ 4688]='h00000dd8;  wr_data_rom[ 4688]='h00000000;
    rd_cycle[ 4689] = 1'b1;  wr_cycle[ 4689] = 1'b0;  addr_rom[ 4689]='h00001b0c;  wr_data_rom[ 4689]='h00000000;
    rd_cycle[ 4690] = 1'b0;  wr_cycle[ 4690] = 1'b1;  addr_rom[ 4690]='h000000e8;  wr_data_rom[ 4690]='h0000197a;
    rd_cycle[ 4691] = 1'b0;  wr_cycle[ 4691] = 1'b1;  addr_rom[ 4691]='h00001d0c;  wr_data_rom[ 4691]='h00000b29;
    rd_cycle[ 4692] = 1'b1;  wr_cycle[ 4692] = 1'b0;  addr_rom[ 4692]='h000002fc;  wr_data_rom[ 4692]='h00000000;
    rd_cycle[ 4693] = 1'b1;  wr_cycle[ 4693] = 1'b0;  addr_rom[ 4693]='h000007dc;  wr_data_rom[ 4693]='h00000000;
    rd_cycle[ 4694] = 1'b0;  wr_cycle[ 4694] = 1'b1;  addr_rom[ 4694]='h000002e0;  wr_data_rom[ 4694]='h0000140c;
    rd_cycle[ 4695] = 1'b1;  wr_cycle[ 4695] = 1'b0;  addr_rom[ 4695]='h00000214;  wr_data_rom[ 4695]='h00000000;
    rd_cycle[ 4696] = 1'b1;  wr_cycle[ 4696] = 1'b0;  addr_rom[ 4696]='h00001420;  wr_data_rom[ 4696]='h00000000;
    rd_cycle[ 4697] = 1'b1;  wr_cycle[ 4697] = 1'b0;  addr_rom[ 4697]='h0000010c;  wr_data_rom[ 4697]='h00000000;
    rd_cycle[ 4698] = 1'b0;  wr_cycle[ 4698] = 1'b1;  addr_rom[ 4698]='h00001b54;  wr_data_rom[ 4698]='h0000032b;
    rd_cycle[ 4699] = 1'b0;  wr_cycle[ 4699] = 1'b1;  addr_rom[ 4699]='h00000c88;  wr_data_rom[ 4699]='h0000012d;
    rd_cycle[ 4700] = 1'b0;  wr_cycle[ 4700] = 1'b1;  addr_rom[ 4700]='h00001eac;  wr_data_rom[ 4700]='h000002e1;
    rd_cycle[ 4701] = 1'b1;  wr_cycle[ 4701] = 1'b0;  addr_rom[ 4701]='h00001c4c;  wr_data_rom[ 4701]='h00000000;
    rd_cycle[ 4702] = 1'b1;  wr_cycle[ 4702] = 1'b0;  addr_rom[ 4702]='h000001b4;  wr_data_rom[ 4702]='h00000000;
    rd_cycle[ 4703] = 1'b0;  wr_cycle[ 4703] = 1'b1;  addr_rom[ 4703]='h00000c0c;  wr_data_rom[ 4703]='h00000ef3;
    rd_cycle[ 4704] = 1'b1;  wr_cycle[ 4704] = 1'b0;  addr_rom[ 4704]='h000011b0;  wr_data_rom[ 4704]='h00000000;
    rd_cycle[ 4705] = 1'b0;  wr_cycle[ 4705] = 1'b1;  addr_rom[ 4705]='h00000cf4;  wr_data_rom[ 4705]='h00000f98;
    rd_cycle[ 4706] = 1'b1;  wr_cycle[ 4706] = 1'b0;  addr_rom[ 4706]='h0000066c;  wr_data_rom[ 4706]='h00000000;
    rd_cycle[ 4707] = 1'b1;  wr_cycle[ 4707] = 1'b0;  addr_rom[ 4707]='h00001e24;  wr_data_rom[ 4707]='h00000000;
    rd_cycle[ 4708] = 1'b0;  wr_cycle[ 4708] = 1'b1;  addr_rom[ 4708]='h0000063c;  wr_data_rom[ 4708]='h00001ed2;
    rd_cycle[ 4709] = 1'b1;  wr_cycle[ 4709] = 1'b0;  addr_rom[ 4709]='h000015b4;  wr_data_rom[ 4709]='h00000000;
    rd_cycle[ 4710] = 1'b0;  wr_cycle[ 4710] = 1'b1;  addr_rom[ 4710]='h00000c9c;  wr_data_rom[ 4710]='h00000077;
    rd_cycle[ 4711] = 1'b1;  wr_cycle[ 4711] = 1'b0;  addr_rom[ 4711]='h00000540;  wr_data_rom[ 4711]='h00000000;
    rd_cycle[ 4712] = 1'b1;  wr_cycle[ 4712] = 1'b0;  addr_rom[ 4712]='h000004c8;  wr_data_rom[ 4712]='h00000000;
    rd_cycle[ 4713] = 1'b1;  wr_cycle[ 4713] = 1'b0;  addr_rom[ 4713]='h00000458;  wr_data_rom[ 4713]='h00000000;
    rd_cycle[ 4714] = 1'b0;  wr_cycle[ 4714] = 1'b1;  addr_rom[ 4714]='h00001e40;  wr_data_rom[ 4714]='h00000254;
    rd_cycle[ 4715] = 1'b1;  wr_cycle[ 4715] = 1'b0;  addr_rom[ 4715]='h00001004;  wr_data_rom[ 4715]='h00000000;
    rd_cycle[ 4716] = 1'b0;  wr_cycle[ 4716] = 1'b1;  addr_rom[ 4716]='h00001350;  wr_data_rom[ 4716]='h00001a21;
    rd_cycle[ 4717] = 1'b0;  wr_cycle[ 4717] = 1'b1;  addr_rom[ 4717]='h00001b74;  wr_data_rom[ 4717]='h000007ce;
    rd_cycle[ 4718] = 1'b0;  wr_cycle[ 4718] = 1'b1;  addr_rom[ 4718]='h000018ac;  wr_data_rom[ 4718]='h00001468;
    rd_cycle[ 4719] = 1'b1;  wr_cycle[ 4719] = 1'b0;  addr_rom[ 4719]='h000013c8;  wr_data_rom[ 4719]='h00000000;
    rd_cycle[ 4720] = 1'b1;  wr_cycle[ 4720] = 1'b0;  addr_rom[ 4720]='h00000d90;  wr_data_rom[ 4720]='h00000000;
    rd_cycle[ 4721] = 1'b1;  wr_cycle[ 4721] = 1'b0;  addr_rom[ 4721]='h0000180c;  wr_data_rom[ 4721]='h00000000;
    rd_cycle[ 4722] = 1'b1;  wr_cycle[ 4722] = 1'b0;  addr_rom[ 4722]='h000008d0;  wr_data_rom[ 4722]='h00000000;
    rd_cycle[ 4723] = 1'b1;  wr_cycle[ 4723] = 1'b0;  addr_rom[ 4723]='h00001d4c;  wr_data_rom[ 4723]='h00000000;
    rd_cycle[ 4724] = 1'b1;  wr_cycle[ 4724] = 1'b0;  addr_rom[ 4724]='h00001eb8;  wr_data_rom[ 4724]='h00000000;
    rd_cycle[ 4725] = 1'b0;  wr_cycle[ 4725] = 1'b1;  addr_rom[ 4725]='h00001000;  wr_data_rom[ 4725]='h00000f40;
    rd_cycle[ 4726] = 1'b0;  wr_cycle[ 4726] = 1'b1;  addr_rom[ 4726]='h00001d74;  wr_data_rom[ 4726]='h0000060b;
    rd_cycle[ 4727] = 1'b1;  wr_cycle[ 4727] = 1'b0;  addr_rom[ 4727]='h00000ed4;  wr_data_rom[ 4727]='h00000000;
    rd_cycle[ 4728] = 1'b1;  wr_cycle[ 4728] = 1'b0;  addr_rom[ 4728]='h000006e0;  wr_data_rom[ 4728]='h00000000;
    rd_cycle[ 4729] = 1'b1;  wr_cycle[ 4729] = 1'b0;  addr_rom[ 4729]='h00000c1c;  wr_data_rom[ 4729]='h00000000;
    rd_cycle[ 4730] = 1'b1;  wr_cycle[ 4730] = 1'b0;  addr_rom[ 4730]='h0000099c;  wr_data_rom[ 4730]='h00000000;
    rd_cycle[ 4731] = 1'b1;  wr_cycle[ 4731] = 1'b0;  addr_rom[ 4731]='h00000434;  wr_data_rom[ 4731]='h00000000;
    rd_cycle[ 4732] = 1'b0;  wr_cycle[ 4732] = 1'b1;  addr_rom[ 4732]='h00000544;  wr_data_rom[ 4732]='h0000061d;
    rd_cycle[ 4733] = 1'b1;  wr_cycle[ 4733] = 1'b0;  addr_rom[ 4733]='h000010c4;  wr_data_rom[ 4733]='h00000000;
    rd_cycle[ 4734] = 1'b0;  wr_cycle[ 4734] = 1'b1;  addr_rom[ 4734]='h00001a54;  wr_data_rom[ 4734]='h00001054;
    rd_cycle[ 4735] = 1'b0;  wr_cycle[ 4735] = 1'b1;  addr_rom[ 4735]='h00001f14;  wr_data_rom[ 4735]='h000018ba;
    rd_cycle[ 4736] = 1'b1;  wr_cycle[ 4736] = 1'b0;  addr_rom[ 4736]='h00001040;  wr_data_rom[ 4736]='h00000000;
    rd_cycle[ 4737] = 1'b0;  wr_cycle[ 4737] = 1'b1;  addr_rom[ 4737]='h0000037c;  wr_data_rom[ 4737]='h0000079f;
    rd_cycle[ 4738] = 1'b0;  wr_cycle[ 4738] = 1'b1;  addr_rom[ 4738]='h000018dc;  wr_data_rom[ 4738]='h00000bcf;
    rd_cycle[ 4739] = 1'b0;  wr_cycle[ 4739] = 1'b1;  addr_rom[ 4739]='h000009d0;  wr_data_rom[ 4739]='h00001030;
    rd_cycle[ 4740] = 1'b1;  wr_cycle[ 4740] = 1'b0;  addr_rom[ 4740]='h00000bd0;  wr_data_rom[ 4740]='h00000000;
    rd_cycle[ 4741] = 1'b0;  wr_cycle[ 4741] = 1'b1;  addr_rom[ 4741]='h000018b4;  wr_data_rom[ 4741]='h0000062c;
    rd_cycle[ 4742] = 1'b1;  wr_cycle[ 4742] = 1'b0;  addr_rom[ 4742]='h00000f34;  wr_data_rom[ 4742]='h00000000;
    rd_cycle[ 4743] = 1'b0;  wr_cycle[ 4743] = 1'b1;  addr_rom[ 4743]='h000016fc;  wr_data_rom[ 4743]='h00001859;
    rd_cycle[ 4744] = 1'b1;  wr_cycle[ 4744] = 1'b0;  addr_rom[ 4744]='h00000e2c;  wr_data_rom[ 4744]='h00000000;
    rd_cycle[ 4745] = 1'b1;  wr_cycle[ 4745] = 1'b0;  addr_rom[ 4745]='h00000c60;  wr_data_rom[ 4745]='h00000000;
    rd_cycle[ 4746] = 1'b0;  wr_cycle[ 4746] = 1'b1;  addr_rom[ 4746]='h00001ab8;  wr_data_rom[ 4746]='h00000ca8;
    rd_cycle[ 4747] = 1'b1;  wr_cycle[ 4747] = 1'b0;  addr_rom[ 4747]='h00000a64;  wr_data_rom[ 4747]='h00000000;
    rd_cycle[ 4748] = 1'b1;  wr_cycle[ 4748] = 1'b0;  addr_rom[ 4748]='h0000003c;  wr_data_rom[ 4748]='h00000000;
    rd_cycle[ 4749] = 1'b1;  wr_cycle[ 4749] = 1'b0;  addr_rom[ 4749]='h00000ed8;  wr_data_rom[ 4749]='h00000000;
    rd_cycle[ 4750] = 1'b0;  wr_cycle[ 4750] = 1'b1;  addr_rom[ 4750]='h00000da8;  wr_data_rom[ 4750]='h0000127a;
    rd_cycle[ 4751] = 1'b1;  wr_cycle[ 4751] = 1'b0;  addr_rom[ 4751]='h000010f8;  wr_data_rom[ 4751]='h00000000;
    rd_cycle[ 4752] = 1'b1;  wr_cycle[ 4752] = 1'b0;  addr_rom[ 4752]='h00000be0;  wr_data_rom[ 4752]='h00000000;
    rd_cycle[ 4753] = 1'b1;  wr_cycle[ 4753] = 1'b0;  addr_rom[ 4753]='h00001cdc;  wr_data_rom[ 4753]='h00000000;
    rd_cycle[ 4754] = 1'b1;  wr_cycle[ 4754] = 1'b0;  addr_rom[ 4754]='h00000698;  wr_data_rom[ 4754]='h00000000;
    rd_cycle[ 4755] = 1'b0;  wr_cycle[ 4755] = 1'b1;  addr_rom[ 4755]='h00000074;  wr_data_rom[ 4755]='h000008cf;
    rd_cycle[ 4756] = 1'b1;  wr_cycle[ 4756] = 1'b0;  addr_rom[ 4756]='h00000a7c;  wr_data_rom[ 4756]='h00000000;
    rd_cycle[ 4757] = 1'b0;  wr_cycle[ 4757] = 1'b1;  addr_rom[ 4757]='h00001b3c;  wr_data_rom[ 4757]='h00000a28;
    rd_cycle[ 4758] = 1'b0;  wr_cycle[ 4758] = 1'b1;  addr_rom[ 4758]='h00000664;  wr_data_rom[ 4758]='h000009f6;
    rd_cycle[ 4759] = 1'b1;  wr_cycle[ 4759] = 1'b0;  addr_rom[ 4759]='h000011a4;  wr_data_rom[ 4759]='h00000000;
    rd_cycle[ 4760] = 1'b1;  wr_cycle[ 4760] = 1'b0;  addr_rom[ 4760]='h00001cc8;  wr_data_rom[ 4760]='h00000000;
    rd_cycle[ 4761] = 1'b1;  wr_cycle[ 4761] = 1'b0;  addr_rom[ 4761]='h00001304;  wr_data_rom[ 4761]='h00000000;
    rd_cycle[ 4762] = 1'b0;  wr_cycle[ 4762] = 1'b1;  addr_rom[ 4762]='h00001f20;  wr_data_rom[ 4762]='h00000496;
    rd_cycle[ 4763] = 1'b1;  wr_cycle[ 4763] = 1'b0;  addr_rom[ 4763]='h000003fc;  wr_data_rom[ 4763]='h00000000;
    rd_cycle[ 4764] = 1'b0;  wr_cycle[ 4764] = 1'b1;  addr_rom[ 4764]='h0000195c;  wr_data_rom[ 4764]='h00001cae;
    rd_cycle[ 4765] = 1'b1;  wr_cycle[ 4765] = 1'b0;  addr_rom[ 4765]='h0000129c;  wr_data_rom[ 4765]='h00000000;
    rd_cycle[ 4766] = 1'b0;  wr_cycle[ 4766] = 1'b1;  addr_rom[ 4766]='h000004c8;  wr_data_rom[ 4766]='h0000193a;
    rd_cycle[ 4767] = 1'b0;  wr_cycle[ 4767] = 1'b1;  addr_rom[ 4767]='h0000030c;  wr_data_rom[ 4767]='h000003db;
    rd_cycle[ 4768] = 1'b1;  wr_cycle[ 4768] = 1'b0;  addr_rom[ 4768]='h0000141c;  wr_data_rom[ 4768]='h00000000;
    rd_cycle[ 4769] = 1'b0;  wr_cycle[ 4769] = 1'b1;  addr_rom[ 4769]='h00001588;  wr_data_rom[ 4769]='h00001841;
    rd_cycle[ 4770] = 1'b0;  wr_cycle[ 4770] = 1'b1;  addr_rom[ 4770]='h00001974;  wr_data_rom[ 4770]='h00001d1d;
    rd_cycle[ 4771] = 1'b1;  wr_cycle[ 4771] = 1'b0;  addr_rom[ 4771]='h00001748;  wr_data_rom[ 4771]='h00000000;
    rd_cycle[ 4772] = 1'b0;  wr_cycle[ 4772] = 1'b1;  addr_rom[ 4772]='h0000037c;  wr_data_rom[ 4772]='h00000a9e;
    rd_cycle[ 4773] = 1'b0;  wr_cycle[ 4773] = 1'b1;  addr_rom[ 4773]='h00000cf4;  wr_data_rom[ 4773]='h000004f6;
    rd_cycle[ 4774] = 1'b0;  wr_cycle[ 4774] = 1'b1;  addr_rom[ 4774]='h0000113c;  wr_data_rom[ 4774]='h00000159;
    rd_cycle[ 4775] = 1'b0;  wr_cycle[ 4775] = 1'b1;  addr_rom[ 4775]='h000007d8;  wr_data_rom[ 4775]='h0000144d;
    rd_cycle[ 4776] = 1'b1;  wr_cycle[ 4776] = 1'b0;  addr_rom[ 4776]='h00001b90;  wr_data_rom[ 4776]='h00000000;
    rd_cycle[ 4777] = 1'b0;  wr_cycle[ 4777] = 1'b1;  addr_rom[ 4777]='h00001910;  wr_data_rom[ 4777]='h00000926;
    rd_cycle[ 4778] = 1'b1;  wr_cycle[ 4778] = 1'b0;  addr_rom[ 4778]='h00000598;  wr_data_rom[ 4778]='h00000000;
    rd_cycle[ 4779] = 1'b0;  wr_cycle[ 4779] = 1'b1;  addr_rom[ 4779]='h000009cc;  wr_data_rom[ 4779]='h00001970;
    rd_cycle[ 4780] = 1'b1;  wr_cycle[ 4780] = 1'b0;  addr_rom[ 4780]='h00000c04;  wr_data_rom[ 4780]='h00000000;
    rd_cycle[ 4781] = 1'b0;  wr_cycle[ 4781] = 1'b1;  addr_rom[ 4781]='h000007ac;  wr_data_rom[ 4781]='h00000171;
    rd_cycle[ 4782] = 1'b1;  wr_cycle[ 4782] = 1'b0;  addr_rom[ 4782]='h00001c6c;  wr_data_rom[ 4782]='h00000000;
    rd_cycle[ 4783] = 1'b1;  wr_cycle[ 4783] = 1'b0;  addr_rom[ 4783]='h00001eb4;  wr_data_rom[ 4783]='h00000000;
    rd_cycle[ 4784] = 1'b0;  wr_cycle[ 4784] = 1'b1;  addr_rom[ 4784]='h00001c20;  wr_data_rom[ 4784]='h00000bee;
    rd_cycle[ 4785] = 1'b0;  wr_cycle[ 4785] = 1'b1;  addr_rom[ 4785]='h000015ac;  wr_data_rom[ 4785]='h000001be;
    rd_cycle[ 4786] = 1'b1;  wr_cycle[ 4786] = 1'b0;  addr_rom[ 4786]='h00001ec4;  wr_data_rom[ 4786]='h00000000;
    rd_cycle[ 4787] = 1'b0;  wr_cycle[ 4787] = 1'b1;  addr_rom[ 4787]='h000016a8;  wr_data_rom[ 4787]='h00000ae2;
    rd_cycle[ 4788] = 1'b1;  wr_cycle[ 4788] = 1'b0;  addr_rom[ 4788]='h00001104;  wr_data_rom[ 4788]='h00000000;
    rd_cycle[ 4789] = 1'b0;  wr_cycle[ 4789] = 1'b1;  addr_rom[ 4789]='h00000f84;  wr_data_rom[ 4789]='h00001053;
    rd_cycle[ 4790] = 1'b1;  wr_cycle[ 4790] = 1'b0;  addr_rom[ 4790]='h000010f0;  wr_data_rom[ 4790]='h00000000;
    rd_cycle[ 4791] = 1'b1;  wr_cycle[ 4791] = 1'b0;  addr_rom[ 4791]='h000011dc;  wr_data_rom[ 4791]='h00000000;
    rd_cycle[ 4792] = 1'b1;  wr_cycle[ 4792] = 1'b0;  addr_rom[ 4792]='h000010e8;  wr_data_rom[ 4792]='h00000000;
    rd_cycle[ 4793] = 1'b1;  wr_cycle[ 4793] = 1'b0;  addr_rom[ 4793]='h00001468;  wr_data_rom[ 4793]='h00000000;
    rd_cycle[ 4794] = 1'b1;  wr_cycle[ 4794] = 1'b0;  addr_rom[ 4794]='h00000ba4;  wr_data_rom[ 4794]='h00000000;
    rd_cycle[ 4795] = 1'b1;  wr_cycle[ 4795] = 1'b0;  addr_rom[ 4795]='h00000be8;  wr_data_rom[ 4795]='h00000000;
    rd_cycle[ 4796] = 1'b0;  wr_cycle[ 4796] = 1'b1;  addr_rom[ 4796]='h00000638;  wr_data_rom[ 4796]='h00001387;
    rd_cycle[ 4797] = 1'b0;  wr_cycle[ 4797] = 1'b1;  addr_rom[ 4797]='h00000f78;  wr_data_rom[ 4797]='h00001970;
    rd_cycle[ 4798] = 1'b1;  wr_cycle[ 4798] = 1'b0;  addr_rom[ 4798]='h00001594;  wr_data_rom[ 4798]='h00000000;
    rd_cycle[ 4799] = 1'b0;  wr_cycle[ 4799] = 1'b1;  addr_rom[ 4799]='h00000f78;  wr_data_rom[ 4799]='h00000f6d;
    rd_cycle[ 4800] = 1'b1;  wr_cycle[ 4800] = 1'b0;  addr_rom[ 4800]='h00000848;  wr_data_rom[ 4800]='h00000000;
    rd_cycle[ 4801] = 1'b1;  wr_cycle[ 4801] = 1'b0;  addr_rom[ 4801]='h00000964;  wr_data_rom[ 4801]='h00000000;
    rd_cycle[ 4802] = 1'b1;  wr_cycle[ 4802] = 1'b0;  addr_rom[ 4802]='h00001cd4;  wr_data_rom[ 4802]='h00000000;
    rd_cycle[ 4803] = 1'b0;  wr_cycle[ 4803] = 1'b1;  addr_rom[ 4803]='h00000ef8;  wr_data_rom[ 4803]='h00001d87;
    rd_cycle[ 4804] = 1'b1;  wr_cycle[ 4804] = 1'b0;  addr_rom[ 4804]='h00000ce8;  wr_data_rom[ 4804]='h00000000;
    rd_cycle[ 4805] = 1'b0;  wr_cycle[ 4805] = 1'b1;  addr_rom[ 4805]='h00001630;  wr_data_rom[ 4805]='h00000daa;
    rd_cycle[ 4806] = 1'b1;  wr_cycle[ 4806] = 1'b0;  addr_rom[ 4806]='h00001598;  wr_data_rom[ 4806]='h00000000;
    rd_cycle[ 4807] = 1'b0;  wr_cycle[ 4807] = 1'b1;  addr_rom[ 4807]='h000002d4;  wr_data_rom[ 4807]='h00001770;
    rd_cycle[ 4808] = 1'b0;  wr_cycle[ 4808] = 1'b1;  addr_rom[ 4808]='h000008e4;  wr_data_rom[ 4808]='h00001e72;
    rd_cycle[ 4809] = 1'b0;  wr_cycle[ 4809] = 1'b1;  addr_rom[ 4809]='h00000268;  wr_data_rom[ 4809]='h000019ab;
    rd_cycle[ 4810] = 1'b1;  wr_cycle[ 4810] = 1'b0;  addr_rom[ 4810]='h00001244;  wr_data_rom[ 4810]='h00000000;
    rd_cycle[ 4811] = 1'b1;  wr_cycle[ 4811] = 1'b0;  addr_rom[ 4811]='h00001724;  wr_data_rom[ 4811]='h00000000;
    rd_cycle[ 4812] = 1'b1;  wr_cycle[ 4812] = 1'b0;  addr_rom[ 4812]='h00000e30;  wr_data_rom[ 4812]='h00000000;
    rd_cycle[ 4813] = 1'b0;  wr_cycle[ 4813] = 1'b1;  addr_rom[ 4813]='h00001600;  wr_data_rom[ 4813]='h000010ac;
    rd_cycle[ 4814] = 1'b0;  wr_cycle[ 4814] = 1'b1;  addr_rom[ 4814]='h00001400;  wr_data_rom[ 4814]='h000007dd;
    rd_cycle[ 4815] = 1'b0;  wr_cycle[ 4815] = 1'b1;  addr_rom[ 4815]='h00000314;  wr_data_rom[ 4815]='h00000c12;
    rd_cycle[ 4816] = 1'b1;  wr_cycle[ 4816] = 1'b0;  addr_rom[ 4816]='h00000e10;  wr_data_rom[ 4816]='h00000000;
    rd_cycle[ 4817] = 1'b0;  wr_cycle[ 4817] = 1'b1;  addr_rom[ 4817]='h000002ac;  wr_data_rom[ 4817]='h00000cea;
    rd_cycle[ 4818] = 1'b1;  wr_cycle[ 4818] = 1'b0;  addr_rom[ 4818]='h000014c0;  wr_data_rom[ 4818]='h00000000;
    rd_cycle[ 4819] = 1'b0;  wr_cycle[ 4819] = 1'b1;  addr_rom[ 4819]='h000012f0;  wr_data_rom[ 4819]='h000000bc;
    rd_cycle[ 4820] = 1'b0;  wr_cycle[ 4820] = 1'b1;  addr_rom[ 4820]='h00001540;  wr_data_rom[ 4820]='h00001b66;
    rd_cycle[ 4821] = 1'b0;  wr_cycle[ 4821] = 1'b1;  addr_rom[ 4821]='h00000318;  wr_data_rom[ 4821]='h00000f40;
    rd_cycle[ 4822] = 1'b1;  wr_cycle[ 4822] = 1'b0;  addr_rom[ 4822]='h0000073c;  wr_data_rom[ 4822]='h00000000;
    rd_cycle[ 4823] = 1'b1;  wr_cycle[ 4823] = 1'b0;  addr_rom[ 4823]='h00001738;  wr_data_rom[ 4823]='h00000000;
    rd_cycle[ 4824] = 1'b1;  wr_cycle[ 4824] = 1'b0;  addr_rom[ 4824]='h00001324;  wr_data_rom[ 4824]='h00000000;
    rd_cycle[ 4825] = 1'b0;  wr_cycle[ 4825] = 1'b1;  addr_rom[ 4825]='h00001920;  wr_data_rom[ 4825]='h00001341;
    rd_cycle[ 4826] = 1'b1;  wr_cycle[ 4826] = 1'b0;  addr_rom[ 4826]='h000014c8;  wr_data_rom[ 4826]='h00000000;
    rd_cycle[ 4827] = 1'b0;  wr_cycle[ 4827] = 1'b1;  addr_rom[ 4827]='h00000748;  wr_data_rom[ 4827]='h0000132d;
    rd_cycle[ 4828] = 1'b1;  wr_cycle[ 4828] = 1'b0;  addr_rom[ 4828]='h000005f8;  wr_data_rom[ 4828]='h00000000;
    rd_cycle[ 4829] = 1'b1;  wr_cycle[ 4829] = 1'b0;  addr_rom[ 4829]='h00001468;  wr_data_rom[ 4829]='h00000000;
    rd_cycle[ 4830] = 1'b1;  wr_cycle[ 4830] = 1'b0;  addr_rom[ 4830]='h00001988;  wr_data_rom[ 4830]='h00000000;
    rd_cycle[ 4831] = 1'b1;  wr_cycle[ 4831] = 1'b0;  addr_rom[ 4831]='h00001bb8;  wr_data_rom[ 4831]='h00000000;
    rd_cycle[ 4832] = 1'b1;  wr_cycle[ 4832] = 1'b0;  addr_rom[ 4832]='h00000d4c;  wr_data_rom[ 4832]='h00000000;
    rd_cycle[ 4833] = 1'b0;  wr_cycle[ 4833] = 1'b1;  addr_rom[ 4833]='h00000ec0;  wr_data_rom[ 4833]='h00000625;
    rd_cycle[ 4834] = 1'b0;  wr_cycle[ 4834] = 1'b1;  addr_rom[ 4834]='h00001288;  wr_data_rom[ 4834]='h00000763;
    rd_cycle[ 4835] = 1'b1;  wr_cycle[ 4835] = 1'b0;  addr_rom[ 4835]='h00000e00;  wr_data_rom[ 4835]='h00000000;
    rd_cycle[ 4836] = 1'b0;  wr_cycle[ 4836] = 1'b1;  addr_rom[ 4836]='h00000bb4;  wr_data_rom[ 4836]='h00001393;
    rd_cycle[ 4837] = 1'b0;  wr_cycle[ 4837] = 1'b1;  addr_rom[ 4837]='h00001cac;  wr_data_rom[ 4837]='h000017d8;
    rd_cycle[ 4838] = 1'b0;  wr_cycle[ 4838] = 1'b1;  addr_rom[ 4838]='h00001900;  wr_data_rom[ 4838]='h000019c9;
    rd_cycle[ 4839] = 1'b1;  wr_cycle[ 4839] = 1'b0;  addr_rom[ 4839]='h000015d8;  wr_data_rom[ 4839]='h00000000;
    rd_cycle[ 4840] = 1'b1;  wr_cycle[ 4840] = 1'b0;  addr_rom[ 4840]='h000014f0;  wr_data_rom[ 4840]='h00000000;
    rd_cycle[ 4841] = 1'b1;  wr_cycle[ 4841] = 1'b0;  addr_rom[ 4841]='h0000021c;  wr_data_rom[ 4841]='h00000000;
    rd_cycle[ 4842] = 1'b0;  wr_cycle[ 4842] = 1'b1;  addr_rom[ 4842]='h00001c88;  wr_data_rom[ 4842]='h000005d6;
    rd_cycle[ 4843] = 1'b1;  wr_cycle[ 4843] = 1'b0;  addr_rom[ 4843]='h0000072c;  wr_data_rom[ 4843]='h00000000;
    rd_cycle[ 4844] = 1'b1;  wr_cycle[ 4844] = 1'b0;  addr_rom[ 4844]='h00001a08;  wr_data_rom[ 4844]='h00000000;
    rd_cycle[ 4845] = 1'b1;  wr_cycle[ 4845] = 1'b0;  addr_rom[ 4845]='h00001a34;  wr_data_rom[ 4845]='h00000000;
    rd_cycle[ 4846] = 1'b0;  wr_cycle[ 4846] = 1'b1;  addr_rom[ 4846]='h00001b2c;  wr_data_rom[ 4846]='h00000a35;
    rd_cycle[ 4847] = 1'b1;  wr_cycle[ 4847] = 1'b0;  addr_rom[ 4847]='h00000e70;  wr_data_rom[ 4847]='h00000000;
    rd_cycle[ 4848] = 1'b1;  wr_cycle[ 4848] = 1'b0;  addr_rom[ 4848]='h00000430;  wr_data_rom[ 4848]='h00000000;
    rd_cycle[ 4849] = 1'b1;  wr_cycle[ 4849] = 1'b0;  addr_rom[ 4849]='h00001bdc;  wr_data_rom[ 4849]='h00000000;
    rd_cycle[ 4850] = 1'b0;  wr_cycle[ 4850] = 1'b1;  addr_rom[ 4850]='h00000a88;  wr_data_rom[ 4850]='h00001776;
    rd_cycle[ 4851] = 1'b1;  wr_cycle[ 4851] = 1'b0;  addr_rom[ 4851]='h00001160;  wr_data_rom[ 4851]='h00000000;
    rd_cycle[ 4852] = 1'b1;  wr_cycle[ 4852] = 1'b0;  addr_rom[ 4852]='h00001078;  wr_data_rom[ 4852]='h00000000;
    rd_cycle[ 4853] = 1'b0;  wr_cycle[ 4853] = 1'b1;  addr_rom[ 4853]='h000002d8;  wr_data_rom[ 4853]='h00001035;
    rd_cycle[ 4854] = 1'b1;  wr_cycle[ 4854] = 1'b0;  addr_rom[ 4854]='h00000478;  wr_data_rom[ 4854]='h00000000;
    rd_cycle[ 4855] = 1'b0;  wr_cycle[ 4855] = 1'b1;  addr_rom[ 4855]='h00000280;  wr_data_rom[ 4855]='h00001da0;
    rd_cycle[ 4856] = 1'b1;  wr_cycle[ 4856] = 1'b0;  addr_rom[ 4856]='h00001de8;  wr_data_rom[ 4856]='h00000000;
    rd_cycle[ 4857] = 1'b1;  wr_cycle[ 4857] = 1'b0;  addr_rom[ 4857]='h00001cb0;  wr_data_rom[ 4857]='h00000000;
    rd_cycle[ 4858] = 1'b1;  wr_cycle[ 4858] = 1'b0;  addr_rom[ 4858]='h000015b0;  wr_data_rom[ 4858]='h00000000;
    rd_cycle[ 4859] = 1'b0;  wr_cycle[ 4859] = 1'b1;  addr_rom[ 4859]='h00001c7c;  wr_data_rom[ 4859]='h00001984;
    rd_cycle[ 4860] = 1'b1;  wr_cycle[ 4860] = 1'b0;  addr_rom[ 4860]='h000006bc;  wr_data_rom[ 4860]='h00000000;
    rd_cycle[ 4861] = 1'b0;  wr_cycle[ 4861] = 1'b1;  addr_rom[ 4861]='h000011c0;  wr_data_rom[ 4861]='h000005b4;
    rd_cycle[ 4862] = 1'b1;  wr_cycle[ 4862] = 1'b0;  addr_rom[ 4862]='h00000228;  wr_data_rom[ 4862]='h00000000;
    rd_cycle[ 4863] = 1'b1;  wr_cycle[ 4863] = 1'b0;  addr_rom[ 4863]='h00001f18;  wr_data_rom[ 4863]='h00000000;
    rd_cycle[ 4864] = 1'b1;  wr_cycle[ 4864] = 1'b0;  addr_rom[ 4864]='h000015d8;  wr_data_rom[ 4864]='h00000000;
    rd_cycle[ 4865] = 1'b1;  wr_cycle[ 4865] = 1'b0;  addr_rom[ 4865]='h00000004;  wr_data_rom[ 4865]='h00000000;
    rd_cycle[ 4866] = 1'b0;  wr_cycle[ 4866] = 1'b1;  addr_rom[ 4866]='h00000ba8;  wr_data_rom[ 4866]='h00001d69;
    rd_cycle[ 4867] = 1'b0;  wr_cycle[ 4867] = 1'b1;  addr_rom[ 4867]='h00001580;  wr_data_rom[ 4867]='h00001815;
    rd_cycle[ 4868] = 1'b1;  wr_cycle[ 4868] = 1'b0;  addr_rom[ 4868]='h0000186c;  wr_data_rom[ 4868]='h00000000;
    rd_cycle[ 4869] = 1'b1;  wr_cycle[ 4869] = 1'b0;  addr_rom[ 4869]='h000003e8;  wr_data_rom[ 4869]='h00000000;
    rd_cycle[ 4870] = 1'b0;  wr_cycle[ 4870] = 1'b1;  addr_rom[ 4870]='h00001d10;  wr_data_rom[ 4870]='h000011b8;
    rd_cycle[ 4871] = 1'b0;  wr_cycle[ 4871] = 1'b1;  addr_rom[ 4871]='h00001d3c;  wr_data_rom[ 4871]='h00000529;
    rd_cycle[ 4872] = 1'b0;  wr_cycle[ 4872] = 1'b1;  addr_rom[ 4872]='h00000f18;  wr_data_rom[ 4872]='h000003b4;
    rd_cycle[ 4873] = 1'b1;  wr_cycle[ 4873] = 1'b0;  addr_rom[ 4873]='h0000132c;  wr_data_rom[ 4873]='h00000000;
    rd_cycle[ 4874] = 1'b0;  wr_cycle[ 4874] = 1'b1;  addr_rom[ 4874]='h00001bd0;  wr_data_rom[ 4874]='h00001c8b;
    rd_cycle[ 4875] = 1'b0;  wr_cycle[ 4875] = 1'b1;  addr_rom[ 4875]='h00001078;  wr_data_rom[ 4875]='h00000119;
    rd_cycle[ 4876] = 1'b0;  wr_cycle[ 4876] = 1'b1;  addr_rom[ 4876]='h0000180c;  wr_data_rom[ 4876]='h00000ab6;
    rd_cycle[ 4877] = 1'b1;  wr_cycle[ 4877] = 1'b0;  addr_rom[ 4877]='h000005b0;  wr_data_rom[ 4877]='h00000000;
    rd_cycle[ 4878] = 1'b1;  wr_cycle[ 4878] = 1'b0;  addr_rom[ 4878]='h00000698;  wr_data_rom[ 4878]='h00000000;
    rd_cycle[ 4879] = 1'b0;  wr_cycle[ 4879] = 1'b1;  addr_rom[ 4879]='h00000bd0;  wr_data_rom[ 4879]='h0000013f;
    rd_cycle[ 4880] = 1'b1;  wr_cycle[ 4880] = 1'b0;  addr_rom[ 4880]='h00000714;  wr_data_rom[ 4880]='h00000000;
    rd_cycle[ 4881] = 1'b1;  wr_cycle[ 4881] = 1'b0;  addr_rom[ 4881]='h0000177c;  wr_data_rom[ 4881]='h00000000;
    rd_cycle[ 4882] = 1'b1;  wr_cycle[ 4882] = 1'b0;  addr_rom[ 4882]='h0000171c;  wr_data_rom[ 4882]='h00000000;
    rd_cycle[ 4883] = 1'b1;  wr_cycle[ 4883] = 1'b0;  addr_rom[ 4883]='h000003dc;  wr_data_rom[ 4883]='h00000000;
    rd_cycle[ 4884] = 1'b0;  wr_cycle[ 4884] = 1'b1;  addr_rom[ 4884]='h00001ad4;  wr_data_rom[ 4884]='h000009f8;
    rd_cycle[ 4885] = 1'b0;  wr_cycle[ 4885] = 1'b1;  addr_rom[ 4885]='h000011c8;  wr_data_rom[ 4885]='h00000f65;
    rd_cycle[ 4886] = 1'b1;  wr_cycle[ 4886] = 1'b0;  addr_rom[ 4886]='h00000a20;  wr_data_rom[ 4886]='h00000000;
    rd_cycle[ 4887] = 1'b0;  wr_cycle[ 4887] = 1'b1;  addr_rom[ 4887]='h00000f58;  wr_data_rom[ 4887]='h00001164;
    rd_cycle[ 4888] = 1'b1;  wr_cycle[ 4888] = 1'b0;  addr_rom[ 4888]='h00000ccc;  wr_data_rom[ 4888]='h00000000;
    rd_cycle[ 4889] = 1'b0;  wr_cycle[ 4889] = 1'b1;  addr_rom[ 4889]='h00000ff8;  wr_data_rom[ 4889]='h00000df4;
    rd_cycle[ 4890] = 1'b1;  wr_cycle[ 4890] = 1'b0;  addr_rom[ 4890]='h00000010;  wr_data_rom[ 4890]='h00000000;
    rd_cycle[ 4891] = 1'b1;  wr_cycle[ 4891] = 1'b0;  addr_rom[ 4891]='h00000720;  wr_data_rom[ 4891]='h00000000;
    rd_cycle[ 4892] = 1'b0;  wr_cycle[ 4892] = 1'b1;  addr_rom[ 4892]='h000011d8;  wr_data_rom[ 4892]='h00000862;
    rd_cycle[ 4893] = 1'b0;  wr_cycle[ 4893] = 1'b1;  addr_rom[ 4893]='h00000128;  wr_data_rom[ 4893]='h00001a2e;
    rd_cycle[ 4894] = 1'b1;  wr_cycle[ 4894] = 1'b0;  addr_rom[ 4894]='h000001cc;  wr_data_rom[ 4894]='h00000000;
    rd_cycle[ 4895] = 1'b1;  wr_cycle[ 4895] = 1'b0;  addr_rom[ 4895]='h000005c4;  wr_data_rom[ 4895]='h00000000;
    rd_cycle[ 4896] = 1'b0;  wr_cycle[ 4896] = 1'b1;  addr_rom[ 4896]='h0000057c;  wr_data_rom[ 4896]='h00001581;
    rd_cycle[ 4897] = 1'b1;  wr_cycle[ 4897] = 1'b0;  addr_rom[ 4897]='h000002c8;  wr_data_rom[ 4897]='h00000000;
    rd_cycle[ 4898] = 1'b0;  wr_cycle[ 4898] = 1'b1;  addr_rom[ 4898]='h00001360;  wr_data_rom[ 4898]='h000011cc;
    rd_cycle[ 4899] = 1'b1;  wr_cycle[ 4899] = 1'b0;  addr_rom[ 4899]='h00001ed4;  wr_data_rom[ 4899]='h00000000;
    rd_cycle[ 4900] = 1'b1;  wr_cycle[ 4900] = 1'b0;  addr_rom[ 4900]='h00000c04;  wr_data_rom[ 4900]='h00000000;
    rd_cycle[ 4901] = 1'b0;  wr_cycle[ 4901] = 1'b1;  addr_rom[ 4901]='h000007e8;  wr_data_rom[ 4901]='h000001c4;
    rd_cycle[ 4902] = 1'b0;  wr_cycle[ 4902] = 1'b1;  addr_rom[ 4902]='h000011bc;  wr_data_rom[ 4902]='h0000157b;
    rd_cycle[ 4903] = 1'b1;  wr_cycle[ 4903] = 1'b0;  addr_rom[ 4903]='h00000320;  wr_data_rom[ 4903]='h00000000;
    rd_cycle[ 4904] = 1'b0;  wr_cycle[ 4904] = 1'b1;  addr_rom[ 4904]='h000003e0;  wr_data_rom[ 4904]='h00000578;
    rd_cycle[ 4905] = 1'b1;  wr_cycle[ 4905] = 1'b0;  addr_rom[ 4905]='h0000189c;  wr_data_rom[ 4905]='h00000000;
    rd_cycle[ 4906] = 1'b0;  wr_cycle[ 4906] = 1'b1;  addr_rom[ 4906]='h00001134;  wr_data_rom[ 4906]='h00001b44;
    rd_cycle[ 4907] = 1'b0;  wr_cycle[ 4907] = 1'b1;  addr_rom[ 4907]='h000004c0;  wr_data_rom[ 4907]='h00000f02;
    rd_cycle[ 4908] = 1'b1;  wr_cycle[ 4908] = 1'b0;  addr_rom[ 4908]='h00000708;  wr_data_rom[ 4908]='h00000000;
    rd_cycle[ 4909] = 1'b0;  wr_cycle[ 4909] = 1'b1;  addr_rom[ 4909]='h00001ac0;  wr_data_rom[ 4909]='h00001c0e;
    rd_cycle[ 4910] = 1'b0;  wr_cycle[ 4910] = 1'b1;  addr_rom[ 4910]='h00001d70;  wr_data_rom[ 4910]='h00000508;
    rd_cycle[ 4911] = 1'b0;  wr_cycle[ 4911] = 1'b1;  addr_rom[ 4911]='h0000100c;  wr_data_rom[ 4911]='h00000ccb;
    rd_cycle[ 4912] = 1'b0;  wr_cycle[ 4912] = 1'b1;  addr_rom[ 4912]='h00000ce8;  wr_data_rom[ 4912]='h00000bf3;
    rd_cycle[ 4913] = 1'b1;  wr_cycle[ 4913] = 1'b0;  addr_rom[ 4913]='h00000344;  wr_data_rom[ 4913]='h00000000;
    rd_cycle[ 4914] = 1'b1;  wr_cycle[ 4914] = 1'b0;  addr_rom[ 4914]='h00001abc;  wr_data_rom[ 4914]='h00000000;
    rd_cycle[ 4915] = 1'b1;  wr_cycle[ 4915] = 1'b0;  addr_rom[ 4915]='h00000afc;  wr_data_rom[ 4915]='h00000000;
    rd_cycle[ 4916] = 1'b1;  wr_cycle[ 4916] = 1'b0;  addr_rom[ 4916]='h00000ab4;  wr_data_rom[ 4916]='h00000000;
    rd_cycle[ 4917] = 1'b0;  wr_cycle[ 4917] = 1'b1;  addr_rom[ 4917]='h000001bc;  wr_data_rom[ 4917]='h0000023d;
    rd_cycle[ 4918] = 1'b1;  wr_cycle[ 4918] = 1'b0;  addr_rom[ 4918]='h000005e4;  wr_data_rom[ 4918]='h00000000;
    rd_cycle[ 4919] = 1'b1;  wr_cycle[ 4919] = 1'b0;  addr_rom[ 4919]='h00001404;  wr_data_rom[ 4919]='h00000000;
    rd_cycle[ 4920] = 1'b0;  wr_cycle[ 4920] = 1'b1;  addr_rom[ 4920]='h00000960;  wr_data_rom[ 4920]='h000013f9;
    rd_cycle[ 4921] = 1'b0;  wr_cycle[ 4921] = 1'b1;  addr_rom[ 4921]='h00000ae0;  wr_data_rom[ 4921]='h000007fb;
    rd_cycle[ 4922] = 1'b0;  wr_cycle[ 4922] = 1'b1;  addr_rom[ 4922]='h00001e1c;  wr_data_rom[ 4922]='h00000559;
    rd_cycle[ 4923] = 1'b1;  wr_cycle[ 4923] = 1'b0;  addr_rom[ 4923]='h00001aa0;  wr_data_rom[ 4923]='h00000000;
    rd_cycle[ 4924] = 1'b0;  wr_cycle[ 4924] = 1'b1;  addr_rom[ 4924]='h00000d24;  wr_data_rom[ 4924]='h000003cf;
    rd_cycle[ 4925] = 1'b0;  wr_cycle[ 4925] = 1'b1;  addr_rom[ 4925]='h00000644;  wr_data_rom[ 4925]='h000011fb;
    rd_cycle[ 4926] = 1'b0;  wr_cycle[ 4926] = 1'b1;  addr_rom[ 4926]='h00001b80;  wr_data_rom[ 4926]='h00001671;
    rd_cycle[ 4927] = 1'b1;  wr_cycle[ 4927] = 1'b0;  addr_rom[ 4927]='h000011fc;  wr_data_rom[ 4927]='h00000000;
    rd_cycle[ 4928] = 1'b1;  wr_cycle[ 4928] = 1'b0;  addr_rom[ 4928]='h00001410;  wr_data_rom[ 4928]='h00000000;
    rd_cycle[ 4929] = 1'b1;  wr_cycle[ 4929] = 1'b0;  addr_rom[ 4929]='h00001814;  wr_data_rom[ 4929]='h00000000;
    rd_cycle[ 4930] = 1'b0;  wr_cycle[ 4930] = 1'b1;  addr_rom[ 4930]='h0000068c;  wr_data_rom[ 4930]='h00000b0d;
    rd_cycle[ 4931] = 1'b0;  wr_cycle[ 4931] = 1'b1;  addr_rom[ 4931]='h00001b68;  wr_data_rom[ 4931]='h000005c1;
    rd_cycle[ 4932] = 1'b1;  wr_cycle[ 4932] = 1'b0;  addr_rom[ 4932]='h00000344;  wr_data_rom[ 4932]='h00000000;
    rd_cycle[ 4933] = 1'b1;  wr_cycle[ 4933] = 1'b0;  addr_rom[ 4933]='h00001c6c;  wr_data_rom[ 4933]='h00000000;
    rd_cycle[ 4934] = 1'b0;  wr_cycle[ 4934] = 1'b1;  addr_rom[ 4934]='h00001190;  wr_data_rom[ 4934]='h00001a11;
    rd_cycle[ 4935] = 1'b1;  wr_cycle[ 4935] = 1'b0;  addr_rom[ 4935]='h000012cc;  wr_data_rom[ 4935]='h00000000;
    rd_cycle[ 4936] = 1'b0;  wr_cycle[ 4936] = 1'b1;  addr_rom[ 4936]='h00000090;  wr_data_rom[ 4936]='h00001425;
    rd_cycle[ 4937] = 1'b1;  wr_cycle[ 4937] = 1'b0;  addr_rom[ 4937]='h00000518;  wr_data_rom[ 4937]='h00000000;
    rd_cycle[ 4938] = 1'b1;  wr_cycle[ 4938] = 1'b0;  addr_rom[ 4938]='h000014b0;  wr_data_rom[ 4938]='h00000000;
    rd_cycle[ 4939] = 1'b0;  wr_cycle[ 4939] = 1'b1;  addr_rom[ 4939]='h00000a50;  wr_data_rom[ 4939]='h00001183;
    rd_cycle[ 4940] = 1'b0;  wr_cycle[ 4940] = 1'b1;  addr_rom[ 4940]='h00001428;  wr_data_rom[ 4940]='h00001864;
    rd_cycle[ 4941] = 1'b0;  wr_cycle[ 4941] = 1'b1;  addr_rom[ 4941]='h000008a0;  wr_data_rom[ 4941]='h00000663;
    rd_cycle[ 4942] = 1'b1;  wr_cycle[ 4942] = 1'b0;  addr_rom[ 4942]='h00001268;  wr_data_rom[ 4942]='h00000000;
    rd_cycle[ 4943] = 1'b1;  wr_cycle[ 4943] = 1'b0;  addr_rom[ 4943]='h00001d98;  wr_data_rom[ 4943]='h00000000;
    rd_cycle[ 4944] = 1'b1;  wr_cycle[ 4944] = 1'b0;  addr_rom[ 4944]='h00001d3c;  wr_data_rom[ 4944]='h00000000;
    rd_cycle[ 4945] = 1'b0;  wr_cycle[ 4945] = 1'b1;  addr_rom[ 4945]='h00001348;  wr_data_rom[ 4945]='h0000169d;
    rd_cycle[ 4946] = 1'b0;  wr_cycle[ 4946] = 1'b1;  addr_rom[ 4946]='h00001d10;  wr_data_rom[ 4946]='h00001864;
    rd_cycle[ 4947] = 1'b1;  wr_cycle[ 4947] = 1'b0;  addr_rom[ 4947]='h000009d0;  wr_data_rom[ 4947]='h00000000;
    rd_cycle[ 4948] = 1'b0;  wr_cycle[ 4948] = 1'b1;  addr_rom[ 4948]='h000013ec;  wr_data_rom[ 4948]='h0000174d;
    rd_cycle[ 4949] = 1'b0;  wr_cycle[ 4949] = 1'b1;  addr_rom[ 4949]='h0000143c;  wr_data_rom[ 4949]='h000004aa;
    rd_cycle[ 4950] = 1'b1;  wr_cycle[ 4950] = 1'b0;  addr_rom[ 4950]='h00000558;  wr_data_rom[ 4950]='h00000000;
    rd_cycle[ 4951] = 1'b1;  wr_cycle[ 4951] = 1'b0;  addr_rom[ 4951]='h00000124;  wr_data_rom[ 4951]='h00000000;
    rd_cycle[ 4952] = 1'b1;  wr_cycle[ 4952] = 1'b0;  addr_rom[ 4952]='h0000165c;  wr_data_rom[ 4952]='h00000000;
    rd_cycle[ 4953] = 1'b1;  wr_cycle[ 4953] = 1'b0;  addr_rom[ 4953]='h000004a4;  wr_data_rom[ 4953]='h00000000;
    rd_cycle[ 4954] = 1'b0;  wr_cycle[ 4954] = 1'b1;  addr_rom[ 4954]='h00000d84;  wr_data_rom[ 4954]='h00000e79;
    rd_cycle[ 4955] = 1'b0;  wr_cycle[ 4955] = 1'b1;  addr_rom[ 4955]='h00000fd0;  wr_data_rom[ 4955]='h000011f5;
    rd_cycle[ 4956] = 1'b1;  wr_cycle[ 4956] = 1'b0;  addr_rom[ 4956]='h00000848;  wr_data_rom[ 4956]='h00000000;
    rd_cycle[ 4957] = 1'b0;  wr_cycle[ 4957] = 1'b1;  addr_rom[ 4957]='h00000f78;  wr_data_rom[ 4957]='h00000b96;
    rd_cycle[ 4958] = 1'b1;  wr_cycle[ 4958] = 1'b0;  addr_rom[ 4958]='h00000638;  wr_data_rom[ 4958]='h00000000;
    rd_cycle[ 4959] = 1'b0;  wr_cycle[ 4959] = 1'b1;  addr_rom[ 4959]='h00001d78;  wr_data_rom[ 4959]='h00001815;
    rd_cycle[ 4960] = 1'b1;  wr_cycle[ 4960] = 1'b0;  addr_rom[ 4960]='h000008b8;  wr_data_rom[ 4960]='h00000000;
    rd_cycle[ 4961] = 1'b0;  wr_cycle[ 4961] = 1'b1;  addr_rom[ 4961]='h000014c0;  wr_data_rom[ 4961]='h000013d8;
    rd_cycle[ 4962] = 1'b0;  wr_cycle[ 4962] = 1'b1;  addr_rom[ 4962]='h00001d7c;  wr_data_rom[ 4962]='h00000a19;
    rd_cycle[ 4963] = 1'b0;  wr_cycle[ 4963] = 1'b1;  addr_rom[ 4963]='h00001a40;  wr_data_rom[ 4963]='h00001776;
    rd_cycle[ 4964] = 1'b0;  wr_cycle[ 4964] = 1'b1;  addr_rom[ 4964]='h00001974;  wr_data_rom[ 4964]='h0000083e;
    rd_cycle[ 4965] = 1'b0;  wr_cycle[ 4965] = 1'b1;  addr_rom[ 4965]='h00001c9c;  wr_data_rom[ 4965]='h00000c4b;
    rd_cycle[ 4966] = 1'b1;  wr_cycle[ 4966] = 1'b0;  addr_rom[ 4966]='h0000041c;  wr_data_rom[ 4966]='h00000000;
    rd_cycle[ 4967] = 1'b0;  wr_cycle[ 4967] = 1'b1;  addr_rom[ 4967]='h00000274;  wr_data_rom[ 4967]='h000008ba;
    rd_cycle[ 4968] = 1'b1;  wr_cycle[ 4968] = 1'b0;  addr_rom[ 4968]='h00001c10;  wr_data_rom[ 4968]='h00000000;
    rd_cycle[ 4969] = 1'b1;  wr_cycle[ 4969] = 1'b0;  addr_rom[ 4969]='h00001324;  wr_data_rom[ 4969]='h00000000;
    rd_cycle[ 4970] = 1'b0;  wr_cycle[ 4970] = 1'b1;  addr_rom[ 4970]='h00001cb8;  wr_data_rom[ 4970]='h000008df;
    rd_cycle[ 4971] = 1'b1;  wr_cycle[ 4971] = 1'b0;  addr_rom[ 4971]='h00000bb4;  wr_data_rom[ 4971]='h00000000;
    rd_cycle[ 4972] = 1'b1;  wr_cycle[ 4972] = 1'b0;  addr_rom[ 4972]='h00001724;  wr_data_rom[ 4972]='h00000000;
    rd_cycle[ 4973] = 1'b0;  wr_cycle[ 4973] = 1'b1;  addr_rom[ 4973]='h000006c4;  wr_data_rom[ 4973]='h00001bd3;
    rd_cycle[ 4974] = 1'b1;  wr_cycle[ 4974] = 1'b0;  addr_rom[ 4974]='h000009dc;  wr_data_rom[ 4974]='h00000000;
    rd_cycle[ 4975] = 1'b1;  wr_cycle[ 4975] = 1'b0;  addr_rom[ 4975]='h00001524;  wr_data_rom[ 4975]='h00000000;
    rd_cycle[ 4976] = 1'b0;  wr_cycle[ 4976] = 1'b1;  addr_rom[ 4976]='h0000154c;  wr_data_rom[ 4976]='h00000e8d;
    rd_cycle[ 4977] = 1'b0;  wr_cycle[ 4977] = 1'b1;  addr_rom[ 4977]='h00001a78;  wr_data_rom[ 4977]='h00000284;
    rd_cycle[ 4978] = 1'b1;  wr_cycle[ 4978] = 1'b0;  addr_rom[ 4978]='h000000fc;  wr_data_rom[ 4978]='h00000000;
    rd_cycle[ 4979] = 1'b0;  wr_cycle[ 4979] = 1'b1;  addr_rom[ 4979]='h00001060;  wr_data_rom[ 4979]='h00000d72;
    rd_cycle[ 4980] = 1'b1;  wr_cycle[ 4980] = 1'b0;  addr_rom[ 4980]='h000012c8;  wr_data_rom[ 4980]='h00000000;
    rd_cycle[ 4981] = 1'b1;  wr_cycle[ 4981] = 1'b0;  addr_rom[ 4981]='h00001a9c;  wr_data_rom[ 4981]='h00000000;
    rd_cycle[ 4982] = 1'b1;  wr_cycle[ 4982] = 1'b0;  addr_rom[ 4982]='h000012a4;  wr_data_rom[ 4982]='h00000000;
    rd_cycle[ 4983] = 1'b0;  wr_cycle[ 4983] = 1'b1;  addr_rom[ 4983]='h0000135c;  wr_data_rom[ 4983]='h00000e3c;
    rd_cycle[ 4984] = 1'b1;  wr_cycle[ 4984] = 1'b0;  addr_rom[ 4984]='h000016dc;  wr_data_rom[ 4984]='h00000000;
    rd_cycle[ 4985] = 1'b0;  wr_cycle[ 4985] = 1'b1;  addr_rom[ 4985]='h00001af0;  wr_data_rom[ 4985]='h00001702;
    rd_cycle[ 4986] = 1'b1;  wr_cycle[ 4986] = 1'b0;  addr_rom[ 4986]='h00001140;  wr_data_rom[ 4986]='h00000000;
    rd_cycle[ 4987] = 1'b1;  wr_cycle[ 4987] = 1'b0;  addr_rom[ 4987]='h000007e4;  wr_data_rom[ 4987]='h00000000;
    rd_cycle[ 4988] = 1'b1;  wr_cycle[ 4988] = 1'b0;  addr_rom[ 4988]='h000000bc;  wr_data_rom[ 4988]='h00000000;
    rd_cycle[ 4989] = 1'b1;  wr_cycle[ 4989] = 1'b0;  addr_rom[ 4989]='h00001e40;  wr_data_rom[ 4989]='h00000000;
    rd_cycle[ 4990] = 1'b0;  wr_cycle[ 4990] = 1'b1;  addr_rom[ 4990]='h000009b4;  wr_data_rom[ 4990]='h0000119b;
    rd_cycle[ 4991] = 1'b1;  wr_cycle[ 4991] = 1'b0;  addr_rom[ 4991]='h00000674;  wr_data_rom[ 4991]='h00000000;
    rd_cycle[ 4992] = 1'b0;  wr_cycle[ 4992] = 1'b1;  addr_rom[ 4992]='h00000b40;  wr_data_rom[ 4992]='h00000740;
    rd_cycle[ 4993] = 1'b0;  wr_cycle[ 4993] = 1'b1;  addr_rom[ 4993]='h000011c4;  wr_data_rom[ 4993]='h00000a25;
    rd_cycle[ 4994] = 1'b0;  wr_cycle[ 4994] = 1'b1;  addr_rom[ 4994]='h0000178c;  wr_data_rom[ 4994]='h00001d7f;
    rd_cycle[ 4995] = 1'b0;  wr_cycle[ 4995] = 1'b1;  addr_rom[ 4995]='h00001a10;  wr_data_rom[ 4995]='h000009a4;
    rd_cycle[ 4996] = 1'b0;  wr_cycle[ 4996] = 1'b1;  addr_rom[ 4996]='h000019e4;  wr_data_rom[ 4996]='h000010e8;
    rd_cycle[ 4997] = 1'b0;  wr_cycle[ 4997] = 1'b1;  addr_rom[ 4997]='h00000518;  wr_data_rom[ 4997]='h00000b2f;
    rd_cycle[ 4998] = 1'b0;  wr_cycle[ 4998] = 1'b1;  addr_rom[ 4998]='h000001dc;  wr_data_rom[ 4998]='h0000060f;
    rd_cycle[ 4999] = 1'b1;  wr_cycle[ 4999] = 1'b0;  addr_rom[ 4999]='h00000e94;  wr_data_rom[ 4999]='h00000000;
    rd_cycle[ 5000] = 1'b0;  wr_cycle[ 5000] = 1'b1;  addr_rom[ 5000]='h00001b9c;  wr_data_rom[ 5000]='h00001e8f;
    rd_cycle[ 5001] = 1'b1;  wr_cycle[ 5001] = 1'b0;  addr_rom[ 5001]='h00000054;  wr_data_rom[ 5001]='h00000000;
    rd_cycle[ 5002] = 1'b1;  wr_cycle[ 5002] = 1'b0;  addr_rom[ 5002]='h00001228;  wr_data_rom[ 5002]='h00000000;
    rd_cycle[ 5003] = 1'b1;  wr_cycle[ 5003] = 1'b0;  addr_rom[ 5003]='h000012ec;  wr_data_rom[ 5003]='h00000000;
    rd_cycle[ 5004] = 1'b0;  wr_cycle[ 5004] = 1'b1;  addr_rom[ 5004]='h00000dc0;  wr_data_rom[ 5004]='h000003a9;
    rd_cycle[ 5005] = 1'b1;  wr_cycle[ 5005] = 1'b0;  addr_rom[ 5005]='h00000f9c;  wr_data_rom[ 5005]='h00000000;
    rd_cycle[ 5006] = 1'b0;  wr_cycle[ 5006] = 1'b1;  addr_rom[ 5006]='h00000580;  wr_data_rom[ 5006]='h0000105b;
    rd_cycle[ 5007] = 1'b0;  wr_cycle[ 5007] = 1'b1;  addr_rom[ 5007]='h000012f4;  wr_data_rom[ 5007]='h00000cff;
    rd_cycle[ 5008] = 1'b0;  wr_cycle[ 5008] = 1'b1;  addr_rom[ 5008]='h00001284;  wr_data_rom[ 5008]='h00000301;
    rd_cycle[ 5009] = 1'b0;  wr_cycle[ 5009] = 1'b1;  addr_rom[ 5009]='h000006c0;  wr_data_rom[ 5009]='h00001783;
    rd_cycle[ 5010] = 1'b0;  wr_cycle[ 5010] = 1'b1;  addr_rom[ 5010]='h000019c4;  wr_data_rom[ 5010]='h0000063d;
    rd_cycle[ 5011] = 1'b0;  wr_cycle[ 5011] = 1'b1;  addr_rom[ 5011]='h0000015c;  wr_data_rom[ 5011]='h000010ca;
    rd_cycle[ 5012] = 1'b0;  wr_cycle[ 5012] = 1'b1;  addr_rom[ 5012]='h000014d4;  wr_data_rom[ 5012]='h00000ade;
    rd_cycle[ 5013] = 1'b1;  wr_cycle[ 5013] = 1'b0;  addr_rom[ 5013]='h00001ee8;  wr_data_rom[ 5013]='h00000000;
    rd_cycle[ 5014] = 1'b0;  wr_cycle[ 5014] = 1'b1;  addr_rom[ 5014]='h0000030c;  wr_data_rom[ 5014]='h00000aff;
    rd_cycle[ 5015] = 1'b1;  wr_cycle[ 5015] = 1'b0;  addr_rom[ 5015]='h00001268;  wr_data_rom[ 5015]='h00000000;
    rd_cycle[ 5016] = 1'b1;  wr_cycle[ 5016] = 1'b0;  addr_rom[ 5016]='h000018ac;  wr_data_rom[ 5016]='h00000000;
    rd_cycle[ 5017] = 1'b1;  wr_cycle[ 5017] = 1'b0;  addr_rom[ 5017]='h0000125c;  wr_data_rom[ 5017]='h00000000;
    rd_cycle[ 5018] = 1'b1;  wr_cycle[ 5018] = 1'b0;  addr_rom[ 5018]='h0000081c;  wr_data_rom[ 5018]='h00000000;
    rd_cycle[ 5019] = 1'b0;  wr_cycle[ 5019] = 1'b1;  addr_rom[ 5019]='h000017ec;  wr_data_rom[ 5019]='h0000137b;
    rd_cycle[ 5020] = 1'b0;  wr_cycle[ 5020] = 1'b1;  addr_rom[ 5020]='h000012fc;  wr_data_rom[ 5020]='h00000732;
    rd_cycle[ 5021] = 1'b1;  wr_cycle[ 5021] = 1'b0;  addr_rom[ 5021]='h00001c28;  wr_data_rom[ 5021]='h00000000;
    rd_cycle[ 5022] = 1'b1;  wr_cycle[ 5022] = 1'b0;  addr_rom[ 5022]='h00000c3c;  wr_data_rom[ 5022]='h00000000;
    rd_cycle[ 5023] = 1'b1;  wr_cycle[ 5023] = 1'b0;  addr_rom[ 5023]='h00001a54;  wr_data_rom[ 5023]='h00000000;
    rd_cycle[ 5024] = 1'b0;  wr_cycle[ 5024] = 1'b1;  addr_rom[ 5024]='h00001280;  wr_data_rom[ 5024]='h000018cd;
    rd_cycle[ 5025] = 1'b0;  wr_cycle[ 5025] = 1'b1;  addr_rom[ 5025]='h0000039c;  wr_data_rom[ 5025]='h000002c4;
    rd_cycle[ 5026] = 1'b1;  wr_cycle[ 5026] = 1'b0;  addr_rom[ 5026]='h000006b8;  wr_data_rom[ 5026]='h00000000;
    rd_cycle[ 5027] = 1'b1;  wr_cycle[ 5027] = 1'b0;  addr_rom[ 5027]='h00000460;  wr_data_rom[ 5027]='h00000000;
    rd_cycle[ 5028] = 1'b0;  wr_cycle[ 5028] = 1'b1;  addr_rom[ 5028]='h00001858;  wr_data_rom[ 5028]='h000006f4;
    rd_cycle[ 5029] = 1'b1;  wr_cycle[ 5029] = 1'b0;  addr_rom[ 5029]='h00001690;  wr_data_rom[ 5029]='h00000000;
    rd_cycle[ 5030] = 1'b0;  wr_cycle[ 5030] = 1'b1;  addr_rom[ 5030]='h000014d4;  wr_data_rom[ 5030]='h000016bc;
    rd_cycle[ 5031] = 1'b1;  wr_cycle[ 5031] = 1'b0;  addr_rom[ 5031]='h000009dc;  wr_data_rom[ 5031]='h00000000;
    rd_cycle[ 5032] = 1'b0;  wr_cycle[ 5032] = 1'b1;  addr_rom[ 5032]='h000005c4;  wr_data_rom[ 5032]='h00000d8f;
    rd_cycle[ 5033] = 1'b0;  wr_cycle[ 5033] = 1'b1;  addr_rom[ 5033]='h000004b0;  wr_data_rom[ 5033]='h00001d05;
    rd_cycle[ 5034] = 1'b0;  wr_cycle[ 5034] = 1'b1;  addr_rom[ 5034]='h00000e0c;  wr_data_rom[ 5034]='h00001189;
    rd_cycle[ 5035] = 1'b1;  wr_cycle[ 5035] = 1'b0;  addr_rom[ 5035]='h000011fc;  wr_data_rom[ 5035]='h00000000;
    rd_cycle[ 5036] = 1'b1;  wr_cycle[ 5036] = 1'b0;  addr_rom[ 5036]='h00001140;  wr_data_rom[ 5036]='h00000000;
    rd_cycle[ 5037] = 1'b1;  wr_cycle[ 5037] = 1'b0;  addr_rom[ 5037]='h000005ec;  wr_data_rom[ 5037]='h00000000;
    rd_cycle[ 5038] = 1'b0;  wr_cycle[ 5038] = 1'b1;  addr_rom[ 5038]='h00000a60;  wr_data_rom[ 5038]='h00001b33;
    rd_cycle[ 5039] = 1'b1;  wr_cycle[ 5039] = 1'b0;  addr_rom[ 5039]='h00001c8c;  wr_data_rom[ 5039]='h00000000;
    rd_cycle[ 5040] = 1'b0;  wr_cycle[ 5040] = 1'b1;  addr_rom[ 5040]='h000011dc;  wr_data_rom[ 5040]='h00000561;
    rd_cycle[ 5041] = 1'b0;  wr_cycle[ 5041] = 1'b1;  addr_rom[ 5041]='h000014e0;  wr_data_rom[ 5041]='h00001d2c;
    rd_cycle[ 5042] = 1'b1;  wr_cycle[ 5042] = 1'b0;  addr_rom[ 5042]='h00000abc;  wr_data_rom[ 5042]='h00000000;
    rd_cycle[ 5043] = 1'b1;  wr_cycle[ 5043] = 1'b0;  addr_rom[ 5043]='h000006c0;  wr_data_rom[ 5043]='h00000000;
    rd_cycle[ 5044] = 1'b1;  wr_cycle[ 5044] = 1'b0;  addr_rom[ 5044]='h00001cf4;  wr_data_rom[ 5044]='h00000000;
    rd_cycle[ 5045] = 1'b1;  wr_cycle[ 5045] = 1'b0;  addr_rom[ 5045]='h00000e48;  wr_data_rom[ 5045]='h00000000;
    rd_cycle[ 5046] = 1'b1;  wr_cycle[ 5046] = 1'b0;  addr_rom[ 5046]='h00001334;  wr_data_rom[ 5046]='h00000000;
    rd_cycle[ 5047] = 1'b0;  wr_cycle[ 5047] = 1'b1;  addr_rom[ 5047]='h00001194;  wr_data_rom[ 5047]='h000005ac;
    rd_cycle[ 5048] = 1'b0;  wr_cycle[ 5048] = 1'b1;  addr_rom[ 5048]='h000016e4;  wr_data_rom[ 5048]='h0000039f;
    rd_cycle[ 5049] = 1'b0;  wr_cycle[ 5049] = 1'b1;  addr_rom[ 5049]='h000007fc;  wr_data_rom[ 5049]='h00001327;
    rd_cycle[ 5050] = 1'b0;  wr_cycle[ 5050] = 1'b1;  addr_rom[ 5050]='h00000f30;  wr_data_rom[ 5050]='h00000a3a;
    rd_cycle[ 5051] = 1'b1;  wr_cycle[ 5051] = 1'b0;  addr_rom[ 5051]='h00000aac;  wr_data_rom[ 5051]='h00000000;
    rd_cycle[ 5052] = 1'b0;  wr_cycle[ 5052] = 1'b1;  addr_rom[ 5052]='h00000b88;  wr_data_rom[ 5052]='h000012d3;
    rd_cycle[ 5053] = 1'b1;  wr_cycle[ 5053] = 1'b0;  addr_rom[ 5053]='h00000e5c;  wr_data_rom[ 5053]='h00000000;
    rd_cycle[ 5054] = 1'b0;  wr_cycle[ 5054] = 1'b1;  addr_rom[ 5054]='h00001a90;  wr_data_rom[ 5054]='h000001e9;
    rd_cycle[ 5055] = 1'b0;  wr_cycle[ 5055] = 1'b1;  addr_rom[ 5055]='h000008a0;  wr_data_rom[ 5055]='h00000b88;
    rd_cycle[ 5056] = 1'b0;  wr_cycle[ 5056] = 1'b1;  addr_rom[ 5056]='h00000a3c;  wr_data_rom[ 5056]='h000015f9;
    rd_cycle[ 5057] = 1'b0;  wr_cycle[ 5057] = 1'b1;  addr_rom[ 5057]='h000007cc;  wr_data_rom[ 5057]='h000015c4;
    rd_cycle[ 5058] = 1'b1;  wr_cycle[ 5058] = 1'b0;  addr_rom[ 5058]='h000004d4;  wr_data_rom[ 5058]='h00000000;
    rd_cycle[ 5059] = 1'b1;  wr_cycle[ 5059] = 1'b0;  addr_rom[ 5059]='h00001128;  wr_data_rom[ 5059]='h00000000;
    rd_cycle[ 5060] = 1'b1;  wr_cycle[ 5060] = 1'b0;  addr_rom[ 5060]='h00001f30;  wr_data_rom[ 5060]='h00000000;
    rd_cycle[ 5061] = 1'b0;  wr_cycle[ 5061] = 1'b1;  addr_rom[ 5061]='h000015e0;  wr_data_rom[ 5061]='h000014ce;
    rd_cycle[ 5062] = 1'b1;  wr_cycle[ 5062] = 1'b0;  addr_rom[ 5062]='h0000133c;  wr_data_rom[ 5062]='h00000000;
    rd_cycle[ 5063] = 1'b0;  wr_cycle[ 5063] = 1'b1;  addr_rom[ 5063]='h000008d0;  wr_data_rom[ 5063]='h00000a59;
    rd_cycle[ 5064] = 1'b0;  wr_cycle[ 5064] = 1'b1;  addr_rom[ 5064]='h00001bd8;  wr_data_rom[ 5064]='h00000d62;
    rd_cycle[ 5065] = 1'b1;  wr_cycle[ 5065] = 1'b0;  addr_rom[ 5065]='h00001ce4;  wr_data_rom[ 5065]='h00000000;
    rd_cycle[ 5066] = 1'b0;  wr_cycle[ 5066] = 1'b1;  addr_rom[ 5066]='h00001914;  wr_data_rom[ 5066]='h00001ebf;
    rd_cycle[ 5067] = 1'b0;  wr_cycle[ 5067] = 1'b1;  addr_rom[ 5067]='h000008c4;  wr_data_rom[ 5067]='h00001483;
    rd_cycle[ 5068] = 1'b1;  wr_cycle[ 5068] = 1'b0;  addr_rom[ 5068]='h0000152c;  wr_data_rom[ 5068]='h00000000;
    rd_cycle[ 5069] = 1'b1;  wr_cycle[ 5069] = 1'b0;  addr_rom[ 5069]='h00000110;  wr_data_rom[ 5069]='h00000000;
    rd_cycle[ 5070] = 1'b0;  wr_cycle[ 5070] = 1'b1;  addr_rom[ 5070]='h00001114;  wr_data_rom[ 5070]='h0000098d;
    rd_cycle[ 5071] = 1'b0;  wr_cycle[ 5071] = 1'b1;  addr_rom[ 5071]='h00001700;  wr_data_rom[ 5071]='h0000095f;
    rd_cycle[ 5072] = 1'b1;  wr_cycle[ 5072] = 1'b0;  addr_rom[ 5072]='h00001a60;  wr_data_rom[ 5072]='h00000000;
    rd_cycle[ 5073] = 1'b0;  wr_cycle[ 5073] = 1'b1;  addr_rom[ 5073]='h0000052c;  wr_data_rom[ 5073]='h0000173c;
    rd_cycle[ 5074] = 1'b1;  wr_cycle[ 5074] = 1'b0;  addr_rom[ 5074]='h000000c4;  wr_data_rom[ 5074]='h00000000;
    rd_cycle[ 5075] = 1'b1;  wr_cycle[ 5075] = 1'b0;  addr_rom[ 5075]='h00001d6c;  wr_data_rom[ 5075]='h00000000;
    rd_cycle[ 5076] = 1'b1;  wr_cycle[ 5076] = 1'b0;  addr_rom[ 5076]='h000006ac;  wr_data_rom[ 5076]='h00000000;
    rd_cycle[ 5077] = 1'b1;  wr_cycle[ 5077] = 1'b0;  addr_rom[ 5077]='h00001920;  wr_data_rom[ 5077]='h00000000;
    rd_cycle[ 5078] = 1'b0;  wr_cycle[ 5078] = 1'b1;  addr_rom[ 5078]='h00001e58;  wr_data_rom[ 5078]='h00001de9;
    rd_cycle[ 5079] = 1'b0;  wr_cycle[ 5079] = 1'b1;  addr_rom[ 5079]='h00000d2c;  wr_data_rom[ 5079]='h00000a2d;
    rd_cycle[ 5080] = 1'b0;  wr_cycle[ 5080] = 1'b1;  addr_rom[ 5080]='h00001590;  wr_data_rom[ 5080]='h0000113d;
    rd_cycle[ 5081] = 1'b0;  wr_cycle[ 5081] = 1'b1;  addr_rom[ 5081]='h00001794;  wr_data_rom[ 5081]='h00000810;
    rd_cycle[ 5082] = 1'b1;  wr_cycle[ 5082] = 1'b0;  addr_rom[ 5082]='h00001ad8;  wr_data_rom[ 5082]='h00000000;
    rd_cycle[ 5083] = 1'b1;  wr_cycle[ 5083] = 1'b0;  addr_rom[ 5083]='h000008c4;  wr_data_rom[ 5083]='h00000000;
    rd_cycle[ 5084] = 1'b1;  wr_cycle[ 5084] = 1'b0;  addr_rom[ 5084]='h00000320;  wr_data_rom[ 5084]='h00000000;
    rd_cycle[ 5085] = 1'b1;  wr_cycle[ 5085] = 1'b0;  addr_rom[ 5085]='h000005a0;  wr_data_rom[ 5085]='h00000000;
    rd_cycle[ 5086] = 1'b1;  wr_cycle[ 5086] = 1'b0;  addr_rom[ 5086]='h00001680;  wr_data_rom[ 5086]='h00000000;
    rd_cycle[ 5087] = 1'b1;  wr_cycle[ 5087] = 1'b0;  addr_rom[ 5087]='h00001214;  wr_data_rom[ 5087]='h00000000;
    rd_cycle[ 5088] = 1'b0;  wr_cycle[ 5088] = 1'b1;  addr_rom[ 5088]='h00001260;  wr_data_rom[ 5088]='h0000068b;
    rd_cycle[ 5089] = 1'b0;  wr_cycle[ 5089] = 1'b1;  addr_rom[ 5089]='h0000092c;  wr_data_rom[ 5089]='h00000fa5;
    rd_cycle[ 5090] = 1'b0;  wr_cycle[ 5090] = 1'b1;  addr_rom[ 5090]='h00001c04;  wr_data_rom[ 5090]='h000018fe;
    rd_cycle[ 5091] = 1'b0;  wr_cycle[ 5091] = 1'b1;  addr_rom[ 5091]='h00000450;  wr_data_rom[ 5091]='h00001d1c;
    rd_cycle[ 5092] = 1'b1;  wr_cycle[ 5092] = 1'b0;  addr_rom[ 5092]='h00000de0;  wr_data_rom[ 5092]='h00000000;
    rd_cycle[ 5093] = 1'b1;  wr_cycle[ 5093] = 1'b0;  addr_rom[ 5093]='h00001944;  wr_data_rom[ 5093]='h00000000;
    rd_cycle[ 5094] = 1'b0;  wr_cycle[ 5094] = 1'b1;  addr_rom[ 5094]='h0000045c;  wr_data_rom[ 5094]='h00001be4;
    rd_cycle[ 5095] = 1'b1;  wr_cycle[ 5095] = 1'b0;  addr_rom[ 5095]='h0000095c;  wr_data_rom[ 5095]='h00000000;
    rd_cycle[ 5096] = 1'b0;  wr_cycle[ 5096] = 1'b1;  addr_rom[ 5096]='h00000f2c;  wr_data_rom[ 5096]='h00000810;
    rd_cycle[ 5097] = 1'b0;  wr_cycle[ 5097] = 1'b1;  addr_rom[ 5097]='h00000184;  wr_data_rom[ 5097]='h000017c5;
    rd_cycle[ 5098] = 1'b0;  wr_cycle[ 5098] = 1'b1;  addr_rom[ 5098]='h000002c0;  wr_data_rom[ 5098]='h00000e4a;
    rd_cycle[ 5099] = 1'b1;  wr_cycle[ 5099] = 1'b0;  addr_rom[ 5099]='h000017d0;  wr_data_rom[ 5099]='h00000000;
    rd_cycle[ 5100] = 1'b1;  wr_cycle[ 5100] = 1'b0;  addr_rom[ 5100]='h00000c90;  wr_data_rom[ 5100]='h00000000;
    rd_cycle[ 5101] = 1'b1;  wr_cycle[ 5101] = 1'b0;  addr_rom[ 5101]='h000008b0;  wr_data_rom[ 5101]='h00000000;
    rd_cycle[ 5102] = 1'b0;  wr_cycle[ 5102] = 1'b1;  addr_rom[ 5102]='h00001768;  wr_data_rom[ 5102]='h000011d1;
    rd_cycle[ 5103] = 1'b1;  wr_cycle[ 5103] = 1'b0;  addr_rom[ 5103]='h000019cc;  wr_data_rom[ 5103]='h00000000;
    rd_cycle[ 5104] = 1'b0;  wr_cycle[ 5104] = 1'b1;  addr_rom[ 5104]='h00001238;  wr_data_rom[ 5104]='h00000113;
    rd_cycle[ 5105] = 1'b1;  wr_cycle[ 5105] = 1'b0;  addr_rom[ 5105]='h00000584;  wr_data_rom[ 5105]='h00000000;
    rd_cycle[ 5106] = 1'b1;  wr_cycle[ 5106] = 1'b0;  addr_rom[ 5106]='h00001a8c;  wr_data_rom[ 5106]='h00000000;
    rd_cycle[ 5107] = 1'b0;  wr_cycle[ 5107] = 1'b1;  addr_rom[ 5107]='h000010f4;  wr_data_rom[ 5107]='h000015ca;
    rd_cycle[ 5108] = 1'b1;  wr_cycle[ 5108] = 1'b0;  addr_rom[ 5108]='h00000104;  wr_data_rom[ 5108]='h00000000;
    rd_cycle[ 5109] = 1'b0;  wr_cycle[ 5109] = 1'b1;  addr_rom[ 5109]='h00000258;  wr_data_rom[ 5109]='h00000c6d;
    rd_cycle[ 5110] = 1'b1;  wr_cycle[ 5110] = 1'b0;  addr_rom[ 5110]='h000003c4;  wr_data_rom[ 5110]='h00000000;
    rd_cycle[ 5111] = 1'b0;  wr_cycle[ 5111] = 1'b1;  addr_rom[ 5111]='h00000050;  wr_data_rom[ 5111]='h00000b8a;
    rd_cycle[ 5112] = 1'b0;  wr_cycle[ 5112] = 1'b1;  addr_rom[ 5112]='h0000138c;  wr_data_rom[ 5112]='h000001b7;
    rd_cycle[ 5113] = 1'b1;  wr_cycle[ 5113] = 1'b0;  addr_rom[ 5113]='h0000039c;  wr_data_rom[ 5113]='h00000000;
    rd_cycle[ 5114] = 1'b0;  wr_cycle[ 5114] = 1'b1;  addr_rom[ 5114]='h00001308;  wr_data_rom[ 5114]='h000010a5;
    rd_cycle[ 5115] = 1'b1;  wr_cycle[ 5115] = 1'b0;  addr_rom[ 5115]='h00001c4c;  wr_data_rom[ 5115]='h00000000;
    rd_cycle[ 5116] = 1'b0;  wr_cycle[ 5116] = 1'b1;  addr_rom[ 5116]='h000003e8;  wr_data_rom[ 5116]='h00001803;
    rd_cycle[ 5117] = 1'b1;  wr_cycle[ 5117] = 1'b0;  addr_rom[ 5117]='h000000d8;  wr_data_rom[ 5117]='h00000000;
    rd_cycle[ 5118] = 1'b0;  wr_cycle[ 5118] = 1'b1;  addr_rom[ 5118]='h0000154c;  wr_data_rom[ 5118]='h00001da9;
    rd_cycle[ 5119] = 1'b1;  wr_cycle[ 5119] = 1'b0;  addr_rom[ 5119]='h000018c0;  wr_data_rom[ 5119]='h00000000;
    rd_cycle[ 5120] = 1'b1;  wr_cycle[ 5120] = 1'b0;  addr_rom[ 5120]='h00001a54;  wr_data_rom[ 5120]='h00000000;
    rd_cycle[ 5121] = 1'b1;  wr_cycle[ 5121] = 1'b0;  addr_rom[ 5121]='h00001c28;  wr_data_rom[ 5121]='h00000000;
    rd_cycle[ 5122] = 1'b1;  wr_cycle[ 5122] = 1'b0;  addr_rom[ 5122]='h000013d0;  wr_data_rom[ 5122]='h00000000;
    rd_cycle[ 5123] = 1'b0;  wr_cycle[ 5123] = 1'b1;  addr_rom[ 5123]='h00001ca8;  wr_data_rom[ 5123]='h00001f39;
    rd_cycle[ 5124] = 1'b0;  wr_cycle[ 5124] = 1'b1;  addr_rom[ 5124]='h00001888;  wr_data_rom[ 5124]='h000000a9;
    rd_cycle[ 5125] = 1'b0;  wr_cycle[ 5125] = 1'b1;  addr_rom[ 5125]='h00001e3c;  wr_data_rom[ 5125]='h00000785;
    rd_cycle[ 5126] = 1'b0;  wr_cycle[ 5126] = 1'b1;  addr_rom[ 5126]='h000005f8;  wr_data_rom[ 5126]='h00000692;
    rd_cycle[ 5127] = 1'b1;  wr_cycle[ 5127] = 1'b0;  addr_rom[ 5127]='h00000b50;  wr_data_rom[ 5127]='h00000000;
    rd_cycle[ 5128] = 1'b1;  wr_cycle[ 5128] = 1'b0;  addr_rom[ 5128]='h00001808;  wr_data_rom[ 5128]='h00000000;
    rd_cycle[ 5129] = 1'b1;  wr_cycle[ 5129] = 1'b0;  addr_rom[ 5129]='h00001a14;  wr_data_rom[ 5129]='h00000000;
    rd_cycle[ 5130] = 1'b0;  wr_cycle[ 5130] = 1'b1;  addr_rom[ 5130]='h000003f0;  wr_data_rom[ 5130]='h000002c5;
    rd_cycle[ 5131] = 1'b1;  wr_cycle[ 5131] = 1'b0;  addr_rom[ 5131]='h00000b2c;  wr_data_rom[ 5131]='h00000000;
    rd_cycle[ 5132] = 1'b1;  wr_cycle[ 5132] = 1'b0;  addr_rom[ 5132]='h00000670;  wr_data_rom[ 5132]='h00000000;
    rd_cycle[ 5133] = 1'b1;  wr_cycle[ 5133] = 1'b0;  addr_rom[ 5133]='h00001284;  wr_data_rom[ 5133]='h00000000;
    rd_cycle[ 5134] = 1'b1;  wr_cycle[ 5134] = 1'b0;  addr_rom[ 5134]='h000001dc;  wr_data_rom[ 5134]='h00000000;
    rd_cycle[ 5135] = 1'b0;  wr_cycle[ 5135] = 1'b1;  addr_rom[ 5135]='h00001068;  wr_data_rom[ 5135]='h0000064b;
    rd_cycle[ 5136] = 1'b0;  wr_cycle[ 5136] = 1'b1;  addr_rom[ 5136]='h00001af8;  wr_data_rom[ 5136]='h00000feb;
    rd_cycle[ 5137] = 1'b0;  wr_cycle[ 5137] = 1'b1;  addr_rom[ 5137]='h000019fc;  wr_data_rom[ 5137]='h00000e5f;
    rd_cycle[ 5138] = 1'b1;  wr_cycle[ 5138] = 1'b0;  addr_rom[ 5138]='h00000740;  wr_data_rom[ 5138]='h00000000;
    rd_cycle[ 5139] = 1'b0;  wr_cycle[ 5139] = 1'b1;  addr_rom[ 5139]='h00000410;  wr_data_rom[ 5139]='h000004ab;
    rd_cycle[ 5140] = 1'b1;  wr_cycle[ 5140] = 1'b0;  addr_rom[ 5140]='h00000214;  wr_data_rom[ 5140]='h00000000;
    rd_cycle[ 5141] = 1'b0;  wr_cycle[ 5141] = 1'b1;  addr_rom[ 5141]='h00001324;  wr_data_rom[ 5141]='h00001cd1;
    rd_cycle[ 5142] = 1'b1;  wr_cycle[ 5142] = 1'b0;  addr_rom[ 5142]='h00001e50;  wr_data_rom[ 5142]='h00000000;
    rd_cycle[ 5143] = 1'b1;  wr_cycle[ 5143] = 1'b0;  addr_rom[ 5143]='h00001254;  wr_data_rom[ 5143]='h00000000;
    rd_cycle[ 5144] = 1'b1;  wr_cycle[ 5144] = 1'b0;  addr_rom[ 5144]='h00000b34;  wr_data_rom[ 5144]='h00000000;
    rd_cycle[ 5145] = 1'b0;  wr_cycle[ 5145] = 1'b1;  addr_rom[ 5145]='h00000618;  wr_data_rom[ 5145]='h00000591;
    rd_cycle[ 5146] = 1'b1;  wr_cycle[ 5146] = 1'b0;  addr_rom[ 5146]='h00001bb8;  wr_data_rom[ 5146]='h00000000;
    rd_cycle[ 5147] = 1'b1;  wr_cycle[ 5147] = 1'b0;  addr_rom[ 5147]='h00000e4c;  wr_data_rom[ 5147]='h00000000;
    rd_cycle[ 5148] = 1'b0;  wr_cycle[ 5148] = 1'b1;  addr_rom[ 5148]='h00001b2c;  wr_data_rom[ 5148]='h00000c57;
    rd_cycle[ 5149] = 1'b1;  wr_cycle[ 5149] = 1'b0;  addr_rom[ 5149]='h00000910;  wr_data_rom[ 5149]='h00000000;
    rd_cycle[ 5150] = 1'b0;  wr_cycle[ 5150] = 1'b1;  addr_rom[ 5150]='h00000254;  wr_data_rom[ 5150]='h00001067;
    rd_cycle[ 5151] = 1'b0;  wr_cycle[ 5151] = 1'b1;  addr_rom[ 5151]='h00001734;  wr_data_rom[ 5151]='h00000cfe;
    rd_cycle[ 5152] = 1'b1;  wr_cycle[ 5152] = 1'b0;  addr_rom[ 5152]='h00000870;  wr_data_rom[ 5152]='h00000000;
    rd_cycle[ 5153] = 1'b1;  wr_cycle[ 5153] = 1'b0;  addr_rom[ 5153]='h000010c4;  wr_data_rom[ 5153]='h00000000;
    rd_cycle[ 5154] = 1'b1;  wr_cycle[ 5154] = 1'b0;  addr_rom[ 5154]='h0000000c;  wr_data_rom[ 5154]='h00000000;
    rd_cycle[ 5155] = 1'b0;  wr_cycle[ 5155] = 1'b1;  addr_rom[ 5155]='h00000a58;  wr_data_rom[ 5155]='h00000359;
    rd_cycle[ 5156] = 1'b0;  wr_cycle[ 5156] = 1'b1;  addr_rom[ 5156]='h000004a8;  wr_data_rom[ 5156]='h00001b11;
    rd_cycle[ 5157] = 1'b0;  wr_cycle[ 5157] = 1'b1;  addr_rom[ 5157]='h000002a4;  wr_data_rom[ 5157]='h0000107f;
    rd_cycle[ 5158] = 1'b0;  wr_cycle[ 5158] = 1'b1;  addr_rom[ 5158]='h00001b38;  wr_data_rom[ 5158]='h000001ae;
    rd_cycle[ 5159] = 1'b0;  wr_cycle[ 5159] = 1'b1;  addr_rom[ 5159]='h00001078;  wr_data_rom[ 5159]='h0000041c;
    rd_cycle[ 5160] = 1'b1;  wr_cycle[ 5160] = 1'b0;  addr_rom[ 5160]='h00001848;  wr_data_rom[ 5160]='h00000000;
    rd_cycle[ 5161] = 1'b1;  wr_cycle[ 5161] = 1'b0;  addr_rom[ 5161]='h00000f08;  wr_data_rom[ 5161]='h00000000;
    rd_cycle[ 5162] = 1'b1;  wr_cycle[ 5162] = 1'b0;  addr_rom[ 5162]='h00000484;  wr_data_rom[ 5162]='h00000000;
    rd_cycle[ 5163] = 1'b1;  wr_cycle[ 5163] = 1'b0;  addr_rom[ 5163]='h0000033c;  wr_data_rom[ 5163]='h00000000;
    rd_cycle[ 5164] = 1'b1;  wr_cycle[ 5164] = 1'b0;  addr_rom[ 5164]='h000014a4;  wr_data_rom[ 5164]='h00000000;
    rd_cycle[ 5165] = 1'b1;  wr_cycle[ 5165] = 1'b0;  addr_rom[ 5165]='h00000eb8;  wr_data_rom[ 5165]='h00000000;
    rd_cycle[ 5166] = 1'b1;  wr_cycle[ 5166] = 1'b0;  addr_rom[ 5166]='h00000214;  wr_data_rom[ 5166]='h00000000;
    rd_cycle[ 5167] = 1'b1;  wr_cycle[ 5167] = 1'b0;  addr_rom[ 5167]='h000005b8;  wr_data_rom[ 5167]='h00000000;
    rd_cycle[ 5168] = 1'b0;  wr_cycle[ 5168] = 1'b1;  addr_rom[ 5168]='h00000a38;  wr_data_rom[ 5168]='h0000197c;
    rd_cycle[ 5169] = 1'b1;  wr_cycle[ 5169] = 1'b0;  addr_rom[ 5169]='h000004a0;  wr_data_rom[ 5169]='h00000000;
    rd_cycle[ 5170] = 1'b0;  wr_cycle[ 5170] = 1'b1;  addr_rom[ 5170]='h000008f8;  wr_data_rom[ 5170]='h00001096;
    rd_cycle[ 5171] = 1'b1;  wr_cycle[ 5171] = 1'b0;  addr_rom[ 5171]='h00001754;  wr_data_rom[ 5171]='h00000000;
    rd_cycle[ 5172] = 1'b1;  wr_cycle[ 5172] = 1'b0;  addr_rom[ 5172]='h00001c98;  wr_data_rom[ 5172]='h00000000;
    rd_cycle[ 5173] = 1'b0;  wr_cycle[ 5173] = 1'b1;  addr_rom[ 5173]='h000004d8;  wr_data_rom[ 5173]='h00000bc3;
    rd_cycle[ 5174] = 1'b0;  wr_cycle[ 5174] = 1'b1;  addr_rom[ 5174]='h0000076c;  wr_data_rom[ 5174]='h0000158b;
    rd_cycle[ 5175] = 1'b1;  wr_cycle[ 5175] = 1'b0;  addr_rom[ 5175]='h00000f30;  wr_data_rom[ 5175]='h00000000;
    rd_cycle[ 5176] = 1'b0;  wr_cycle[ 5176] = 1'b1;  addr_rom[ 5176]='h00000cb4;  wr_data_rom[ 5176]='h00001c84;
    rd_cycle[ 5177] = 1'b1;  wr_cycle[ 5177] = 1'b0;  addr_rom[ 5177]='h00001dd4;  wr_data_rom[ 5177]='h00000000;
    rd_cycle[ 5178] = 1'b0;  wr_cycle[ 5178] = 1'b1;  addr_rom[ 5178]='h00001524;  wr_data_rom[ 5178]='h0000020e;
    rd_cycle[ 5179] = 1'b1;  wr_cycle[ 5179] = 1'b0;  addr_rom[ 5179]='h00001594;  wr_data_rom[ 5179]='h00000000;
    rd_cycle[ 5180] = 1'b1;  wr_cycle[ 5180] = 1'b0;  addr_rom[ 5180]='h00000614;  wr_data_rom[ 5180]='h00000000;
    rd_cycle[ 5181] = 1'b1;  wr_cycle[ 5181] = 1'b0;  addr_rom[ 5181]='h00001ab8;  wr_data_rom[ 5181]='h00000000;
    rd_cycle[ 5182] = 1'b0;  wr_cycle[ 5182] = 1'b1;  addr_rom[ 5182]='h00001ac8;  wr_data_rom[ 5182]='h00001e80;
    rd_cycle[ 5183] = 1'b0;  wr_cycle[ 5183] = 1'b1;  addr_rom[ 5183]='h000019a8;  wr_data_rom[ 5183]='h00000db8;
    rd_cycle[ 5184] = 1'b0;  wr_cycle[ 5184] = 1'b1;  addr_rom[ 5184]='h0000198c;  wr_data_rom[ 5184]='h000000fe;
    rd_cycle[ 5185] = 1'b1;  wr_cycle[ 5185] = 1'b0;  addr_rom[ 5185]='h00001368;  wr_data_rom[ 5185]='h00000000;
    rd_cycle[ 5186] = 1'b1;  wr_cycle[ 5186] = 1'b0;  addr_rom[ 5186]='h000018b4;  wr_data_rom[ 5186]='h00000000;
    rd_cycle[ 5187] = 1'b0;  wr_cycle[ 5187] = 1'b1;  addr_rom[ 5187]='h000010bc;  wr_data_rom[ 5187]='h00001b0e;
    rd_cycle[ 5188] = 1'b1;  wr_cycle[ 5188] = 1'b0;  addr_rom[ 5188]='h000009cc;  wr_data_rom[ 5188]='h00000000;
    rd_cycle[ 5189] = 1'b0;  wr_cycle[ 5189] = 1'b1;  addr_rom[ 5189]='h00001eb8;  wr_data_rom[ 5189]='h00001770;
    rd_cycle[ 5190] = 1'b1;  wr_cycle[ 5190] = 1'b0;  addr_rom[ 5190]='h000008d4;  wr_data_rom[ 5190]='h00000000;
    rd_cycle[ 5191] = 1'b0;  wr_cycle[ 5191] = 1'b1;  addr_rom[ 5191]='h000005e0;  wr_data_rom[ 5191]='h00000682;
    rd_cycle[ 5192] = 1'b0;  wr_cycle[ 5192] = 1'b1;  addr_rom[ 5192]='h00001de0;  wr_data_rom[ 5192]='h00000b3e;
    rd_cycle[ 5193] = 1'b0;  wr_cycle[ 5193] = 1'b1;  addr_rom[ 5193]='h00000e64;  wr_data_rom[ 5193]='h000015e8;
    rd_cycle[ 5194] = 1'b1;  wr_cycle[ 5194] = 1'b0;  addr_rom[ 5194]='h00001720;  wr_data_rom[ 5194]='h00000000;
    rd_cycle[ 5195] = 1'b0;  wr_cycle[ 5195] = 1'b1;  addr_rom[ 5195]='h0000140c;  wr_data_rom[ 5195]='h00001e60;
    rd_cycle[ 5196] = 1'b1;  wr_cycle[ 5196] = 1'b0;  addr_rom[ 5196]='h00001e50;  wr_data_rom[ 5196]='h00000000;
    rd_cycle[ 5197] = 1'b1;  wr_cycle[ 5197] = 1'b0;  addr_rom[ 5197]='h00001c38;  wr_data_rom[ 5197]='h00000000;
    rd_cycle[ 5198] = 1'b0;  wr_cycle[ 5198] = 1'b1;  addr_rom[ 5198]='h00000ff0;  wr_data_rom[ 5198]='h000011fb;
    rd_cycle[ 5199] = 1'b0;  wr_cycle[ 5199] = 1'b1;  addr_rom[ 5199]='h000000ac;  wr_data_rom[ 5199]='h00000068;
    rd_cycle[ 5200] = 1'b1;  wr_cycle[ 5200] = 1'b0;  addr_rom[ 5200]='h000011d0;  wr_data_rom[ 5200]='h00000000;
    rd_cycle[ 5201] = 1'b0;  wr_cycle[ 5201] = 1'b1;  addr_rom[ 5201]='h0000155c;  wr_data_rom[ 5201]='h000014b5;
    rd_cycle[ 5202] = 1'b1;  wr_cycle[ 5202] = 1'b0;  addr_rom[ 5202]='h00001b6c;  wr_data_rom[ 5202]='h00000000;
    rd_cycle[ 5203] = 1'b0;  wr_cycle[ 5203] = 1'b1;  addr_rom[ 5203]='h0000086c;  wr_data_rom[ 5203]='h00000f47;
    rd_cycle[ 5204] = 1'b1;  wr_cycle[ 5204] = 1'b0;  addr_rom[ 5204]='h00000d34;  wr_data_rom[ 5204]='h00000000;
    rd_cycle[ 5205] = 1'b1;  wr_cycle[ 5205] = 1'b0;  addr_rom[ 5205]='h00000140;  wr_data_rom[ 5205]='h00000000;
    rd_cycle[ 5206] = 1'b0;  wr_cycle[ 5206] = 1'b1;  addr_rom[ 5206]='h00001980;  wr_data_rom[ 5206]='h00001cfe;
    rd_cycle[ 5207] = 1'b0;  wr_cycle[ 5207] = 1'b1;  addr_rom[ 5207]='h000000f8;  wr_data_rom[ 5207]='h00001969;
    rd_cycle[ 5208] = 1'b1;  wr_cycle[ 5208] = 1'b0;  addr_rom[ 5208]='h00000ea4;  wr_data_rom[ 5208]='h00000000;
    rd_cycle[ 5209] = 1'b0;  wr_cycle[ 5209] = 1'b1;  addr_rom[ 5209]='h00000210;  wr_data_rom[ 5209]='h00000e3b;
    rd_cycle[ 5210] = 1'b1;  wr_cycle[ 5210] = 1'b0;  addr_rom[ 5210]='h00000b0c;  wr_data_rom[ 5210]='h00000000;
    rd_cycle[ 5211] = 1'b0;  wr_cycle[ 5211] = 1'b1;  addr_rom[ 5211]='h00000808;  wr_data_rom[ 5211]='h000009e2;
    rd_cycle[ 5212] = 1'b0;  wr_cycle[ 5212] = 1'b1;  addr_rom[ 5212]='h000005ac;  wr_data_rom[ 5212]='h0000187f;
    rd_cycle[ 5213] = 1'b1;  wr_cycle[ 5213] = 1'b0;  addr_rom[ 5213]='h00000134;  wr_data_rom[ 5213]='h00000000;
    rd_cycle[ 5214] = 1'b0;  wr_cycle[ 5214] = 1'b1;  addr_rom[ 5214]='h000015b0;  wr_data_rom[ 5214]='h00000054;
    rd_cycle[ 5215] = 1'b0;  wr_cycle[ 5215] = 1'b1;  addr_rom[ 5215]='h000009a4;  wr_data_rom[ 5215]='h00000fef;
    rd_cycle[ 5216] = 1'b1;  wr_cycle[ 5216] = 1'b0;  addr_rom[ 5216]='h00001184;  wr_data_rom[ 5216]='h00000000;
    rd_cycle[ 5217] = 1'b0;  wr_cycle[ 5217] = 1'b1;  addr_rom[ 5217]='h00000234;  wr_data_rom[ 5217]='h00001b0f;
    rd_cycle[ 5218] = 1'b1;  wr_cycle[ 5218] = 1'b0;  addr_rom[ 5218]='h00000fb8;  wr_data_rom[ 5218]='h00000000;
    rd_cycle[ 5219] = 1'b1;  wr_cycle[ 5219] = 1'b0;  addr_rom[ 5219]='h00001e04;  wr_data_rom[ 5219]='h00000000;
    rd_cycle[ 5220] = 1'b1;  wr_cycle[ 5220] = 1'b0;  addr_rom[ 5220]='h00001d08;  wr_data_rom[ 5220]='h00000000;
    rd_cycle[ 5221] = 1'b0;  wr_cycle[ 5221] = 1'b1;  addr_rom[ 5221]='h000019a0;  wr_data_rom[ 5221]='h00000622;
    rd_cycle[ 5222] = 1'b1;  wr_cycle[ 5222] = 1'b0;  addr_rom[ 5222]='h0000139c;  wr_data_rom[ 5222]='h00000000;
    rd_cycle[ 5223] = 1'b1;  wr_cycle[ 5223] = 1'b0;  addr_rom[ 5223]='h00000c94;  wr_data_rom[ 5223]='h00000000;
    rd_cycle[ 5224] = 1'b0;  wr_cycle[ 5224] = 1'b1;  addr_rom[ 5224]='h00000c5c;  wr_data_rom[ 5224]='h00001bcc;
    rd_cycle[ 5225] = 1'b0;  wr_cycle[ 5225] = 1'b1;  addr_rom[ 5225]='h00001120;  wr_data_rom[ 5225]='h00000984;
    rd_cycle[ 5226] = 1'b0;  wr_cycle[ 5226] = 1'b1;  addr_rom[ 5226]='h000011c0;  wr_data_rom[ 5226]='h000009f1;
    rd_cycle[ 5227] = 1'b1;  wr_cycle[ 5227] = 1'b0;  addr_rom[ 5227]='h00000c3c;  wr_data_rom[ 5227]='h00000000;
    rd_cycle[ 5228] = 1'b1;  wr_cycle[ 5228] = 1'b0;  addr_rom[ 5228]='h00000ed8;  wr_data_rom[ 5228]='h00000000;
    rd_cycle[ 5229] = 1'b0;  wr_cycle[ 5229] = 1'b1;  addr_rom[ 5229]='h000012e8;  wr_data_rom[ 5229]='h0000159b;
    rd_cycle[ 5230] = 1'b1;  wr_cycle[ 5230] = 1'b0;  addr_rom[ 5230]='h0000168c;  wr_data_rom[ 5230]='h00000000;
    rd_cycle[ 5231] = 1'b1;  wr_cycle[ 5231] = 1'b0;  addr_rom[ 5231]='h00000dfc;  wr_data_rom[ 5231]='h00000000;
    rd_cycle[ 5232] = 1'b1;  wr_cycle[ 5232] = 1'b0;  addr_rom[ 5232]='h00001334;  wr_data_rom[ 5232]='h00000000;
    rd_cycle[ 5233] = 1'b1;  wr_cycle[ 5233] = 1'b0;  addr_rom[ 5233]='h00001a74;  wr_data_rom[ 5233]='h00000000;
    rd_cycle[ 5234] = 1'b1;  wr_cycle[ 5234] = 1'b0;  addr_rom[ 5234]='h00001d7c;  wr_data_rom[ 5234]='h00000000;
    rd_cycle[ 5235] = 1'b1;  wr_cycle[ 5235] = 1'b0;  addr_rom[ 5235]='h0000010c;  wr_data_rom[ 5235]='h00000000;
    rd_cycle[ 5236] = 1'b1;  wr_cycle[ 5236] = 1'b0;  addr_rom[ 5236]='h00001074;  wr_data_rom[ 5236]='h00000000;
    rd_cycle[ 5237] = 1'b1;  wr_cycle[ 5237] = 1'b0;  addr_rom[ 5237]='h00000f34;  wr_data_rom[ 5237]='h00000000;
    rd_cycle[ 5238] = 1'b1;  wr_cycle[ 5238] = 1'b0;  addr_rom[ 5238]='h000009d0;  wr_data_rom[ 5238]='h00000000;
    rd_cycle[ 5239] = 1'b0;  wr_cycle[ 5239] = 1'b1;  addr_rom[ 5239]='h00000824;  wr_data_rom[ 5239]='h000003cf;
    rd_cycle[ 5240] = 1'b0;  wr_cycle[ 5240] = 1'b1;  addr_rom[ 5240]='h00000fb8;  wr_data_rom[ 5240]='h000008bb;
    rd_cycle[ 5241] = 1'b0;  wr_cycle[ 5241] = 1'b1;  addr_rom[ 5241]='h000008a0;  wr_data_rom[ 5241]='h00001b33;
    rd_cycle[ 5242] = 1'b1;  wr_cycle[ 5242] = 1'b0;  addr_rom[ 5242]='h00001adc;  wr_data_rom[ 5242]='h00000000;
    rd_cycle[ 5243] = 1'b1;  wr_cycle[ 5243] = 1'b0;  addr_rom[ 5243]='h0000045c;  wr_data_rom[ 5243]='h00000000;
    rd_cycle[ 5244] = 1'b1;  wr_cycle[ 5244] = 1'b0;  addr_rom[ 5244]='h00000f68;  wr_data_rom[ 5244]='h00000000;
    rd_cycle[ 5245] = 1'b1;  wr_cycle[ 5245] = 1'b0;  addr_rom[ 5245]='h00000840;  wr_data_rom[ 5245]='h00000000;
    rd_cycle[ 5246] = 1'b1;  wr_cycle[ 5246] = 1'b0;  addr_rom[ 5246]='h000005cc;  wr_data_rom[ 5246]='h00000000;
    rd_cycle[ 5247] = 1'b1;  wr_cycle[ 5247] = 1'b0;  addr_rom[ 5247]='h00000d68;  wr_data_rom[ 5247]='h00000000;
    rd_cycle[ 5248] = 1'b0;  wr_cycle[ 5248] = 1'b1;  addr_rom[ 5248]='h00001528;  wr_data_rom[ 5248]='h00001af6;
    rd_cycle[ 5249] = 1'b1;  wr_cycle[ 5249] = 1'b0;  addr_rom[ 5249]='h00001b70;  wr_data_rom[ 5249]='h00000000;
    rd_cycle[ 5250] = 1'b0;  wr_cycle[ 5250] = 1'b1;  addr_rom[ 5250]='h00000ebc;  wr_data_rom[ 5250]='h00001344;
    rd_cycle[ 5251] = 1'b0;  wr_cycle[ 5251] = 1'b1;  addr_rom[ 5251]='h000018f8;  wr_data_rom[ 5251]='h00001a93;
    rd_cycle[ 5252] = 1'b0;  wr_cycle[ 5252] = 1'b1;  addr_rom[ 5252]='h00001468;  wr_data_rom[ 5252]='h00000f51;
    rd_cycle[ 5253] = 1'b1;  wr_cycle[ 5253] = 1'b0;  addr_rom[ 5253]='h0000112c;  wr_data_rom[ 5253]='h00000000;
    rd_cycle[ 5254] = 1'b1;  wr_cycle[ 5254] = 1'b0;  addr_rom[ 5254]='h00001950;  wr_data_rom[ 5254]='h00000000;
    rd_cycle[ 5255] = 1'b1;  wr_cycle[ 5255] = 1'b0;  addr_rom[ 5255]='h00000200;  wr_data_rom[ 5255]='h00000000;
    rd_cycle[ 5256] = 1'b1;  wr_cycle[ 5256] = 1'b0;  addr_rom[ 5256]='h00000e04;  wr_data_rom[ 5256]='h00000000;
    rd_cycle[ 5257] = 1'b1;  wr_cycle[ 5257] = 1'b0;  addr_rom[ 5257]='h000001dc;  wr_data_rom[ 5257]='h00000000;
    rd_cycle[ 5258] = 1'b0;  wr_cycle[ 5258] = 1'b1;  addr_rom[ 5258]='h00000cd8;  wr_data_rom[ 5258]='h000012fb;
    rd_cycle[ 5259] = 1'b1;  wr_cycle[ 5259] = 1'b0;  addr_rom[ 5259]='h00001d94;  wr_data_rom[ 5259]='h00000000;
    rd_cycle[ 5260] = 1'b0;  wr_cycle[ 5260] = 1'b1;  addr_rom[ 5260]='h00001924;  wr_data_rom[ 5260]='h00001200;
    rd_cycle[ 5261] = 1'b0;  wr_cycle[ 5261] = 1'b1;  addr_rom[ 5261]='h00000e00;  wr_data_rom[ 5261]='h0000174f;
    rd_cycle[ 5262] = 1'b1;  wr_cycle[ 5262] = 1'b0;  addr_rom[ 5262]='h000018f8;  wr_data_rom[ 5262]='h00000000;
    rd_cycle[ 5263] = 1'b0;  wr_cycle[ 5263] = 1'b1;  addr_rom[ 5263]='h00001880;  wr_data_rom[ 5263]='h00001bda;
    rd_cycle[ 5264] = 1'b0;  wr_cycle[ 5264] = 1'b1;  addr_rom[ 5264]='h00000ea8;  wr_data_rom[ 5264]='h000014d5;
    rd_cycle[ 5265] = 1'b0;  wr_cycle[ 5265] = 1'b1;  addr_rom[ 5265]='h000016c8;  wr_data_rom[ 5265]='h000009e3;
    rd_cycle[ 5266] = 1'b0;  wr_cycle[ 5266] = 1'b1;  addr_rom[ 5266]='h000019c8;  wr_data_rom[ 5266]='h000004ad;
    rd_cycle[ 5267] = 1'b0;  wr_cycle[ 5267] = 1'b1;  addr_rom[ 5267]='h00000640;  wr_data_rom[ 5267]='h000008c8;
    rd_cycle[ 5268] = 1'b0;  wr_cycle[ 5268] = 1'b1;  addr_rom[ 5268]='h000015e4;  wr_data_rom[ 5268]='h000016f8;
    rd_cycle[ 5269] = 1'b0;  wr_cycle[ 5269] = 1'b1;  addr_rom[ 5269]='h00001894;  wr_data_rom[ 5269]='h00001b27;
    rd_cycle[ 5270] = 1'b1;  wr_cycle[ 5270] = 1'b0;  addr_rom[ 5270]='h000008bc;  wr_data_rom[ 5270]='h00000000;
    rd_cycle[ 5271] = 1'b0;  wr_cycle[ 5271] = 1'b1;  addr_rom[ 5271]='h00000488;  wr_data_rom[ 5271]='h00001b8a;
    rd_cycle[ 5272] = 1'b0;  wr_cycle[ 5272] = 1'b1;  addr_rom[ 5272]='h00000764;  wr_data_rom[ 5272]='h00001646;
    rd_cycle[ 5273] = 1'b0;  wr_cycle[ 5273] = 1'b1;  addr_rom[ 5273]='h000006f4;  wr_data_rom[ 5273]='h00001d7d;
    rd_cycle[ 5274] = 1'b0;  wr_cycle[ 5274] = 1'b1;  addr_rom[ 5274]='h00001908;  wr_data_rom[ 5274]='h00001dcf;
    rd_cycle[ 5275] = 1'b0;  wr_cycle[ 5275] = 1'b1;  addr_rom[ 5275]='h000013cc;  wr_data_rom[ 5275]='h000017cf;
    rd_cycle[ 5276] = 1'b0;  wr_cycle[ 5276] = 1'b1;  addr_rom[ 5276]='h00000ddc;  wr_data_rom[ 5276]='h000014f2;
    rd_cycle[ 5277] = 1'b1;  wr_cycle[ 5277] = 1'b0;  addr_rom[ 5277]='h00000108;  wr_data_rom[ 5277]='h00000000;
    rd_cycle[ 5278] = 1'b0;  wr_cycle[ 5278] = 1'b1;  addr_rom[ 5278]='h00001e88;  wr_data_rom[ 5278]='h00000131;
    rd_cycle[ 5279] = 1'b0;  wr_cycle[ 5279] = 1'b1;  addr_rom[ 5279]='h0000177c;  wr_data_rom[ 5279]='h000012da;
    rd_cycle[ 5280] = 1'b1;  wr_cycle[ 5280] = 1'b0;  addr_rom[ 5280]='h00001a54;  wr_data_rom[ 5280]='h00000000;
    rd_cycle[ 5281] = 1'b1;  wr_cycle[ 5281] = 1'b0;  addr_rom[ 5281]='h00000418;  wr_data_rom[ 5281]='h00000000;
    rd_cycle[ 5282] = 1'b0;  wr_cycle[ 5282] = 1'b1;  addr_rom[ 5282]='h000010dc;  wr_data_rom[ 5282]='h0000128b;
    rd_cycle[ 5283] = 1'b1;  wr_cycle[ 5283] = 1'b0;  addr_rom[ 5283]='h00001d10;  wr_data_rom[ 5283]='h00000000;
    rd_cycle[ 5284] = 1'b1;  wr_cycle[ 5284] = 1'b0;  addr_rom[ 5284]='h000002e4;  wr_data_rom[ 5284]='h00000000;
    rd_cycle[ 5285] = 1'b1;  wr_cycle[ 5285] = 1'b0;  addr_rom[ 5285]='h00000ff0;  wr_data_rom[ 5285]='h00000000;
    rd_cycle[ 5286] = 1'b1;  wr_cycle[ 5286] = 1'b0;  addr_rom[ 5286]='h000006fc;  wr_data_rom[ 5286]='h00000000;
    rd_cycle[ 5287] = 1'b1;  wr_cycle[ 5287] = 1'b0;  addr_rom[ 5287]='h00001cb4;  wr_data_rom[ 5287]='h00000000;
    rd_cycle[ 5288] = 1'b1;  wr_cycle[ 5288] = 1'b0;  addr_rom[ 5288]='h0000170c;  wr_data_rom[ 5288]='h00000000;
    rd_cycle[ 5289] = 1'b0;  wr_cycle[ 5289] = 1'b1;  addr_rom[ 5289]='h00000cb8;  wr_data_rom[ 5289]='h0000122c;
    rd_cycle[ 5290] = 1'b1;  wr_cycle[ 5290] = 1'b0;  addr_rom[ 5290]='h00001754;  wr_data_rom[ 5290]='h00000000;
    rd_cycle[ 5291] = 1'b1;  wr_cycle[ 5291] = 1'b0;  addr_rom[ 5291]='h00000d28;  wr_data_rom[ 5291]='h00000000;
    rd_cycle[ 5292] = 1'b1;  wr_cycle[ 5292] = 1'b0;  addr_rom[ 5292]='h00001d00;  wr_data_rom[ 5292]='h00000000;
    rd_cycle[ 5293] = 1'b1;  wr_cycle[ 5293] = 1'b0;  addr_rom[ 5293]='h00001634;  wr_data_rom[ 5293]='h00000000;
    rd_cycle[ 5294] = 1'b0;  wr_cycle[ 5294] = 1'b1;  addr_rom[ 5294]='h000015c8;  wr_data_rom[ 5294]='h000006ba;
    rd_cycle[ 5295] = 1'b1;  wr_cycle[ 5295] = 1'b0;  addr_rom[ 5295]='h00001910;  wr_data_rom[ 5295]='h00000000;
    rd_cycle[ 5296] = 1'b0;  wr_cycle[ 5296] = 1'b1;  addr_rom[ 5296]='h00000904;  wr_data_rom[ 5296]='h00001558;
    rd_cycle[ 5297] = 1'b1;  wr_cycle[ 5297] = 1'b0;  addr_rom[ 5297]='h000019f8;  wr_data_rom[ 5297]='h00000000;
    rd_cycle[ 5298] = 1'b1;  wr_cycle[ 5298] = 1'b0;  addr_rom[ 5298]='h00001c04;  wr_data_rom[ 5298]='h00000000;
    rd_cycle[ 5299] = 1'b1;  wr_cycle[ 5299] = 1'b0;  addr_rom[ 5299]='h00000e4c;  wr_data_rom[ 5299]='h00000000;
    rd_cycle[ 5300] = 1'b0;  wr_cycle[ 5300] = 1'b1;  addr_rom[ 5300]='h0000020c;  wr_data_rom[ 5300]='h00000326;
    rd_cycle[ 5301] = 1'b0;  wr_cycle[ 5301] = 1'b1;  addr_rom[ 5301]='h00001690;  wr_data_rom[ 5301]='h00000936;
    rd_cycle[ 5302] = 1'b1;  wr_cycle[ 5302] = 1'b0;  addr_rom[ 5302]='h00001b90;  wr_data_rom[ 5302]='h00000000;
    rd_cycle[ 5303] = 1'b0;  wr_cycle[ 5303] = 1'b1;  addr_rom[ 5303]='h000006d8;  wr_data_rom[ 5303]='h00000afc;
    rd_cycle[ 5304] = 1'b1;  wr_cycle[ 5304] = 1'b0;  addr_rom[ 5304]='h00001ecc;  wr_data_rom[ 5304]='h00000000;
    rd_cycle[ 5305] = 1'b1;  wr_cycle[ 5305] = 1'b0;  addr_rom[ 5305]='h00000920;  wr_data_rom[ 5305]='h00000000;
    rd_cycle[ 5306] = 1'b1;  wr_cycle[ 5306] = 1'b0;  addr_rom[ 5306]='h00000678;  wr_data_rom[ 5306]='h00000000;
    rd_cycle[ 5307] = 1'b0;  wr_cycle[ 5307] = 1'b1;  addr_rom[ 5307]='h00000ca4;  wr_data_rom[ 5307]='h00001dc1;
    rd_cycle[ 5308] = 1'b1;  wr_cycle[ 5308] = 1'b0;  addr_rom[ 5308]='h00001844;  wr_data_rom[ 5308]='h00000000;
    rd_cycle[ 5309] = 1'b0;  wr_cycle[ 5309] = 1'b1;  addr_rom[ 5309]='h00000ddc;  wr_data_rom[ 5309]='h0000093c;
    rd_cycle[ 5310] = 1'b1;  wr_cycle[ 5310] = 1'b0;  addr_rom[ 5310]='h00001440;  wr_data_rom[ 5310]='h00000000;
    rd_cycle[ 5311] = 1'b0;  wr_cycle[ 5311] = 1'b1;  addr_rom[ 5311]='h00000948;  wr_data_rom[ 5311]='h00001851;
    rd_cycle[ 5312] = 1'b1;  wr_cycle[ 5312] = 1'b0;  addr_rom[ 5312]='h00000bcc;  wr_data_rom[ 5312]='h00000000;
    rd_cycle[ 5313] = 1'b0;  wr_cycle[ 5313] = 1'b1;  addr_rom[ 5313]='h00001ee4;  wr_data_rom[ 5313]='h00000f9e;
    rd_cycle[ 5314] = 1'b0;  wr_cycle[ 5314] = 1'b1;  addr_rom[ 5314]='h0000086c;  wr_data_rom[ 5314]='h00001b9c;
    rd_cycle[ 5315] = 1'b1;  wr_cycle[ 5315] = 1'b0;  addr_rom[ 5315]='h0000076c;  wr_data_rom[ 5315]='h00000000;
    rd_cycle[ 5316] = 1'b1;  wr_cycle[ 5316] = 1'b0;  addr_rom[ 5316]='h00001c98;  wr_data_rom[ 5316]='h00000000;
    rd_cycle[ 5317] = 1'b0;  wr_cycle[ 5317] = 1'b1;  addr_rom[ 5317]='h00000518;  wr_data_rom[ 5317]='h00001e3e;
    rd_cycle[ 5318] = 1'b1;  wr_cycle[ 5318] = 1'b0;  addr_rom[ 5318]='h00001198;  wr_data_rom[ 5318]='h00000000;
    rd_cycle[ 5319] = 1'b1;  wr_cycle[ 5319] = 1'b0;  addr_rom[ 5319]='h00001a08;  wr_data_rom[ 5319]='h00000000;
    rd_cycle[ 5320] = 1'b0;  wr_cycle[ 5320] = 1'b1;  addr_rom[ 5320]='h00000e08;  wr_data_rom[ 5320]='h0000075f;
    rd_cycle[ 5321] = 1'b1;  wr_cycle[ 5321] = 1'b0;  addr_rom[ 5321]='h00001904;  wr_data_rom[ 5321]='h00000000;
    rd_cycle[ 5322] = 1'b1;  wr_cycle[ 5322] = 1'b0;  addr_rom[ 5322]='h000010f0;  wr_data_rom[ 5322]='h00000000;
    rd_cycle[ 5323] = 1'b1;  wr_cycle[ 5323] = 1'b0;  addr_rom[ 5323]='h00000914;  wr_data_rom[ 5323]='h00000000;
    rd_cycle[ 5324] = 1'b1;  wr_cycle[ 5324] = 1'b0;  addr_rom[ 5324]='h00000958;  wr_data_rom[ 5324]='h00000000;
    rd_cycle[ 5325] = 1'b0;  wr_cycle[ 5325] = 1'b1;  addr_rom[ 5325]='h00001af4;  wr_data_rom[ 5325]='h0000101b;
    rd_cycle[ 5326] = 1'b1;  wr_cycle[ 5326] = 1'b0;  addr_rom[ 5326]='h00000430;  wr_data_rom[ 5326]='h00000000;
    rd_cycle[ 5327] = 1'b0;  wr_cycle[ 5327] = 1'b1;  addr_rom[ 5327]='h00000d94;  wr_data_rom[ 5327]='h0000195d;
    rd_cycle[ 5328] = 1'b1;  wr_cycle[ 5328] = 1'b0;  addr_rom[ 5328]='h00000408;  wr_data_rom[ 5328]='h00000000;
    rd_cycle[ 5329] = 1'b1;  wr_cycle[ 5329] = 1'b0;  addr_rom[ 5329]='h00001ad0;  wr_data_rom[ 5329]='h00000000;
    rd_cycle[ 5330] = 1'b0;  wr_cycle[ 5330] = 1'b1;  addr_rom[ 5330]='h0000007c;  wr_data_rom[ 5330]='h00001f06;
    rd_cycle[ 5331] = 1'b1;  wr_cycle[ 5331] = 1'b0;  addr_rom[ 5331]='h00001e50;  wr_data_rom[ 5331]='h00000000;
    rd_cycle[ 5332] = 1'b0;  wr_cycle[ 5332] = 1'b1;  addr_rom[ 5332]='h0000065c;  wr_data_rom[ 5332]='h00001957;
    rd_cycle[ 5333] = 1'b1;  wr_cycle[ 5333] = 1'b0;  addr_rom[ 5333]='h000016e4;  wr_data_rom[ 5333]='h00000000;
    rd_cycle[ 5334] = 1'b0;  wr_cycle[ 5334] = 1'b1;  addr_rom[ 5334]='h00001d14;  wr_data_rom[ 5334]='h0000130c;
    rd_cycle[ 5335] = 1'b0;  wr_cycle[ 5335] = 1'b1;  addr_rom[ 5335]='h000015cc;  wr_data_rom[ 5335]='h00001ed6;
    rd_cycle[ 5336] = 1'b0;  wr_cycle[ 5336] = 1'b1;  addr_rom[ 5336]='h000012a0;  wr_data_rom[ 5336]='h00000731;
    rd_cycle[ 5337] = 1'b1;  wr_cycle[ 5337] = 1'b0;  addr_rom[ 5337]='h0000141c;  wr_data_rom[ 5337]='h00000000;
    rd_cycle[ 5338] = 1'b0;  wr_cycle[ 5338] = 1'b1;  addr_rom[ 5338]='h00000540;  wr_data_rom[ 5338]='h00000d22;
    rd_cycle[ 5339] = 1'b1;  wr_cycle[ 5339] = 1'b0;  addr_rom[ 5339]='h00000960;  wr_data_rom[ 5339]='h00000000;
    rd_cycle[ 5340] = 1'b0;  wr_cycle[ 5340] = 1'b1;  addr_rom[ 5340]='h000011b4;  wr_data_rom[ 5340]='h00001c84;
    rd_cycle[ 5341] = 1'b1;  wr_cycle[ 5341] = 1'b0;  addr_rom[ 5341]='h00001024;  wr_data_rom[ 5341]='h00000000;
    rd_cycle[ 5342] = 1'b0;  wr_cycle[ 5342] = 1'b1;  addr_rom[ 5342]='h00000460;  wr_data_rom[ 5342]='h00000cc5;
    rd_cycle[ 5343] = 1'b1;  wr_cycle[ 5343] = 1'b0;  addr_rom[ 5343]='h00001408;  wr_data_rom[ 5343]='h00000000;
    rd_cycle[ 5344] = 1'b0;  wr_cycle[ 5344] = 1'b1;  addr_rom[ 5344]='h00001db8;  wr_data_rom[ 5344]='h000005bc;
    rd_cycle[ 5345] = 1'b0;  wr_cycle[ 5345] = 1'b1;  addr_rom[ 5345]='h00001848;  wr_data_rom[ 5345]='h00001763;
    rd_cycle[ 5346] = 1'b0;  wr_cycle[ 5346] = 1'b1;  addr_rom[ 5346]='h000005fc;  wr_data_rom[ 5346]='h000002e6;
    rd_cycle[ 5347] = 1'b0;  wr_cycle[ 5347] = 1'b1;  addr_rom[ 5347]='h000008cc;  wr_data_rom[ 5347]='h000014e2;
    rd_cycle[ 5348] = 1'b1;  wr_cycle[ 5348] = 1'b0;  addr_rom[ 5348]='h00000d78;  wr_data_rom[ 5348]='h00000000;
    rd_cycle[ 5349] = 1'b1;  wr_cycle[ 5349] = 1'b0;  addr_rom[ 5349]='h00001d38;  wr_data_rom[ 5349]='h00000000;
    rd_cycle[ 5350] = 1'b0;  wr_cycle[ 5350] = 1'b1;  addr_rom[ 5350]='h00000064;  wr_data_rom[ 5350]='h0000156c;
    rd_cycle[ 5351] = 1'b1;  wr_cycle[ 5351] = 1'b0;  addr_rom[ 5351]='h000012c8;  wr_data_rom[ 5351]='h00000000;
    rd_cycle[ 5352] = 1'b0;  wr_cycle[ 5352] = 1'b1;  addr_rom[ 5352]='h00001188;  wr_data_rom[ 5352]='h00000519;
    rd_cycle[ 5353] = 1'b1;  wr_cycle[ 5353] = 1'b0;  addr_rom[ 5353]='h0000127c;  wr_data_rom[ 5353]='h00000000;
    rd_cycle[ 5354] = 1'b0;  wr_cycle[ 5354] = 1'b1;  addr_rom[ 5354]='h00000b04;  wr_data_rom[ 5354]='h00000ec7;
    rd_cycle[ 5355] = 1'b1;  wr_cycle[ 5355] = 1'b0;  addr_rom[ 5355]='h00000f08;  wr_data_rom[ 5355]='h00000000;
    rd_cycle[ 5356] = 1'b0;  wr_cycle[ 5356] = 1'b1;  addr_rom[ 5356]='h0000162c;  wr_data_rom[ 5356]='h00001404;
    rd_cycle[ 5357] = 1'b0;  wr_cycle[ 5357] = 1'b1;  addr_rom[ 5357]='h00001784;  wr_data_rom[ 5357]='h00001dbf;
    rd_cycle[ 5358] = 1'b0;  wr_cycle[ 5358] = 1'b1;  addr_rom[ 5358]='h000009f0;  wr_data_rom[ 5358]='h0000101b;
    rd_cycle[ 5359] = 1'b0;  wr_cycle[ 5359] = 1'b1;  addr_rom[ 5359]='h00000204;  wr_data_rom[ 5359]='h000014f8;
    rd_cycle[ 5360] = 1'b1;  wr_cycle[ 5360] = 1'b0;  addr_rom[ 5360]='h000002f8;  wr_data_rom[ 5360]='h00000000;
    rd_cycle[ 5361] = 1'b1;  wr_cycle[ 5361] = 1'b0;  addr_rom[ 5361]='h00000b40;  wr_data_rom[ 5361]='h00000000;
    rd_cycle[ 5362] = 1'b0;  wr_cycle[ 5362] = 1'b1;  addr_rom[ 5362]='h000012b8;  wr_data_rom[ 5362]='h00001450;
    rd_cycle[ 5363] = 1'b1;  wr_cycle[ 5363] = 1'b0;  addr_rom[ 5363]='h00000a38;  wr_data_rom[ 5363]='h00000000;
    rd_cycle[ 5364] = 1'b1;  wr_cycle[ 5364] = 1'b0;  addr_rom[ 5364]='h00001520;  wr_data_rom[ 5364]='h00000000;
    rd_cycle[ 5365] = 1'b1;  wr_cycle[ 5365] = 1'b0;  addr_rom[ 5365]='h000011dc;  wr_data_rom[ 5365]='h00000000;
    rd_cycle[ 5366] = 1'b1;  wr_cycle[ 5366] = 1'b0;  addr_rom[ 5366]='h00001124;  wr_data_rom[ 5366]='h00000000;
    rd_cycle[ 5367] = 1'b1;  wr_cycle[ 5367] = 1'b0;  addr_rom[ 5367]='h0000148c;  wr_data_rom[ 5367]='h00000000;
    rd_cycle[ 5368] = 1'b0;  wr_cycle[ 5368] = 1'b1;  addr_rom[ 5368]='h00000dd8;  wr_data_rom[ 5368]='h00001017;
    rd_cycle[ 5369] = 1'b1;  wr_cycle[ 5369] = 1'b0;  addr_rom[ 5369]='h00001130;  wr_data_rom[ 5369]='h00000000;
    rd_cycle[ 5370] = 1'b1;  wr_cycle[ 5370] = 1'b0;  addr_rom[ 5370]='h000005a4;  wr_data_rom[ 5370]='h00000000;
    rd_cycle[ 5371] = 1'b0;  wr_cycle[ 5371] = 1'b1;  addr_rom[ 5371]='h000019dc;  wr_data_rom[ 5371]='h000013df;
    rd_cycle[ 5372] = 1'b0;  wr_cycle[ 5372] = 1'b1;  addr_rom[ 5372]='h00000090;  wr_data_rom[ 5372]='h00001632;
    rd_cycle[ 5373] = 1'b0;  wr_cycle[ 5373] = 1'b1;  addr_rom[ 5373]='h000010a4;  wr_data_rom[ 5373]='h00000ff1;
    rd_cycle[ 5374] = 1'b1;  wr_cycle[ 5374] = 1'b0;  addr_rom[ 5374]='h00000434;  wr_data_rom[ 5374]='h00000000;
    rd_cycle[ 5375] = 1'b1;  wr_cycle[ 5375] = 1'b0;  addr_rom[ 5375]='h00000514;  wr_data_rom[ 5375]='h00000000;
    rd_cycle[ 5376] = 1'b1;  wr_cycle[ 5376] = 1'b0;  addr_rom[ 5376]='h00001b08;  wr_data_rom[ 5376]='h00000000;
    rd_cycle[ 5377] = 1'b1;  wr_cycle[ 5377] = 1'b0;  addr_rom[ 5377]='h00000224;  wr_data_rom[ 5377]='h00000000;
    rd_cycle[ 5378] = 1'b0;  wr_cycle[ 5378] = 1'b1;  addr_rom[ 5378]='h00000984;  wr_data_rom[ 5378]='h000001e6;
    rd_cycle[ 5379] = 1'b1;  wr_cycle[ 5379] = 1'b0;  addr_rom[ 5379]='h00001f0c;  wr_data_rom[ 5379]='h00000000;
    rd_cycle[ 5380] = 1'b1;  wr_cycle[ 5380] = 1'b0;  addr_rom[ 5380]='h00000700;  wr_data_rom[ 5380]='h00000000;
    rd_cycle[ 5381] = 1'b0;  wr_cycle[ 5381] = 1'b1;  addr_rom[ 5381]='h00001ee4;  wr_data_rom[ 5381]='h00000817;
    rd_cycle[ 5382] = 1'b1;  wr_cycle[ 5382] = 1'b0;  addr_rom[ 5382]='h00000498;  wr_data_rom[ 5382]='h00000000;
    rd_cycle[ 5383] = 1'b0;  wr_cycle[ 5383] = 1'b1;  addr_rom[ 5383]='h0000199c;  wr_data_rom[ 5383]='h00000be7;
    rd_cycle[ 5384] = 1'b0;  wr_cycle[ 5384] = 1'b1;  addr_rom[ 5384]='h00001d70;  wr_data_rom[ 5384]='h00000f54;
    rd_cycle[ 5385] = 1'b1;  wr_cycle[ 5385] = 1'b0;  addr_rom[ 5385]='h00001260;  wr_data_rom[ 5385]='h00000000;
    rd_cycle[ 5386] = 1'b0;  wr_cycle[ 5386] = 1'b1;  addr_rom[ 5386]='h00001db4;  wr_data_rom[ 5386]='h00000e4e;
    rd_cycle[ 5387] = 1'b0;  wr_cycle[ 5387] = 1'b1;  addr_rom[ 5387]='h0000009c;  wr_data_rom[ 5387]='h0000131c;
    rd_cycle[ 5388] = 1'b1;  wr_cycle[ 5388] = 1'b0;  addr_rom[ 5388]='h00000c68;  wr_data_rom[ 5388]='h00000000;
    rd_cycle[ 5389] = 1'b0;  wr_cycle[ 5389] = 1'b1;  addr_rom[ 5389]='h000013d0;  wr_data_rom[ 5389]='h000012d4;
    rd_cycle[ 5390] = 1'b1;  wr_cycle[ 5390] = 1'b0;  addr_rom[ 5390]='h00000f34;  wr_data_rom[ 5390]='h00000000;
    rd_cycle[ 5391] = 1'b1;  wr_cycle[ 5391] = 1'b0;  addr_rom[ 5391]='h00000a28;  wr_data_rom[ 5391]='h00000000;
    rd_cycle[ 5392] = 1'b0;  wr_cycle[ 5392] = 1'b1;  addr_rom[ 5392]='h00000b40;  wr_data_rom[ 5392]='h000003f1;
    rd_cycle[ 5393] = 1'b0;  wr_cycle[ 5393] = 1'b1;  addr_rom[ 5393]='h0000190c;  wr_data_rom[ 5393]='h0000013d;
    rd_cycle[ 5394] = 1'b1;  wr_cycle[ 5394] = 1'b0;  addr_rom[ 5394]='h000009e4;  wr_data_rom[ 5394]='h00000000;
    rd_cycle[ 5395] = 1'b1;  wr_cycle[ 5395] = 1'b0;  addr_rom[ 5395]='h000000ec;  wr_data_rom[ 5395]='h00000000;
    rd_cycle[ 5396] = 1'b1;  wr_cycle[ 5396] = 1'b0;  addr_rom[ 5396]='h00000380;  wr_data_rom[ 5396]='h00000000;
    rd_cycle[ 5397] = 1'b0;  wr_cycle[ 5397] = 1'b1;  addr_rom[ 5397]='h000012a0;  wr_data_rom[ 5397]='h00000ac2;
    rd_cycle[ 5398] = 1'b0;  wr_cycle[ 5398] = 1'b1;  addr_rom[ 5398]='h000006a8;  wr_data_rom[ 5398]='h00001979;
    rd_cycle[ 5399] = 1'b1;  wr_cycle[ 5399] = 1'b0;  addr_rom[ 5399]='h00000e4c;  wr_data_rom[ 5399]='h00000000;
    rd_cycle[ 5400] = 1'b1;  wr_cycle[ 5400] = 1'b0;  addr_rom[ 5400]='h000007fc;  wr_data_rom[ 5400]='h00000000;
    rd_cycle[ 5401] = 1'b1;  wr_cycle[ 5401] = 1'b0;  addr_rom[ 5401]='h00001648;  wr_data_rom[ 5401]='h00000000;
    rd_cycle[ 5402] = 1'b0;  wr_cycle[ 5402] = 1'b1;  addr_rom[ 5402]='h00001660;  wr_data_rom[ 5402]='h00000e8b;
    rd_cycle[ 5403] = 1'b1;  wr_cycle[ 5403] = 1'b0;  addr_rom[ 5403]='h000002bc;  wr_data_rom[ 5403]='h00000000;
    rd_cycle[ 5404] = 1'b1;  wr_cycle[ 5404] = 1'b0;  addr_rom[ 5404]='h00000dbc;  wr_data_rom[ 5404]='h00000000;
    rd_cycle[ 5405] = 1'b0;  wr_cycle[ 5405] = 1'b1;  addr_rom[ 5405]='h00001354;  wr_data_rom[ 5405]='h0000021a;
    rd_cycle[ 5406] = 1'b1;  wr_cycle[ 5406] = 1'b0;  addr_rom[ 5406]='h000009b8;  wr_data_rom[ 5406]='h00000000;
    rd_cycle[ 5407] = 1'b0;  wr_cycle[ 5407] = 1'b1;  addr_rom[ 5407]='h000010c4;  wr_data_rom[ 5407]='h00001991;
    rd_cycle[ 5408] = 1'b0;  wr_cycle[ 5408] = 1'b1;  addr_rom[ 5408]='h00001320;  wr_data_rom[ 5408]='h00000077;
    rd_cycle[ 5409] = 1'b1;  wr_cycle[ 5409] = 1'b0;  addr_rom[ 5409]='h000016a0;  wr_data_rom[ 5409]='h00000000;
    rd_cycle[ 5410] = 1'b0;  wr_cycle[ 5410] = 1'b1;  addr_rom[ 5410]='h000008c8;  wr_data_rom[ 5410]='h00001bbc;
    rd_cycle[ 5411] = 1'b1;  wr_cycle[ 5411] = 1'b0;  addr_rom[ 5411]='h0000072c;  wr_data_rom[ 5411]='h00000000;
    rd_cycle[ 5412] = 1'b1;  wr_cycle[ 5412] = 1'b0;  addr_rom[ 5412]='h000017bc;  wr_data_rom[ 5412]='h00000000;
    rd_cycle[ 5413] = 1'b1;  wr_cycle[ 5413] = 1'b0;  addr_rom[ 5413]='h000014e0;  wr_data_rom[ 5413]='h00000000;
    rd_cycle[ 5414] = 1'b0;  wr_cycle[ 5414] = 1'b1;  addr_rom[ 5414]='h00001d10;  wr_data_rom[ 5414]='h00000f0b;
    rd_cycle[ 5415] = 1'b0;  wr_cycle[ 5415] = 1'b1;  addr_rom[ 5415]='h00001164;  wr_data_rom[ 5415]='h00000753;
    rd_cycle[ 5416] = 1'b0;  wr_cycle[ 5416] = 1'b1;  addr_rom[ 5416]='h000018e8;  wr_data_rom[ 5416]='h00001b18;
    rd_cycle[ 5417] = 1'b1;  wr_cycle[ 5417] = 1'b0;  addr_rom[ 5417]='h00000ac8;  wr_data_rom[ 5417]='h00000000;
    rd_cycle[ 5418] = 1'b1;  wr_cycle[ 5418] = 1'b0;  addr_rom[ 5418]='h00000b8c;  wr_data_rom[ 5418]='h00000000;
    rd_cycle[ 5419] = 1'b1;  wr_cycle[ 5419] = 1'b0;  addr_rom[ 5419]='h000007c8;  wr_data_rom[ 5419]='h00000000;
    rd_cycle[ 5420] = 1'b1;  wr_cycle[ 5420] = 1'b0;  addr_rom[ 5420]='h00001cc8;  wr_data_rom[ 5420]='h00000000;
    rd_cycle[ 5421] = 1'b0;  wr_cycle[ 5421] = 1'b1;  addr_rom[ 5421]='h0000061c;  wr_data_rom[ 5421]='h0000092d;
    rd_cycle[ 5422] = 1'b0;  wr_cycle[ 5422] = 1'b1;  addr_rom[ 5422]='h00001c88;  wr_data_rom[ 5422]='h00001c04;
    rd_cycle[ 5423] = 1'b0;  wr_cycle[ 5423] = 1'b1;  addr_rom[ 5423]='h00001764;  wr_data_rom[ 5423]='h00001ce9;
    rd_cycle[ 5424] = 1'b1;  wr_cycle[ 5424] = 1'b0;  addr_rom[ 5424]='h00001388;  wr_data_rom[ 5424]='h00000000;
    rd_cycle[ 5425] = 1'b1;  wr_cycle[ 5425] = 1'b0;  addr_rom[ 5425]='h00000e80;  wr_data_rom[ 5425]='h00000000;
    rd_cycle[ 5426] = 1'b0;  wr_cycle[ 5426] = 1'b1;  addr_rom[ 5426]='h0000120c;  wr_data_rom[ 5426]='h000019db;
    rd_cycle[ 5427] = 1'b1;  wr_cycle[ 5427] = 1'b0;  addr_rom[ 5427]='h00000810;  wr_data_rom[ 5427]='h00000000;
    rd_cycle[ 5428] = 1'b1;  wr_cycle[ 5428] = 1'b0;  addr_rom[ 5428]='h000007d8;  wr_data_rom[ 5428]='h00000000;
    rd_cycle[ 5429] = 1'b0;  wr_cycle[ 5429] = 1'b1;  addr_rom[ 5429]='h00001044;  wr_data_rom[ 5429]='h00000b2c;
    rd_cycle[ 5430] = 1'b1;  wr_cycle[ 5430] = 1'b0;  addr_rom[ 5430]='h00001398;  wr_data_rom[ 5430]='h00000000;
    rd_cycle[ 5431] = 1'b0;  wr_cycle[ 5431] = 1'b1;  addr_rom[ 5431]='h0000157c;  wr_data_rom[ 5431]='h000018fd;
    rd_cycle[ 5432] = 1'b1;  wr_cycle[ 5432] = 1'b0;  addr_rom[ 5432]='h000004c0;  wr_data_rom[ 5432]='h00000000;
    rd_cycle[ 5433] = 1'b1;  wr_cycle[ 5433] = 1'b0;  addr_rom[ 5433]='h00000d9c;  wr_data_rom[ 5433]='h00000000;
    rd_cycle[ 5434] = 1'b1;  wr_cycle[ 5434] = 1'b0;  addr_rom[ 5434]='h0000070c;  wr_data_rom[ 5434]='h00000000;
    rd_cycle[ 5435] = 1'b0;  wr_cycle[ 5435] = 1'b1;  addr_rom[ 5435]='h000010d4;  wr_data_rom[ 5435]='h00000c82;
    rd_cycle[ 5436] = 1'b0;  wr_cycle[ 5436] = 1'b1;  addr_rom[ 5436]='h00001308;  wr_data_rom[ 5436]='h0000188f;
    rd_cycle[ 5437] = 1'b1;  wr_cycle[ 5437] = 1'b0;  addr_rom[ 5437]='h00001884;  wr_data_rom[ 5437]='h00000000;
    rd_cycle[ 5438] = 1'b1;  wr_cycle[ 5438] = 1'b0;  addr_rom[ 5438]='h0000111c;  wr_data_rom[ 5438]='h00000000;
    rd_cycle[ 5439] = 1'b1;  wr_cycle[ 5439] = 1'b0;  addr_rom[ 5439]='h00000c94;  wr_data_rom[ 5439]='h00000000;
    rd_cycle[ 5440] = 1'b0;  wr_cycle[ 5440] = 1'b1;  addr_rom[ 5440]='h0000070c;  wr_data_rom[ 5440]='h0000056c;
    rd_cycle[ 5441] = 1'b0;  wr_cycle[ 5441] = 1'b1;  addr_rom[ 5441]='h00001548;  wr_data_rom[ 5441]='h00000015;
    rd_cycle[ 5442] = 1'b0;  wr_cycle[ 5442] = 1'b1;  addr_rom[ 5442]='h00001540;  wr_data_rom[ 5442]='h000013e5;
    rd_cycle[ 5443] = 1'b0;  wr_cycle[ 5443] = 1'b1;  addr_rom[ 5443]='h00000054;  wr_data_rom[ 5443]='h000008b8;
    rd_cycle[ 5444] = 1'b1;  wr_cycle[ 5444] = 1'b0;  addr_rom[ 5444]='h00001104;  wr_data_rom[ 5444]='h00000000;
    rd_cycle[ 5445] = 1'b1;  wr_cycle[ 5445] = 1'b0;  addr_rom[ 5445]='h00000560;  wr_data_rom[ 5445]='h00000000;
    rd_cycle[ 5446] = 1'b1;  wr_cycle[ 5446] = 1'b0;  addr_rom[ 5446]='h00001030;  wr_data_rom[ 5446]='h00000000;
    rd_cycle[ 5447] = 1'b1;  wr_cycle[ 5447] = 1'b0;  addr_rom[ 5447]='h00000f98;  wr_data_rom[ 5447]='h00000000;
    rd_cycle[ 5448] = 1'b0;  wr_cycle[ 5448] = 1'b1;  addr_rom[ 5448]='h00001488;  wr_data_rom[ 5448]='h00000a80;
    rd_cycle[ 5449] = 1'b1;  wr_cycle[ 5449] = 1'b0;  addr_rom[ 5449]='h00001078;  wr_data_rom[ 5449]='h00000000;
    rd_cycle[ 5450] = 1'b1;  wr_cycle[ 5450] = 1'b0;  addr_rom[ 5450]='h00000394;  wr_data_rom[ 5450]='h00000000;
    rd_cycle[ 5451] = 1'b1;  wr_cycle[ 5451] = 1'b0;  addr_rom[ 5451]='h00000b64;  wr_data_rom[ 5451]='h00000000;
    rd_cycle[ 5452] = 1'b1;  wr_cycle[ 5452] = 1'b0;  addr_rom[ 5452]='h00000584;  wr_data_rom[ 5452]='h00000000;
    rd_cycle[ 5453] = 1'b1;  wr_cycle[ 5453] = 1'b0;  addr_rom[ 5453]='h0000099c;  wr_data_rom[ 5453]='h00000000;
    rd_cycle[ 5454] = 1'b1;  wr_cycle[ 5454] = 1'b0;  addr_rom[ 5454]='h000007e4;  wr_data_rom[ 5454]='h00000000;
    rd_cycle[ 5455] = 1'b0;  wr_cycle[ 5455] = 1'b1;  addr_rom[ 5455]='h00000d80;  wr_data_rom[ 5455]='h0000020b;
    rd_cycle[ 5456] = 1'b0;  wr_cycle[ 5456] = 1'b1;  addr_rom[ 5456]='h000011a8;  wr_data_rom[ 5456]='h00000cb2;
    rd_cycle[ 5457] = 1'b0;  wr_cycle[ 5457] = 1'b1;  addr_rom[ 5457]='h00000ea0;  wr_data_rom[ 5457]='h000005ec;
    rd_cycle[ 5458] = 1'b1;  wr_cycle[ 5458] = 1'b0;  addr_rom[ 5458]='h00000f98;  wr_data_rom[ 5458]='h00000000;
    rd_cycle[ 5459] = 1'b0;  wr_cycle[ 5459] = 1'b1;  addr_rom[ 5459]='h0000124c;  wr_data_rom[ 5459]='h00000bdb;
    rd_cycle[ 5460] = 1'b0;  wr_cycle[ 5460] = 1'b1;  addr_rom[ 5460]='h00001124;  wr_data_rom[ 5460]='h000019b1;
    rd_cycle[ 5461] = 1'b1;  wr_cycle[ 5461] = 1'b0;  addr_rom[ 5461]='h00001838;  wr_data_rom[ 5461]='h00000000;
    rd_cycle[ 5462] = 1'b1;  wr_cycle[ 5462] = 1'b0;  addr_rom[ 5462]='h00000cbc;  wr_data_rom[ 5462]='h00000000;
    rd_cycle[ 5463] = 1'b0;  wr_cycle[ 5463] = 1'b1;  addr_rom[ 5463]='h000012c4;  wr_data_rom[ 5463]='h00000a1b;
    rd_cycle[ 5464] = 1'b0;  wr_cycle[ 5464] = 1'b1;  addr_rom[ 5464]='h000006b0;  wr_data_rom[ 5464]='h00001119;
    rd_cycle[ 5465] = 1'b1;  wr_cycle[ 5465] = 1'b0;  addr_rom[ 5465]='h000001f4;  wr_data_rom[ 5465]='h00000000;
    rd_cycle[ 5466] = 1'b0;  wr_cycle[ 5466] = 1'b1;  addr_rom[ 5466]='h000001a8;  wr_data_rom[ 5466]='h00001c77;
    rd_cycle[ 5467] = 1'b0;  wr_cycle[ 5467] = 1'b1;  addr_rom[ 5467]='h000011e0;  wr_data_rom[ 5467]='h000002da;
    rd_cycle[ 5468] = 1'b0;  wr_cycle[ 5468] = 1'b1;  addr_rom[ 5468]='h00001328;  wr_data_rom[ 5468]='h00000a79;
    rd_cycle[ 5469] = 1'b0;  wr_cycle[ 5469] = 1'b1;  addr_rom[ 5469]='h00001638;  wr_data_rom[ 5469]='h0000111f;
    rd_cycle[ 5470] = 1'b0;  wr_cycle[ 5470] = 1'b1;  addr_rom[ 5470]='h00001840;  wr_data_rom[ 5470]='h00000285;
    rd_cycle[ 5471] = 1'b0;  wr_cycle[ 5471] = 1'b1;  addr_rom[ 5471]='h00001ec4;  wr_data_rom[ 5471]='h00001339;
    rd_cycle[ 5472] = 1'b1;  wr_cycle[ 5472] = 1'b0;  addr_rom[ 5472]='h000002c0;  wr_data_rom[ 5472]='h00000000;
    rd_cycle[ 5473] = 1'b0;  wr_cycle[ 5473] = 1'b1;  addr_rom[ 5473]='h00001d80;  wr_data_rom[ 5473]='h00001712;
    rd_cycle[ 5474] = 1'b1;  wr_cycle[ 5474] = 1'b0;  addr_rom[ 5474]='h00001088;  wr_data_rom[ 5474]='h00000000;
    rd_cycle[ 5475] = 1'b0;  wr_cycle[ 5475] = 1'b1;  addr_rom[ 5475]='h00001634;  wr_data_rom[ 5475]='h0000005a;
    rd_cycle[ 5476] = 1'b1;  wr_cycle[ 5476] = 1'b0;  addr_rom[ 5476]='h00000354;  wr_data_rom[ 5476]='h00000000;
    rd_cycle[ 5477] = 1'b1;  wr_cycle[ 5477] = 1'b0;  addr_rom[ 5477]='h000013e8;  wr_data_rom[ 5477]='h00000000;
    rd_cycle[ 5478] = 1'b1;  wr_cycle[ 5478] = 1'b0;  addr_rom[ 5478]='h000015a4;  wr_data_rom[ 5478]='h00000000;
    rd_cycle[ 5479] = 1'b1;  wr_cycle[ 5479] = 1'b0;  addr_rom[ 5479]='h00000e60;  wr_data_rom[ 5479]='h00000000;
    rd_cycle[ 5480] = 1'b0;  wr_cycle[ 5480] = 1'b1;  addr_rom[ 5480]='h0000083c;  wr_data_rom[ 5480]='h00000989;
    rd_cycle[ 5481] = 1'b1;  wr_cycle[ 5481] = 1'b0;  addr_rom[ 5481]='h00001224;  wr_data_rom[ 5481]='h00000000;
    rd_cycle[ 5482] = 1'b1;  wr_cycle[ 5482] = 1'b0;  addr_rom[ 5482]='h00001668;  wr_data_rom[ 5482]='h00000000;
    rd_cycle[ 5483] = 1'b0;  wr_cycle[ 5483] = 1'b1;  addr_rom[ 5483]='h0000193c;  wr_data_rom[ 5483]='h000019ba;
    rd_cycle[ 5484] = 1'b1;  wr_cycle[ 5484] = 1'b0;  addr_rom[ 5484]='h00000d5c;  wr_data_rom[ 5484]='h00000000;
    rd_cycle[ 5485] = 1'b1;  wr_cycle[ 5485] = 1'b0;  addr_rom[ 5485]='h00001914;  wr_data_rom[ 5485]='h00000000;
    rd_cycle[ 5486] = 1'b1;  wr_cycle[ 5486] = 1'b0;  addr_rom[ 5486]='h00000090;  wr_data_rom[ 5486]='h00000000;
    rd_cycle[ 5487] = 1'b1;  wr_cycle[ 5487] = 1'b0;  addr_rom[ 5487]='h00001b54;  wr_data_rom[ 5487]='h00000000;
    rd_cycle[ 5488] = 1'b1;  wr_cycle[ 5488] = 1'b0;  addr_rom[ 5488]='h00001c80;  wr_data_rom[ 5488]='h00000000;
    rd_cycle[ 5489] = 1'b0;  wr_cycle[ 5489] = 1'b1;  addr_rom[ 5489]='h00001004;  wr_data_rom[ 5489]='h00001006;
    rd_cycle[ 5490] = 1'b0;  wr_cycle[ 5490] = 1'b1;  addr_rom[ 5490]='h000008f0;  wr_data_rom[ 5490]='h000016ca;
    rd_cycle[ 5491] = 1'b1;  wr_cycle[ 5491] = 1'b0;  addr_rom[ 5491]='h00001674;  wr_data_rom[ 5491]='h00000000;
    rd_cycle[ 5492] = 1'b1;  wr_cycle[ 5492] = 1'b0;  addr_rom[ 5492]='h00000ec8;  wr_data_rom[ 5492]='h00000000;
    rd_cycle[ 5493] = 1'b1;  wr_cycle[ 5493] = 1'b0;  addr_rom[ 5493]='h0000177c;  wr_data_rom[ 5493]='h00000000;
    rd_cycle[ 5494] = 1'b0;  wr_cycle[ 5494] = 1'b1;  addr_rom[ 5494]='h000015f8;  wr_data_rom[ 5494]='h00000a80;
    rd_cycle[ 5495] = 1'b0;  wr_cycle[ 5495] = 1'b1;  addr_rom[ 5495]='h000003c8;  wr_data_rom[ 5495]='h00000462;
    rd_cycle[ 5496] = 1'b0;  wr_cycle[ 5496] = 1'b1;  addr_rom[ 5496]='h00001020;  wr_data_rom[ 5496]='h00000779;
    rd_cycle[ 5497] = 1'b0;  wr_cycle[ 5497] = 1'b1;  addr_rom[ 5497]='h000017e8;  wr_data_rom[ 5497]='h000012e3;
    rd_cycle[ 5498] = 1'b1;  wr_cycle[ 5498] = 1'b0;  addr_rom[ 5498]='h00001e6c;  wr_data_rom[ 5498]='h00000000;
    rd_cycle[ 5499] = 1'b1;  wr_cycle[ 5499] = 1'b0;  addr_rom[ 5499]='h0000022c;  wr_data_rom[ 5499]='h00000000;
    rd_cycle[ 5500] = 1'b0;  wr_cycle[ 5500] = 1'b1;  addr_rom[ 5500]='h000013ac;  wr_data_rom[ 5500]='h00001b07;
    rd_cycle[ 5501] = 1'b0;  wr_cycle[ 5501] = 1'b1;  addr_rom[ 5501]='h0000011c;  wr_data_rom[ 5501]='h00000fd5;
    rd_cycle[ 5502] = 1'b0;  wr_cycle[ 5502] = 1'b1;  addr_rom[ 5502]='h00001be8;  wr_data_rom[ 5502]='h00000ac4;
    rd_cycle[ 5503] = 1'b0;  wr_cycle[ 5503] = 1'b1;  addr_rom[ 5503]='h00001c24;  wr_data_rom[ 5503]='h00000068;
    rd_cycle[ 5504] = 1'b1;  wr_cycle[ 5504] = 1'b0;  addr_rom[ 5504]='h000011e0;  wr_data_rom[ 5504]='h00000000;
    rd_cycle[ 5505] = 1'b0;  wr_cycle[ 5505] = 1'b1;  addr_rom[ 5505]='h0000085c;  wr_data_rom[ 5505]='h00000eb8;
    rd_cycle[ 5506] = 1'b0;  wr_cycle[ 5506] = 1'b1;  addr_rom[ 5506]='h000003b0;  wr_data_rom[ 5506]='h000008d8;
    rd_cycle[ 5507] = 1'b0;  wr_cycle[ 5507] = 1'b1;  addr_rom[ 5507]='h0000049c;  wr_data_rom[ 5507]='h000010a4;
    rd_cycle[ 5508] = 1'b1;  wr_cycle[ 5508] = 1'b0;  addr_rom[ 5508]='h000010d8;  wr_data_rom[ 5508]='h00000000;
    rd_cycle[ 5509] = 1'b1;  wr_cycle[ 5509] = 1'b0;  addr_rom[ 5509]='h00000a40;  wr_data_rom[ 5509]='h00000000;
    rd_cycle[ 5510] = 1'b1;  wr_cycle[ 5510] = 1'b0;  addr_rom[ 5510]='h00001108;  wr_data_rom[ 5510]='h00000000;
    rd_cycle[ 5511] = 1'b0;  wr_cycle[ 5511] = 1'b1;  addr_rom[ 5511]='h000002bc;  wr_data_rom[ 5511]='h00000684;
    rd_cycle[ 5512] = 1'b1;  wr_cycle[ 5512] = 1'b0;  addr_rom[ 5512]='h00000404;  wr_data_rom[ 5512]='h00000000;
    rd_cycle[ 5513] = 1'b0;  wr_cycle[ 5513] = 1'b1;  addr_rom[ 5513]='h000001d0;  wr_data_rom[ 5513]='h00001599;
    rd_cycle[ 5514] = 1'b0;  wr_cycle[ 5514] = 1'b1;  addr_rom[ 5514]='h000012a0;  wr_data_rom[ 5514]='h000019be;
    rd_cycle[ 5515] = 1'b1;  wr_cycle[ 5515] = 1'b0;  addr_rom[ 5515]='h0000114c;  wr_data_rom[ 5515]='h00000000;
    rd_cycle[ 5516] = 1'b0;  wr_cycle[ 5516] = 1'b1;  addr_rom[ 5516]='h00001984;  wr_data_rom[ 5516]='h0000174e;
    rd_cycle[ 5517] = 1'b0;  wr_cycle[ 5517] = 1'b1;  addr_rom[ 5517]='h00001538;  wr_data_rom[ 5517]='h00000b6f;
    rd_cycle[ 5518] = 1'b0;  wr_cycle[ 5518] = 1'b1;  addr_rom[ 5518]='h00001e78;  wr_data_rom[ 5518]='h00001426;
    rd_cycle[ 5519] = 1'b0;  wr_cycle[ 5519] = 1'b1;  addr_rom[ 5519]='h000006f0;  wr_data_rom[ 5519]='h000016ad;
    rd_cycle[ 5520] = 1'b1;  wr_cycle[ 5520] = 1'b0;  addr_rom[ 5520]='h00000b20;  wr_data_rom[ 5520]='h00000000;
    rd_cycle[ 5521] = 1'b0;  wr_cycle[ 5521] = 1'b1;  addr_rom[ 5521]='h000004c4;  wr_data_rom[ 5521]='h00001cc3;
    rd_cycle[ 5522] = 1'b0;  wr_cycle[ 5522] = 1'b1;  addr_rom[ 5522]='h00000fb0;  wr_data_rom[ 5522]='h000003cf;
    rd_cycle[ 5523] = 1'b1;  wr_cycle[ 5523] = 1'b0;  addr_rom[ 5523]='h00001d10;  wr_data_rom[ 5523]='h00000000;
    rd_cycle[ 5524] = 1'b0;  wr_cycle[ 5524] = 1'b1;  addr_rom[ 5524]='h00001d6c;  wr_data_rom[ 5524]='h00001828;
    rd_cycle[ 5525] = 1'b1;  wr_cycle[ 5525] = 1'b0;  addr_rom[ 5525]='h00001510;  wr_data_rom[ 5525]='h00000000;
    rd_cycle[ 5526] = 1'b0;  wr_cycle[ 5526] = 1'b1;  addr_rom[ 5526]='h00000dd4;  wr_data_rom[ 5526]='h000008ec;
    rd_cycle[ 5527] = 1'b0;  wr_cycle[ 5527] = 1'b1;  addr_rom[ 5527]='h00001710;  wr_data_rom[ 5527]='h00001ef8;
    rd_cycle[ 5528] = 1'b0;  wr_cycle[ 5528] = 1'b1;  addr_rom[ 5528]='h00001e50;  wr_data_rom[ 5528]='h00001c70;
    rd_cycle[ 5529] = 1'b1;  wr_cycle[ 5529] = 1'b0;  addr_rom[ 5529]='h00000204;  wr_data_rom[ 5529]='h00000000;
    rd_cycle[ 5530] = 1'b1;  wr_cycle[ 5530] = 1'b0;  addr_rom[ 5530]='h000011e8;  wr_data_rom[ 5530]='h00000000;
    rd_cycle[ 5531] = 1'b0;  wr_cycle[ 5531] = 1'b1;  addr_rom[ 5531]='h00000a04;  wr_data_rom[ 5531]='h00000aee;
    rd_cycle[ 5532] = 1'b1;  wr_cycle[ 5532] = 1'b0;  addr_rom[ 5532]='h000017c0;  wr_data_rom[ 5532]='h00000000;
    rd_cycle[ 5533] = 1'b0;  wr_cycle[ 5533] = 1'b1;  addr_rom[ 5533]='h00000b78;  wr_data_rom[ 5533]='h0000147e;
    rd_cycle[ 5534] = 1'b0;  wr_cycle[ 5534] = 1'b1;  addr_rom[ 5534]='h00001618;  wr_data_rom[ 5534]='h00000755;
    rd_cycle[ 5535] = 1'b0;  wr_cycle[ 5535] = 1'b1;  addr_rom[ 5535]='h00001060;  wr_data_rom[ 5535]='h000018de;
    rd_cycle[ 5536] = 1'b1;  wr_cycle[ 5536] = 1'b0;  addr_rom[ 5536]='h00001a28;  wr_data_rom[ 5536]='h00000000;
    rd_cycle[ 5537] = 1'b1;  wr_cycle[ 5537] = 1'b0;  addr_rom[ 5537]='h00001f1c;  wr_data_rom[ 5537]='h00000000;
    rd_cycle[ 5538] = 1'b1;  wr_cycle[ 5538] = 1'b0;  addr_rom[ 5538]='h00000998;  wr_data_rom[ 5538]='h00000000;
    rd_cycle[ 5539] = 1'b1;  wr_cycle[ 5539] = 1'b0;  addr_rom[ 5539]='h00001d30;  wr_data_rom[ 5539]='h00000000;
    rd_cycle[ 5540] = 1'b0;  wr_cycle[ 5540] = 1'b1;  addr_rom[ 5540]='h00000d24;  wr_data_rom[ 5540]='h00000ae8;
    rd_cycle[ 5541] = 1'b0;  wr_cycle[ 5541] = 1'b1;  addr_rom[ 5541]='h00001484;  wr_data_rom[ 5541]='h00000536;
    rd_cycle[ 5542] = 1'b0;  wr_cycle[ 5542] = 1'b1;  addr_rom[ 5542]='h00001730;  wr_data_rom[ 5542]='h00001391;
    rd_cycle[ 5543] = 1'b1;  wr_cycle[ 5543] = 1'b0;  addr_rom[ 5543]='h00000994;  wr_data_rom[ 5543]='h00000000;
    rd_cycle[ 5544] = 1'b1;  wr_cycle[ 5544] = 1'b0;  addr_rom[ 5544]='h00000a30;  wr_data_rom[ 5544]='h00000000;
    rd_cycle[ 5545] = 1'b0;  wr_cycle[ 5545] = 1'b1;  addr_rom[ 5545]='h00001460;  wr_data_rom[ 5545]='h00000192;
    rd_cycle[ 5546] = 1'b1;  wr_cycle[ 5546] = 1'b0;  addr_rom[ 5546]='h00001bd4;  wr_data_rom[ 5546]='h00000000;
    rd_cycle[ 5547] = 1'b1;  wr_cycle[ 5547] = 1'b0;  addr_rom[ 5547]='h00001a40;  wr_data_rom[ 5547]='h00000000;
    rd_cycle[ 5548] = 1'b1;  wr_cycle[ 5548] = 1'b0;  addr_rom[ 5548]='h0000092c;  wr_data_rom[ 5548]='h00000000;
    rd_cycle[ 5549] = 1'b0;  wr_cycle[ 5549] = 1'b1;  addr_rom[ 5549]='h00000bc8;  wr_data_rom[ 5549]='h00001e30;
    rd_cycle[ 5550] = 1'b1;  wr_cycle[ 5550] = 1'b0;  addr_rom[ 5550]='h0000191c;  wr_data_rom[ 5550]='h00000000;
    rd_cycle[ 5551] = 1'b0;  wr_cycle[ 5551] = 1'b1;  addr_rom[ 5551]='h00001b7c;  wr_data_rom[ 5551]='h000013c8;
    rd_cycle[ 5552] = 1'b0;  wr_cycle[ 5552] = 1'b1;  addr_rom[ 5552]='h00001ae4;  wr_data_rom[ 5552]='h000017d3;
    rd_cycle[ 5553] = 1'b1;  wr_cycle[ 5553] = 1'b0;  addr_rom[ 5553]='h0000192c;  wr_data_rom[ 5553]='h00000000;
    rd_cycle[ 5554] = 1'b0;  wr_cycle[ 5554] = 1'b1;  addr_rom[ 5554]='h000019b4;  wr_data_rom[ 5554]='h00000d7f;
    rd_cycle[ 5555] = 1'b0;  wr_cycle[ 5555] = 1'b1;  addr_rom[ 5555]='h000016b4;  wr_data_rom[ 5555]='h00000ac9;
    rd_cycle[ 5556] = 1'b0;  wr_cycle[ 5556] = 1'b1;  addr_rom[ 5556]='h000013bc;  wr_data_rom[ 5556]='h000000b7;
    rd_cycle[ 5557] = 1'b0;  wr_cycle[ 5557] = 1'b1;  addr_rom[ 5557]='h000019c4;  wr_data_rom[ 5557]='h000005f5;
    rd_cycle[ 5558] = 1'b0;  wr_cycle[ 5558] = 1'b1;  addr_rom[ 5558]='h00001e5c;  wr_data_rom[ 5558]='h000006fa;
    rd_cycle[ 5559] = 1'b0;  wr_cycle[ 5559] = 1'b1;  addr_rom[ 5559]='h00001e3c;  wr_data_rom[ 5559]='h0000031d;
    rd_cycle[ 5560] = 1'b0;  wr_cycle[ 5560] = 1'b1;  addr_rom[ 5560]='h00001b9c;  wr_data_rom[ 5560]='h00001cea;
    rd_cycle[ 5561] = 1'b1;  wr_cycle[ 5561] = 1'b0;  addr_rom[ 5561]='h00001b94;  wr_data_rom[ 5561]='h00000000;
    rd_cycle[ 5562] = 1'b1;  wr_cycle[ 5562] = 1'b0;  addr_rom[ 5562]='h00000764;  wr_data_rom[ 5562]='h00000000;
    rd_cycle[ 5563] = 1'b1;  wr_cycle[ 5563] = 1'b0;  addr_rom[ 5563]='h00000228;  wr_data_rom[ 5563]='h00000000;
    rd_cycle[ 5564] = 1'b1;  wr_cycle[ 5564] = 1'b0;  addr_rom[ 5564]='h000005f8;  wr_data_rom[ 5564]='h00000000;
    rd_cycle[ 5565] = 1'b0;  wr_cycle[ 5565] = 1'b1;  addr_rom[ 5565]='h00000fec;  wr_data_rom[ 5565]='h000015a8;
    rd_cycle[ 5566] = 1'b0;  wr_cycle[ 5566] = 1'b1;  addr_rom[ 5566]='h0000144c;  wr_data_rom[ 5566]='h000019a6;
    rd_cycle[ 5567] = 1'b1;  wr_cycle[ 5567] = 1'b0;  addr_rom[ 5567]='h00000acc;  wr_data_rom[ 5567]='h00000000;
    rd_cycle[ 5568] = 1'b1;  wr_cycle[ 5568] = 1'b0;  addr_rom[ 5568]='h00000074;  wr_data_rom[ 5568]='h00000000;
    rd_cycle[ 5569] = 1'b1;  wr_cycle[ 5569] = 1'b0;  addr_rom[ 5569]='h00001240;  wr_data_rom[ 5569]='h00000000;
    rd_cycle[ 5570] = 1'b1;  wr_cycle[ 5570] = 1'b0;  addr_rom[ 5570]='h000017e4;  wr_data_rom[ 5570]='h00000000;
    rd_cycle[ 5571] = 1'b1;  wr_cycle[ 5571] = 1'b0;  addr_rom[ 5571]='h00001e20;  wr_data_rom[ 5571]='h00000000;
    rd_cycle[ 5572] = 1'b1;  wr_cycle[ 5572] = 1'b0;  addr_rom[ 5572]='h000000f0;  wr_data_rom[ 5572]='h00000000;
    rd_cycle[ 5573] = 1'b0;  wr_cycle[ 5573] = 1'b1;  addr_rom[ 5573]='h000015f8;  wr_data_rom[ 5573]='h0000061a;
    rd_cycle[ 5574] = 1'b0;  wr_cycle[ 5574] = 1'b1;  addr_rom[ 5574]='h00001b24;  wr_data_rom[ 5574]='h000011f2;
    rd_cycle[ 5575] = 1'b1;  wr_cycle[ 5575] = 1'b0;  addr_rom[ 5575]='h00001140;  wr_data_rom[ 5575]='h00000000;
    rd_cycle[ 5576] = 1'b0;  wr_cycle[ 5576] = 1'b1;  addr_rom[ 5576]='h00000eec;  wr_data_rom[ 5576]='h0000082a;
    rd_cycle[ 5577] = 1'b1;  wr_cycle[ 5577] = 1'b0;  addr_rom[ 5577]='h000000cc;  wr_data_rom[ 5577]='h00000000;
    rd_cycle[ 5578] = 1'b0;  wr_cycle[ 5578] = 1'b1;  addr_rom[ 5578]='h00001974;  wr_data_rom[ 5578]='h00001d95;
    rd_cycle[ 5579] = 1'b0;  wr_cycle[ 5579] = 1'b1;  addr_rom[ 5579]='h000001c0;  wr_data_rom[ 5579]='h000009ec;
    rd_cycle[ 5580] = 1'b1;  wr_cycle[ 5580] = 1'b0;  addr_rom[ 5580]='h00001724;  wr_data_rom[ 5580]='h00000000;
    rd_cycle[ 5581] = 1'b0;  wr_cycle[ 5581] = 1'b1;  addr_rom[ 5581]='h000010d4;  wr_data_rom[ 5581]='h00001ccd;
    rd_cycle[ 5582] = 1'b0;  wr_cycle[ 5582] = 1'b1;  addr_rom[ 5582]='h00001008;  wr_data_rom[ 5582]='h00001e2f;
    rd_cycle[ 5583] = 1'b1;  wr_cycle[ 5583] = 1'b0;  addr_rom[ 5583]='h00000f0c;  wr_data_rom[ 5583]='h00000000;
    rd_cycle[ 5584] = 1'b0;  wr_cycle[ 5584] = 1'b1;  addr_rom[ 5584]='h000010f0;  wr_data_rom[ 5584]='h00000c8a;
    rd_cycle[ 5585] = 1'b1;  wr_cycle[ 5585] = 1'b0;  addr_rom[ 5585]='h00000a98;  wr_data_rom[ 5585]='h00000000;
    rd_cycle[ 5586] = 1'b0;  wr_cycle[ 5586] = 1'b1;  addr_rom[ 5586]='h00001af0;  wr_data_rom[ 5586]='h00001dcf;
    rd_cycle[ 5587] = 1'b0;  wr_cycle[ 5587] = 1'b1;  addr_rom[ 5587]='h0000163c;  wr_data_rom[ 5587]='h0000084b;
    rd_cycle[ 5588] = 1'b1;  wr_cycle[ 5588] = 1'b0;  addr_rom[ 5588]='h0000149c;  wr_data_rom[ 5588]='h00000000;
    rd_cycle[ 5589] = 1'b1;  wr_cycle[ 5589] = 1'b0;  addr_rom[ 5589]='h0000000c;  wr_data_rom[ 5589]='h00000000;
    rd_cycle[ 5590] = 1'b0;  wr_cycle[ 5590] = 1'b1;  addr_rom[ 5590]='h00000bf0;  wr_data_rom[ 5590]='h00000779;
    rd_cycle[ 5591] = 1'b1;  wr_cycle[ 5591] = 1'b0;  addr_rom[ 5591]='h000003d4;  wr_data_rom[ 5591]='h00000000;
    rd_cycle[ 5592] = 1'b1;  wr_cycle[ 5592] = 1'b0;  addr_rom[ 5592]='h00001ef8;  wr_data_rom[ 5592]='h00000000;
    rd_cycle[ 5593] = 1'b0;  wr_cycle[ 5593] = 1'b1;  addr_rom[ 5593]='h000014c0;  wr_data_rom[ 5593]='h000010bb;
    rd_cycle[ 5594] = 1'b1;  wr_cycle[ 5594] = 1'b0;  addr_rom[ 5594]='h000002bc;  wr_data_rom[ 5594]='h00000000;
    rd_cycle[ 5595] = 1'b1;  wr_cycle[ 5595] = 1'b0;  addr_rom[ 5595]='h00000818;  wr_data_rom[ 5595]='h00000000;
    rd_cycle[ 5596] = 1'b1;  wr_cycle[ 5596] = 1'b0;  addr_rom[ 5596]='h000018a8;  wr_data_rom[ 5596]='h00000000;
    rd_cycle[ 5597] = 1'b0;  wr_cycle[ 5597] = 1'b1;  addr_rom[ 5597]='h00000ecc;  wr_data_rom[ 5597]='h0000018b;
    rd_cycle[ 5598] = 1'b1;  wr_cycle[ 5598] = 1'b0;  addr_rom[ 5598]='h00000a34;  wr_data_rom[ 5598]='h00000000;
    rd_cycle[ 5599] = 1'b0;  wr_cycle[ 5599] = 1'b1;  addr_rom[ 5599]='h00001a88;  wr_data_rom[ 5599]='h0000022a;
    rd_cycle[ 5600] = 1'b0;  wr_cycle[ 5600] = 1'b1;  addr_rom[ 5600]='h00001424;  wr_data_rom[ 5600]='h000009dc;
    rd_cycle[ 5601] = 1'b0;  wr_cycle[ 5601] = 1'b1;  addr_rom[ 5601]='h000014cc;  wr_data_rom[ 5601]='h00000f9a;
    rd_cycle[ 5602] = 1'b0;  wr_cycle[ 5602] = 1'b1;  addr_rom[ 5602]='h00001ecc;  wr_data_rom[ 5602]='h00001793;
    rd_cycle[ 5603] = 1'b0;  wr_cycle[ 5603] = 1'b1;  addr_rom[ 5603]='h00001970;  wr_data_rom[ 5603]='h00000319;
    rd_cycle[ 5604] = 1'b0;  wr_cycle[ 5604] = 1'b1;  addr_rom[ 5604]='h00001bd8;  wr_data_rom[ 5604]='h0000149e;
    rd_cycle[ 5605] = 1'b1;  wr_cycle[ 5605] = 1'b0;  addr_rom[ 5605]='h00000cc8;  wr_data_rom[ 5605]='h00000000;
    rd_cycle[ 5606] = 1'b0;  wr_cycle[ 5606] = 1'b1;  addr_rom[ 5606]='h00001864;  wr_data_rom[ 5606]='h00000b33;
    rd_cycle[ 5607] = 1'b0;  wr_cycle[ 5607] = 1'b1;  addr_rom[ 5607]='h00000cdc;  wr_data_rom[ 5607]='h000010ba;
    rd_cycle[ 5608] = 1'b1;  wr_cycle[ 5608] = 1'b0;  addr_rom[ 5608]='h0000021c;  wr_data_rom[ 5608]='h00000000;
    rd_cycle[ 5609] = 1'b0;  wr_cycle[ 5609] = 1'b1;  addr_rom[ 5609]='h00001c50;  wr_data_rom[ 5609]='h00000ff7;
    rd_cycle[ 5610] = 1'b0;  wr_cycle[ 5610] = 1'b1;  addr_rom[ 5610]='h00000700;  wr_data_rom[ 5610]='h00001dbd;
    rd_cycle[ 5611] = 1'b0;  wr_cycle[ 5611] = 1'b1;  addr_rom[ 5611]='h00001188;  wr_data_rom[ 5611]='h0000101d;
    rd_cycle[ 5612] = 1'b1;  wr_cycle[ 5612] = 1'b0;  addr_rom[ 5612]='h00000a9c;  wr_data_rom[ 5612]='h00000000;
    rd_cycle[ 5613] = 1'b1;  wr_cycle[ 5613] = 1'b0;  addr_rom[ 5613]='h00000c70;  wr_data_rom[ 5613]='h00000000;
    rd_cycle[ 5614] = 1'b0;  wr_cycle[ 5614] = 1'b1;  addr_rom[ 5614]='h00001290;  wr_data_rom[ 5614]='h000010d3;
    rd_cycle[ 5615] = 1'b1;  wr_cycle[ 5615] = 1'b0;  addr_rom[ 5615]='h00000944;  wr_data_rom[ 5615]='h00000000;
    rd_cycle[ 5616] = 1'b0;  wr_cycle[ 5616] = 1'b1;  addr_rom[ 5616]='h0000109c;  wr_data_rom[ 5616]='h00001a2b;
    rd_cycle[ 5617] = 1'b1;  wr_cycle[ 5617] = 1'b0;  addr_rom[ 5617]='h00001b50;  wr_data_rom[ 5617]='h00000000;
    rd_cycle[ 5618] = 1'b1;  wr_cycle[ 5618] = 1'b0;  addr_rom[ 5618]='h00001ed0;  wr_data_rom[ 5618]='h00000000;
    rd_cycle[ 5619] = 1'b1;  wr_cycle[ 5619] = 1'b0;  addr_rom[ 5619]='h000012b8;  wr_data_rom[ 5619]='h00000000;
    rd_cycle[ 5620] = 1'b0;  wr_cycle[ 5620] = 1'b1;  addr_rom[ 5620]='h00001a88;  wr_data_rom[ 5620]='h00000f8e;
    rd_cycle[ 5621] = 1'b1;  wr_cycle[ 5621] = 1'b0;  addr_rom[ 5621]='h00000154;  wr_data_rom[ 5621]='h00000000;
    rd_cycle[ 5622] = 1'b0;  wr_cycle[ 5622] = 1'b1;  addr_rom[ 5622]='h00000d58;  wr_data_rom[ 5622]='h00000237;
    rd_cycle[ 5623] = 1'b1;  wr_cycle[ 5623] = 1'b0;  addr_rom[ 5623]='h000001fc;  wr_data_rom[ 5623]='h00000000;
    rd_cycle[ 5624] = 1'b0;  wr_cycle[ 5624] = 1'b1;  addr_rom[ 5624]='h00000200;  wr_data_rom[ 5624]='h00000003;
    rd_cycle[ 5625] = 1'b1;  wr_cycle[ 5625] = 1'b0;  addr_rom[ 5625]='h0000124c;  wr_data_rom[ 5625]='h00000000;
    rd_cycle[ 5626] = 1'b0;  wr_cycle[ 5626] = 1'b1;  addr_rom[ 5626]='h0000140c;  wr_data_rom[ 5626]='h000008e3;
    rd_cycle[ 5627] = 1'b0;  wr_cycle[ 5627] = 1'b1;  addr_rom[ 5627]='h000010c8;  wr_data_rom[ 5627]='h00000195;
    rd_cycle[ 5628] = 1'b1;  wr_cycle[ 5628] = 1'b0;  addr_rom[ 5628]='h00001578;  wr_data_rom[ 5628]='h00000000;
    rd_cycle[ 5629] = 1'b1;  wr_cycle[ 5629] = 1'b0;  addr_rom[ 5629]='h00000728;  wr_data_rom[ 5629]='h00000000;
    rd_cycle[ 5630] = 1'b0;  wr_cycle[ 5630] = 1'b1;  addr_rom[ 5630]='h00001978;  wr_data_rom[ 5630]='h00001c32;
    rd_cycle[ 5631] = 1'b0;  wr_cycle[ 5631] = 1'b1;  addr_rom[ 5631]='h00001860;  wr_data_rom[ 5631]='h00000028;
    rd_cycle[ 5632] = 1'b1;  wr_cycle[ 5632] = 1'b0;  addr_rom[ 5632]='h000003f8;  wr_data_rom[ 5632]='h00000000;
    rd_cycle[ 5633] = 1'b0;  wr_cycle[ 5633] = 1'b1;  addr_rom[ 5633]='h00000f28;  wr_data_rom[ 5633]='h00000c66;
    rd_cycle[ 5634] = 1'b0;  wr_cycle[ 5634] = 1'b1;  addr_rom[ 5634]='h00000b2c;  wr_data_rom[ 5634]='h000007b1;
    rd_cycle[ 5635] = 1'b0;  wr_cycle[ 5635] = 1'b1;  addr_rom[ 5635]='h000001b4;  wr_data_rom[ 5635]='h0000058b;
    rd_cycle[ 5636] = 1'b0;  wr_cycle[ 5636] = 1'b1;  addr_rom[ 5636]='h000011c8;  wr_data_rom[ 5636]='h000006db;
    rd_cycle[ 5637] = 1'b1;  wr_cycle[ 5637] = 1'b0;  addr_rom[ 5637]='h00000e88;  wr_data_rom[ 5637]='h00000000;
    rd_cycle[ 5638] = 1'b1;  wr_cycle[ 5638] = 1'b0;  addr_rom[ 5638]='h000003bc;  wr_data_rom[ 5638]='h00000000;
    rd_cycle[ 5639] = 1'b1;  wr_cycle[ 5639] = 1'b0;  addr_rom[ 5639]='h00000ec0;  wr_data_rom[ 5639]='h00000000;
    rd_cycle[ 5640] = 1'b1;  wr_cycle[ 5640] = 1'b0;  addr_rom[ 5640]='h000015e4;  wr_data_rom[ 5640]='h00000000;
    rd_cycle[ 5641] = 1'b1;  wr_cycle[ 5641] = 1'b0;  addr_rom[ 5641]='h000010a8;  wr_data_rom[ 5641]='h00000000;
    rd_cycle[ 5642] = 1'b0;  wr_cycle[ 5642] = 1'b1;  addr_rom[ 5642]='h00001ee8;  wr_data_rom[ 5642]='h000000c5;
    rd_cycle[ 5643] = 1'b0;  wr_cycle[ 5643] = 1'b1;  addr_rom[ 5643]='h00000c4c;  wr_data_rom[ 5643]='h000011b4;
    rd_cycle[ 5644] = 1'b1;  wr_cycle[ 5644] = 1'b0;  addr_rom[ 5644]='h000013e0;  wr_data_rom[ 5644]='h00000000;
    rd_cycle[ 5645] = 1'b0;  wr_cycle[ 5645] = 1'b1;  addr_rom[ 5645]='h00000d28;  wr_data_rom[ 5645]='h0000169d;
    rd_cycle[ 5646] = 1'b1;  wr_cycle[ 5646] = 1'b0;  addr_rom[ 5646]='h00001af8;  wr_data_rom[ 5646]='h00000000;
    rd_cycle[ 5647] = 1'b0;  wr_cycle[ 5647] = 1'b1;  addr_rom[ 5647]='h000019b0;  wr_data_rom[ 5647]='h00001f0c;
    rd_cycle[ 5648] = 1'b1;  wr_cycle[ 5648] = 1'b0;  addr_rom[ 5648]='h00000e2c;  wr_data_rom[ 5648]='h00000000;
    rd_cycle[ 5649] = 1'b1;  wr_cycle[ 5649] = 1'b0;  addr_rom[ 5649]='h000012a0;  wr_data_rom[ 5649]='h00000000;
    rd_cycle[ 5650] = 1'b0;  wr_cycle[ 5650] = 1'b1;  addr_rom[ 5650]='h00001090;  wr_data_rom[ 5650]='h00001559;
    rd_cycle[ 5651] = 1'b1;  wr_cycle[ 5651] = 1'b0;  addr_rom[ 5651]='h000011dc;  wr_data_rom[ 5651]='h00000000;
    rd_cycle[ 5652] = 1'b1;  wr_cycle[ 5652] = 1'b0;  addr_rom[ 5652]='h00001730;  wr_data_rom[ 5652]='h00000000;
    rd_cycle[ 5653] = 1'b0;  wr_cycle[ 5653] = 1'b1;  addr_rom[ 5653]='h00001400;  wr_data_rom[ 5653]='h00001ddd;
    rd_cycle[ 5654] = 1'b1;  wr_cycle[ 5654] = 1'b0;  addr_rom[ 5654]='h00001848;  wr_data_rom[ 5654]='h00000000;
    rd_cycle[ 5655] = 1'b0;  wr_cycle[ 5655] = 1'b1;  addr_rom[ 5655]='h00001904;  wr_data_rom[ 5655]='h00001590;
    rd_cycle[ 5656] = 1'b1;  wr_cycle[ 5656] = 1'b0;  addr_rom[ 5656]='h00000678;  wr_data_rom[ 5656]='h00000000;
    rd_cycle[ 5657] = 1'b0;  wr_cycle[ 5657] = 1'b1;  addr_rom[ 5657]='h00000d94;  wr_data_rom[ 5657]='h00000786;
    rd_cycle[ 5658] = 1'b0;  wr_cycle[ 5658] = 1'b1;  addr_rom[ 5658]='h00001630;  wr_data_rom[ 5658]='h00001878;
    rd_cycle[ 5659] = 1'b1;  wr_cycle[ 5659] = 1'b0;  addr_rom[ 5659]='h000010c0;  wr_data_rom[ 5659]='h00000000;
    rd_cycle[ 5660] = 1'b1;  wr_cycle[ 5660] = 1'b0;  addr_rom[ 5660]='h00001cdc;  wr_data_rom[ 5660]='h00000000;
    rd_cycle[ 5661] = 1'b0;  wr_cycle[ 5661] = 1'b1;  addr_rom[ 5661]='h000000dc;  wr_data_rom[ 5661]='h00000107;
    rd_cycle[ 5662] = 1'b0;  wr_cycle[ 5662] = 1'b1;  addr_rom[ 5662]='h00000478;  wr_data_rom[ 5662]='h00000f1c;
    rd_cycle[ 5663] = 1'b0;  wr_cycle[ 5663] = 1'b1;  addr_rom[ 5663]='h00001a9c;  wr_data_rom[ 5663]='h00001249;
    rd_cycle[ 5664] = 1'b1;  wr_cycle[ 5664] = 1'b0;  addr_rom[ 5664]='h0000089c;  wr_data_rom[ 5664]='h00000000;
    rd_cycle[ 5665] = 1'b1;  wr_cycle[ 5665] = 1'b0;  addr_rom[ 5665]='h00000e74;  wr_data_rom[ 5665]='h00000000;
    rd_cycle[ 5666] = 1'b0;  wr_cycle[ 5666] = 1'b1;  addr_rom[ 5666]='h00001448;  wr_data_rom[ 5666]='h000012b0;
    rd_cycle[ 5667] = 1'b0;  wr_cycle[ 5667] = 1'b1;  addr_rom[ 5667]='h000011a8;  wr_data_rom[ 5667]='h00000dbc;
    rd_cycle[ 5668] = 1'b0;  wr_cycle[ 5668] = 1'b1;  addr_rom[ 5668]='h00001758;  wr_data_rom[ 5668]='h00000021;
    rd_cycle[ 5669] = 1'b1;  wr_cycle[ 5669] = 1'b0;  addr_rom[ 5669]='h00000c98;  wr_data_rom[ 5669]='h00000000;
    rd_cycle[ 5670] = 1'b1;  wr_cycle[ 5670] = 1'b0;  addr_rom[ 5670]='h00000854;  wr_data_rom[ 5670]='h00000000;
    rd_cycle[ 5671] = 1'b0;  wr_cycle[ 5671] = 1'b1;  addr_rom[ 5671]='h000012c4;  wr_data_rom[ 5671]='h00001e2c;
    rd_cycle[ 5672] = 1'b0;  wr_cycle[ 5672] = 1'b1;  addr_rom[ 5672]='h0000072c;  wr_data_rom[ 5672]='h0000146e;
    rd_cycle[ 5673] = 1'b0;  wr_cycle[ 5673] = 1'b1;  addr_rom[ 5673]='h00000f18;  wr_data_rom[ 5673]='h00000c9c;
    rd_cycle[ 5674] = 1'b1;  wr_cycle[ 5674] = 1'b0;  addr_rom[ 5674]='h00000808;  wr_data_rom[ 5674]='h00000000;
    rd_cycle[ 5675] = 1'b1;  wr_cycle[ 5675] = 1'b0;  addr_rom[ 5675]='h00000dec;  wr_data_rom[ 5675]='h00000000;
    rd_cycle[ 5676] = 1'b1;  wr_cycle[ 5676] = 1'b0;  addr_rom[ 5676]='h00000048;  wr_data_rom[ 5676]='h00000000;
    rd_cycle[ 5677] = 1'b0;  wr_cycle[ 5677] = 1'b1;  addr_rom[ 5677]='h0000037c;  wr_data_rom[ 5677]='h00000f7b;
    rd_cycle[ 5678] = 1'b1;  wr_cycle[ 5678] = 1'b0;  addr_rom[ 5678]='h00000704;  wr_data_rom[ 5678]='h00000000;
    rd_cycle[ 5679] = 1'b1;  wr_cycle[ 5679] = 1'b0;  addr_rom[ 5679]='h00001dc0;  wr_data_rom[ 5679]='h00000000;
    rd_cycle[ 5680] = 1'b0;  wr_cycle[ 5680] = 1'b1;  addr_rom[ 5680]='h000019f4;  wr_data_rom[ 5680]='h00000e6b;
    rd_cycle[ 5681] = 1'b1;  wr_cycle[ 5681] = 1'b0;  addr_rom[ 5681]='h00000724;  wr_data_rom[ 5681]='h00000000;
    rd_cycle[ 5682] = 1'b0;  wr_cycle[ 5682] = 1'b1;  addr_rom[ 5682]='h00000ef0;  wr_data_rom[ 5682]='h000011b9;
    rd_cycle[ 5683] = 1'b1;  wr_cycle[ 5683] = 1'b0;  addr_rom[ 5683]='h00000250;  wr_data_rom[ 5683]='h00000000;
    rd_cycle[ 5684] = 1'b1;  wr_cycle[ 5684] = 1'b0;  addr_rom[ 5684]='h00000448;  wr_data_rom[ 5684]='h00000000;
    rd_cycle[ 5685] = 1'b1;  wr_cycle[ 5685] = 1'b0;  addr_rom[ 5685]='h000005a4;  wr_data_rom[ 5685]='h00000000;
    rd_cycle[ 5686] = 1'b1;  wr_cycle[ 5686] = 1'b0;  addr_rom[ 5686]='h00001444;  wr_data_rom[ 5686]='h00000000;
    rd_cycle[ 5687] = 1'b0;  wr_cycle[ 5687] = 1'b1;  addr_rom[ 5687]='h00001ee4;  wr_data_rom[ 5687]='h00001c91;
    rd_cycle[ 5688] = 1'b1;  wr_cycle[ 5688] = 1'b0;  addr_rom[ 5688]='h00001d5c;  wr_data_rom[ 5688]='h00000000;
    rd_cycle[ 5689] = 1'b1;  wr_cycle[ 5689] = 1'b0;  addr_rom[ 5689]='h00000f04;  wr_data_rom[ 5689]='h00000000;
    rd_cycle[ 5690] = 1'b0;  wr_cycle[ 5690] = 1'b1;  addr_rom[ 5690]='h00000a1c;  wr_data_rom[ 5690]='h0000125d;
    rd_cycle[ 5691] = 1'b1;  wr_cycle[ 5691] = 1'b0;  addr_rom[ 5691]='h000000f0;  wr_data_rom[ 5691]='h00000000;
    rd_cycle[ 5692] = 1'b1;  wr_cycle[ 5692] = 1'b0;  addr_rom[ 5692]='h0000147c;  wr_data_rom[ 5692]='h00000000;
    rd_cycle[ 5693] = 1'b1;  wr_cycle[ 5693] = 1'b0;  addr_rom[ 5693]='h00001164;  wr_data_rom[ 5693]='h00000000;
    rd_cycle[ 5694] = 1'b0;  wr_cycle[ 5694] = 1'b1;  addr_rom[ 5694]='h00001af0;  wr_data_rom[ 5694]='h000013d9;
    rd_cycle[ 5695] = 1'b0;  wr_cycle[ 5695] = 1'b1;  addr_rom[ 5695]='h00000624;  wr_data_rom[ 5695]='h000002cf;
    rd_cycle[ 5696] = 1'b1;  wr_cycle[ 5696] = 1'b0;  addr_rom[ 5696]='h00000380;  wr_data_rom[ 5696]='h00000000;
    rd_cycle[ 5697] = 1'b0;  wr_cycle[ 5697] = 1'b1;  addr_rom[ 5697]='h00001944;  wr_data_rom[ 5697]='h00000878;
    rd_cycle[ 5698] = 1'b0;  wr_cycle[ 5698] = 1'b1;  addr_rom[ 5698]='h000004b4;  wr_data_rom[ 5698]='h00000cff;
    rd_cycle[ 5699] = 1'b1;  wr_cycle[ 5699] = 1'b0;  addr_rom[ 5699]='h00000834;  wr_data_rom[ 5699]='h00000000;
    rd_cycle[ 5700] = 1'b1;  wr_cycle[ 5700] = 1'b0;  addr_rom[ 5700]='h00001870;  wr_data_rom[ 5700]='h00000000;
    rd_cycle[ 5701] = 1'b1;  wr_cycle[ 5701] = 1'b0;  addr_rom[ 5701]='h00000b8c;  wr_data_rom[ 5701]='h00000000;
    rd_cycle[ 5702] = 1'b1;  wr_cycle[ 5702] = 1'b0;  addr_rom[ 5702]='h00000c88;  wr_data_rom[ 5702]='h00000000;
    rd_cycle[ 5703] = 1'b0;  wr_cycle[ 5703] = 1'b1;  addr_rom[ 5703]='h00001eb0;  wr_data_rom[ 5703]='h00000e3a;
    rd_cycle[ 5704] = 1'b1;  wr_cycle[ 5704] = 1'b0;  addr_rom[ 5704]='h000002b0;  wr_data_rom[ 5704]='h00000000;
    rd_cycle[ 5705] = 1'b1;  wr_cycle[ 5705] = 1'b0;  addr_rom[ 5705]='h00001454;  wr_data_rom[ 5705]='h00000000;
    rd_cycle[ 5706] = 1'b1;  wr_cycle[ 5706] = 1'b0;  addr_rom[ 5706]='h0000053c;  wr_data_rom[ 5706]='h00000000;
    rd_cycle[ 5707] = 1'b0;  wr_cycle[ 5707] = 1'b1;  addr_rom[ 5707]='h00000c28;  wr_data_rom[ 5707]='h00000af9;
    rd_cycle[ 5708] = 1'b0;  wr_cycle[ 5708] = 1'b1;  addr_rom[ 5708]='h0000116c;  wr_data_rom[ 5708]='h00000b49;
    rd_cycle[ 5709] = 1'b1;  wr_cycle[ 5709] = 1'b0;  addr_rom[ 5709]='h00001640;  wr_data_rom[ 5709]='h00000000;
    rd_cycle[ 5710] = 1'b0;  wr_cycle[ 5710] = 1'b1;  addr_rom[ 5710]='h00001820;  wr_data_rom[ 5710]='h00000557;
    rd_cycle[ 5711] = 1'b1;  wr_cycle[ 5711] = 1'b0;  addr_rom[ 5711]='h000005c4;  wr_data_rom[ 5711]='h00000000;
    rd_cycle[ 5712] = 1'b1;  wr_cycle[ 5712] = 1'b0;  addr_rom[ 5712]='h00000fd0;  wr_data_rom[ 5712]='h00000000;
    rd_cycle[ 5713] = 1'b1;  wr_cycle[ 5713] = 1'b0;  addr_rom[ 5713]='h00000bc8;  wr_data_rom[ 5713]='h00000000;
    rd_cycle[ 5714] = 1'b1;  wr_cycle[ 5714] = 1'b0;  addr_rom[ 5714]='h00000508;  wr_data_rom[ 5714]='h00000000;
    rd_cycle[ 5715] = 1'b1;  wr_cycle[ 5715] = 1'b0;  addr_rom[ 5715]='h000011c8;  wr_data_rom[ 5715]='h00000000;
    rd_cycle[ 5716] = 1'b1;  wr_cycle[ 5716] = 1'b0;  addr_rom[ 5716]='h00000378;  wr_data_rom[ 5716]='h00000000;
    rd_cycle[ 5717] = 1'b0;  wr_cycle[ 5717] = 1'b1;  addr_rom[ 5717]='h0000128c;  wr_data_rom[ 5717]='h00001718;
    rd_cycle[ 5718] = 1'b0;  wr_cycle[ 5718] = 1'b1;  addr_rom[ 5718]='h00000540;  wr_data_rom[ 5718]='h00001092;
    rd_cycle[ 5719] = 1'b0;  wr_cycle[ 5719] = 1'b1;  addr_rom[ 5719]='h000003a4;  wr_data_rom[ 5719]='h00000fb5;
    rd_cycle[ 5720] = 1'b1;  wr_cycle[ 5720] = 1'b0;  addr_rom[ 5720]='h00001ac0;  wr_data_rom[ 5720]='h00000000;
    rd_cycle[ 5721] = 1'b0;  wr_cycle[ 5721] = 1'b1;  addr_rom[ 5721]='h000005d8;  wr_data_rom[ 5721]='h00001df7;
    rd_cycle[ 5722] = 1'b1;  wr_cycle[ 5722] = 1'b0;  addr_rom[ 5722]='h00000060;  wr_data_rom[ 5722]='h00000000;
    rd_cycle[ 5723] = 1'b0;  wr_cycle[ 5723] = 1'b1;  addr_rom[ 5723]='h000016a4;  wr_data_rom[ 5723]='h00000bf2;
    rd_cycle[ 5724] = 1'b1;  wr_cycle[ 5724] = 1'b0;  addr_rom[ 5724]='h000012ac;  wr_data_rom[ 5724]='h00000000;
    rd_cycle[ 5725] = 1'b1;  wr_cycle[ 5725] = 1'b0;  addr_rom[ 5725]='h00001e50;  wr_data_rom[ 5725]='h00000000;
    rd_cycle[ 5726] = 1'b1;  wr_cycle[ 5726] = 1'b0;  addr_rom[ 5726]='h0000059c;  wr_data_rom[ 5726]='h00000000;
    rd_cycle[ 5727] = 1'b1;  wr_cycle[ 5727] = 1'b0;  addr_rom[ 5727]='h0000025c;  wr_data_rom[ 5727]='h00000000;
    rd_cycle[ 5728] = 1'b1;  wr_cycle[ 5728] = 1'b0;  addr_rom[ 5728]='h00000540;  wr_data_rom[ 5728]='h00000000;
    rd_cycle[ 5729] = 1'b1;  wr_cycle[ 5729] = 1'b0;  addr_rom[ 5729]='h00001b2c;  wr_data_rom[ 5729]='h00000000;
    rd_cycle[ 5730] = 1'b0;  wr_cycle[ 5730] = 1'b1;  addr_rom[ 5730]='h000014f8;  wr_data_rom[ 5730]='h000009fa;
    rd_cycle[ 5731] = 1'b0;  wr_cycle[ 5731] = 1'b1;  addr_rom[ 5731]='h00001d30;  wr_data_rom[ 5731]='h000019af;
    rd_cycle[ 5732] = 1'b1;  wr_cycle[ 5732] = 1'b0;  addr_rom[ 5732]='h00001518;  wr_data_rom[ 5732]='h00000000;
    rd_cycle[ 5733] = 1'b0;  wr_cycle[ 5733] = 1'b1;  addr_rom[ 5733]='h000007d8;  wr_data_rom[ 5733]='h000009e5;
    rd_cycle[ 5734] = 1'b1;  wr_cycle[ 5734] = 1'b0;  addr_rom[ 5734]='h000009e0;  wr_data_rom[ 5734]='h00000000;
    rd_cycle[ 5735] = 1'b1;  wr_cycle[ 5735] = 1'b0;  addr_rom[ 5735]='h00001070;  wr_data_rom[ 5735]='h00000000;
    rd_cycle[ 5736] = 1'b0;  wr_cycle[ 5736] = 1'b1;  addr_rom[ 5736]='h00001018;  wr_data_rom[ 5736]='h000013e2;
    rd_cycle[ 5737] = 1'b1;  wr_cycle[ 5737] = 1'b0;  addr_rom[ 5737]='h00000c78;  wr_data_rom[ 5737]='h00000000;
    rd_cycle[ 5738] = 1'b0;  wr_cycle[ 5738] = 1'b1;  addr_rom[ 5738]='h00000d64;  wr_data_rom[ 5738]='h00001d32;
    rd_cycle[ 5739] = 1'b1;  wr_cycle[ 5739] = 1'b0;  addr_rom[ 5739]='h000002ac;  wr_data_rom[ 5739]='h00000000;
    rd_cycle[ 5740] = 1'b0;  wr_cycle[ 5740] = 1'b1;  addr_rom[ 5740]='h00001ce4;  wr_data_rom[ 5740]='h00001040;
    rd_cycle[ 5741] = 1'b1;  wr_cycle[ 5741] = 1'b0;  addr_rom[ 5741]='h00001e90;  wr_data_rom[ 5741]='h00000000;
    rd_cycle[ 5742] = 1'b1;  wr_cycle[ 5742] = 1'b0;  addr_rom[ 5742]='h0000111c;  wr_data_rom[ 5742]='h00000000;
    rd_cycle[ 5743] = 1'b0;  wr_cycle[ 5743] = 1'b1;  addr_rom[ 5743]='h00001440;  wr_data_rom[ 5743]='h00001252;
    rd_cycle[ 5744] = 1'b0;  wr_cycle[ 5744] = 1'b1;  addr_rom[ 5744]='h000011f0;  wr_data_rom[ 5744]='h000013a8;
    rd_cycle[ 5745] = 1'b0;  wr_cycle[ 5745] = 1'b1;  addr_rom[ 5745]='h00001b18;  wr_data_rom[ 5745]='h0000116c;
    rd_cycle[ 5746] = 1'b0;  wr_cycle[ 5746] = 1'b1;  addr_rom[ 5746]='h00000c70;  wr_data_rom[ 5746]='h000005ce;
    rd_cycle[ 5747] = 1'b0;  wr_cycle[ 5747] = 1'b1;  addr_rom[ 5747]='h00001da4;  wr_data_rom[ 5747]='h00000625;
    rd_cycle[ 5748] = 1'b0;  wr_cycle[ 5748] = 1'b1;  addr_rom[ 5748]='h00000fa0;  wr_data_rom[ 5748]='h0000196a;
    rd_cycle[ 5749] = 1'b1;  wr_cycle[ 5749] = 1'b0;  addr_rom[ 5749]='h00001400;  wr_data_rom[ 5749]='h00000000;
    rd_cycle[ 5750] = 1'b1;  wr_cycle[ 5750] = 1'b0;  addr_rom[ 5750]='h00000424;  wr_data_rom[ 5750]='h00000000;
    rd_cycle[ 5751] = 1'b0;  wr_cycle[ 5751] = 1'b1;  addr_rom[ 5751]='h0000133c;  wr_data_rom[ 5751]='h00000a09;
    rd_cycle[ 5752] = 1'b0;  wr_cycle[ 5752] = 1'b1;  addr_rom[ 5752]='h0000174c;  wr_data_rom[ 5752]='h0000052f;
    rd_cycle[ 5753] = 1'b1;  wr_cycle[ 5753] = 1'b0;  addr_rom[ 5753]='h000014f4;  wr_data_rom[ 5753]='h00000000;
    rd_cycle[ 5754] = 1'b0;  wr_cycle[ 5754] = 1'b1;  addr_rom[ 5754]='h00001764;  wr_data_rom[ 5754]='h0000172d;
    rd_cycle[ 5755] = 1'b0;  wr_cycle[ 5755] = 1'b1;  addr_rom[ 5755]='h00000d74;  wr_data_rom[ 5755]='h000011d5;
    rd_cycle[ 5756] = 1'b1;  wr_cycle[ 5756] = 1'b0;  addr_rom[ 5756]='h0000139c;  wr_data_rom[ 5756]='h00000000;
    rd_cycle[ 5757] = 1'b0;  wr_cycle[ 5757] = 1'b1;  addr_rom[ 5757]='h000010ac;  wr_data_rom[ 5757]='h00000252;
    rd_cycle[ 5758] = 1'b0;  wr_cycle[ 5758] = 1'b1;  addr_rom[ 5758]='h00001a48;  wr_data_rom[ 5758]='h000013cd;
    rd_cycle[ 5759] = 1'b1;  wr_cycle[ 5759] = 1'b0;  addr_rom[ 5759]='h00000070;  wr_data_rom[ 5759]='h00000000;
    rd_cycle[ 5760] = 1'b0;  wr_cycle[ 5760] = 1'b1;  addr_rom[ 5760]='h00000130;  wr_data_rom[ 5760]='h00000ad2;
    rd_cycle[ 5761] = 1'b0;  wr_cycle[ 5761] = 1'b1;  addr_rom[ 5761]='h00000890;  wr_data_rom[ 5761]='h00000661;
    rd_cycle[ 5762] = 1'b0;  wr_cycle[ 5762] = 1'b1;  addr_rom[ 5762]='h0000181c;  wr_data_rom[ 5762]='h00001b94;
    rd_cycle[ 5763] = 1'b1;  wr_cycle[ 5763] = 1'b0;  addr_rom[ 5763]='h00001794;  wr_data_rom[ 5763]='h00000000;
    rd_cycle[ 5764] = 1'b0;  wr_cycle[ 5764] = 1'b1;  addr_rom[ 5764]='h00000a40;  wr_data_rom[ 5764]='h0000083e;
    rd_cycle[ 5765] = 1'b0;  wr_cycle[ 5765] = 1'b1;  addr_rom[ 5765]='h00001154;  wr_data_rom[ 5765]='h00000902;
    rd_cycle[ 5766] = 1'b1;  wr_cycle[ 5766] = 1'b0;  addr_rom[ 5766]='h000017b0;  wr_data_rom[ 5766]='h00000000;
    rd_cycle[ 5767] = 1'b0;  wr_cycle[ 5767] = 1'b1;  addr_rom[ 5767]='h00001b64;  wr_data_rom[ 5767]='h00001253;
    rd_cycle[ 5768] = 1'b0;  wr_cycle[ 5768] = 1'b1;  addr_rom[ 5768]='h000004f0;  wr_data_rom[ 5768]='h00001c35;
    rd_cycle[ 5769] = 1'b1;  wr_cycle[ 5769] = 1'b0;  addr_rom[ 5769]='h000003fc;  wr_data_rom[ 5769]='h00000000;
    rd_cycle[ 5770] = 1'b1;  wr_cycle[ 5770] = 1'b0;  addr_rom[ 5770]='h000001b0;  wr_data_rom[ 5770]='h00000000;
    rd_cycle[ 5771] = 1'b0;  wr_cycle[ 5771] = 1'b1;  addr_rom[ 5771]='h00001dcc;  wr_data_rom[ 5771]='h00000a72;
    rd_cycle[ 5772] = 1'b1;  wr_cycle[ 5772] = 1'b0;  addr_rom[ 5772]='h000003b4;  wr_data_rom[ 5772]='h00000000;
    rd_cycle[ 5773] = 1'b0;  wr_cycle[ 5773] = 1'b1;  addr_rom[ 5773]='h0000128c;  wr_data_rom[ 5773]='h00001345;
    rd_cycle[ 5774] = 1'b1;  wr_cycle[ 5774] = 1'b0;  addr_rom[ 5774]='h00001214;  wr_data_rom[ 5774]='h00000000;
    rd_cycle[ 5775] = 1'b1;  wr_cycle[ 5775] = 1'b0;  addr_rom[ 5775]='h00001b40;  wr_data_rom[ 5775]='h00000000;
    rd_cycle[ 5776] = 1'b1;  wr_cycle[ 5776] = 1'b0;  addr_rom[ 5776]='h00001b14;  wr_data_rom[ 5776]='h00000000;
    rd_cycle[ 5777] = 1'b0;  wr_cycle[ 5777] = 1'b1;  addr_rom[ 5777]='h00000c24;  wr_data_rom[ 5777]='h000015b1;
    rd_cycle[ 5778] = 1'b0;  wr_cycle[ 5778] = 1'b1;  addr_rom[ 5778]='h00001794;  wr_data_rom[ 5778]='h00000c64;
    rd_cycle[ 5779] = 1'b0;  wr_cycle[ 5779] = 1'b1;  addr_rom[ 5779]='h000014ac;  wr_data_rom[ 5779]='h00000954;
    rd_cycle[ 5780] = 1'b1;  wr_cycle[ 5780] = 1'b0;  addr_rom[ 5780]='h0000156c;  wr_data_rom[ 5780]='h00000000;
    rd_cycle[ 5781] = 1'b1;  wr_cycle[ 5781] = 1'b0;  addr_rom[ 5781]='h00000f20;  wr_data_rom[ 5781]='h00000000;
    rd_cycle[ 5782] = 1'b0;  wr_cycle[ 5782] = 1'b1;  addr_rom[ 5782]='h000009f0;  wr_data_rom[ 5782]='h00000e4f;
    rd_cycle[ 5783] = 1'b0;  wr_cycle[ 5783] = 1'b1;  addr_rom[ 5783]='h00001b58;  wr_data_rom[ 5783]='h0000015e;
    rd_cycle[ 5784] = 1'b0;  wr_cycle[ 5784] = 1'b1;  addr_rom[ 5784]='h00000d74;  wr_data_rom[ 5784]='h00000186;
    rd_cycle[ 5785] = 1'b0;  wr_cycle[ 5785] = 1'b1;  addr_rom[ 5785]='h00001f18;  wr_data_rom[ 5785]='h000006ba;
    rd_cycle[ 5786] = 1'b0;  wr_cycle[ 5786] = 1'b1;  addr_rom[ 5786]='h00001a34;  wr_data_rom[ 5786]='h00001f2a;
    rd_cycle[ 5787] = 1'b0;  wr_cycle[ 5787] = 1'b1;  addr_rom[ 5787]='h00000084;  wr_data_rom[ 5787]='h00001a32;
    rd_cycle[ 5788] = 1'b0;  wr_cycle[ 5788] = 1'b1;  addr_rom[ 5788]='h00001e5c;  wr_data_rom[ 5788]='h00001bd6;
    rd_cycle[ 5789] = 1'b1;  wr_cycle[ 5789] = 1'b0;  addr_rom[ 5789]='h00000520;  wr_data_rom[ 5789]='h00000000;
    rd_cycle[ 5790] = 1'b0;  wr_cycle[ 5790] = 1'b1;  addr_rom[ 5790]='h00000e3c;  wr_data_rom[ 5790]='h0000004f;
    rd_cycle[ 5791] = 1'b0;  wr_cycle[ 5791] = 1'b1;  addr_rom[ 5791]='h00000b48;  wr_data_rom[ 5791]='h00001047;
    rd_cycle[ 5792] = 1'b0;  wr_cycle[ 5792] = 1'b1;  addr_rom[ 5792]='h00000554;  wr_data_rom[ 5792]='h00001bd2;
    rd_cycle[ 5793] = 1'b1;  wr_cycle[ 5793] = 1'b0;  addr_rom[ 5793]='h00000340;  wr_data_rom[ 5793]='h00000000;
    rd_cycle[ 5794] = 1'b0;  wr_cycle[ 5794] = 1'b1;  addr_rom[ 5794]='h00000910;  wr_data_rom[ 5794]='h000016ac;
    rd_cycle[ 5795] = 1'b1;  wr_cycle[ 5795] = 1'b0;  addr_rom[ 5795]='h00001820;  wr_data_rom[ 5795]='h00000000;
    rd_cycle[ 5796] = 1'b1;  wr_cycle[ 5796] = 1'b0;  addr_rom[ 5796]='h000009f8;  wr_data_rom[ 5796]='h00000000;
    rd_cycle[ 5797] = 1'b0;  wr_cycle[ 5797] = 1'b1;  addr_rom[ 5797]='h00000438;  wr_data_rom[ 5797]='h00001abd;
    rd_cycle[ 5798] = 1'b0;  wr_cycle[ 5798] = 1'b1;  addr_rom[ 5798]='h000003f8;  wr_data_rom[ 5798]='h00001cc6;
    rd_cycle[ 5799] = 1'b0;  wr_cycle[ 5799] = 1'b1;  addr_rom[ 5799]='h000001b4;  wr_data_rom[ 5799]='h00000743;
    rd_cycle[ 5800] = 1'b1;  wr_cycle[ 5800] = 1'b0;  addr_rom[ 5800]='h000006b4;  wr_data_rom[ 5800]='h00000000;
    rd_cycle[ 5801] = 1'b0;  wr_cycle[ 5801] = 1'b1;  addr_rom[ 5801]='h00000fb8;  wr_data_rom[ 5801]='h00001cbf;
    rd_cycle[ 5802] = 1'b0;  wr_cycle[ 5802] = 1'b1;  addr_rom[ 5802]='h000013d4;  wr_data_rom[ 5802]='h00001b24;
    rd_cycle[ 5803] = 1'b0;  wr_cycle[ 5803] = 1'b1;  addr_rom[ 5803]='h00000320;  wr_data_rom[ 5803]='h00001a9f;
    rd_cycle[ 5804] = 1'b0;  wr_cycle[ 5804] = 1'b1;  addr_rom[ 5804]='h000007d8;  wr_data_rom[ 5804]='h0000062c;
    rd_cycle[ 5805] = 1'b1;  wr_cycle[ 5805] = 1'b0;  addr_rom[ 5805]='h00001b7c;  wr_data_rom[ 5805]='h00000000;
    rd_cycle[ 5806] = 1'b1;  wr_cycle[ 5806] = 1'b0;  addr_rom[ 5806]='h00000680;  wr_data_rom[ 5806]='h00000000;
    rd_cycle[ 5807] = 1'b0;  wr_cycle[ 5807] = 1'b1;  addr_rom[ 5807]='h00001950;  wr_data_rom[ 5807]='h00000254;
    rd_cycle[ 5808] = 1'b1;  wr_cycle[ 5808] = 1'b0;  addr_rom[ 5808]='h0000031c;  wr_data_rom[ 5808]='h00000000;
    rd_cycle[ 5809] = 1'b1;  wr_cycle[ 5809] = 1'b0;  addr_rom[ 5809]='h00000694;  wr_data_rom[ 5809]='h00000000;
    rd_cycle[ 5810] = 1'b0;  wr_cycle[ 5810] = 1'b1;  addr_rom[ 5810]='h00000980;  wr_data_rom[ 5810]='h00001c2b;
    rd_cycle[ 5811] = 1'b0;  wr_cycle[ 5811] = 1'b1;  addr_rom[ 5811]='h00001940;  wr_data_rom[ 5811]='h00001801;
    rd_cycle[ 5812] = 1'b1;  wr_cycle[ 5812] = 1'b0;  addr_rom[ 5812]='h00000100;  wr_data_rom[ 5812]='h00000000;
    rd_cycle[ 5813] = 1'b0;  wr_cycle[ 5813] = 1'b1;  addr_rom[ 5813]='h00000a14;  wr_data_rom[ 5813]='h000003e9;
    rd_cycle[ 5814] = 1'b1;  wr_cycle[ 5814] = 1'b0;  addr_rom[ 5814]='h000012e0;  wr_data_rom[ 5814]='h00000000;
    rd_cycle[ 5815] = 1'b0;  wr_cycle[ 5815] = 1'b1;  addr_rom[ 5815]='h00000840;  wr_data_rom[ 5815]='h00001d0d;
    rd_cycle[ 5816] = 1'b0;  wr_cycle[ 5816] = 1'b1;  addr_rom[ 5816]='h0000075c;  wr_data_rom[ 5816]='h0000101a;
    rd_cycle[ 5817] = 1'b1;  wr_cycle[ 5817] = 1'b0;  addr_rom[ 5817]='h00000368;  wr_data_rom[ 5817]='h00000000;
    rd_cycle[ 5818] = 1'b0;  wr_cycle[ 5818] = 1'b1;  addr_rom[ 5818]='h00001958;  wr_data_rom[ 5818]='h00000452;
    rd_cycle[ 5819] = 1'b0;  wr_cycle[ 5819] = 1'b1;  addr_rom[ 5819]='h00000f10;  wr_data_rom[ 5819]='h00001045;
    rd_cycle[ 5820] = 1'b1;  wr_cycle[ 5820] = 1'b0;  addr_rom[ 5820]='h00000634;  wr_data_rom[ 5820]='h00000000;
    rd_cycle[ 5821] = 1'b1;  wr_cycle[ 5821] = 1'b0;  addr_rom[ 5821]='h00001948;  wr_data_rom[ 5821]='h00000000;
    rd_cycle[ 5822] = 1'b1;  wr_cycle[ 5822] = 1'b0;  addr_rom[ 5822]='h00000c94;  wr_data_rom[ 5822]='h00000000;
    rd_cycle[ 5823] = 1'b1;  wr_cycle[ 5823] = 1'b0;  addr_rom[ 5823]='h00000d48;  wr_data_rom[ 5823]='h00000000;
    rd_cycle[ 5824] = 1'b0;  wr_cycle[ 5824] = 1'b1;  addr_rom[ 5824]='h000012f8;  wr_data_rom[ 5824]='h00000b58;
    rd_cycle[ 5825] = 1'b1;  wr_cycle[ 5825] = 1'b0;  addr_rom[ 5825]='h00000c8c;  wr_data_rom[ 5825]='h00000000;
    rd_cycle[ 5826] = 1'b1;  wr_cycle[ 5826] = 1'b0;  addr_rom[ 5826]='h00000528;  wr_data_rom[ 5826]='h00000000;
    rd_cycle[ 5827] = 1'b0;  wr_cycle[ 5827] = 1'b1;  addr_rom[ 5827]='h00000404;  wr_data_rom[ 5827]='h00000dd6;
    rd_cycle[ 5828] = 1'b0;  wr_cycle[ 5828] = 1'b1;  addr_rom[ 5828]='h000008b8;  wr_data_rom[ 5828]='h00000013;
    rd_cycle[ 5829] = 1'b0;  wr_cycle[ 5829] = 1'b1;  addr_rom[ 5829]='h00001a80;  wr_data_rom[ 5829]='h0000047b;
    rd_cycle[ 5830] = 1'b1;  wr_cycle[ 5830] = 1'b0;  addr_rom[ 5830]='h0000012c;  wr_data_rom[ 5830]='h00000000;
    rd_cycle[ 5831] = 1'b0;  wr_cycle[ 5831] = 1'b1;  addr_rom[ 5831]='h00001bc8;  wr_data_rom[ 5831]='h000009fb;
    rd_cycle[ 5832] = 1'b1;  wr_cycle[ 5832] = 1'b0;  addr_rom[ 5832]='h00000ce4;  wr_data_rom[ 5832]='h00000000;
    rd_cycle[ 5833] = 1'b1;  wr_cycle[ 5833] = 1'b0;  addr_rom[ 5833]='h000012d8;  wr_data_rom[ 5833]='h00000000;
    rd_cycle[ 5834] = 1'b0;  wr_cycle[ 5834] = 1'b1;  addr_rom[ 5834]='h00001164;  wr_data_rom[ 5834]='h000013a8;
    rd_cycle[ 5835] = 1'b1;  wr_cycle[ 5835] = 1'b0;  addr_rom[ 5835]='h00001748;  wr_data_rom[ 5835]='h00000000;
    rd_cycle[ 5836] = 1'b0;  wr_cycle[ 5836] = 1'b1;  addr_rom[ 5836]='h00001e18;  wr_data_rom[ 5836]='h00000f22;
    rd_cycle[ 5837] = 1'b1;  wr_cycle[ 5837] = 1'b0;  addr_rom[ 5837]='h00001c2c;  wr_data_rom[ 5837]='h00000000;
    rd_cycle[ 5838] = 1'b0;  wr_cycle[ 5838] = 1'b1;  addr_rom[ 5838]='h000000c0;  wr_data_rom[ 5838]='h00000deb;
    rd_cycle[ 5839] = 1'b1;  wr_cycle[ 5839] = 1'b0;  addr_rom[ 5839]='h00000f8c;  wr_data_rom[ 5839]='h00000000;
    rd_cycle[ 5840] = 1'b0;  wr_cycle[ 5840] = 1'b1;  addr_rom[ 5840]='h000010ec;  wr_data_rom[ 5840]='h00001b35;
    rd_cycle[ 5841] = 1'b1;  wr_cycle[ 5841] = 1'b0;  addr_rom[ 5841]='h000010d0;  wr_data_rom[ 5841]='h00000000;
    rd_cycle[ 5842] = 1'b1;  wr_cycle[ 5842] = 1'b0;  addr_rom[ 5842]='h00000ecc;  wr_data_rom[ 5842]='h00000000;
    rd_cycle[ 5843] = 1'b1;  wr_cycle[ 5843] = 1'b0;  addr_rom[ 5843]='h00001a8c;  wr_data_rom[ 5843]='h00000000;
    rd_cycle[ 5844] = 1'b0;  wr_cycle[ 5844] = 1'b1;  addr_rom[ 5844]='h000014f4;  wr_data_rom[ 5844]='h00001083;
    rd_cycle[ 5845] = 1'b0;  wr_cycle[ 5845] = 1'b1;  addr_rom[ 5845]='h00001d24;  wr_data_rom[ 5845]='h000011eb;
    rd_cycle[ 5846] = 1'b0;  wr_cycle[ 5846] = 1'b1;  addr_rom[ 5846]='h000014b4;  wr_data_rom[ 5846]='h00001b34;
    rd_cycle[ 5847] = 1'b0;  wr_cycle[ 5847] = 1'b1;  addr_rom[ 5847]='h00000fa8;  wr_data_rom[ 5847]='h000019ed;
    rd_cycle[ 5848] = 1'b1;  wr_cycle[ 5848] = 1'b0;  addr_rom[ 5848]='h000018b0;  wr_data_rom[ 5848]='h00000000;
    rd_cycle[ 5849] = 1'b1;  wr_cycle[ 5849] = 1'b0;  addr_rom[ 5849]='h0000088c;  wr_data_rom[ 5849]='h00000000;
    rd_cycle[ 5850] = 1'b1;  wr_cycle[ 5850] = 1'b0;  addr_rom[ 5850]='h00000034;  wr_data_rom[ 5850]='h00000000;
    rd_cycle[ 5851] = 1'b1;  wr_cycle[ 5851] = 1'b0;  addr_rom[ 5851]='h000000b0;  wr_data_rom[ 5851]='h00000000;
    rd_cycle[ 5852] = 1'b1;  wr_cycle[ 5852] = 1'b0;  addr_rom[ 5852]='h00001730;  wr_data_rom[ 5852]='h00000000;
    rd_cycle[ 5853] = 1'b1;  wr_cycle[ 5853] = 1'b0;  addr_rom[ 5853]='h00000e7c;  wr_data_rom[ 5853]='h00000000;
    rd_cycle[ 5854] = 1'b0;  wr_cycle[ 5854] = 1'b1;  addr_rom[ 5854]='h000013ac;  wr_data_rom[ 5854]='h00001bd1;
    rd_cycle[ 5855] = 1'b0;  wr_cycle[ 5855] = 1'b1;  addr_rom[ 5855]='h00001724;  wr_data_rom[ 5855]='h0000004f;
    rd_cycle[ 5856] = 1'b0;  wr_cycle[ 5856] = 1'b1;  addr_rom[ 5856]='h00000a88;  wr_data_rom[ 5856]='h00001c8a;
    rd_cycle[ 5857] = 1'b0;  wr_cycle[ 5857] = 1'b1;  addr_rom[ 5857]='h00000bc8;  wr_data_rom[ 5857]='h000019d7;
    rd_cycle[ 5858] = 1'b0;  wr_cycle[ 5858] = 1'b1;  addr_rom[ 5858]='h000014c8;  wr_data_rom[ 5858]='h0000047f;
    rd_cycle[ 5859] = 1'b0;  wr_cycle[ 5859] = 1'b1;  addr_rom[ 5859]='h00000284;  wr_data_rom[ 5859]='h00001a56;
    rd_cycle[ 5860] = 1'b1;  wr_cycle[ 5860] = 1'b0;  addr_rom[ 5860]='h00001648;  wr_data_rom[ 5860]='h00000000;
    rd_cycle[ 5861] = 1'b0;  wr_cycle[ 5861] = 1'b1;  addr_rom[ 5861]='h000014e4;  wr_data_rom[ 5861]='h00001015;
    rd_cycle[ 5862] = 1'b0;  wr_cycle[ 5862] = 1'b1;  addr_rom[ 5862]='h00000398;  wr_data_rom[ 5862]='h00000212;
    rd_cycle[ 5863] = 1'b1;  wr_cycle[ 5863] = 1'b0;  addr_rom[ 5863]='h00000128;  wr_data_rom[ 5863]='h00000000;
    rd_cycle[ 5864] = 1'b1;  wr_cycle[ 5864] = 1'b0;  addr_rom[ 5864]='h00000a04;  wr_data_rom[ 5864]='h00000000;
    rd_cycle[ 5865] = 1'b1;  wr_cycle[ 5865] = 1'b0;  addr_rom[ 5865]='h000007c0;  wr_data_rom[ 5865]='h00000000;
    rd_cycle[ 5866] = 1'b1;  wr_cycle[ 5866] = 1'b0;  addr_rom[ 5866]='h000000b8;  wr_data_rom[ 5866]='h00000000;
    rd_cycle[ 5867] = 1'b0;  wr_cycle[ 5867] = 1'b1;  addr_rom[ 5867]='h000016f8;  wr_data_rom[ 5867]='h000000a0;
    rd_cycle[ 5868] = 1'b0;  wr_cycle[ 5868] = 1'b1;  addr_rom[ 5868]='h00001394;  wr_data_rom[ 5868]='h000000eb;
    rd_cycle[ 5869] = 1'b0;  wr_cycle[ 5869] = 1'b1;  addr_rom[ 5869]='h00001d0c;  wr_data_rom[ 5869]='h000012a5;
    rd_cycle[ 5870] = 1'b1;  wr_cycle[ 5870] = 1'b0;  addr_rom[ 5870]='h0000144c;  wr_data_rom[ 5870]='h00000000;
    rd_cycle[ 5871] = 1'b0;  wr_cycle[ 5871] = 1'b1;  addr_rom[ 5871]='h00001d4c;  wr_data_rom[ 5871]='h000011a1;
    rd_cycle[ 5872] = 1'b1;  wr_cycle[ 5872] = 1'b0;  addr_rom[ 5872]='h00000428;  wr_data_rom[ 5872]='h00000000;
    rd_cycle[ 5873] = 1'b0;  wr_cycle[ 5873] = 1'b1;  addr_rom[ 5873]='h00001a24;  wr_data_rom[ 5873]='h000012c5;
    rd_cycle[ 5874] = 1'b1;  wr_cycle[ 5874] = 1'b0;  addr_rom[ 5874]='h0000100c;  wr_data_rom[ 5874]='h00000000;
    rd_cycle[ 5875] = 1'b0;  wr_cycle[ 5875] = 1'b1;  addr_rom[ 5875]='h00000124;  wr_data_rom[ 5875]='h000019bc;
    rd_cycle[ 5876] = 1'b1;  wr_cycle[ 5876] = 1'b0;  addr_rom[ 5876]='h0000115c;  wr_data_rom[ 5876]='h00000000;
    rd_cycle[ 5877] = 1'b0;  wr_cycle[ 5877] = 1'b1;  addr_rom[ 5877]='h0000104c;  wr_data_rom[ 5877]='h000014f1;
    rd_cycle[ 5878] = 1'b0;  wr_cycle[ 5878] = 1'b1;  addr_rom[ 5878]='h00000bac;  wr_data_rom[ 5878]='h0000131a;
    rd_cycle[ 5879] = 1'b1;  wr_cycle[ 5879] = 1'b0;  addr_rom[ 5879]='h00000b5c;  wr_data_rom[ 5879]='h00000000;
    rd_cycle[ 5880] = 1'b0;  wr_cycle[ 5880] = 1'b1;  addr_rom[ 5880]='h00001e48;  wr_data_rom[ 5880]='h0000177f;
    rd_cycle[ 5881] = 1'b0;  wr_cycle[ 5881] = 1'b1;  addr_rom[ 5881]='h00001508;  wr_data_rom[ 5881]='h00001355;
    rd_cycle[ 5882] = 1'b0;  wr_cycle[ 5882] = 1'b1;  addr_rom[ 5882]='h00000014;  wr_data_rom[ 5882]='h000004fb;
    rd_cycle[ 5883] = 1'b0;  wr_cycle[ 5883] = 1'b1;  addr_rom[ 5883]='h00001650;  wr_data_rom[ 5883]='h00001f3b;
    rd_cycle[ 5884] = 1'b1;  wr_cycle[ 5884] = 1'b0;  addr_rom[ 5884]='h00000418;  wr_data_rom[ 5884]='h00000000;
    rd_cycle[ 5885] = 1'b1;  wr_cycle[ 5885] = 1'b0;  addr_rom[ 5885]='h00000440;  wr_data_rom[ 5885]='h00000000;
    rd_cycle[ 5886] = 1'b1;  wr_cycle[ 5886] = 1'b0;  addr_rom[ 5886]='h00000fb8;  wr_data_rom[ 5886]='h00000000;
    rd_cycle[ 5887] = 1'b0;  wr_cycle[ 5887] = 1'b1;  addr_rom[ 5887]='h00000460;  wr_data_rom[ 5887]='h00001d5e;
    rd_cycle[ 5888] = 1'b0;  wr_cycle[ 5888] = 1'b1;  addr_rom[ 5888]='h00000f04;  wr_data_rom[ 5888]='h0000096c;
    rd_cycle[ 5889] = 1'b1;  wr_cycle[ 5889] = 1'b0;  addr_rom[ 5889]='h0000008c;  wr_data_rom[ 5889]='h00000000;
    rd_cycle[ 5890] = 1'b0;  wr_cycle[ 5890] = 1'b1;  addr_rom[ 5890]='h00001ee0;  wr_data_rom[ 5890]='h00000785;
    rd_cycle[ 5891] = 1'b1;  wr_cycle[ 5891] = 1'b0;  addr_rom[ 5891]='h00001198;  wr_data_rom[ 5891]='h00000000;
    rd_cycle[ 5892] = 1'b1;  wr_cycle[ 5892] = 1'b0;  addr_rom[ 5892]='h00001c14;  wr_data_rom[ 5892]='h00000000;
    rd_cycle[ 5893] = 1'b0;  wr_cycle[ 5893] = 1'b1;  addr_rom[ 5893]='h00001748;  wr_data_rom[ 5893]='h0000042c;
    rd_cycle[ 5894] = 1'b1;  wr_cycle[ 5894] = 1'b0;  addr_rom[ 5894]='h00000974;  wr_data_rom[ 5894]='h00000000;
    rd_cycle[ 5895] = 1'b1;  wr_cycle[ 5895] = 1'b0;  addr_rom[ 5895]='h000014cc;  wr_data_rom[ 5895]='h00000000;
    rd_cycle[ 5896] = 1'b1;  wr_cycle[ 5896] = 1'b0;  addr_rom[ 5896]='h00000d54;  wr_data_rom[ 5896]='h00000000;
    rd_cycle[ 5897] = 1'b1;  wr_cycle[ 5897] = 1'b0;  addr_rom[ 5897]='h00001d2c;  wr_data_rom[ 5897]='h00000000;
    rd_cycle[ 5898] = 1'b0;  wr_cycle[ 5898] = 1'b1;  addr_rom[ 5898]='h00001550;  wr_data_rom[ 5898]='h00000efa;
    rd_cycle[ 5899] = 1'b0;  wr_cycle[ 5899] = 1'b1;  addr_rom[ 5899]='h000014e8;  wr_data_rom[ 5899]='h00000eee;
    rd_cycle[ 5900] = 1'b0;  wr_cycle[ 5900] = 1'b1;  addr_rom[ 5900]='h0000109c;  wr_data_rom[ 5900]='h00001b0a;
    rd_cycle[ 5901] = 1'b1;  wr_cycle[ 5901] = 1'b0;  addr_rom[ 5901]='h00001858;  wr_data_rom[ 5901]='h00000000;
    rd_cycle[ 5902] = 1'b1;  wr_cycle[ 5902] = 1'b0;  addr_rom[ 5902]='h00000568;  wr_data_rom[ 5902]='h00000000;
    rd_cycle[ 5903] = 1'b1;  wr_cycle[ 5903] = 1'b0;  addr_rom[ 5903]='h000019c8;  wr_data_rom[ 5903]='h00000000;
    rd_cycle[ 5904] = 1'b1;  wr_cycle[ 5904] = 1'b0;  addr_rom[ 5904]='h000005bc;  wr_data_rom[ 5904]='h00000000;
    rd_cycle[ 5905] = 1'b1;  wr_cycle[ 5905] = 1'b0;  addr_rom[ 5905]='h00000108;  wr_data_rom[ 5905]='h00000000;
    rd_cycle[ 5906] = 1'b0;  wr_cycle[ 5906] = 1'b1;  addr_rom[ 5906]='h00000450;  wr_data_rom[ 5906]='h00001151;
    rd_cycle[ 5907] = 1'b1;  wr_cycle[ 5907] = 1'b0;  addr_rom[ 5907]='h00001b28;  wr_data_rom[ 5907]='h00000000;
    rd_cycle[ 5908] = 1'b0;  wr_cycle[ 5908] = 1'b1;  addr_rom[ 5908]='h000009e4;  wr_data_rom[ 5908]='h00001558;
    rd_cycle[ 5909] = 1'b1;  wr_cycle[ 5909] = 1'b0;  addr_rom[ 5909]='h00000854;  wr_data_rom[ 5909]='h00000000;
    rd_cycle[ 5910] = 1'b0;  wr_cycle[ 5910] = 1'b1;  addr_rom[ 5910]='h00000600;  wr_data_rom[ 5910]='h00001cba;
    rd_cycle[ 5911] = 1'b0;  wr_cycle[ 5911] = 1'b1;  addr_rom[ 5911]='h00000ff0;  wr_data_rom[ 5911]='h00001c9f;
    rd_cycle[ 5912] = 1'b0;  wr_cycle[ 5912] = 1'b1;  addr_rom[ 5912]='h00000f0c;  wr_data_rom[ 5912]='h000002e3;
    rd_cycle[ 5913] = 1'b1;  wr_cycle[ 5913] = 1'b0;  addr_rom[ 5913]='h00001b2c;  wr_data_rom[ 5913]='h00000000;
    rd_cycle[ 5914] = 1'b0;  wr_cycle[ 5914] = 1'b1;  addr_rom[ 5914]='h000012a0;  wr_data_rom[ 5914]='h00001143;
    rd_cycle[ 5915] = 1'b0;  wr_cycle[ 5915] = 1'b1;  addr_rom[ 5915]='h000013a8;  wr_data_rom[ 5915]='h00000139;
    rd_cycle[ 5916] = 1'b0;  wr_cycle[ 5916] = 1'b1;  addr_rom[ 5916]='h00001cf8;  wr_data_rom[ 5916]='h000016b8;
    rd_cycle[ 5917] = 1'b0;  wr_cycle[ 5917] = 1'b1;  addr_rom[ 5917]='h00001154;  wr_data_rom[ 5917]='h00000c96;
    rd_cycle[ 5918] = 1'b0;  wr_cycle[ 5918] = 1'b1;  addr_rom[ 5918]='h00001814;  wr_data_rom[ 5918]='h00001e61;
    rd_cycle[ 5919] = 1'b0;  wr_cycle[ 5919] = 1'b1;  addr_rom[ 5919]='h00001cec;  wr_data_rom[ 5919]='h00001489;
    rd_cycle[ 5920] = 1'b0;  wr_cycle[ 5920] = 1'b1;  addr_rom[ 5920]='h00001d88;  wr_data_rom[ 5920]='h00001afb;
    rd_cycle[ 5921] = 1'b0;  wr_cycle[ 5921] = 1'b1;  addr_rom[ 5921]='h00001ae0;  wr_data_rom[ 5921]='h00001bdc;
    rd_cycle[ 5922] = 1'b0;  wr_cycle[ 5922] = 1'b1;  addr_rom[ 5922]='h00001af0;  wr_data_rom[ 5922]='h00000e64;
    rd_cycle[ 5923] = 1'b1;  wr_cycle[ 5923] = 1'b0;  addr_rom[ 5923]='h0000062c;  wr_data_rom[ 5923]='h00000000;
    rd_cycle[ 5924] = 1'b0;  wr_cycle[ 5924] = 1'b1;  addr_rom[ 5924]='h00000628;  wr_data_rom[ 5924]='h00001227;
    rd_cycle[ 5925] = 1'b1;  wr_cycle[ 5925] = 1'b0;  addr_rom[ 5925]='h000016f8;  wr_data_rom[ 5925]='h00000000;
    rd_cycle[ 5926] = 1'b1;  wr_cycle[ 5926] = 1'b0;  addr_rom[ 5926]='h00000b58;  wr_data_rom[ 5926]='h00000000;
    rd_cycle[ 5927] = 1'b0;  wr_cycle[ 5927] = 1'b1;  addr_rom[ 5927]='h00000224;  wr_data_rom[ 5927]='h00000f51;
    rd_cycle[ 5928] = 1'b1;  wr_cycle[ 5928] = 1'b0;  addr_rom[ 5928]='h00001718;  wr_data_rom[ 5928]='h00000000;
    rd_cycle[ 5929] = 1'b0;  wr_cycle[ 5929] = 1'b1;  addr_rom[ 5929]='h0000102c;  wr_data_rom[ 5929]='h00000075;
    rd_cycle[ 5930] = 1'b0;  wr_cycle[ 5930] = 1'b1;  addr_rom[ 5930]='h00000e68;  wr_data_rom[ 5930]='h000017cb;
    rd_cycle[ 5931] = 1'b0;  wr_cycle[ 5931] = 1'b1;  addr_rom[ 5931]='h00001248;  wr_data_rom[ 5931]='h00001a04;
    rd_cycle[ 5932] = 1'b1;  wr_cycle[ 5932] = 1'b0;  addr_rom[ 5932]='h000004cc;  wr_data_rom[ 5932]='h00000000;
    rd_cycle[ 5933] = 1'b0;  wr_cycle[ 5933] = 1'b1;  addr_rom[ 5933]='h00000acc;  wr_data_rom[ 5933]='h00001ccd;
    rd_cycle[ 5934] = 1'b1;  wr_cycle[ 5934] = 1'b0;  addr_rom[ 5934]='h00001d4c;  wr_data_rom[ 5934]='h00000000;
    rd_cycle[ 5935] = 1'b0;  wr_cycle[ 5935] = 1'b1;  addr_rom[ 5935]='h00000758;  wr_data_rom[ 5935]='h00001820;
    rd_cycle[ 5936] = 1'b1;  wr_cycle[ 5936] = 1'b0;  addr_rom[ 5936]='h00000738;  wr_data_rom[ 5936]='h00000000;
    rd_cycle[ 5937] = 1'b1;  wr_cycle[ 5937] = 1'b0;  addr_rom[ 5937]='h00001d74;  wr_data_rom[ 5937]='h00000000;
    rd_cycle[ 5938] = 1'b1;  wr_cycle[ 5938] = 1'b0;  addr_rom[ 5938]='h000009e8;  wr_data_rom[ 5938]='h00000000;
    rd_cycle[ 5939] = 1'b0;  wr_cycle[ 5939] = 1'b1;  addr_rom[ 5939]='h00000bd0;  wr_data_rom[ 5939]='h00001b24;
    rd_cycle[ 5940] = 1'b0;  wr_cycle[ 5940] = 1'b1;  addr_rom[ 5940]='h00000ee8;  wr_data_rom[ 5940]='h00001f1c;
    rd_cycle[ 5941] = 1'b1;  wr_cycle[ 5941] = 1'b0;  addr_rom[ 5941]='h00001c4c;  wr_data_rom[ 5941]='h00000000;
    rd_cycle[ 5942] = 1'b0;  wr_cycle[ 5942] = 1'b1;  addr_rom[ 5942]='h00000f20;  wr_data_rom[ 5942]='h00000345;
    rd_cycle[ 5943] = 1'b0;  wr_cycle[ 5943] = 1'b1;  addr_rom[ 5943]='h00001b54;  wr_data_rom[ 5943]='h0000199f;
    rd_cycle[ 5944] = 1'b0;  wr_cycle[ 5944] = 1'b1;  addr_rom[ 5944]='h00000fb8;  wr_data_rom[ 5944]='h00000040;
    rd_cycle[ 5945] = 1'b0;  wr_cycle[ 5945] = 1'b1;  addr_rom[ 5945]='h000019b4;  wr_data_rom[ 5945]='h00001188;
    rd_cycle[ 5946] = 1'b0;  wr_cycle[ 5946] = 1'b1;  addr_rom[ 5946]='h00000ae4;  wr_data_rom[ 5946]='h000018f8;
    rd_cycle[ 5947] = 1'b0;  wr_cycle[ 5947] = 1'b1;  addr_rom[ 5947]='h0000136c;  wr_data_rom[ 5947]='h00000613;
    rd_cycle[ 5948] = 1'b0;  wr_cycle[ 5948] = 1'b1;  addr_rom[ 5948]='h00000750;  wr_data_rom[ 5948]='h00000ea4;
    rd_cycle[ 5949] = 1'b1;  wr_cycle[ 5949] = 1'b0;  addr_rom[ 5949]='h00000af4;  wr_data_rom[ 5949]='h00000000;
    rd_cycle[ 5950] = 1'b0;  wr_cycle[ 5950] = 1'b1;  addr_rom[ 5950]='h00000c08;  wr_data_rom[ 5950]='h000014fa;
    rd_cycle[ 5951] = 1'b1;  wr_cycle[ 5951] = 1'b0;  addr_rom[ 5951]='h000014d8;  wr_data_rom[ 5951]='h00000000;
    rd_cycle[ 5952] = 1'b1;  wr_cycle[ 5952] = 1'b0;  addr_rom[ 5952]='h000007f8;  wr_data_rom[ 5952]='h00000000;
    rd_cycle[ 5953] = 1'b1;  wr_cycle[ 5953] = 1'b0;  addr_rom[ 5953]='h00000300;  wr_data_rom[ 5953]='h00000000;
    rd_cycle[ 5954] = 1'b0;  wr_cycle[ 5954] = 1'b1;  addr_rom[ 5954]='h000000c0;  wr_data_rom[ 5954]='h0000107a;
    rd_cycle[ 5955] = 1'b0;  wr_cycle[ 5955] = 1'b1;  addr_rom[ 5955]='h00000674;  wr_data_rom[ 5955]='h00000eba;
    rd_cycle[ 5956] = 1'b1;  wr_cycle[ 5956] = 1'b0;  addr_rom[ 5956]='h00000b80;  wr_data_rom[ 5956]='h00000000;
    rd_cycle[ 5957] = 1'b0;  wr_cycle[ 5957] = 1'b1;  addr_rom[ 5957]='h000003e8;  wr_data_rom[ 5957]='h00000488;
    rd_cycle[ 5958] = 1'b0;  wr_cycle[ 5958] = 1'b1;  addr_rom[ 5958]='h00001b24;  wr_data_rom[ 5958]='h00001015;
    rd_cycle[ 5959] = 1'b0;  wr_cycle[ 5959] = 1'b1;  addr_rom[ 5959]='h00001da0;  wr_data_rom[ 5959]='h000013bd;
    rd_cycle[ 5960] = 1'b0;  wr_cycle[ 5960] = 1'b1;  addr_rom[ 5960]='h00001b18;  wr_data_rom[ 5960]='h00000394;
    rd_cycle[ 5961] = 1'b1;  wr_cycle[ 5961] = 1'b0;  addr_rom[ 5961]='h00000cd8;  wr_data_rom[ 5961]='h00000000;
    rd_cycle[ 5962] = 1'b1;  wr_cycle[ 5962] = 1'b0;  addr_rom[ 5962]='h000017f8;  wr_data_rom[ 5962]='h00000000;
    rd_cycle[ 5963] = 1'b1;  wr_cycle[ 5963] = 1'b0;  addr_rom[ 5963]='h00001a84;  wr_data_rom[ 5963]='h00000000;
    rd_cycle[ 5964] = 1'b1;  wr_cycle[ 5964] = 1'b0;  addr_rom[ 5964]='h00000db0;  wr_data_rom[ 5964]='h00000000;
    rd_cycle[ 5965] = 1'b1;  wr_cycle[ 5965] = 1'b0;  addr_rom[ 5965]='h000012f8;  wr_data_rom[ 5965]='h00000000;
    rd_cycle[ 5966] = 1'b0;  wr_cycle[ 5966] = 1'b1;  addr_rom[ 5966]='h000009e4;  wr_data_rom[ 5966]='h00001256;
    rd_cycle[ 5967] = 1'b1;  wr_cycle[ 5967] = 1'b0;  addr_rom[ 5967]='h00000cf0;  wr_data_rom[ 5967]='h00000000;
    rd_cycle[ 5968] = 1'b0;  wr_cycle[ 5968] = 1'b1;  addr_rom[ 5968]='h00001210;  wr_data_rom[ 5968]='h000019c6;
    rd_cycle[ 5969] = 1'b0;  wr_cycle[ 5969] = 1'b1;  addr_rom[ 5969]='h00000f78;  wr_data_rom[ 5969]='h000010ff;
    rd_cycle[ 5970] = 1'b0;  wr_cycle[ 5970] = 1'b1;  addr_rom[ 5970]='h000015e4;  wr_data_rom[ 5970]='h000013c6;
    rd_cycle[ 5971] = 1'b1;  wr_cycle[ 5971] = 1'b0;  addr_rom[ 5971]='h0000092c;  wr_data_rom[ 5971]='h00000000;
    rd_cycle[ 5972] = 1'b0;  wr_cycle[ 5972] = 1'b1;  addr_rom[ 5972]='h00000110;  wr_data_rom[ 5972]='h0000140c;
    rd_cycle[ 5973] = 1'b0;  wr_cycle[ 5973] = 1'b1;  addr_rom[ 5973]='h00000f64;  wr_data_rom[ 5973]='h0000156f;
    rd_cycle[ 5974] = 1'b1;  wr_cycle[ 5974] = 1'b0;  addr_rom[ 5974]='h00001788;  wr_data_rom[ 5974]='h00000000;
    rd_cycle[ 5975] = 1'b1;  wr_cycle[ 5975] = 1'b0;  addr_rom[ 5975]='h00001860;  wr_data_rom[ 5975]='h00000000;
    rd_cycle[ 5976] = 1'b0;  wr_cycle[ 5976] = 1'b1;  addr_rom[ 5976]='h000011ac;  wr_data_rom[ 5976]='h00000926;
    rd_cycle[ 5977] = 1'b0;  wr_cycle[ 5977] = 1'b1;  addr_rom[ 5977]='h00000da0;  wr_data_rom[ 5977]='h00001dcb;
    rd_cycle[ 5978] = 1'b0;  wr_cycle[ 5978] = 1'b1;  addr_rom[ 5978]='h000015c8;  wr_data_rom[ 5978]='h00001439;
    rd_cycle[ 5979] = 1'b0;  wr_cycle[ 5979] = 1'b1;  addr_rom[ 5979]='h0000175c;  wr_data_rom[ 5979]='h00001b99;
    rd_cycle[ 5980] = 1'b0;  wr_cycle[ 5980] = 1'b1;  addr_rom[ 5980]='h00001ab4;  wr_data_rom[ 5980]='h000011e9;
    rd_cycle[ 5981] = 1'b1;  wr_cycle[ 5981] = 1'b0;  addr_rom[ 5981]='h00000de4;  wr_data_rom[ 5981]='h00000000;
    rd_cycle[ 5982] = 1'b1;  wr_cycle[ 5982] = 1'b0;  addr_rom[ 5982]='h00000bb4;  wr_data_rom[ 5982]='h00000000;
    rd_cycle[ 5983] = 1'b1;  wr_cycle[ 5983] = 1'b0;  addr_rom[ 5983]='h000008e8;  wr_data_rom[ 5983]='h00000000;
    rd_cycle[ 5984] = 1'b0;  wr_cycle[ 5984] = 1'b1;  addr_rom[ 5984]='h00001964;  wr_data_rom[ 5984]='h0000090c;
    rd_cycle[ 5985] = 1'b0;  wr_cycle[ 5985] = 1'b1;  addr_rom[ 5985]='h0000144c;  wr_data_rom[ 5985]='h000014c5;
    rd_cycle[ 5986] = 1'b1;  wr_cycle[ 5986] = 1'b0;  addr_rom[ 5986]='h000006c4;  wr_data_rom[ 5986]='h00000000;
    rd_cycle[ 5987] = 1'b1;  wr_cycle[ 5987] = 1'b0;  addr_rom[ 5987]='h0000034c;  wr_data_rom[ 5987]='h00000000;
    rd_cycle[ 5988] = 1'b0;  wr_cycle[ 5988] = 1'b1;  addr_rom[ 5988]='h000009f4;  wr_data_rom[ 5988]='h0000113b;
    rd_cycle[ 5989] = 1'b1;  wr_cycle[ 5989] = 1'b0;  addr_rom[ 5989]='h00000228;  wr_data_rom[ 5989]='h00000000;
    rd_cycle[ 5990] = 1'b1;  wr_cycle[ 5990] = 1'b0;  addr_rom[ 5990]='h00001434;  wr_data_rom[ 5990]='h00000000;
    rd_cycle[ 5991] = 1'b1;  wr_cycle[ 5991] = 1'b0;  addr_rom[ 5991]='h00000e74;  wr_data_rom[ 5991]='h00000000;
    rd_cycle[ 5992] = 1'b1;  wr_cycle[ 5992] = 1'b0;  addr_rom[ 5992]='h00000c0c;  wr_data_rom[ 5992]='h00000000;
    rd_cycle[ 5993] = 1'b1;  wr_cycle[ 5993] = 1'b0;  addr_rom[ 5993]='h00000458;  wr_data_rom[ 5993]='h00000000;
    rd_cycle[ 5994] = 1'b0;  wr_cycle[ 5994] = 1'b1;  addr_rom[ 5994]='h00000b84;  wr_data_rom[ 5994]='h00000347;
    rd_cycle[ 5995] = 1'b1;  wr_cycle[ 5995] = 1'b0;  addr_rom[ 5995]='h00000dac;  wr_data_rom[ 5995]='h00000000;
    rd_cycle[ 5996] = 1'b1;  wr_cycle[ 5996] = 1'b0;  addr_rom[ 5996]='h000007c0;  wr_data_rom[ 5996]='h00000000;
    rd_cycle[ 5997] = 1'b1;  wr_cycle[ 5997] = 1'b0;  addr_rom[ 5997]='h00001c94;  wr_data_rom[ 5997]='h00000000;
    rd_cycle[ 5998] = 1'b1;  wr_cycle[ 5998] = 1'b0;  addr_rom[ 5998]='h00001704;  wr_data_rom[ 5998]='h00000000;
    rd_cycle[ 5999] = 1'b0;  wr_cycle[ 5999] = 1'b1;  addr_rom[ 5999]='h00001ba4;  wr_data_rom[ 5999]='h00000895;
    rd_cycle[ 6000] = 1'b0;  wr_cycle[ 6000] = 1'b1;  addr_rom[ 6000]='h000001ac;  wr_data_rom[ 6000]='h000015d2;
    rd_cycle[ 6001] = 1'b1;  wr_cycle[ 6001] = 1'b0;  addr_rom[ 6001]='h00001970;  wr_data_rom[ 6001]='h00000000;
    rd_cycle[ 6002] = 1'b0;  wr_cycle[ 6002] = 1'b1;  addr_rom[ 6002]='h000005b4;  wr_data_rom[ 6002]='h0000165b;
    rd_cycle[ 6003] = 1'b1;  wr_cycle[ 6003] = 1'b0;  addr_rom[ 6003]='h00001f20;  wr_data_rom[ 6003]='h00000000;
    rd_cycle[ 6004] = 1'b1;  wr_cycle[ 6004] = 1'b0;  addr_rom[ 6004]='h00001168;  wr_data_rom[ 6004]='h00000000;
    rd_cycle[ 6005] = 1'b0;  wr_cycle[ 6005] = 1'b1;  addr_rom[ 6005]='h000011c8;  wr_data_rom[ 6005]='h00000979;
    rd_cycle[ 6006] = 1'b1;  wr_cycle[ 6006] = 1'b0;  addr_rom[ 6006]='h0000181c;  wr_data_rom[ 6006]='h00000000;
    rd_cycle[ 6007] = 1'b0;  wr_cycle[ 6007] = 1'b1;  addr_rom[ 6007]='h00001a3c;  wr_data_rom[ 6007]='h0000012e;
    rd_cycle[ 6008] = 1'b1;  wr_cycle[ 6008] = 1'b0;  addr_rom[ 6008]='h000016b8;  wr_data_rom[ 6008]='h00000000;
    rd_cycle[ 6009] = 1'b0;  wr_cycle[ 6009] = 1'b1;  addr_rom[ 6009]='h000016d0;  wr_data_rom[ 6009]='h000008fc;
    rd_cycle[ 6010] = 1'b0;  wr_cycle[ 6010] = 1'b1;  addr_rom[ 6010]='h000011d0;  wr_data_rom[ 6010]='h000015ae;
    rd_cycle[ 6011] = 1'b0;  wr_cycle[ 6011] = 1'b1;  addr_rom[ 6011]='h00001ce8;  wr_data_rom[ 6011]='h000000f0;
    rd_cycle[ 6012] = 1'b1;  wr_cycle[ 6012] = 1'b0;  addr_rom[ 6012]='h000006bc;  wr_data_rom[ 6012]='h00000000;
    rd_cycle[ 6013] = 1'b0;  wr_cycle[ 6013] = 1'b1;  addr_rom[ 6013]='h00000148;  wr_data_rom[ 6013]='h00001724;
    rd_cycle[ 6014] = 1'b1;  wr_cycle[ 6014] = 1'b0;  addr_rom[ 6014]='h00001620;  wr_data_rom[ 6014]='h00000000;
    rd_cycle[ 6015] = 1'b1;  wr_cycle[ 6015] = 1'b0;  addr_rom[ 6015]='h000015b8;  wr_data_rom[ 6015]='h00000000;
    rd_cycle[ 6016] = 1'b1;  wr_cycle[ 6016] = 1'b0;  addr_rom[ 6016]='h00000de8;  wr_data_rom[ 6016]='h00000000;
    rd_cycle[ 6017] = 1'b0;  wr_cycle[ 6017] = 1'b1;  addr_rom[ 6017]='h00000130;  wr_data_rom[ 6017]='h00001a60;
    rd_cycle[ 6018] = 1'b1;  wr_cycle[ 6018] = 1'b0;  addr_rom[ 6018]='h00001bd4;  wr_data_rom[ 6018]='h00000000;
    rd_cycle[ 6019] = 1'b0;  wr_cycle[ 6019] = 1'b1;  addr_rom[ 6019]='h00000584;  wr_data_rom[ 6019]='h00001053;
    rd_cycle[ 6020] = 1'b0;  wr_cycle[ 6020] = 1'b1;  addr_rom[ 6020]='h00000e70;  wr_data_rom[ 6020]='h000007ea;
    rd_cycle[ 6021] = 1'b0;  wr_cycle[ 6021] = 1'b1;  addr_rom[ 6021]='h000016dc;  wr_data_rom[ 6021]='h00001a5b;
    rd_cycle[ 6022] = 1'b0;  wr_cycle[ 6022] = 1'b1;  addr_rom[ 6022]='h000010d0;  wr_data_rom[ 6022]='h00000a79;
    rd_cycle[ 6023] = 1'b1;  wr_cycle[ 6023] = 1'b0;  addr_rom[ 6023]='h00000228;  wr_data_rom[ 6023]='h00000000;
    rd_cycle[ 6024] = 1'b0;  wr_cycle[ 6024] = 1'b1;  addr_rom[ 6024]='h00001164;  wr_data_rom[ 6024]='h00000f3d;
    rd_cycle[ 6025] = 1'b1;  wr_cycle[ 6025] = 1'b0;  addr_rom[ 6025]='h000019f4;  wr_data_rom[ 6025]='h00000000;
    rd_cycle[ 6026] = 1'b0;  wr_cycle[ 6026] = 1'b1;  addr_rom[ 6026]='h000011e0;  wr_data_rom[ 6026]='h0000184a;
    rd_cycle[ 6027] = 1'b1;  wr_cycle[ 6027] = 1'b0;  addr_rom[ 6027]='h00001838;  wr_data_rom[ 6027]='h00000000;
    rd_cycle[ 6028] = 1'b0;  wr_cycle[ 6028] = 1'b1;  addr_rom[ 6028]='h00001a9c;  wr_data_rom[ 6028]='h00000778;
    rd_cycle[ 6029] = 1'b1;  wr_cycle[ 6029] = 1'b0;  addr_rom[ 6029]='h00000c04;  wr_data_rom[ 6029]='h00000000;
    rd_cycle[ 6030] = 1'b1;  wr_cycle[ 6030] = 1'b0;  addr_rom[ 6030]='h00000f64;  wr_data_rom[ 6030]='h00000000;
    rd_cycle[ 6031] = 1'b0;  wr_cycle[ 6031] = 1'b1;  addr_rom[ 6031]='h000012b8;  wr_data_rom[ 6031]='h00000e37;
    rd_cycle[ 6032] = 1'b0;  wr_cycle[ 6032] = 1'b1;  addr_rom[ 6032]='h00001344;  wr_data_rom[ 6032]='h0000193b;
    rd_cycle[ 6033] = 1'b0;  wr_cycle[ 6033] = 1'b1;  addr_rom[ 6033]='h0000134c;  wr_data_rom[ 6033]='h00000efc;
    rd_cycle[ 6034] = 1'b1;  wr_cycle[ 6034] = 1'b0;  addr_rom[ 6034]='h00001130;  wr_data_rom[ 6034]='h00000000;
    rd_cycle[ 6035] = 1'b1;  wr_cycle[ 6035] = 1'b0;  addr_rom[ 6035]='h00000dc4;  wr_data_rom[ 6035]='h00000000;
    rd_cycle[ 6036] = 1'b1;  wr_cycle[ 6036] = 1'b0;  addr_rom[ 6036]='h000015f8;  wr_data_rom[ 6036]='h00000000;
    rd_cycle[ 6037] = 1'b0;  wr_cycle[ 6037] = 1'b1;  addr_rom[ 6037]='h00001d28;  wr_data_rom[ 6037]='h00000b8f;
    rd_cycle[ 6038] = 1'b0;  wr_cycle[ 6038] = 1'b1;  addr_rom[ 6038]='h000018e8;  wr_data_rom[ 6038]='h00000a30;
    rd_cycle[ 6039] = 1'b0;  wr_cycle[ 6039] = 1'b1;  addr_rom[ 6039]='h00000a24;  wr_data_rom[ 6039]='h0000155a;
    rd_cycle[ 6040] = 1'b1;  wr_cycle[ 6040] = 1'b0;  addr_rom[ 6040]='h00001a40;  wr_data_rom[ 6040]='h00000000;
    rd_cycle[ 6041] = 1'b1;  wr_cycle[ 6041] = 1'b0;  addr_rom[ 6041]='h00001aec;  wr_data_rom[ 6041]='h00000000;
    rd_cycle[ 6042] = 1'b1;  wr_cycle[ 6042] = 1'b0;  addr_rom[ 6042]='h000006f8;  wr_data_rom[ 6042]='h00000000;
    rd_cycle[ 6043] = 1'b1;  wr_cycle[ 6043] = 1'b0;  addr_rom[ 6043]='h000015b0;  wr_data_rom[ 6043]='h00000000;
    rd_cycle[ 6044] = 1'b1;  wr_cycle[ 6044] = 1'b0;  addr_rom[ 6044]='h00000a78;  wr_data_rom[ 6044]='h00000000;
    rd_cycle[ 6045] = 1'b0;  wr_cycle[ 6045] = 1'b1;  addr_rom[ 6045]='h00000264;  wr_data_rom[ 6045]='h0000009c;
    rd_cycle[ 6046] = 1'b0;  wr_cycle[ 6046] = 1'b1;  addr_rom[ 6046]='h00001e68;  wr_data_rom[ 6046]='h00001b87;
    rd_cycle[ 6047] = 1'b0;  wr_cycle[ 6047] = 1'b1;  addr_rom[ 6047]='h00001c94;  wr_data_rom[ 6047]='h00000f10;
    rd_cycle[ 6048] = 1'b1;  wr_cycle[ 6048] = 1'b0;  addr_rom[ 6048]='h0000076c;  wr_data_rom[ 6048]='h00000000;
    rd_cycle[ 6049] = 1'b1;  wr_cycle[ 6049] = 1'b0;  addr_rom[ 6049]='h000015e4;  wr_data_rom[ 6049]='h00000000;
    rd_cycle[ 6050] = 1'b0;  wr_cycle[ 6050] = 1'b1;  addr_rom[ 6050]='h0000123c;  wr_data_rom[ 6050]='h00001a5a;
    rd_cycle[ 6051] = 1'b1;  wr_cycle[ 6051] = 1'b0;  addr_rom[ 6051]='h00001774;  wr_data_rom[ 6051]='h00000000;
    rd_cycle[ 6052] = 1'b0;  wr_cycle[ 6052] = 1'b1;  addr_rom[ 6052]='h00000bc8;  wr_data_rom[ 6052]='h00001dcd;
    rd_cycle[ 6053] = 1'b0;  wr_cycle[ 6053] = 1'b1;  addr_rom[ 6053]='h00001b20;  wr_data_rom[ 6053]='h00001d6e;
    rd_cycle[ 6054] = 1'b0;  wr_cycle[ 6054] = 1'b1;  addr_rom[ 6054]='h00000374;  wr_data_rom[ 6054]='h00000d02;
    rd_cycle[ 6055] = 1'b0;  wr_cycle[ 6055] = 1'b1;  addr_rom[ 6055]='h00001e70;  wr_data_rom[ 6055]='h0000151e;
    rd_cycle[ 6056] = 1'b1;  wr_cycle[ 6056] = 1'b0;  addr_rom[ 6056]='h000009a4;  wr_data_rom[ 6056]='h00000000;
    rd_cycle[ 6057] = 1'b0;  wr_cycle[ 6057] = 1'b1;  addr_rom[ 6057]='h00000c68;  wr_data_rom[ 6057]='h000014b0;
    rd_cycle[ 6058] = 1'b1;  wr_cycle[ 6058] = 1'b0;  addr_rom[ 6058]='h00001568;  wr_data_rom[ 6058]='h00000000;
    rd_cycle[ 6059] = 1'b0;  wr_cycle[ 6059] = 1'b1;  addr_rom[ 6059]='h0000166c;  wr_data_rom[ 6059]='h00000691;
    rd_cycle[ 6060] = 1'b0;  wr_cycle[ 6060] = 1'b1;  addr_rom[ 6060]='h000002ac;  wr_data_rom[ 6060]='h000006ce;
    rd_cycle[ 6061] = 1'b0;  wr_cycle[ 6061] = 1'b1;  addr_rom[ 6061]='h00001bec;  wr_data_rom[ 6061]='h00001992;
    rd_cycle[ 6062] = 1'b1;  wr_cycle[ 6062] = 1'b0;  addr_rom[ 6062]='h00000c70;  wr_data_rom[ 6062]='h00000000;
    rd_cycle[ 6063] = 1'b0;  wr_cycle[ 6063] = 1'b1;  addr_rom[ 6063]='h00000bc4;  wr_data_rom[ 6063]='h00001b78;
    rd_cycle[ 6064] = 1'b0;  wr_cycle[ 6064] = 1'b1;  addr_rom[ 6064]='h00001624;  wr_data_rom[ 6064]='h000007e0;
    rd_cycle[ 6065] = 1'b0;  wr_cycle[ 6065] = 1'b1;  addr_rom[ 6065]='h000000ec;  wr_data_rom[ 6065]='h000019d1;
    rd_cycle[ 6066] = 1'b1;  wr_cycle[ 6066] = 1'b0;  addr_rom[ 6066]='h00000f38;  wr_data_rom[ 6066]='h00000000;
    rd_cycle[ 6067] = 1'b1;  wr_cycle[ 6067] = 1'b0;  addr_rom[ 6067]='h000001a0;  wr_data_rom[ 6067]='h00000000;
    rd_cycle[ 6068] = 1'b1;  wr_cycle[ 6068] = 1'b0;  addr_rom[ 6068]='h00000cd8;  wr_data_rom[ 6068]='h00000000;
    rd_cycle[ 6069] = 1'b1;  wr_cycle[ 6069] = 1'b0;  addr_rom[ 6069]='h000010c8;  wr_data_rom[ 6069]='h00000000;
    rd_cycle[ 6070] = 1'b1;  wr_cycle[ 6070] = 1'b0;  addr_rom[ 6070]='h000003f4;  wr_data_rom[ 6070]='h00000000;
    rd_cycle[ 6071] = 1'b1;  wr_cycle[ 6071] = 1'b0;  addr_rom[ 6071]='h000002bc;  wr_data_rom[ 6071]='h00000000;
    rd_cycle[ 6072] = 1'b0;  wr_cycle[ 6072] = 1'b1;  addr_rom[ 6072]='h0000116c;  wr_data_rom[ 6072]='h00001b1f;
    rd_cycle[ 6073] = 1'b1;  wr_cycle[ 6073] = 1'b0;  addr_rom[ 6073]='h00001304;  wr_data_rom[ 6073]='h00000000;
    rd_cycle[ 6074] = 1'b0;  wr_cycle[ 6074] = 1'b1;  addr_rom[ 6074]='h00001758;  wr_data_rom[ 6074]='h00000b7e;
    rd_cycle[ 6075] = 1'b1;  wr_cycle[ 6075] = 1'b0;  addr_rom[ 6075]='h00001e6c;  wr_data_rom[ 6075]='h00000000;
    rd_cycle[ 6076] = 1'b1;  wr_cycle[ 6076] = 1'b0;  addr_rom[ 6076]='h000000a0;  wr_data_rom[ 6076]='h00000000;
    rd_cycle[ 6077] = 1'b0;  wr_cycle[ 6077] = 1'b1;  addr_rom[ 6077]='h0000156c;  wr_data_rom[ 6077]='h00001ea5;
    rd_cycle[ 6078] = 1'b0;  wr_cycle[ 6078] = 1'b1;  addr_rom[ 6078]='h000004e8;  wr_data_rom[ 6078]='h00000769;
    rd_cycle[ 6079] = 1'b0;  wr_cycle[ 6079] = 1'b1;  addr_rom[ 6079]='h00000374;  wr_data_rom[ 6079]='h00000702;
    rd_cycle[ 6080] = 1'b1;  wr_cycle[ 6080] = 1'b0;  addr_rom[ 6080]='h00000608;  wr_data_rom[ 6080]='h00000000;
    rd_cycle[ 6081] = 1'b1;  wr_cycle[ 6081] = 1'b0;  addr_rom[ 6081]='h000009c0;  wr_data_rom[ 6081]='h00000000;
    rd_cycle[ 6082] = 1'b1;  wr_cycle[ 6082] = 1'b0;  addr_rom[ 6082]='h00001104;  wr_data_rom[ 6082]='h00000000;
    rd_cycle[ 6083] = 1'b0;  wr_cycle[ 6083] = 1'b1;  addr_rom[ 6083]='h00001cdc;  wr_data_rom[ 6083]='h00000d18;
    rd_cycle[ 6084] = 1'b0;  wr_cycle[ 6084] = 1'b1;  addr_rom[ 6084]='h000002bc;  wr_data_rom[ 6084]='h00000aa4;
    rd_cycle[ 6085] = 1'b0;  wr_cycle[ 6085] = 1'b1;  addr_rom[ 6085]='h00000e88;  wr_data_rom[ 6085]='h00000173;
    rd_cycle[ 6086] = 1'b1;  wr_cycle[ 6086] = 1'b0;  addr_rom[ 6086]='h000006ac;  wr_data_rom[ 6086]='h00000000;
    rd_cycle[ 6087] = 1'b1;  wr_cycle[ 6087] = 1'b0;  addr_rom[ 6087]='h00000444;  wr_data_rom[ 6087]='h00000000;
    rd_cycle[ 6088] = 1'b1;  wr_cycle[ 6088] = 1'b0;  addr_rom[ 6088]='h000015c8;  wr_data_rom[ 6088]='h00000000;
    rd_cycle[ 6089] = 1'b1;  wr_cycle[ 6089] = 1'b0;  addr_rom[ 6089]='h0000078c;  wr_data_rom[ 6089]='h00000000;
    rd_cycle[ 6090] = 1'b0;  wr_cycle[ 6090] = 1'b1;  addr_rom[ 6090]='h00000ac4;  wr_data_rom[ 6090]='h00001eb6;
    rd_cycle[ 6091] = 1'b1;  wr_cycle[ 6091] = 1'b0;  addr_rom[ 6091]='h00000274;  wr_data_rom[ 6091]='h00000000;
    rd_cycle[ 6092] = 1'b1;  wr_cycle[ 6092] = 1'b0;  addr_rom[ 6092]='h00000f90;  wr_data_rom[ 6092]='h00000000;
    rd_cycle[ 6093] = 1'b0;  wr_cycle[ 6093] = 1'b1;  addr_rom[ 6093]='h000018b0;  wr_data_rom[ 6093]='h000010da;
    rd_cycle[ 6094] = 1'b1;  wr_cycle[ 6094] = 1'b0;  addr_rom[ 6094]='h0000178c;  wr_data_rom[ 6094]='h00000000;
    rd_cycle[ 6095] = 1'b0;  wr_cycle[ 6095] = 1'b1;  addr_rom[ 6095]='h00001510;  wr_data_rom[ 6095]='h000003ed;
    rd_cycle[ 6096] = 1'b0;  wr_cycle[ 6096] = 1'b1;  addr_rom[ 6096]='h00000f30;  wr_data_rom[ 6096]='h0000037a;
    rd_cycle[ 6097] = 1'b0;  wr_cycle[ 6097] = 1'b1;  addr_rom[ 6097]='h00001710;  wr_data_rom[ 6097]='h00001d93;
    rd_cycle[ 6098] = 1'b1;  wr_cycle[ 6098] = 1'b0;  addr_rom[ 6098]='h00000f20;  wr_data_rom[ 6098]='h00000000;
    rd_cycle[ 6099] = 1'b1;  wr_cycle[ 6099] = 1'b0;  addr_rom[ 6099]='h00001cd0;  wr_data_rom[ 6099]='h00000000;
    rd_cycle[ 6100] = 1'b1;  wr_cycle[ 6100] = 1'b0;  addr_rom[ 6100]='h00001110;  wr_data_rom[ 6100]='h00000000;
    rd_cycle[ 6101] = 1'b0;  wr_cycle[ 6101] = 1'b1;  addr_rom[ 6101]='h0000053c;  wr_data_rom[ 6101]='h0000153c;
    rd_cycle[ 6102] = 1'b1;  wr_cycle[ 6102] = 1'b0;  addr_rom[ 6102]='h00001394;  wr_data_rom[ 6102]='h00000000;
    rd_cycle[ 6103] = 1'b1;  wr_cycle[ 6103] = 1'b0;  addr_rom[ 6103]='h00000984;  wr_data_rom[ 6103]='h00000000;
    rd_cycle[ 6104] = 1'b0;  wr_cycle[ 6104] = 1'b1;  addr_rom[ 6104]='h000004dc;  wr_data_rom[ 6104]='h0000170a;
    rd_cycle[ 6105] = 1'b1;  wr_cycle[ 6105] = 1'b0;  addr_rom[ 6105]='h00001f28;  wr_data_rom[ 6105]='h00000000;
    rd_cycle[ 6106] = 1'b1;  wr_cycle[ 6106] = 1'b0;  addr_rom[ 6106]='h00001260;  wr_data_rom[ 6106]='h00000000;
    rd_cycle[ 6107] = 1'b0;  wr_cycle[ 6107] = 1'b1;  addr_rom[ 6107]='h00001444;  wr_data_rom[ 6107]='h00001905;
    rd_cycle[ 6108] = 1'b0;  wr_cycle[ 6108] = 1'b1;  addr_rom[ 6108]='h00000de0;  wr_data_rom[ 6108]='h00000175;
    rd_cycle[ 6109] = 1'b1;  wr_cycle[ 6109] = 1'b0;  addr_rom[ 6109]='h000013e8;  wr_data_rom[ 6109]='h00000000;
    rd_cycle[ 6110] = 1'b0;  wr_cycle[ 6110] = 1'b1;  addr_rom[ 6110]='h00000ed4;  wr_data_rom[ 6110]='h000011af;
    rd_cycle[ 6111] = 1'b1;  wr_cycle[ 6111] = 1'b0;  addr_rom[ 6111]='h00001a1c;  wr_data_rom[ 6111]='h00000000;
    rd_cycle[ 6112] = 1'b1;  wr_cycle[ 6112] = 1'b0;  addr_rom[ 6112]='h00000dfc;  wr_data_rom[ 6112]='h00000000;
    rd_cycle[ 6113] = 1'b1;  wr_cycle[ 6113] = 1'b0;  addr_rom[ 6113]='h00000558;  wr_data_rom[ 6113]='h00000000;
    rd_cycle[ 6114] = 1'b1;  wr_cycle[ 6114] = 1'b0;  addr_rom[ 6114]='h00000220;  wr_data_rom[ 6114]='h00000000;
    rd_cycle[ 6115] = 1'b1;  wr_cycle[ 6115] = 1'b0;  addr_rom[ 6115]='h0000092c;  wr_data_rom[ 6115]='h00000000;
    rd_cycle[ 6116] = 1'b1;  wr_cycle[ 6116] = 1'b0;  addr_rom[ 6116]='h0000017c;  wr_data_rom[ 6116]='h00000000;
    rd_cycle[ 6117] = 1'b1;  wr_cycle[ 6117] = 1'b0;  addr_rom[ 6117]='h00000258;  wr_data_rom[ 6117]='h00000000;
    rd_cycle[ 6118] = 1'b0;  wr_cycle[ 6118] = 1'b1;  addr_rom[ 6118]='h00000f58;  wr_data_rom[ 6118]='h000005db;
    rd_cycle[ 6119] = 1'b1;  wr_cycle[ 6119] = 1'b0;  addr_rom[ 6119]='h000016a0;  wr_data_rom[ 6119]='h00000000;
    rd_cycle[ 6120] = 1'b1;  wr_cycle[ 6120] = 1'b0;  addr_rom[ 6120]='h00000f84;  wr_data_rom[ 6120]='h00000000;
    rd_cycle[ 6121] = 1'b0;  wr_cycle[ 6121] = 1'b1;  addr_rom[ 6121]='h000000c8;  wr_data_rom[ 6121]='h000012cb;
    rd_cycle[ 6122] = 1'b0;  wr_cycle[ 6122] = 1'b1;  addr_rom[ 6122]='h000018a0;  wr_data_rom[ 6122]='h00000ace;
    rd_cycle[ 6123] = 1'b1;  wr_cycle[ 6123] = 1'b0;  addr_rom[ 6123]='h00000b10;  wr_data_rom[ 6123]='h00000000;
    rd_cycle[ 6124] = 1'b0;  wr_cycle[ 6124] = 1'b1;  addr_rom[ 6124]='h000006f0;  wr_data_rom[ 6124]='h00000afd;
    rd_cycle[ 6125] = 1'b1;  wr_cycle[ 6125] = 1'b0;  addr_rom[ 6125]='h00000364;  wr_data_rom[ 6125]='h00000000;
    rd_cycle[ 6126] = 1'b1;  wr_cycle[ 6126] = 1'b0;  addr_rom[ 6126]='h000001bc;  wr_data_rom[ 6126]='h00000000;
    rd_cycle[ 6127] = 1'b1;  wr_cycle[ 6127] = 1'b0;  addr_rom[ 6127]='h00001828;  wr_data_rom[ 6127]='h00000000;
    rd_cycle[ 6128] = 1'b0;  wr_cycle[ 6128] = 1'b1;  addr_rom[ 6128]='h00001dbc;  wr_data_rom[ 6128]='h0000124a;
    rd_cycle[ 6129] = 1'b0;  wr_cycle[ 6129] = 1'b1;  addr_rom[ 6129]='h00001b20;  wr_data_rom[ 6129]='h00000e43;
    rd_cycle[ 6130] = 1'b0;  wr_cycle[ 6130] = 1'b1;  addr_rom[ 6130]='h00001188;  wr_data_rom[ 6130]='h00000474;
    rd_cycle[ 6131] = 1'b1;  wr_cycle[ 6131] = 1'b0;  addr_rom[ 6131]='h00001ba8;  wr_data_rom[ 6131]='h00000000;
    rd_cycle[ 6132] = 1'b0;  wr_cycle[ 6132] = 1'b1;  addr_rom[ 6132]='h0000043c;  wr_data_rom[ 6132]='h0000145f;
    rd_cycle[ 6133] = 1'b0;  wr_cycle[ 6133] = 1'b1;  addr_rom[ 6133]='h000015e8;  wr_data_rom[ 6133]='h00000afe;
    rd_cycle[ 6134] = 1'b0;  wr_cycle[ 6134] = 1'b1;  addr_rom[ 6134]='h0000047c;  wr_data_rom[ 6134]='h00001be4;
    rd_cycle[ 6135] = 1'b1;  wr_cycle[ 6135] = 1'b0;  addr_rom[ 6135]='h00000a8c;  wr_data_rom[ 6135]='h00000000;
    rd_cycle[ 6136] = 1'b1;  wr_cycle[ 6136] = 1'b0;  addr_rom[ 6136]='h00001190;  wr_data_rom[ 6136]='h00000000;
    rd_cycle[ 6137] = 1'b0;  wr_cycle[ 6137] = 1'b1;  addr_rom[ 6137]='h00000768;  wr_data_rom[ 6137]='h00001aa1;
    rd_cycle[ 6138] = 1'b0;  wr_cycle[ 6138] = 1'b1;  addr_rom[ 6138]='h00001048;  wr_data_rom[ 6138]='h00001184;
    rd_cycle[ 6139] = 1'b0;  wr_cycle[ 6139] = 1'b1;  addr_rom[ 6139]='h0000135c;  wr_data_rom[ 6139]='h00000dfc;
    rd_cycle[ 6140] = 1'b1;  wr_cycle[ 6140] = 1'b0;  addr_rom[ 6140]='h00000f2c;  wr_data_rom[ 6140]='h00000000;
    rd_cycle[ 6141] = 1'b1;  wr_cycle[ 6141] = 1'b0;  addr_rom[ 6141]='h00001af8;  wr_data_rom[ 6141]='h00000000;
    rd_cycle[ 6142] = 1'b1;  wr_cycle[ 6142] = 1'b0;  addr_rom[ 6142]='h00000cf8;  wr_data_rom[ 6142]='h00000000;
    rd_cycle[ 6143] = 1'b1;  wr_cycle[ 6143] = 1'b0;  addr_rom[ 6143]='h00000e44;  wr_data_rom[ 6143]='h00000000;
    rd_cycle[ 6144] = 1'b0;  wr_cycle[ 6144] = 1'b1;  addr_rom[ 6144]='h000012a8;  wr_data_rom[ 6144]='h000004e4;
    rd_cycle[ 6145] = 1'b0;  wr_cycle[ 6145] = 1'b1;  addr_rom[ 6145]='h000009c8;  wr_data_rom[ 6145]='h00001aa5;
    rd_cycle[ 6146] = 1'b1;  wr_cycle[ 6146] = 1'b0;  addr_rom[ 6146]='h0000016c;  wr_data_rom[ 6146]='h00000000;
    rd_cycle[ 6147] = 1'b1;  wr_cycle[ 6147] = 1'b0;  addr_rom[ 6147]='h00001654;  wr_data_rom[ 6147]='h00000000;
    rd_cycle[ 6148] = 1'b1;  wr_cycle[ 6148] = 1'b0;  addr_rom[ 6148]='h000018d4;  wr_data_rom[ 6148]='h00000000;
    rd_cycle[ 6149] = 1'b0;  wr_cycle[ 6149] = 1'b1;  addr_rom[ 6149]='h00000278;  wr_data_rom[ 6149]='h00001777;
    rd_cycle[ 6150] = 1'b1;  wr_cycle[ 6150] = 1'b0;  addr_rom[ 6150]='h00000cd8;  wr_data_rom[ 6150]='h00000000;
    rd_cycle[ 6151] = 1'b0;  wr_cycle[ 6151] = 1'b1;  addr_rom[ 6151]='h00001504;  wr_data_rom[ 6151]='h000009e0;
    rd_cycle[ 6152] = 1'b1;  wr_cycle[ 6152] = 1'b0;  addr_rom[ 6152]='h00001450;  wr_data_rom[ 6152]='h00000000;
    rd_cycle[ 6153] = 1'b1;  wr_cycle[ 6153] = 1'b0;  addr_rom[ 6153]='h00001584;  wr_data_rom[ 6153]='h00000000;
    rd_cycle[ 6154] = 1'b1;  wr_cycle[ 6154] = 1'b0;  addr_rom[ 6154]='h00000074;  wr_data_rom[ 6154]='h00000000;
    rd_cycle[ 6155] = 1'b0;  wr_cycle[ 6155] = 1'b1;  addr_rom[ 6155]='h00001c7c;  wr_data_rom[ 6155]='h000017c3;
    rd_cycle[ 6156] = 1'b1;  wr_cycle[ 6156] = 1'b0;  addr_rom[ 6156]='h000005c8;  wr_data_rom[ 6156]='h00000000;
    rd_cycle[ 6157] = 1'b1;  wr_cycle[ 6157] = 1'b0;  addr_rom[ 6157]='h000016d4;  wr_data_rom[ 6157]='h00000000;
    rd_cycle[ 6158] = 1'b1;  wr_cycle[ 6158] = 1'b0;  addr_rom[ 6158]='h00000ac0;  wr_data_rom[ 6158]='h00000000;
    rd_cycle[ 6159] = 1'b1;  wr_cycle[ 6159] = 1'b0;  addr_rom[ 6159]='h00000234;  wr_data_rom[ 6159]='h00000000;
    rd_cycle[ 6160] = 1'b0;  wr_cycle[ 6160] = 1'b1;  addr_rom[ 6160]='h00001c5c;  wr_data_rom[ 6160]='h00000b87;
    rd_cycle[ 6161] = 1'b0;  wr_cycle[ 6161] = 1'b1;  addr_rom[ 6161]='h000017d4;  wr_data_rom[ 6161]='h00001713;
    rd_cycle[ 6162] = 1'b1;  wr_cycle[ 6162] = 1'b0;  addr_rom[ 6162]='h00001ad0;  wr_data_rom[ 6162]='h00000000;
    rd_cycle[ 6163] = 1'b1;  wr_cycle[ 6163] = 1'b0;  addr_rom[ 6163]='h00001d30;  wr_data_rom[ 6163]='h00000000;
    rd_cycle[ 6164] = 1'b1;  wr_cycle[ 6164] = 1'b0;  addr_rom[ 6164]='h00001ce8;  wr_data_rom[ 6164]='h00000000;
    rd_cycle[ 6165] = 1'b1;  wr_cycle[ 6165] = 1'b0;  addr_rom[ 6165]='h0000171c;  wr_data_rom[ 6165]='h00000000;
    rd_cycle[ 6166] = 1'b1;  wr_cycle[ 6166] = 1'b0;  addr_rom[ 6166]='h00001454;  wr_data_rom[ 6166]='h00000000;
    rd_cycle[ 6167] = 1'b0;  wr_cycle[ 6167] = 1'b1;  addr_rom[ 6167]='h0000100c;  wr_data_rom[ 6167]='h00000183;
    rd_cycle[ 6168] = 1'b0;  wr_cycle[ 6168] = 1'b1;  addr_rom[ 6168]='h000011f8;  wr_data_rom[ 6168]='h0000184e;
    rd_cycle[ 6169] = 1'b0;  wr_cycle[ 6169] = 1'b1;  addr_rom[ 6169]='h0000133c;  wr_data_rom[ 6169]='h00000389;
    rd_cycle[ 6170] = 1'b0;  wr_cycle[ 6170] = 1'b1;  addr_rom[ 6170]='h000018b0;  wr_data_rom[ 6170]='h0000078a;
    rd_cycle[ 6171] = 1'b0;  wr_cycle[ 6171] = 1'b1;  addr_rom[ 6171]='h0000175c;  wr_data_rom[ 6171]='h000018e2;
    rd_cycle[ 6172] = 1'b0;  wr_cycle[ 6172] = 1'b1;  addr_rom[ 6172]='h000008d8;  wr_data_rom[ 6172]='h00001d16;
    rd_cycle[ 6173] = 1'b0;  wr_cycle[ 6173] = 1'b1;  addr_rom[ 6173]='h00000ddc;  wr_data_rom[ 6173]='h00001ed1;
    rd_cycle[ 6174] = 1'b0;  wr_cycle[ 6174] = 1'b1;  addr_rom[ 6174]='h00000488;  wr_data_rom[ 6174]='h000004a5;
    rd_cycle[ 6175] = 1'b1;  wr_cycle[ 6175] = 1'b0;  addr_rom[ 6175]='h0000136c;  wr_data_rom[ 6175]='h00000000;
    rd_cycle[ 6176] = 1'b0;  wr_cycle[ 6176] = 1'b1;  addr_rom[ 6176]='h00000308;  wr_data_rom[ 6176]='h000008f9;
    rd_cycle[ 6177] = 1'b1;  wr_cycle[ 6177] = 1'b0;  addr_rom[ 6177]='h000018a4;  wr_data_rom[ 6177]='h00000000;
    rd_cycle[ 6178] = 1'b0;  wr_cycle[ 6178] = 1'b1;  addr_rom[ 6178]='h000009ec;  wr_data_rom[ 6178]='h00000c11;
    rd_cycle[ 6179] = 1'b1;  wr_cycle[ 6179] = 1'b0;  addr_rom[ 6179]='h00001070;  wr_data_rom[ 6179]='h00000000;
    rd_cycle[ 6180] = 1'b1;  wr_cycle[ 6180] = 1'b0;  addr_rom[ 6180]='h00001a9c;  wr_data_rom[ 6180]='h00000000;
    rd_cycle[ 6181] = 1'b0;  wr_cycle[ 6181] = 1'b1;  addr_rom[ 6181]='h000010f0;  wr_data_rom[ 6181]='h0000121b;
    rd_cycle[ 6182] = 1'b0;  wr_cycle[ 6182] = 1'b1;  addr_rom[ 6182]='h00000bcc;  wr_data_rom[ 6182]='h00000bc6;
    rd_cycle[ 6183] = 1'b1;  wr_cycle[ 6183] = 1'b0;  addr_rom[ 6183]='h00000574;  wr_data_rom[ 6183]='h00000000;
    rd_cycle[ 6184] = 1'b0;  wr_cycle[ 6184] = 1'b1;  addr_rom[ 6184]='h0000083c;  wr_data_rom[ 6184]='h000010f9;
    rd_cycle[ 6185] = 1'b0;  wr_cycle[ 6185] = 1'b1;  addr_rom[ 6185]='h00001350;  wr_data_rom[ 6185]='h00000fc8;
    rd_cycle[ 6186] = 1'b0;  wr_cycle[ 6186] = 1'b1;  addr_rom[ 6186]='h00000328;  wr_data_rom[ 6186]='h000017f8;
    rd_cycle[ 6187] = 1'b0;  wr_cycle[ 6187] = 1'b1;  addr_rom[ 6187]='h00001690;  wr_data_rom[ 6187]='h0000162a;
    rd_cycle[ 6188] = 1'b0;  wr_cycle[ 6188] = 1'b1;  addr_rom[ 6188]='h000009b0;  wr_data_rom[ 6188]='h00001506;
    rd_cycle[ 6189] = 1'b1;  wr_cycle[ 6189] = 1'b0;  addr_rom[ 6189]='h00000df8;  wr_data_rom[ 6189]='h00000000;
    rd_cycle[ 6190] = 1'b0;  wr_cycle[ 6190] = 1'b1;  addr_rom[ 6190]='h00000980;  wr_data_rom[ 6190]='h000018d2;
    rd_cycle[ 6191] = 1'b0;  wr_cycle[ 6191] = 1'b1;  addr_rom[ 6191]='h00000a40;  wr_data_rom[ 6191]='h0000077a;
    rd_cycle[ 6192] = 1'b0;  wr_cycle[ 6192] = 1'b1;  addr_rom[ 6192]='h00000968;  wr_data_rom[ 6192]='h000019b5;
    rd_cycle[ 6193] = 1'b0;  wr_cycle[ 6193] = 1'b1;  addr_rom[ 6193]='h00000324;  wr_data_rom[ 6193]='h000014fd;
    rd_cycle[ 6194] = 1'b0;  wr_cycle[ 6194] = 1'b1;  addr_rom[ 6194]='h00001434;  wr_data_rom[ 6194]='h0000098d;
    rd_cycle[ 6195] = 1'b0;  wr_cycle[ 6195] = 1'b1;  addr_rom[ 6195]='h00001f18;  wr_data_rom[ 6195]='h00000b99;
    rd_cycle[ 6196] = 1'b1;  wr_cycle[ 6196] = 1'b0;  addr_rom[ 6196]='h0000154c;  wr_data_rom[ 6196]='h00000000;
    rd_cycle[ 6197] = 1'b0;  wr_cycle[ 6197] = 1'b1;  addr_rom[ 6197]='h000016d4;  wr_data_rom[ 6197]='h0000012b;
    rd_cycle[ 6198] = 1'b0;  wr_cycle[ 6198] = 1'b1;  addr_rom[ 6198]='h000003f8;  wr_data_rom[ 6198]='h0000013a;
    rd_cycle[ 6199] = 1'b0;  wr_cycle[ 6199] = 1'b1;  addr_rom[ 6199]='h000000ac;  wr_data_rom[ 6199]='h000011c7;
    rd_cycle[ 6200] = 1'b0;  wr_cycle[ 6200] = 1'b1;  addr_rom[ 6200]='h00001028;  wr_data_rom[ 6200]='h000013aa;
    rd_cycle[ 6201] = 1'b0;  wr_cycle[ 6201] = 1'b1;  addr_rom[ 6201]='h00000d78;  wr_data_rom[ 6201]='h00000dd6;
    rd_cycle[ 6202] = 1'b0;  wr_cycle[ 6202] = 1'b1;  addr_rom[ 6202]='h00001304;  wr_data_rom[ 6202]='h000006c0;
    rd_cycle[ 6203] = 1'b1;  wr_cycle[ 6203] = 1'b0;  addr_rom[ 6203]='h00001924;  wr_data_rom[ 6203]='h00000000;
    rd_cycle[ 6204] = 1'b0;  wr_cycle[ 6204] = 1'b1;  addr_rom[ 6204]='h00000fdc;  wr_data_rom[ 6204]='h00001f03;
    rd_cycle[ 6205] = 1'b0;  wr_cycle[ 6205] = 1'b1;  addr_rom[ 6205]='h00001d70;  wr_data_rom[ 6205]='h00000fef;
    rd_cycle[ 6206] = 1'b1;  wr_cycle[ 6206] = 1'b0;  addr_rom[ 6206]='h00000dfc;  wr_data_rom[ 6206]='h00000000;
    rd_cycle[ 6207] = 1'b1;  wr_cycle[ 6207] = 1'b0;  addr_rom[ 6207]='h0000045c;  wr_data_rom[ 6207]='h00000000;
    rd_cycle[ 6208] = 1'b0;  wr_cycle[ 6208] = 1'b1;  addr_rom[ 6208]='h00000058;  wr_data_rom[ 6208]='h00000858;
    rd_cycle[ 6209] = 1'b0;  wr_cycle[ 6209] = 1'b1;  addr_rom[ 6209]='h00001bec;  wr_data_rom[ 6209]='h000006c1;
    rd_cycle[ 6210] = 1'b0;  wr_cycle[ 6210] = 1'b1;  addr_rom[ 6210]='h000001dc;  wr_data_rom[ 6210]='h000016ac;
    rd_cycle[ 6211] = 1'b1;  wr_cycle[ 6211] = 1'b0;  addr_rom[ 6211]='h00001818;  wr_data_rom[ 6211]='h00000000;
    rd_cycle[ 6212] = 1'b1;  wr_cycle[ 6212] = 1'b0;  addr_rom[ 6212]='h000011f4;  wr_data_rom[ 6212]='h00000000;
    rd_cycle[ 6213] = 1'b0;  wr_cycle[ 6213] = 1'b1;  addr_rom[ 6213]='h00000a58;  wr_data_rom[ 6213]='h0000166f;
    rd_cycle[ 6214] = 1'b0;  wr_cycle[ 6214] = 1'b1;  addr_rom[ 6214]='h00001778;  wr_data_rom[ 6214]='h0000062f;
    rd_cycle[ 6215] = 1'b1;  wr_cycle[ 6215] = 1'b0;  addr_rom[ 6215]='h000013e0;  wr_data_rom[ 6215]='h00000000;
    rd_cycle[ 6216] = 1'b0;  wr_cycle[ 6216] = 1'b1;  addr_rom[ 6216]='h00000724;  wr_data_rom[ 6216]='h00001d03;
    rd_cycle[ 6217] = 1'b1;  wr_cycle[ 6217] = 1'b0;  addr_rom[ 6217]='h0000084c;  wr_data_rom[ 6217]='h00000000;
    rd_cycle[ 6218] = 1'b0;  wr_cycle[ 6218] = 1'b1;  addr_rom[ 6218]='h00000b38;  wr_data_rom[ 6218]='h000000ba;
    rd_cycle[ 6219] = 1'b0;  wr_cycle[ 6219] = 1'b1;  addr_rom[ 6219]='h00001b14;  wr_data_rom[ 6219]='h00000c06;
    rd_cycle[ 6220] = 1'b1;  wr_cycle[ 6220] = 1'b0;  addr_rom[ 6220]='h00000b4c;  wr_data_rom[ 6220]='h00000000;
    rd_cycle[ 6221] = 1'b1;  wr_cycle[ 6221] = 1'b0;  addr_rom[ 6221]='h00000aa8;  wr_data_rom[ 6221]='h00000000;
    rd_cycle[ 6222] = 1'b1;  wr_cycle[ 6222] = 1'b0;  addr_rom[ 6222]='h00001d5c;  wr_data_rom[ 6222]='h00000000;
    rd_cycle[ 6223] = 1'b1;  wr_cycle[ 6223] = 1'b0;  addr_rom[ 6223]='h00000860;  wr_data_rom[ 6223]='h00000000;
    rd_cycle[ 6224] = 1'b0;  wr_cycle[ 6224] = 1'b1;  addr_rom[ 6224]='h000015a0;  wr_data_rom[ 6224]='h000000dc;
    rd_cycle[ 6225] = 1'b0;  wr_cycle[ 6225] = 1'b1;  addr_rom[ 6225]='h000002a8;  wr_data_rom[ 6225]='h00000261;
    rd_cycle[ 6226] = 1'b1;  wr_cycle[ 6226] = 1'b0;  addr_rom[ 6226]='h00000db4;  wr_data_rom[ 6226]='h00000000;
    rd_cycle[ 6227] = 1'b1;  wr_cycle[ 6227] = 1'b0;  addr_rom[ 6227]='h000018b0;  wr_data_rom[ 6227]='h00000000;
    rd_cycle[ 6228] = 1'b1;  wr_cycle[ 6228] = 1'b0;  addr_rom[ 6228]='h00001cfc;  wr_data_rom[ 6228]='h00000000;
    rd_cycle[ 6229] = 1'b1;  wr_cycle[ 6229] = 1'b0;  addr_rom[ 6229]='h00000050;  wr_data_rom[ 6229]='h00000000;
    rd_cycle[ 6230] = 1'b1;  wr_cycle[ 6230] = 1'b0;  addr_rom[ 6230]='h000016b0;  wr_data_rom[ 6230]='h00000000;
    rd_cycle[ 6231] = 1'b0;  wr_cycle[ 6231] = 1'b1;  addr_rom[ 6231]='h00001c38;  wr_data_rom[ 6231]='h00000f17;
    rd_cycle[ 6232] = 1'b0;  wr_cycle[ 6232] = 1'b1;  addr_rom[ 6232]='h00001434;  wr_data_rom[ 6232]='h00001e02;
    rd_cycle[ 6233] = 1'b0;  wr_cycle[ 6233] = 1'b1;  addr_rom[ 6233]='h00000f58;  wr_data_rom[ 6233]='h00000b38;
    rd_cycle[ 6234] = 1'b0;  wr_cycle[ 6234] = 1'b1;  addr_rom[ 6234]='h00001a10;  wr_data_rom[ 6234]='h00000150;
    rd_cycle[ 6235] = 1'b1;  wr_cycle[ 6235] = 1'b0;  addr_rom[ 6235]='h0000185c;  wr_data_rom[ 6235]='h00000000;
    rd_cycle[ 6236] = 1'b0;  wr_cycle[ 6236] = 1'b1;  addr_rom[ 6236]='h0000154c;  wr_data_rom[ 6236]='h000007ea;
    rd_cycle[ 6237] = 1'b0;  wr_cycle[ 6237] = 1'b1;  addr_rom[ 6237]='h00000aac;  wr_data_rom[ 6237]='h00001ac9;
    rd_cycle[ 6238] = 1'b0;  wr_cycle[ 6238] = 1'b1;  addr_rom[ 6238]='h00000220;  wr_data_rom[ 6238]='h000009b8;
    rd_cycle[ 6239] = 1'b0;  wr_cycle[ 6239] = 1'b1;  addr_rom[ 6239]='h000010cc;  wr_data_rom[ 6239]='h00000b1a;
    rd_cycle[ 6240] = 1'b0;  wr_cycle[ 6240] = 1'b1;  addr_rom[ 6240]='h00001e0c;  wr_data_rom[ 6240]='h000000df;
    rd_cycle[ 6241] = 1'b1;  wr_cycle[ 6241] = 1'b0;  addr_rom[ 6241]='h00000c0c;  wr_data_rom[ 6241]='h00000000;
    rd_cycle[ 6242] = 1'b1;  wr_cycle[ 6242] = 1'b0;  addr_rom[ 6242]='h00001898;  wr_data_rom[ 6242]='h00000000;
    rd_cycle[ 6243] = 1'b1;  wr_cycle[ 6243] = 1'b0;  addr_rom[ 6243]='h00001af4;  wr_data_rom[ 6243]='h00000000;
    rd_cycle[ 6244] = 1'b1;  wr_cycle[ 6244] = 1'b0;  addr_rom[ 6244]='h00000f28;  wr_data_rom[ 6244]='h00000000;
    rd_cycle[ 6245] = 1'b0;  wr_cycle[ 6245] = 1'b1;  addr_rom[ 6245]='h00001038;  wr_data_rom[ 6245]='h000018ee;
    rd_cycle[ 6246] = 1'b0;  wr_cycle[ 6246] = 1'b1;  addr_rom[ 6246]='h00001b88;  wr_data_rom[ 6246]='h00001c0d;
    rd_cycle[ 6247] = 1'b0;  wr_cycle[ 6247] = 1'b1;  addr_rom[ 6247]='h00001064;  wr_data_rom[ 6247]='h00000ff7;
    rd_cycle[ 6248] = 1'b1;  wr_cycle[ 6248] = 1'b0;  addr_rom[ 6248]='h00001e78;  wr_data_rom[ 6248]='h00000000;
    rd_cycle[ 6249] = 1'b1;  wr_cycle[ 6249] = 1'b0;  addr_rom[ 6249]='h0000068c;  wr_data_rom[ 6249]='h00000000;
    rd_cycle[ 6250] = 1'b0;  wr_cycle[ 6250] = 1'b1;  addr_rom[ 6250]='h00001944;  wr_data_rom[ 6250]='h00000cba;
    rd_cycle[ 6251] = 1'b0;  wr_cycle[ 6251] = 1'b1;  addr_rom[ 6251]='h00001cb8;  wr_data_rom[ 6251]='h00000fcc;
    rd_cycle[ 6252] = 1'b0;  wr_cycle[ 6252] = 1'b1;  addr_rom[ 6252]='h000001b4;  wr_data_rom[ 6252]='h000012ee;
    rd_cycle[ 6253] = 1'b0;  wr_cycle[ 6253] = 1'b1;  addr_rom[ 6253]='h0000008c;  wr_data_rom[ 6253]='h0000068d;
    rd_cycle[ 6254] = 1'b0;  wr_cycle[ 6254] = 1'b1;  addr_rom[ 6254]='h0000103c;  wr_data_rom[ 6254]='h0000145f;
    rd_cycle[ 6255] = 1'b1;  wr_cycle[ 6255] = 1'b0;  addr_rom[ 6255]='h00001804;  wr_data_rom[ 6255]='h00000000;
    rd_cycle[ 6256] = 1'b0;  wr_cycle[ 6256] = 1'b1;  addr_rom[ 6256]='h00001334;  wr_data_rom[ 6256]='h000019a5;
    rd_cycle[ 6257] = 1'b0;  wr_cycle[ 6257] = 1'b1;  addr_rom[ 6257]='h00000ea8;  wr_data_rom[ 6257]='h000013d1;
    rd_cycle[ 6258] = 1'b1;  wr_cycle[ 6258] = 1'b0;  addr_rom[ 6258]='h000007f4;  wr_data_rom[ 6258]='h00000000;
    rd_cycle[ 6259] = 1'b1;  wr_cycle[ 6259] = 1'b0;  addr_rom[ 6259]='h000002f4;  wr_data_rom[ 6259]='h00000000;
    rd_cycle[ 6260] = 1'b1;  wr_cycle[ 6260] = 1'b0;  addr_rom[ 6260]='h00001168;  wr_data_rom[ 6260]='h00000000;
    rd_cycle[ 6261] = 1'b0;  wr_cycle[ 6261] = 1'b1;  addr_rom[ 6261]='h000018a0;  wr_data_rom[ 6261]='h00000445;
    rd_cycle[ 6262] = 1'b1;  wr_cycle[ 6262] = 1'b0;  addr_rom[ 6262]='h00001454;  wr_data_rom[ 6262]='h00000000;
    rd_cycle[ 6263] = 1'b0;  wr_cycle[ 6263] = 1'b1;  addr_rom[ 6263]='h00000d88;  wr_data_rom[ 6263]='h000001da;
    rd_cycle[ 6264] = 1'b0;  wr_cycle[ 6264] = 1'b1;  addr_rom[ 6264]='h00001a14;  wr_data_rom[ 6264]='h00001a84;
    rd_cycle[ 6265] = 1'b1;  wr_cycle[ 6265] = 1'b0;  addr_rom[ 6265]='h00000780;  wr_data_rom[ 6265]='h00000000;
    rd_cycle[ 6266] = 1'b1;  wr_cycle[ 6266] = 1'b0;  addr_rom[ 6266]='h00001b98;  wr_data_rom[ 6266]='h00000000;
    rd_cycle[ 6267] = 1'b1;  wr_cycle[ 6267] = 1'b0;  addr_rom[ 6267]='h00001734;  wr_data_rom[ 6267]='h00000000;
    rd_cycle[ 6268] = 1'b0;  wr_cycle[ 6268] = 1'b1;  addr_rom[ 6268]='h00000918;  wr_data_rom[ 6268]='h00001d61;
    rd_cycle[ 6269] = 1'b1;  wr_cycle[ 6269] = 1'b0;  addr_rom[ 6269]='h000001fc;  wr_data_rom[ 6269]='h00000000;
    rd_cycle[ 6270] = 1'b0;  wr_cycle[ 6270] = 1'b1;  addr_rom[ 6270]='h000015c8;  wr_data_rom[ 6270]='h00001437;
    rd_cycle[ 6271] = 1'b0;  wr_cycle[ 6271] = 1'b1;  addr_rom[ 6271]='h00001544;  wr_data_rom[ 6271]='h0000192d;
    rd_cycle[ 6272] = 1'b1;  wr_cycle[ 6272] = 1'b0;  addr_rom[ 6272]='h00001af8;  wr_data_rom[ 6272]='h00000000;
    rd_cycle[ 6273] = 1'b0;  wr_cycle[ 6273] = 1'b1;  addr_rom[ 6273]='h00000f94;  wr_data_rom[ 6273]='h0000094d;
    rd_cycle[ 6274] = 1'b1;  wr_cycle[ 6274] = 1'b0;  addr_rom[ 6274]='h00001d7c;  wr_data_rom[ 6274]='h00000000;
    rd_cycle[ 6275] = 1'b1;  wr_cycle[ 6275] = 1'b0;  addr_rom[ 6275]='h00000510;  wr_data_rom[ 6275]='h00000000;
    rd_cycle[ 6276] = 1'b1;  wr_cycle[ 6276] = 1'b0;  addr_rom[ 6276]='h00000930;  wr_data_rom[ 6276]='h00000000;
    rd_cycle[ 6277] = 1'b1;  wr_cycle[ 6277] = 1'b0;  addr_rom[ 6277]='h00001d04;  wr_data_rom[ 6277]='h00000000;
    rd_cycle[ 6278] = 1'b0;  wr_cycle[ 6278] = 1'b1;  addr_rom[ 6278]='h00001c94;  wr_data_rom[ 6278]='h00000b5f;
    rd_cycle[ 6279] = 1'b0;  wr_cycle[ 6279] = 1'b1;  addr_rom[ 6279]='h00000ebc;  wr_data_rom[ 6279]='h0000010f;
    rd_cycle[ 6280] = 1'b1;  wr_cycle[ 6280] = 1'b0;  addr_rom[ 6280]='h00001458;  wr_data_rom[ 6280]='h00000000;
    rd_cycle[ 6281] = 1'b1;  wr_cycle[ 6281] = 1'b0;  addr_rom[ 6281]='h00000a10;  wr_data_rom[ 6281]='h00000000;
    rd_cycle[ 6282] = 1'b1;  wr_cycle[ 6282] = 1'b0;  addr_rom[ 6282]='h00001f30;  wr_data_rom[ 6282]='h00000000;
    rd_cycle[ 6283] = 1'b0;  wr_cycle[ 6283] = 1'b1;  addr_rom[ 6283]='h00000f88;  wr_data_rom[ 6283]='h00000b93;
    rd_cycle[ 6284] = 1'b1;  wr_cycle[ 6284] = 1'b0;  addr_rom[ 6284]='h000007b4;  wr_data_rom[ 6284]='h00000000;
    rd_cycle[ 6285] = 1'b1;  wr_cycle[ 6285] = 1'b0;  addr_rom[ 6285]='h000005c0;  wr_data_rom[ 6285]='h00000000;
    rd_cycle[ 6286] = 1'b0;  wr_cycle[ 6286] = 1'b1;  addr_rom[ 6286]='h0000036c;  wr_data_rom[ 6286]='h00000c0a;
    rd_cycle[ 6287] = 1'b1;  wr_cycle[ 6287] = 1'b0;  addr_rom[ 6287]='h00000578;  wr_data_rom[ 6287]='h00000000;
    rd_cycle[ 6288] = 1'b1;  wr_cycle[ 6288] = 1'b0;  addr_rom[ 6288]='h000004b0;  wr_data_rom[ 6288]='h00000000;
    rd_cycle[ 6289] = 1'b0;  wr_cycle[ 6289] = 1'b1;  addr_rom[ 6289]='h000017a4;  wr_data_rom[ 6289]='h00000baf;
    rd_cycle[ 6290] = 1'b0;  wr_cycle[ 6290] = 1'b1;  addr_rom[ 6290]='h0000143c;  wr_data_rom[ 6290]='h00001c7f;
    rd_cycle[ 6291] = 1'b0;  wr_cycle[ 6291] = 1'b1;  addr_rom[ 6291]='h000014d0;  wr_data_rom[ 6291]='h00000983;
    rd_cycle[ 6292] = 1'b1;  wr_cycle[ 6292] = 1'b0;  addr_rom[ 6292]='h00001040;  wr_data_rom[ 6292]='h00000000;
    rd_cycle[ 6293] = 1'b1;  wr_cycle[ 6293] = 1'b0;  addr_rom[ 6293]='h00000f54;  wr_data_rom[ 6293]='h00000000;
    rd_cycle[ 6294] = 1'b0;  wr_cycle[ 6294] = 1'b1;  addr_rom[ 6294]='h00000e00;  wr_data_rom[ 6294]='h00000a56;
    rd_cycle[ 6295] = 1'b1;  wr_cycle[ 6295] = 1'b0;  addr_rom[ 6295]='h00000504;  wr_data_rom[ 6295]='h00000000;
    rd_cycle[ 6296] = 1'b0;  wr_cycle[ 6296] = 1'b1;  addr_rom[ 6296]='h0000084c;  wr_data_rom[ 6296]='h00000748;
    rd_cycle[ 6297] = 1'b0;  wr_cycle[ 6297] = 1'b1;  addr_rom[ 6297]='h0000023c;  wr_data_rom[ 6297]='h00001d37;
    rd_cycle[ 6298] = 1'b1;  wr_cycle[ 6298] = 1'b0;  addr_rom[ 6298]='h00000ff4;  wr_data_rom[ 6298]='h00000000;
    rd_cycle[ 6299] = 1'b1;  wr_cycle[ 6299] = 1'b0;  addr_rom[ 6299]='h00001ea4;  wr_data_rom[ 6299]='h00000000;
    rd_cycle[ 6300] = 1'b1;  wr_cycle[ 6300] = 1'b0;  addr_rom[ 6300]='h00001e28;  wr_data_rom[ 6300]='h00000000;
    rd_cycle[ 6301] = 1'b0;  wr_cycle[ 6301] = 1'b1;  addr_rom[ 6301]='h00001e78;  wr_data_rom[ 6301]='h000011cd;
    rd_cycle[ 6302] = 1'b0;  wr_cycle[ 6302] = 1'b1;  addr_rom[ 6302]='h0000196c;  wr_data_rom[ 6302]='h000013a8;
    rd_cycle[ 6303] = 1'b0;  wr_cycle[ 6303] = 1'b1;  addr_rom[ 6303]='h00001c88;  wr_data_rom[ 6303]='h00000bae;
    rd_cycle[ 6304] = 1'b1;  wr_cycle[ 6304] = 1'b0;  addr_rom[ 6304]='h00000030;  wr_data_rom[ 6304]='h00000000;
    rd_cycle[ 6305] = 1'b0;  wr_cycle[ 6305] = 1'b1;  addr_rom[ 6305]='h00001b30;  wr_data_rom[ 6305]='h00001bba;
    rd_cycle[ 6306] = 1'b0;  wr_cycle[ 6306] = 1'b1;  addr_rom[ 6306]='h00000c64;  wr_data_rom[ 6306]='h000008c3;
    rd_cycle[ 6307] = 1'b0;  wr_cycle[ 6307] = 1'b1;  addr_rom[ 6307]='h00000434;  wr_data_rom[ 6307]='h000015cb;
    rd_cycle[ 6308] = 1'b1;  wr_cycle[ 6308] = 1'b0;  addr_rom[ 6308]='h000001d8;  wr_data_rom[ 6308]='h00000000;
    rd_cycle[ 6309] = 1'b0;  wr_cycle[ 6309] = 1'b1;  addr_rom[ 6309]='h00000d2c;  wr_data_rom[ 6309]='h0000181a;
    rd_cycle[ 6310] = 1'b1;  wr_cycle[ 6310] = 1'b0;  addr_rom[ 6310]='h00001d88;  wr_data_rom[ 6310]='h00000000;
    rd_cycle[ 6311] = 1'b0;  wr_cycle[ 6311] = 1'b1;  addr_rom[ 6311]='h00001ba4;  wr_data_rom[ 6311]='h00001d5e;
    rd_cycle[ 6312] = 1'b0;  wr_cycle[ 6312] = 1'b1;  addr_rom[ 6312]='h00000898;  wr_data_rom[ 6312]='h00001cbf;
    rd_cycle[ 6313] = 1'b1;  wr_cycle[ 6313] = 1'b0;  addr_rom[ 6313]='h00001e08;  wr_data_rom[ 6313]='h00000000;
    rd_cycle[ 6314] = 1'b1;  wr_cycle[ 6314] = 1'b0;  addr_rom[ 6314]='h00000330;  wr_data_rom[ 6314]='h00000000;
    rd_cycle[ 6315] = 1'b1;  wr_cycle[ 6315] = 1'b0;  addr_rom[ 6315]='h00001534;  wr_data_rom[ 6315]='h00000000;
    rd_cycle[ 6316] = 1'b0;  wr_cycle[ 6316] = 1'b1;  addr_rom[ 6316]='h000018c4;  wr_data_rom[ 6316]='h000012bb;
    rd_cycle[ 6317] = 1'b1;  wr_cycle[ 6317] = 1'b0;  addr_rom[ 6317]='h00001aac;  wr_data_rom[ 6317]='h00000000;
    rd_cycle[ 6318] = 1'b1;  wr_cycle[ 6318] = 1'b0;  addr_rom[ 6318]='h0000125c;  wr_data_rom[ 6318]='h00000000;
    rd_cycle[ 6319] = 1'b1;  wr_cycle[ 6319] = 1'b0;  addr_rom[ 6319]='h00001eec;  wr_data_rom[ 6319]='h00000000;
    rd_cycle[ 6320] = 1'b0;  wr_cycle[ 6320] = 1'b1;  addr_rom[ 6320]='h000000f8;  wr_data_rom[ 6320]='h00000f07;
    rd_cycle[ 6321] = 1'b0;  wr_cycle[ 6321] = 1'b1;  addr_rom[ 6321]='h00000778;  wr_data_rom[ 6321]='h000013d7;
    rd_cycle[ 6322] = 1'b1;  wr_cycle[ 6322] = 1'b0;  addr_rom[ 6322]='h0000054c;  wr_data_rom[ 6322]='h00000000;
    rd_cycle[ 6323] = 1'b1;  wr_cycle[ 6323] = 1'b0;  addr_rom[ 6323]='h00001f1c;  wr_data_rom[ 6323]='h00000000;
    rd_cycle[ 6324] = 1'b0;  wr_cycle[ 6324] = 1'b1;  addr_rom[ 6324]='h000018e4;  wr_data_rom[ 6324]='h00001f03;
    rd_cycle[ 6325] = 1'b1;  wr_cycle[ 6325] = 1'b0;  addr_rom[ 6325]='h00000180;  wr_data_rom[ 6325]='h00000000;
    rd_cycle[ 6326] = 1'b1;  wr_cycle[ 6326] = 1'b0;  addr_rom[ 6326]='h00000f08;  wr_data_rom[ 6326]='h00000000;
    rd_cycle[ 6327] = 1'b0;  wr_cycle[ 6327] = 1'b1;  addr_rom[ 6327]='h00001adc;  wr_data_rom[ 6327]='h000014b8;
    rd_cycle[ 6328] = 1'b0;  wr_cycle[ 6328] = 1'b1;  addr_rom[ 6328]='h0000071c;  wr_data_rom[ 6328]='h00000dfe;
    rd_cycle[ 6329] = 1'b0;  wr_cycle[ 6329] = 1'b1;  addr_rom[ 6329]='h0000176c;  wr_data_rom[ 6329]='h00000c16;
    rd_cycle[ 6330] = 1'b1;  wr_cycle[ 6330] = 1'b0;  addr_rom[ 6330]='h00000f80;  wr_data_rom[ 6330]='h00000000;
    rd_cycle[ 6331] = 1'b1;  wr_cycle[ 6331] = 1'b0;  addr_rom[ 6331]='h00000864;  wr_data_rom[ 6331]='h00000000;
    rd_cycle[ 6332] = 1'b1;  wr_cycle[ 6332] = 1'b0;  addr_rom[ 6332]='h00000d44;  wr_data_rom[ 6332]='h00000000;
    rd_cycle[ 6333] = 1'b0;  wr_cycle[ 6333] = 1'b1;  addr_rom[ 6333]='h00001e64;  wr_data_rom[ 6333]='h00001897;
    rd_cycle[ 6334] = 1'b0;  wr_cycle[ 6334] = 1'b1;  addr_rom[ 6334]='h00001d7c;  wr_data_rom[ 6334]='h000009d6;
    rd_cycle[ 6335] = 1'b1;  wr_cycle[ 6335] = 1'b0;  addr_rom[ 6335]='h00001064;  wr_data_rom[ 6335]='h00000000;
    rd_cycle[ 6336] = 1'b0;  wr_cycle[ 6336] = 1'b1;  addr_rom[ 6336]='h000010e4;  wr_data_rom[ 6336]='h0000157e;
    rd_cycle[ 6337] = 1'b0;  wr_cycle[ 6337] = 1'b1;  addr_rom[ 6337]='h000001fc;  wr_data_rom[ 6337]='h000007d7;
    rd_cycle[ 6338] = 1'b0;  wr_cycle[ 6338] = 1'b1;  addr_rom[ 6338]='h00001b74;  wr_data_rom[ 6338]='h00001ec3;
    rd_cycle[ 6339] = 1'b1;  wr_cycle[ 6339] = 1'b0;  addr_rom[ 6339]='h00001794;  wr_data_rom[ 6339]='h00000000;
    rd_cycle[ 6340] = 1'b1;  wr_cycle[ 6340] = 1'b0;  addr_rom[ 6340]='h00001c98;  wr_data_rom[ 6340]='h00000000;
    rd_cycle[ 6341] = 1'b1;  wr_cycle[ 6341] = 1'b0;  addr_rom[ 6341]='h00001b9c;  wr_data_rom[ 6341]='h00000000;
    rd_cycle[ 6342] = 1'b1;  wr_cycle[ 6342] = 1'b0;  addr_rom[ 6342]='h000008b8;  wr_data_rom[ 6342]='h00000000;
    rd_cycle[ 6343] = 1'b0;  wr_cycle[ 6343] = 1'b1;  addr_rom[ 6343]='h00000170;  wr_data_rom[ 6343]='h00000855;
    rd_cycle[ 6344] = 1'b0;  wr_cycle[ 6344] = 1'b1;  addr_rom[ 6344]='h0000091c;  wr_data_rom[ 6344]='h00000912;
    rd_cycle[ 6345] = 1'b1;  wr_cycle[ 6345] = 1'b0;  addr_rom[ 6345]='h0000068c;  wr_data_rom[ 6345]='h00000000;
    rd_cycle[ 6346] = 1'b0;  wr_cycle[ 6346] = 1'b1;  addr_rom[ 6346]='h000016c8;  wr_data_rom[ 6346]='h00000dc0;
    rd_cycle[ 6347] = 1'b1;  wr_cycle[ 6347] = 1'b0;  addr_rom[ 6347]='h00001b4c;  wr_data_rom[ 6347]='h00000000;
    rd_cycle[ 6348] = 1'b0;  wr_cycle[ 6348] = 1'b1;  addr_rom[ 6348]='h00001dfc;  wr_data_rom[ 6348]='h00000f68;
    rd_cycle[ 6349] = 1'b1;  wr_cycle[ 6349] = 1'b0;  addr_rom[ 6349]='h000013d4;  wr_data_rom[ 6349]='h00000000;
    rd_cycle[ 6350] = 1'b0;  wr_cycle[ 6350] = 1'b1;  addr_rom[ 6350]='h000019d8;  wr_data_rom[ 6350]='h000015b2;
    rd_cycle[ 6351] = 1'b0;  wr_cycle[ 6351] = 1'b1;  addr_rom[ 6351]='h00000c48;  wr_data_rom[ 6351]='h00000553;
    rd_cycle[ 6352] = 1'b0;  wr_cycle[ 6352] = 1'b1;  addr_rom[ 6352]='h00001430;  wr_data_rom[ 6352]='h00001b32;
    rd_cycle[ 6353] = 1'b1;  wr_cycle[ 6353] = 1'b0;  addr_rom[ 6353]='h000009a8;  wr_data_rom[ 6353]='h00000000;
    rd_cycle[ 6354] = 1'b0;  wr_cycle[ 6354] = 1'b1;  addr_rom[ 6354]='h00001140;  wr_data_rom[ 6354]='h00001a85;
    rd_cycle[ 6355] = 1'b0;  wr_cycle[ 6355] = 1'b1;  addr_rom[ 6355]='h00000044;  wr_data_rom[ 6355]='h00001570;
    rd_cycle[ 6356] = 1'b1;  wr_cycle[ 6356] = 1'b0;  addr_rom[ 6356]='h00000704;  wr_data_rom[ 6356]='h00000000;
    rd_cycle[ 6357] = 1'b0;  wr_cycle[ 6357] = 1'b1;  addr_rom[ 6357]='h000011cc;  wr_data_rom[ 6357]='h00001b9a;
    rd_cycle[ 6358] = 1'b0;  wr_cycle[ 6358] = 1'b1;  addr_rom[ 6358]='h00001268;  wr_data_rom[ 6358]='h00000449;
    rd_cycle[ 6359] = 1'b1;  wr_cycle[ 6359] = 1'b0;  addr_rom[ 6359]='h00000a78;  wr_data_rom[ 6359]='h00000000;
    rd_cycle[ 6360] = 1'b1;  wr_cycle[ 6360] = 1'b0;  addr_rom[ 6360]='h00000ab4;  wr_data_rom[ 6360]='h00000000;
    rd_cycle[ 6361] = 1'b1;  wr_cycle[ 6361] = 1'b0;  addr_rom[ 6361]='h000018cc;  wr_data_rom[ 6361]='h00000000;
    rd_cycle[ 6362] = 1'b1;  wr_cycle[ 6362] = 1'b0;  addr_rom[ 6362]='h000013a8;  wr_data_rom[ 6362]='h00000000;
    rd_cycle[ 6363] = 1'b0;  wr_cycle[ 6363] = 1'b1;  addr_rom[ 6363]='h00000df8;  wr_data_rom[ 6363]='h00000c62;
    rd_cycle[ 6364] = 1'b1;  wr_cycle[ 6364] = 1'b0;  addr_rom[ 6364]='h000013e0;  wr_data_rom[ 6364]='h00000000;
    rd_cycle[ 6365] = 1'b1;  wr_cycle[ 6365] = 1'b0;  addr_rom[ 6365]='h00000c20;  wr_data_rom[ 6365]='h00000000;
    rd_cycle[ 6366] = 1'b1;  wr_cycle[ 6366] = 1'b0;  addr_rom[ 6366]='h00001ad0;  wr_data_rom[ 6366]='h00000000;
    rd_cycle[ 6367] = 1'b1;  wr_cycle[ 6367] = 1'b0;  addr_rom[ 6367]='h000003c0;  wr_data_rom[ 6367]='h00000000;
    rd_cycle[ 6368] = 1'b1;  wr_cycle[ 6368] = 1'b0;  addr_rom[ 6368]='h00000064;  wr_data_rom[ 6368]='h00000000;
    rd_cycle[ 6369] = 1'b1;  wr_cycle[ 6369] = 1'b0;  addr_rom[ 6369]='h00000154;  wr_data_rom[ 6369]='h00000000;
    rd_cycle[ 6370] = 1'b0;  wr_cycle[ 6370] = 1'b1;  addr_rom[ 6370]='h00000580;  wr_data_rom[ 6370]='h00000246;
    rd_cycle[ 6371] = 1'b0;  wr_cycle[ 6371] = 1'b1;  addr_rom[ 6371]='h0000129c;  wr_data_rom[ 6371]='h000015f2;
    rd_cycle[ 6372] = 1'b0;  wr_cycle[ 6372] = 1'b1;  addr_rom[ 6372]='h00000e0c;  wr_data_rom[ 6372]='h00000385;
    rd_cycle[ 6373] = 1'b1;  wr_cycle[ 6373] = 1'b0;  addr_rom[ 6373]='h00001dec;  wr_data_rom[ 6373]='h00000000;
    rd_cycle[ 6374] = 1'b1;  wr_cycle[ 6374] = 1'b0;  addr_rom[ 6374]='h000001d0;  wr_data_rom[ 6374]='h00000000;
    rd_cycle[ 6375] = 1'b0;  wr_cycle[ 6375] = 1'b1;  addr_rom[ 6375]='h000003a4;  wr_data_rom[ 6375]='h00001a43;
    rd_cycle[ 6376] = 1'b1;  wr_cycle[ 6376] = 1'b0;  addr_rom[ 6376]='h00001018;  wr_data_rom[ 6376]='h00000000;
    rd_cycle[ 6377] = 1'b0;  wr_cycle[ 6377] = 1'b1;  addr_rom[ 6377]='h00001220;  wr_data_rom[ 6377]='h000016de;
    rd_cycle[ 6378] = 1'b0;  wr_cycle[ 6378] = 1'b1;  addr_rom[ 6378]='h00000004;  wr_data_rom[ 6378]='h0000036c;
    rd_cycle[ 6379] = 1'b1;  wr_cycle[ 6379] = 1'b0;  addr_rom[ 6379]='h0000123c;  wr_data_rom[ 6379]='h00000000;
    rd_cycle[ 6380] = 1'b0;  wr_cycle[ 6380] = 1'b1;  addr_rom[ 6380]='h00001e74;  wr_data_rom[ 6380]='h000016a6;
    rd_cycle[ 6381] = 1'b1;  wr_cycle[ 6381] = 1'b0;  addr_rom[ 6381]='h000014f0;  wr_data_rom[ 6381]='h00000000;
    rd_cycle[ 6382] = 1'b1;  wr_cycle[ 6382] = 1'b0;  addr_rom[ 6382]='h000003bc;  wr_data_rom[ 6382]='h00000000;
    rd_cycle[ 6383] = 1'b0;  wr_cycle[ 6383] = 1'b1;  addr_rom[ 6383]='h00001c78;  wr_data_rom[ 6383]='h000001b5;
    rd_cycle[ 6384] = 1'b1;  wr_cycle[ 6384] = 1'b0;  addr_rom[ 6384]='h00001c48;  wr_data_rom[ 6384]='h00000000;
    rd_cycle[ 6385] = 1'b1;  wr_cycle[ 6385] = 1'b0;  addr_rom[ 6385]='h0000094c;  wr_data_rom[ 6385]='h00000000;
    rd_cycle[ 6386] = 1'b0;  wr_cycle[ 6386] = 1'b1;  addr_rom[ 6386]='h000019e0;  wr_data_rom[ 6386]='h0000155a;
    rd_cycle[ 6387] = 1'b1;  wr_cycle[ 6387] = 1'b0;  addr_rom[ 6387]='h00001d40;  wr_data_rom[ 6387]='h00000000;
    rd_cycle[ 6388] = 1'b1;  wr_cycle[ 6388] = 1'b0;  addr_rom[ 6388]='h000009fc;  wr_data_rom[ 6388]='h00000000;
    rd_cycle[ 6389] = 1'b0;  wr_cycle[ 6389] = 1'b1;  addr_rom[ 6389]='h00001f08;  wr_data_rom[ 6389]='h00000204;
    rd_cycle[ 6390] = 1'b1;  wr_cycle[ 6390] = 1'b0;  addr_rom[ 6390]='h00001a3c;  wr_data_rom[ 6390]='h00000000;
    rd_cycle[ 6391] = 1'b1;  wr_cycle[ 6391] = 1'b0;  addr_rom[ 6391]='h00000a50;  wr_data_rom[ 6391]='h00000000;
    rd_cycle[ 6392] = 1'b1;  wr_cycle[ 6392] = 1'b0;  addr_rom[ 6392]='h0000021c;  wr_data_rom[ 6392]='h00000000;
    rd_cycle[ 6393] = 1'b1;  wr_cycle[ 6393] = 1'b0;  addr_rom[ 6393]='h00001f0c;  wr_data_rom[ 6393]='h00000000;
    rd_cycle[ 6394] = 1'b1;  wr_cycle[ 6394] = 1'b0;  addr_rom[ 6394]='h00001a18;  wr_data_rom[ 6394]='h00000000;
    rd_cycle[ 6395] = 1'b0;  wr_cycle[ 6395] = 1'b1;  addr_rom[ 6395]='h00001010;  wr_data_rom[ 6395]='h000010f8;
    rd_cycle[ 6396] = 1'b0;  wr_cycle[ 6396] = 1'b1;  addr_rom[ 6396]='h00000240;  wr_data_rom[ 6396]='h000012ce;
    rd_cycle[ 6397] = 1'b0;  wr_cycle[ 6397] = 1'b1;  addr_rom[ 6397]='h00001980;  wr_data_rom[ 6397]='h00000470;
    rd_cycle[ 6398] = 1'b1;  wr_cycle[ 6398] = 1'b0;  addr_rom[ 6398]='h00000674;  wr_data_rom[ 6398]='h00000000;
    rd_cycle[ 6399] = 1'b0;  wr_cycle[ 6399] = 1'b1;  addr_rom[ 6399]='h00000510;  wr_data_rom[ 6399]='h00000020;
    rd_cycle[ 6400] = 1'b0;  wr_cycle[ 6400] = 1'b1;  addr_rom[ 6400]='h00000938;  wr_data_rom[ 6400]='h0000109e;
    rd_cycle[ 6401] = 1'b1;  wr_cycle[ 6401] = 1'b0;  addr_rom[ 6401]='h00000e58;  wr_data_rom[ 6401]='h00000000;
    rd_cycle[ 6402] = 1'b0;  wr_cycle[ 6402] = 1'b1;  addr_rom[ 6402]='h00000e68;  wr_data_rom[ 6402]='h00000174;
    rd_cycle[ 6403] = 1'b0;  wr_cycle[ 6403] = 1'b1;  addr_rom[ 6403]='h00001494;  wr_data_rom[ 6403]='h00001215;
    rd_cycle[ 6404] = 1'b1;  wr_cycle[ 6404] = 1'b0;  addr_rom[ 6404]='h00000ed4;  wr_data_rom[ 6404]='h00000000;
    rd_cycle[ 6405] = 1'b1;  wr_cycle[ 6405] = 1'b0;  addr_rom[ 6405]='h0000064c;  wr_data_rom[ 6405]='h00000000;
    rd_cycle[ 6406] = 1'b0;  wr_cycle[ 6406] = 1'b1;  addr_rom[ 6406]='h00000488;  wr_data_rom[ 6406]='h00000de2;
    rd_cycle[ 6407] = 1'b1;  wr_cycle[ 6407] = 1'b0;  addr_rom[ 6407]='h00001a74;  wr_data_rom[ 6407]='h00000000;
    rd_cycle[ 6408] = 1'b0;  wr_cycle[ 6408] = 1'b1;  addr_rom[ 6408]='h00001478;  wr_data_rom[ 6408]='h00001c91;
    rd_cycle[ 6409] = 1'b1;  wr_cycle[ 6409] = 1'b0;  addr_rom[ 6409]='h000001d4;  wr_data_rom[ 6409]='h00000000;
    rd_cycle[ 6410] = 1'b0;  wr_cycle[ 6410] = 1'b1;  addr_rom[ 6410]='h00000bd8;  wr_data_rom[ 6410]='h00000da3;
    rd_cycle[ 6411] = 1'b1;  wr_cycle[ 6411] = 1'b0;  addr_rom[ 6411]='h00001244;  wr_data_rom[ 6411]='h00000000;
    rd_cycle[ 6412] = 1'b1;  wr_cycle[ 6412] = 1'b0;  addr_rom[ 6412]='h00001978;  wr_data_rom[ 6412]='h00000000;
    rd_cycle[ 6413] = 1'b1;  wr_cycle[ 6413] = 1'b0;  addr_rom[ 6413]='h00000a80;  wr_data_rom[ 6413]='h00000000;
    rd_cycle[ 6414] = 1'b1;  wr_cycle[ 6414] = 1'b0;  addr_rom[ 6414]='h000017a8;  wr_data_rom[ 6414]='h00000000;
    rd_cycle[ 6415] = 1'b1;  wr_cycle[ 6415] = 1'b0;  addr_rom[ 6415]='h00001b5c;  wr_data_rom[ 6415]='h00000000;
    rd_cycle[ 6416] = 1'b1;  wr_cycle[ 6416] = 1'b0;  addr_rom[ 6416]='h000018f0;  wr_data_rom[ 6416]='h00000000;
    rd_cycle[ 6417] = 1'b0;  wr_cycle[ 6417] = 1'b1;  addr_rom[ 6417]='h00000808;  wr_data_rom[ 6417]='h000007f7;
    rd_cycle[ 6418] = 1'b1;  wr_cycle[ 6418] = 1'b0;  addr_rom[ 6418]='h00001858;  wr_data_rom[ 6418]='h00000000;
    rd_cycle[ 6419] = 1'b0;  wr_cycle[ 6419] = 1'b1;  addr_rom[ 6419]='h00001bf0;  wr_data_rom[ 6419]='h000012bc;
    rd_cycle[ 6420] = 1'b0;  wr_cycle[ 6420] = 1'b1;  addr_rom[ 6420]='h00000944;  wr_data_rom[ 6420]='h0000005c;
    rd_cycle[ 6421] = 1'b0;  wr_cycle[ 6421] = 1'b1;  addr_rom[ 6421]='h00000630;  wr_data_rom[ 6421]='h00001861;
    rd_cycle[ 6422] = 1'b0;  wr_cycle[ 6422] = 1'b1;  addr_rom[ 6422]='h00001238;  wr_data_rom[ 6422]='h000018a2;
    rd_cycle[ 6423] = 1'b0;  wr_cycle[ 6423] = 1'b1;  addr_rom[ 6423]='h000016d0;  wr_data_rom[ 6423]='h00001673;
    rd_cycle[ 6424] = 1'b1;  wr_cycle[ 6424] = 1'b0;  addr_rom[ 6424]='h00001404;  wr_data_rom[ 6424]='h00000000;
    rd_cycle[ 6425] = 1'b1;  wr_cycle[ 6425] = 1'b0;  addr_rom[ 6425]='h00001dcc;  wr_data_rom[ 6425]='h00000000;
    rd_cycle[ 6426] = 1'b1;  wr_cycle[ 6426] = 1'b0;  addr_rom[ 6426]='h00001840;  wr_data_rom[ 6426]='h00000000;
    rd_cycle[ 6427] = 1'b0;  wr_cycle[ 6427] = 1'b1;  addr_rom[ 6427]='h00001a44;  wr_data_rom[ 6427]='h00000a54;
    rd_cycle[ 6428] = 1'b0;  wr_cycle[ 6428] = 1'b1;  addr_rom[ 6428]='h00000f28;  wr_data_rom[ 6428]='h00001460;
    rd_cycle[ 6429] = 1'b0;  wr_cycle[ 6429] = 1'b1;  addr_rom[ 6429]='h000000cc;  wr_data_rom[ 6429]='h000010b6;
    rd_cycle[ 6430] = 1'b0;  wr_cycle[ 6430] = 1'b1;  addr_rom[ 6430]='h00000288;  wr_data_rom[ 6430]='h000000ff;
    rd_cycle[ 6431] = 1'b1;  wr_cycle[ 6431] = 1'b0;  addr_rom[ 6431]='h00000768;  wr_data_rom[ 6431]='h00000000;
    rd_cycle[ 6432] = 1'b0;  wr_cycle[ 6432] = 1'b1;  addr_rom[ 6432]='h00001e0c;  wr_data_rom[ 6432]='h00001b54;
    rd_cycle[ 6433] = 1'b1;  wr_cycle[ 6433] = 1'b0;  addr_rom[ 6433]='h000007c8;  wr_data_rom[ 6433]='h00000000;
    rd_cycle[ 6434] = 1'b1;  wr_cycle[ 6434] = 1'b0;  addr_rom[ 6434]='h00000a98;  wr_data_rom[ 6434]='h00000000;
    rd_cycle[ 6435] = 1'b0;  wr_cycle[ 6435] = 1'b1;  addr_rom[ 6435]='h00000254;  wr_data_rom[ 6435]='h00000c37;
    rd_cycle[ 6436] = 1'b1;  wr_cycle[ 6436] = 1'b0;  addr_rom[ 6436]='h000007fc;  wr_data_rom[ 6436]='h00000000;
    rd_cycle[ 6437] = 1'b0;  wr_cycle[ 6437] = 1'b1;  addr_rom[ 6437]='h000003d8;  wr_data_rom[ 6437]='h00000e78;
    rd_cycle[ 6438] = 1'b0;  wr_cycle[ 6438] = 1'b1;  addr_rom[ 6438]='h00001960;  wr_data_rom[ 6438]='h0000068f;
    rd_cycle[ 6439] = 1'b0;  wr_cycle[ 6439] = 1'b1;  addr_rom[ 6439]='h000012ac;  wr_data_rom[ 6439]='h0000156e;
    rd_cycle[ 6440] = 1'b0;  wr_cycle[ 6440] = 1'b1;  addr_rom[ 6440]='h00001f14;  wr_data_rom[ 6440]='h00000523;
    rd_cycle[ 6441] = 1'b1;  wr_cycle[ 6441] = 1'b0;  addr_rom[ 6441]='h000005bc;  wr_data_rom[ 6441]='h00000000;
    rd_cycle[ 6442] = 1'b0;  wr_cycle[ 6442] = 1'b1;  addr_rom[ 6442]='h00001468;  wr_data_rom[ 6442]='h00000a01;
    rd_cycle[ 6443] = 1'b0;  wr_cycle[ 6443] = 1'b1;  addr_rom[ 6443]='h00001904;  wr_data_rom[ 6443]='h00001bbd;
    rd_cycle[ 6444] = 1'b0;  wr_cycle[ 6444] = 1'b1;  addr_rom[ 6444]='h000008b0;  wr_data_rom[ 6444]='h00001463;
    rd_cycle[ 6445] = 1'b0;  wr_cycle[ 6445] = 1'b1;  addr_rom[ 6445]='h00000a28;  wr_data_rom[ 6445]='h000014d8;
    rd_cycle[ 6446] = 1'b1;  wr_cycle[ 6446] = 1'b0;  addr_rom[ 6446]='h000016fc;  wr_data_rom[ 6446]='h00000000;
    rd_cycle[ 6447] = 1'b1;  wr_cycle[ 6447] = 1'b0;  addr_rom[ 6447]='h00000404;  wr_data_rom[ 6447]='h00000000;
    rd_cycle[ 6448] = 1'b1;  wr_cycle[ 6448] = 1'b0;  addr_rom[ 6448]='h00000b44;  wr_data_rom[ 6448]='h00000000;
    rd_cycle[ 6449] = 1'b1;  wr_cycle[ 6449] = 1'b0;  addr_rom[ 6449]='h00001650;  wr_data_rom[ 6449]='h00000000;
    rd_cycle[ 6450] = 1'b1;  wr_cycle[ 6450] = 1'b0;  addr_rom[ 6450]='h0000016c;  wr_data_rom[ 6450]='h00000000;
    rd_cycle[ 6451] = 1'b1;  wr_cycle[ 6451] = 1'b0;  addr_rom[ 6451]='h000005fc;  wr_data_rom[ 6451]='h00000000;
    rd_cycle[ 6452] = 1'b0;  wr_cycle[ 6452] = 1'b1;  addr_rom[ 6452]='h000014a8;  wr_data_rom[ 6452]='h00001b89;
    rd_cycle[ 6453] = 1'b1;  wr_cycle[ 6453] = 1'b0;  addr_rom[ 6453]='h00000890;  wr_data_rom[ 6453]='h00000000;
    rd_cycle[ 6454] = 1'b0;  wr_cycle[ 6454] = 1'b1;  addr_rom[ 6454]='h000001a8;  wr_data_rom[ 6454]='h000017e0;
    rd_cycle[ 6455] = 1'b0;  wr_cycle[ 6455] = 1'b1;  addr_rom[ 6455]='h00001f28;  wr_data_rom[ 6455]='h00001810;
    rd_cycle[ 6456] = 1'b1;  wr_cycle[ 6456] = 1'b0;  addr_rom[ 6456]='h000016ec;  wr_data_rom[ 6456]='h00000000;
    rd_cycle[ 6457] = 1'b1;  wr_cycle[ 6457] = 1'b0;  addr_rom[ 6457]='h00001580;  wr_data_rom[ 6457]='h00000000;
    rd_cycle[ 6458] = 1'b0;  wr_cycle[ 6458] = 1'b1;  addr_rom[ 6458]='h00001998;  wr_data_rom[ 6458]='h00000ca3;
    rd_cycle[ 6459] = 1'b0;  wr_cycle[ 6459] = 1'b1;  addr_rom[ 6459]='h00001290;  wr_data_rom[ 6459]='h00000864;
    rd_cycle[ 6460] = 1'b1;  wr_cycle[ 6460] = 1'b0;  addr_rom[ 6460]='h00000e80;  wr_data_rom[ 6460]='h00000000;
    rd_cycle[ 6461] = 1'b0;  wr_cycle[ 6461] = 1'b1;  addr_rom[ 6461]='h000015b8;  wr_data_rom[ 6461]='h000008f3;
    rd_cycle[ 6462] = 1'b0;  wr_cycle[ 6462] = 1'b1;  addr_rom[ 6462]='h000019e0;  wr_data_rom[ 6462]='h0000096e;
    rd_cycle[ 6463] = 1'b1;  wr_cycle[ 6463] = 1'b0;  addr_rom[ 6463]='h000002ec;  wr_data_rom[ 6463]='h00000000;
    rd_cycle[ 6464] = 1'b1;  wr_cycle[ 6464] = 1'b0;  addr_rom[ 6464]='h0000156c;  wr_data_rom[ 6464]='h00000000;
    rd_cycle[ 6465] = 1'b0;  wr_cycle[ 6465] = 1'b1;  addr_rom[ 6465]='h00000004;  wr_data_rom[ 6465]='h0000161a;
    rd_cycle[ 6466] = 1'b0;  wr_cycle[ 6466] = 1'b1;  addr_rom[ 6466]='h0000139c;  wr_data_rom[ 6466]='h0000066d;
    rd_cycle[ 6467] = 1'b0;  wr_cycle[ 6467] = 1'b1;  addr_rom[ 6467]='h00000cb0;  wr_data_rom[ 6467]='h00001d92;
    rd_cycle[ 6468] = 1'b0;  wr_cycle[ 6468] = 1'b1;  addr_rom[ 6468]='h00001858;  wr_data_rom[ 6468]='h00001072;
    rd_cycle[ 6469] = 1'b0;  wr_cycle[ 6469] = 1'b1;  addr_rom[ 6469]='h00001708;  wr_data_rom[ 6469]='h00000a8d;
    rd_cycle[ 6470] = 1'b0;  wr_cycle[ 6470] = 1'b1;  addr_rom[ 6470]='h00000c24;  wr_data_rom[ 6470]='h000004b4;
    rd_cycle[ 6471] = 1'b1;  wr_cycle[ 6471] = 1'b0;  addr_rom[ 6471]='h00001be0;  wr_data_rom[ 6471]='h00000000;
    rd_cycle[ 6472] = 1'b0;  wr_cycle[ 6472] = 1'b1;  addr_rom[ 6472]='h00001858;  wr_data_rom[ 6472]='h00000ec7;
    rd_cycle[ 6473] = 1'b1;  wr_cycle[ 6473] = 1'b0;  addr_rom[ 6473]='h0000015c;  wr_data_rom[ 6473]='h00000000;
    rd_cycle[ 6474] = 1'b0;  wr_cycle[ 6474] = 1'b1;  addr_rom[ 6474]='h00001d78;  wr_data_rom[ 6474]='h00000fa7;
    rd_cycle[ 6475] = 1'b1;  wr_cycle[ 6475] = 1'b0;  addr_rom[ 6475]='h00001a44;  wr_data_rom[ 6475]='h00000000;
    rd_cycle[ 6476] = 1'b1;  wr_cycle[ 6476] = 1'b0;  addr_rom[ 6476]='h000016b8;  wr_data_rom[ 6476]='h00000000;
    rd_cycle[ 6477] = 1'b1;  wr_cycle[ 6477] = 1'b0;  addr_rom[ 6477]='h00001004;  wr_data_rom[ 6477]='h00000000;
    rd_cycle[ 6478] = 1'b0;  wr_cycle[ 6478] = 1'b1;  addr_rom[ 6478]='h000017d8;  wr_data_rom[ 6478]='h000011b0;
    rd_cycle[ 6479] = 1'b1;  wr_cycle[ 6479] = 1'b0;  addr_rom[ 6479]='h00000108;  wr_data_rom[ 6479]='h00000000;
    rd_cycle[ 6480] = 1'b0;  wr_cycle[ 6480] = 1'b1;  addr_rom[ 6480]='h00001a94;  wr_data_rom[ 6480]='h00001933;
    rd_cycle[ 6481] = 1'b0;  wr_cycle[ 6481] = 1'b1;  addr_rom[ 6481]='h0000114c;  wr_data_rom[ 6481]='h000004ee;
    rd_cycle[ 6482] = 1'b1;  wr_cycle[ 6482] = 1'b0;  addr_rom[ 6482]='h00001d70;  wr_data_rom[ 6482]='h00000000;
    rd_cycle[ 6483] = 1'b1;  wr_cycle[ 6483] = 1'b0;  addr_rom[ 6483]='h00001d90;  wr_data_rom[ 6483]='h00000000;
    rd_cycle[ 6484] = 1'b0;  wr_cycle[ 6484] = 1'b1;  addr_rom[ 6484]='h00001814;  wr_data_rom[ 6484]='h00000196;
    rd_cycle[ 6485] = 1'b1;  wr_cycle[ 6485] = 1'b0;  addr_rom[ 6485]='h0000164c;  wr_data_rom[ 6485]='h00000000;
    rd_cycle[ 6486] = 1'b0;  wr_cycle[ 6486] = 1'b1;  addr_rom[ 6486]='h0000137c;  wr_data_rom[ 6486]='h0000117d;
    rd_cycle[ 6487] = 1'b0;  wr_cycle[ 6487] = 1'b1;  addr_rom[ 6487]='h0000087c;  wr_data_rom[ 6487]='h000001cf;
    rd_cycle[ 6488] = 1'b1;  wr_cycle[ 6488] = 1'b0;  addr_rom[ 6488]='h00001e3c;  wr_data_rom[ 6488]='h00000000;
    rd_cycle[ 6489] = 1'b1;  wr_cycle[ 6489] = 1'b0;  addr_rom[ 6489]='h000002f4;  wr_data_rom[ 6489]='h00000000;
    rd_cycle[ 6490] = 1'b1;  wr_cycle[ 6490] = 1'b0;  addr_rom[ 6490]='h0000180c;  wr_data_rom[ 6490]='h00000000;
    rd_cycle[ 6491] = 1'b1;  wr_cycle[ 6491] = 1'b0;  addr_rom[ 6491]='h00001084;  wr_data_rom[ 6491]='h00000000;
    rd_cycle[ 6492] = 1'b0;  wr_cycle[ 6492] = 1'b1;  addr_rom[ 6492]='h000008f8;  wr_data_rom[ 6492]='h000018fc;
    rd_cycle[ 6493] = 1'b0;  wr_cycle[ 6493] = 1'b1;  addr_rom[ 6493]='h000011b8;  wr_data_rom[ 6493]='h00000e52;
    rd_cycle[ 6494] = 1'b0;  wr_cycle[ 6494] = 1'b1;  addr_rom[ 6494]='h00000bfc;  wr_data_rom[ 6494]='h00000634;
    rd_cycle[ 6495] = 1'b0;  wr_cycle[ 6495] = 1'b1;  addr_rom[ 6495]='h00000250;  wr_data_rom[ 6495]='h00000bc1;
    rd_cycle[ 6496] = 1'b1;  wr_cycle[ 6496] = 1'b0;  addr_rom[ 6496]='h00000d2c;  wr_data_rom[ 6496]='h00000000;
    rd_cycle[ 6497] = 1'b0;  wr_cycle[ 6497] = 1'b1;  addr_rom[ 6497]='h00000fc8;  wr_data_rom[ 6497]='h00001f3a;
    rd_cycle[ 6498] = 1'b0;  wr_cycle[ 6498] = 1'b1;  addr_rom[ 6498]='h00000ce8;  wr_data_rom[ 6498]='h00001c5f;
    rd_cycle[ 6499] = 1'b1;  wr_cycle[ 6499] = 1'b0;  addr_rom[ 6499]='h00001bc8;  wr_data_rom[ 6499]='h00000000;
    rd_cycle[ 6500] = 1'b1;  wr_cycle[ 6500] = 1'b0;  addr_rom[ 6500]='h000016c0;  wr_data_rom[ 6500]='h00000000;
    rd_cycle[ 6501] = 1'b0;  wr_cycle[ 6501] = 1'b1;  addr_rom[ 6501]='h000003dc;  wr_data_rom[ 6501]='h00000304;
    rd_cycle[ 6502] = 1'b1;  wr_cycle[ 6502] = 1'b0;  addr_rom[ 6502]='h000003a0;  wr_data_rom[ 6502]='h00000000;
    rd_cycle[ 6503] = 1'b1;  wr_cycle[ 6503] = 1'b0;  addr_rom[ 6503]='h00001684;  wr_data_rom[ 6503]='h00000000;
    rd_cycle[ 6504] = 1'b0;  wr_cycle[ 6504] = 1'b1;  addr_rom[ 6504]='h0000011c;  wr_data_rom[ 6504]='h00001126;
    rd_cycle[ 6505] = 1'b1;  wr_cycle[ 6505] = 1'b0;  addr_rom[ 6505]='h000014fc;  wr_data_rom[ 6505]='h00000000;
    rd_cycle[ 6506] = 1'b1;  wr_cycle[ 6506] = 1'b0;  addr_rom[ 6506]='h00001a60;  wr_data_rom[ 6506]='h00000000;
    rd_cycle[ 6507] = 1'b1;  wr_cycle[ 6507] = 1'b0;  addr_rom[ 6507]='h00000754;  wr_data_rom[ 6507]='h00000000;
    rd_cycle[ 6508] = 1'b0;  wr_cycle[ 6508] = 1'b1;  addr_rom[ 6508]='h0000153c;  wr_data_rom[ 6508]='h0000038d;
    rd_cycle[ 6509] = 1'b0;  wr_cycle[ 6509] = 1'b1;  addr_rom[ 6509]='h000006ac;  wr_data_rom[ 6509]='h000013fe;
    rd_cycle[ 6510] = 1'b0;  wr_cycle[ 6510] = 1'b1;  addr_rom[ 6510]='h000008ac;  wr_data_rom[ 6510]='h00001a47;
    rd_cycle[ 6511] = 1'b0;  wr_cycle[ 6511] = 1'b1;  addr_rom[ 6511]='h00000760;  wr_data_rom[ 6511]='h000007ef;
    rd_cycle[ 6512] = 1'b0;  wr_cycle[ 6512] = 1'b1;  addr_rom[ 6512]='h00000a6c;  wr_data_rom[ 6512]='h00001758;
    rd_cycle[ 6513] = 1'b1;  wr_cycle[ 6513] = 1'b0;  addr_rom[ 6513]='h00001868;  wr_data_rom[ 6513]='h00000000;
    rd_cycle[ 6514] = 1'b0;  wr_cycle[ 6514] = 1'b1;  addr_rom[ 6514]='h00001048;  wr_data_rom[ 6514]='h00000258;
    rd_cycle[ 6515] = 1'b0;  wr_cycle[ 6515] = 1'b1;  addr_rom[ 6515]='h0000172c;  wr_data_rom[ 6515]='h00000ac8;
    rd_cycle[ 6516] = 1'b0;  wr_cycle[ 6516] = 1'b1;  addr_rom[ 6516]='h00001f08;  wr_data_rom[ 6516]='h0000008d;
    rd_cycle[ 6517] = 1'b1;  wr_cycle[ 6517] = 1'b0;  addr_rom[ 6517]='h00001b20;  wr_data_rom[ 6517]='h00000000;
    rd_cycle[ 6518] = 1'b1;  wr_cycle[ 6518] = 1'b0;  addr_rom[ 6518]='h0000033c;  wr_data_rom[ 6518]='h00000000;
    rd_cycle[ 6519] = 1'b1;  wr_cycle[ 6519] = 1'b0;  addr_rom[ 6519]='h00001b38;  wr_data_rom[ 6519]='h00000000;
    rd_cycle[ 6520] = 1'b1;  wr_cycle[ 6520] = 1'b0;  addr_rom[ 6520]='h00001b00;  wr_data_rom[ 6520]='h00000000;
    rd_cycle[ 6521] = 1'b0;  wr_cycle[ 6521] = 1'b1;  addr_rom[ 6521]='h00000c14;  wr_data_rom[ 6521]='h0000044c;
    rd_cycle[ 6522] = 1'b0;  wr_cycle[ 6522] = 1'b1;  addr_rom[ 6522]='h00000f3c;  wr_data_rom[ 6522]='h00000923;
    rd_cycle[ 6523] = 1'b0;  wr_cycle[ 6523] = 1'b1;  addr_rom[ 6523]='h0000110c;  wr_data_rom[ 6523]='h00000bd2;
    rd_cycle[ 6524] = 1'b1;  wr_cycle[ 6524] = 1'b0;  addr_rom[ 6524]='h00000d40;  wr_data_rom[ 6524]='h00000000;
    rd_cycle[ 6525] = 1'b1;  wr_cycle[ 6525] = 1'b0;  addr_rom[ 6525]='h00001234;  wr_data_rom[ 6525]='h00000000;
    rd_cycle[ 6526] = 1'b0;  wr_cycle[ 6526] = 1'b1;  addr_rom[ 6526]='h00000460;  wr_data_rom[ 6526]='h0000136d;
    rd_cycle[ 6527] = 1'b1;  wr_cycle[ 6527] = 1'b0;  addr_rom[ 6527]='h000004cc;  wr_data_rom[ 6527]='h00000000;
    rd_cycle[ 6528] = 1'b1;  wr_cycle[ 6528] = 1'b0;  addr_rom[ 6528]='h00001434;  wr_data_rom[ 6528]='h00000000;
    rd_cycle[ 6529] = 1'b1;  wr_cycle[ 6529] = 1'b0;  addr_rom[ 6529]='h0000060c;  wr_data_rom[ 6529]='h00000000;
    rd_cycle[ 6530] = 1'b1;  wr_cycle[ 6530] = 1'b0;  addr_rom[ 6530]='h00001144;  wr_data_rom[ 6530]='h00000000;
    rd_cycle[ 6531] = 1'b1;  wr_cycle[ 6531] = 1'b0;  addr_rom[ 6531]='h00000cd0;  wr_data_rom[ 6531]='h00000000;
    rd_cycle[ 6532] = 1'b1;  wr_cycle[ 6532] = 1'b0;  addr_rom[ 6532]='h00001d50;  wr_data_rom[ 6532]='h00000000;
    rd_cycle[ 6533] = 1'b0;  wr_cycle[ 6533] = 1'b1;  addr_rom[ 6533]='h00001c78;  wr_data_rom[ 6533]='h00000bd2;
    rd_cycle[ 6534] = 1'b1;  wr_cycle[ 6534] = 1'b0;  addr_rom[ 6534]='h000012c0;  wr_data_rom[ 6534]='h00000000;
    rd_cycle[ 6535] = 1'b0;  wr_cycle[ 6535] = 1'b1;  addr_rom[ 6535]='h00000404;  wr_data_rom[ 6535]='h00001c2a;
    rd_cycle[ 6536] = 1'b1;  wr_cycle[ 6536] = 1'b0;  addr_rom[ 6536]='h00001490;  wr_data_rom[ 6536]='h00000000;
    rd_cycle[ 6537] = 1'b0;  wr_cycle[ 6537] = 1'b1;  addr_rom[ 6537]='h00000204;  wr_data_rom[ 6537]='h000004a1;
    rd_cycle[ 6538] = 1'b1;  wr_cycle[ 6538] = 1'b0;  addr_rom[ 6538]='h000008c4;  wr_data_rom[ 6538]='h00000000;
    rd_cycle[ 6539] = 1'b0;  wr_cycle[ 6539] = 1'b1;  addr_rom[ 6539]='h00000b18;  wr_data_rom[ 6539]='h00000805;
    rd_cycle[ 6540] = 1'b1;  wr_cycle[ 6540] = 1'b0;  addr_rom[ 6540]='h00000e20;  wr_data_rom[ 6540]='h00000000;
    rd_cycle[ 6541] = 1'b1;  wr_cycle[ 6541] = 1'b0;  addr_rom[ 6541]='h00001404;  wr_data_rom[ 6541]='h00000000;
    rd_cycle[ 6542] = 1'b0;  wr_cycle[ 6542] = 1'b1;  addr_rom[ 6542]='h00001640;  wr_data_rom[ 6542]='h00001e30;
    rd_cycle[ 6543] = 1'b0;  wr_cycle[ 6543] = 1'b1;  addr_rom[ 6543]='h00001a50;  wr_data_rom[ 6543]='h0000137d;
    rd_cycle[ 6544] = 1'b1;  wr_cycle[ 6544] = 1'b0;  addr_rom[ 6544]='h000014e8;  wr_data_rom[ 6544]='h00000000;
    rd_cycle[ 6545] = 1'b1;  wr_cycle[ 6545] = 1'b0;  addr_rom[ 6545]='h00001e88;  wr_data_rom[ 6545]='h00000000;
    rd_cycle[ 6546] = 1'b1;  wr_cycle[ 6546] = 1'b0;  addr_rom[ 6546]='h00001450;  wr_data_rom[ 6546]='h00000000;
    rd_cycle[ 6547] = 1'b1;  wr_cycle[ 6547] = 1'b0;  addr_rom[ 6547]='h00000994;  wr_data_rom[ 6547]='h00000000;
    rd_cycle[ 6548] = 1'b1;  wr_cycle[ 6548] = 1'b0;  addr_rom[ 6548]='h00000d68;  wr_data_rom[ 6548]='h00000000;
    rd_cycle[ 6549] = 1'b0;  wr_cycle[ 6549] = 1'b1;  addr_rom[ 6549]='h000001ec;  wr_data_rom[ 6549]='h0000180b;
    rd_cycle[ 6550] = 1'b1;  wr_cycle[ 6550] = 1'b0;  addr_rom[ 6550]='h00000a98;  wr_data_rom[ 6550]='h00000000;
    rd_cycle[ 6551] = 1'b0;  wr_cycle[ 6551] = 1'b1;  addr_rom[ 6551]='h00001a50;  wr_data_rom[ 6551]='h0000176a;
    rd_cycle[ 6552] = 1'b1;  wr_cycle[ 6552] = 1'b0;  addr_rom[ 6552]='h0000035c;  wr_data_rom[ 6552]='h00000000;
    rd_cycle[ 6553] = 1'b1;  wr_cycle[ 6553] = 1'b0;  addr_rom[ 6553]='h000001ec;  wr_data_rom[ 6553]='h00000000;
    rd_cycle[ 6554] = 1'b1;  wr_cycle[ 6554] = 1'b0;  addr_rom[ 6554]='h00000090;  wr_data_rom[ 6554]='h00000000;
    rd_cycle[ 6555] = 1'b1;  wr_cycle[ 6555] = 1'b0;  addr_rom[ 6555]='h000019ac;  wr_data_rom[ 6555]='h00000000;
    rd_cycle[ 6556] = 1'b1;  wr_cycle[ 6556] = 1'b0;  addr_rom[ 6556]='h00000758;  wr_data_rom[ 6556]='h00000000;
    rd_cycle[ 6557] = 1'b0;  wr_cycle[ 6557] = 1'b1;  addr_rom[ 6557]='h000013b8;  wr_data_rom[ 6557]='h00000f47;
    rd_cycle[ 6558] = 1'b0;  wr_cycle[ 6558] = 1'b1;  addr_rom[ 6558]='h00000d64;  wr_data_rom[ 6558]='h00001392;
    rd_cycle[ 6559] = 1'b1;  wr_cycle[ 6559] = 1'b0;  addr_rom[ 6559]='h00001908;  wr_data_rom[ 6559]='h00000000;
    rd_cycle[ 6560] = 1'b1;  wr_cycle[ 6560] = 1'b0;  addr_rom[ 6560]='h00001554;  wr_data_rom[ 6560]='h00000000;
    rd_cycle[ 6561] = 1'b1;  wr_cycle[ 6561] = 1'b0;  addr_rom[ 6561]='h00001784;  wr_data_rom[ 6561]='h00000000;
    rd_cycle[ 6562] = 1'b1;  wr_cycle[ 6562] = 1'b0;  addr_rom[ 6562]='h00000ad4;  wr_data_rom[ 6562]='h00000000;
    rd_cycle[ 6563] = 1'b1;  wr_cycle[ 6563] = 1'b0;  addr_rom[ 6563]='h00001394;  wr_data_rom[ 6563]='h00000000;
    rd_cycle[ 6564] = 1'b1;  wr_cycle[ 6564] = 1'b0;  addr_rom[ 6564]='h00001df0;  wr_data_rom[ 6564]='h00000000;
    rd_cycle[ 6565] = 1'b0;  wr_cycle[ 6565] = 1'b1;  addr_rom[ 6565]='h00000388;  wr_data_rom[ 6565]='h000013c7;
    rd_cycle[ 6566] = 1'b0;  wr_cycle[ 6566] = 1'b1;  addr_rom[ 6566]='h00000cd8;  wr_data_rom[ 6566]='h00000b14;
    rd_cycle[ 6567] = 1'b0;  wr_cycle[ 6567] = 1'b1;  addr_rom[ 6567]='h00001864;  wr_data_rom[ 6567]='h0000142a;
    rd_cycle[ 6568] = 1'b1;  wr_cycle[ 6568] = 1'b0;  addr_rom[ 6568]='h00001388;  wr_data_rom[ 6568]='h00000000;
    rd_cycle[ 6569] = 1'b1;  wr_cycle[ 6569] = 1'b0;  addr_rom[ 6569]='h0000071c;  wr_data_rom[ 6569]='h00000000;
    rd_cycle[ 6570] = 1'b1;  wr_cycle[ 6570] = 1'b0;  addr_rom[ 6570]='h00000594;  wr_data_rom[ 6570]='h00000000;
    rd_cycle[ 6571] = 1'b0;  wr_cycle[ 6571] = 1'b1;  addr_rom[ 6571]='h00000b70;  wr_data_rom[ 6571]='h00000b59;
    rd_cycle[ 6572] = 1'b1;  wr_cycle[ 6572] = 1'b0;  addr_rom[ 6572]='h00001220;  wr_data_rom[ 6572]='h00000000;
    rd_cycle[ 6573] = 1'b1;  wr_cycle[ 6573] = 1'b0;  addr_rom[ 6573]='h000010a4;  wr_data_rom[ 6573]='h00000000;
    rd_cycle[ 6574] = 1'b0;  wr_cycle[ 6574] = 1'b1;  addr_rom[ 6574]='h00001628;  wr_data_rom[ 6574]='h00001117;
    rd_cycle[ 6575] = 1'b0;  wr_cycle[ 6575] = 1'b1;  addr_rom[ 6575]='h00000614;  wr_data_rom[ 6575]='h00001c8b;
    rd_cycle[ 6576] = 1'b1;  wr_cycle[ 6576] = 1'b0;  addr_rom[ 6576]='h00000a68;  wr_data_rom[ 6576]='h00000000;
    rd_cycle[ 6577] = 1'b0;  wr_cycle[ 6577] = 1'b1;  addr_rom[ 6577]='h00001ee8;  wr_data_rom[ 6577]='h0000157a;
    rd_cycle[ 6578] = 1'b1;  wr_cycle[ 6578] = 1'b0;  addr_rom[ 6578]='h00000120;  wr_data_rom[ 6578]='h00000000;
    rd_cycle[ 6579] = 1'b0;  wr_cycle[ 6579] = 1'b1;  addr_rom[ 6579]='h00001188;  wr_data_rom[ 6579]='h0000076b;
    rd_cycle[ 6580] = 1'b1;  wr_cycle[ 6580] = 1'b0;  addr_rom[ 6580]='h00000204;  wr_data_rom[ 6580]='h00000000;
    rd_cycle[ 6581] = 1'b0;  wr_cycle[ 6581] = 1'b1;  addr_rom[ 6581]='h00001770;  wr_data_rom[ 6581]='h00000d38;
    rd_cycle[ 6582] = 1'b1;  wr_cycle[ 6582] = 1'b0;  addr_rom[ 6582]='h00000f84;  wr_data_rom[ 6582]='h00000000;
    rd_cycle[ 6583] = 1'b0;  wr_cycle[ 6583] = 1'b1;  addr_rom[ 6583]='h00001414;  wr_data_rom[ 6583]='h00000c4a;
    rd_cycle[ 6584] = 1'b1;  wr_cycle[ 6584] = 1'b0;  addr_rom[ 6584]='h00001ab8;  wr_data_rom[ 6584]='h00000000;
    rd_cycle[ 6585] = 1'b1;  wr_cycle[ 6585] = 1'b0;  addr_rom[ 6585]='h000003c8;  wr_data_rom[ 6585]='h00000000;
    rd_cycle[ 6586] = 1'b1;  wr_cycle[ 6586] = 1'b0;  addr_rom[ 6586]='h000011fc;  wr_data_rom[ 6586]='h00000000;
    rd_cycle[ 6587] = 1'b1;  wr_cycle[ 6587] = 1'b0;  addr_rom[ 6587]='h0000018c;  wr_data_rom[ 6587]='h00000000;
    rd_cycle[ 6588] = 1'b1;  wr_cycle[ 6588] = 1'b0;  addr_rom[ 6588]='h000012b8;  wr_data_rom[ 6588]='h00000000;
    rd_cycle[ 6589] = 1'b0;  wr_cycle[ 6589] = 1'b1;  addr_rom[ 6589]='h000014cc;  wr_data_rom[ 6589]='h000014d6;
    rd_cycle[ 6590] = 1'b1;  wr_cycle[ 6590] = 1'b0;  addr_rom[ 6590]='h00001afc;  wr_data_rom[ 6590]='h00000000;
    rd_cycle[ 6591] = 1'b0;  wr_cycle[ 6591] = 1'b1;  addr_rom[ 6591]='h00000ab4;  wr_data_rom[ 6591]='h00001def;
    rd_cycle[ 6592] = 1'b0;  wr_cycle[ 6592] = 1'b1;  addr_rom[ 6592]='h000005d8;  wr_data_rom[ 6592]='h00001db3;
    rd_cycle[ 6593] = 1'b1;  wr_cycle[ 6593] = 1'b0;  addr_rom[ 6593]='h0000080c;  wr_data_rom[ 6593]='h00000000;
    rd_cycle[ 6594] = 1'b1;  wr_cycle[ 6594] = 1'b0;  addr_rom[ 6594]='h00000de8;  wr_data_rom[ 6594]='h00000000;
    rd_cycle[ 6595] = 1'b0;  wr_cycle[ 6595] = 1'b1;  addr_rom[ 6595]='h000018a4;  wr_data_rom[ 6595]='h00001e8d;
    rd_cycle[ 6596] = 1'b1;  wr_cycle[ 6596] = 1'b0;  addr_rom[ 6596]='h00001a10;  wr_data_rom[ 6596]='h00000000;
    rd_cycle[ 6597] = 1'b1;  wr_cycle[ 6597] = 1'b0;  addr_rom[ 6597]='h00000438;  wr_data_rom[ 6597]='h00000000;
    rd_cycle[ 6598] = 1'b1;  wr_cycle[ 6598] = 1'b0;  addr_rom[ 6598]='h00000e38;  wr_data_rom[ 6598]='h00000000;
    rd_cycle[ 6599] = 1'b0;  wr_cycle[ 6599] = 1'b1;  addr_rom[ 6599]='h00000928;  wr_data_rom[ 6599]='h00000389;
    rd_cycle[ 6600] = 1'b1;  wr_cycle[ 6600] = 1'b0;  addr_rom[ 6600]='h00000524;  wr_data_rom[ 6600]='h00000000;
    rd_cycle[ 6601] = 1'b0;  wr_cycle[ 6601] = 1'b1;  addr_rom[ 6601]='h00001790;  wr_data_rom[ 6601]='h00001a59;
    rd_cycle[ 6602] = 1'b0;  wr_cycle[ 6602] = 1'b1;  addr_rom[ 6602]='h00001148;  wr_data_rom[ 6602]='h00000958;
    rd_cycle[ 6603] = 1'b1;  wr_cycle[ 6603] = 1'b0;  addr_rom[ 6603]='h0000176c;  wr_data_rom[ 6603]='h00000000;
    rd_cycle[ 6604] = 1'b0;  wr_cycle[ 6604] = 1'b1;  addr_rom[ 6604]='h000003ec;  wr_data_rom[ 6604]='h00000f56;
    rd_cycle[ 6605] = 1'b1;  wr_cycle[ 6605] = 1'b0;  addr_rom[ 6605]='h00001844;  wr_data_rom[ 6605]='h00000000;
    rd_cycle[ 6606] = 1'b1;  wr_cycle[ 6606] = 1'b0;  addr_rom[ 6606]='h00001750;  wr_data_rom[ 6606]='h00000000;
    rd_cycle[ 6607] = 1'b0;  wr_cycle[ 6607] = 1'b1;  addr_rom[ 6607]='h000016c0;  wr_data_rom[ 6607]='h0000111b;
    rd_cycle[ 6608] = 1'b0;  wr_cycle[ 6608] = 1'b1;  addr_rom[ 6608]='h00000c90;  wr_data_rom[ 6608]='h000011d8;
    rd_cycle[ 6609] = 1'b0;  wr_cycle[ 6609] = 1'b1;  addr_rom[ 6609]='h00000504;  wr_data_rom[ 6609]='h000007f6;
    rd_cycle[ 6610] = 1'b1;  wr_cycle[ 6610] = 1'b0;  addr_rom[ 6610]='h00000120;  wr_data_rom[ 6610]='h00000000;
    rd_cycle[ 6611] = 1'b0;  wr_cycle[ 6611] = 1'b1;  addr_rom[ 6611]='h00000aa4;  wr_data_rom[ 6611]='h00001675;
    rd_cycle[ 6612] = 1'b0;  wr_cycle[ 6612] = 1'b1;  addr_rom[ 6612]='h00001d0c;  wr_data_rom[ 6612]='h000017ab;
    rd_cycle[ 6613] = 1'b0;  wr_cycle[ 6613] = 1'b1;  addr_rom[ 6613]='h0000105c;  wr_data_rom[ 6613]='h00001d31;
    rd_cycle[ 6614] = 1'b1;  wr_cycle[ 6614] = 1'b0;  addr_rom[ 6614]='h00001db0;  wr_data_rom[ 6614]='h00000000;
    rd_cycle[ 6615] = 1'b0;  wr_cycle[ 6615] = 1'b1;  addr_rom[ 6615]='h00001778;  wr_data_rom[ 6615]='h000015e5;
    rd_cycle[ 6616] = 1'b1;  wr_cycle[ 6616] = 1'b0;  addr_rom[ 6616]='h000015a8;  wr_data_rom[ 6616]='h00000000;
    rd_cycle[ 6617] = 1'b1;  wr_cycle[ 6617] = 1'b0;  addr_rom[ 6617]='h00001140;  wr_data_rom[ 6617]='h00000000;
    rd_cycle[ 6618] = 1'b1;  wr_cycle[ 6618] = 1'b0;  addr_rom[ 6618]='h00000de0;  wr_data_rom[ 6618]='h00000000;
    rd_cycle[ 6619] = 1'b0;  wr_cycle[ 6619] = 1'b1;  addr_rom[ 6619]='h00001488;  wr_data_rom[ 6619]='h00001985;
    rd_cycle[ 6620] = 1'b1;  wr_cycle[ 6620] = 1'b0;  addr_rom[ 6620]='h000015ac;  wr_data_rom[ 6620]='h00000000;
    rd_cycle[ 6621] = 1'b1;  wr_cycle[ 6621] = 1'b0;  addr_rom[ 6621]='h00001d20;  wr_data_rom[ 6621]='h00000000;
    rd_cycle[ 6622] = 1'b1;  wr_cycle[ 6622] = 1'b0;  addr_rom[ 6622]='h00000e44;  wr_data_rom[ 6622]='h00000000;
    rd_cycle[ 6623] = 1'b0;  wr_cycle[ 6623] = 1'b1;  addr_rom[ 6623]='h00001744;  wr_data_rom[ 6623]='h0000046c;
    rd_cycle[ 6624] = 1'b1;  wr_cycle[ 6624] = 1'b0;  addr_rom[ 6624]='h000000dc;  wr_data_rom[ 6624]='h00000000;
    rd_cycle[ 6625] = 1'b0;  wr_cycle[ 6625] = 1'b1;  addr_rom[ 6625]='h00001794;  wr_data_rom[ 6625]='h00000811;
    rd_cycle[ 6626] = 1'b1;  wr_cycle[ 6626] = 1'b0;  addr_rom[ 6626]='h00001138;  wr_data_rom[ 6626]='h00000000;
    rd_cycle[ 6627] = 1'b0;  wr_cycle[ 6627] = 1'b1;  addr_rom[ 6627]='h00000838;  wr_data_rom[ 6627]='h00000b92;
    rd_cycle[ 6628] = 1'b0;  wr_cycle[ 6628] = 1'b1;  addr_rom[ 6628]='h00000f44;  wr_data_rom[ 6628]='h00000748;
    rd_cycle[ 6629] = 1'b1;  wr_cycle[ 6629] = 1'b0;  addr_rom[ 6629]='h00001e74;  wr_data_rom[ 6629]='h00000000;
    rd_cycle[ 6630] = 1'b0;  wr_cycle[ 6630] = 1'b1;  addr_rom[ 6630]='h00000690;  wr_data_rom[ 6630]='h00001c73;
    rd_cycle[ 6631] = 1'b0;  wr_cycle[ 6631] = 1'b1;  addr_rom[ 6631]='h00000f2c;  wr_data_rom[ 6631]='h00001108;
    rd_cycle[ 6632] = 1'b0;  wr_cycle[ 6632] = 1'b1;  addr_rom[ 6632]='h0000054c;  wr_data_rom[ 6632]='h00001838;
    rd_cycle[ 6633] = 1'b1;  wr_cycle[ 6633] = 1'b0;  addr_rom[ 6633]='h00000370;  wr_data_rom[ 6633]='h00000000;
    rd_cycle[ 6634] = 1'b0;  wr_cycle[ 6634] = 1'b1;  addr_rom[ 6634]='h0000028c;  wr_data_rom[ 6634]='h0000066a;
    rd_cycle[ 6635] = 1'b1;  wr_cycle[ 6635] = 1'b0;  addr_rom[ 6635]='h00000d90;  wr_data_rom[ 6635]='h00000000;
    rd_cycle[ 6636] = 1'b1;  wr_cycle[ 6636] = 1'b0;  addr_rom[ 6636]='h000013c0;  wr_data_rom[ 6636]='h00000000;
    rd_cycle[ 6637] = 1'b0;  wr_cycle[ 6637] = 1'b1;  addr_rom[ 6637]='h000001cc;  wr_data_rom[ 6637]='h00001dd3;
    rd_cycle[ 6638] = 1'b0;  wr_cycle[ 6638] = 1'b1;  addr_rom[ 6638]='h00000a84;  wr_data_rom[ 6638]='h00000022;
    rd_cycle[ 6639] = 1'b0;  wr_cycle[ 6639] = 1'b1;  addr_rom[ 6639]='h000008f8;  wr_data_rom[ 6639]='h00000e89;
    rd_cycle[ 6640] = 1'b1;  wr_cycle[ 6640] = 1'b0;  addr_rom[ 6640]='h00001b10;  wr_data_rom[ 6640]='h00000000;
    rd_cycle[ 6641] = 1'b1;  wr_cycle[ 6641] = 1'b0;  addr_rom[ 6641]='h00001704;  wr_data_rom[ 6641]='h00000000;
    rd_cycle[ 6642] = 1'b0;  wr_cycle[ 6642] = 1'b1;  addr_rom[ 6642]='h000006a0;  wr_data_rom[ 6642]='h000012ce;
    rd_cycle[ 6643] = 1'b0;  wr_cycle[ 6643] = 1'b1;  addr_rom[ 6643]='h000016d0;  wr_data_rom[ 6643]='h000015aa;
    rd_cycle[ 6644] = 1'b1;  wr_cycle[ 6644] = 1'b0;  addr_rom[ 6644]='h000018a8;  wr_data_rom[ 6644]='h00000000;
    rd_cycle[ 6645] = 1'b0;  wr_cycle[ 6645] = 1'b1;  addr_rom[ 6645]='h00001c90;  wr_data_rom[ 6645]='h000010d9;
    rd_cycle[ 6646] = 1'b1;  wr_cycle[ 6646] = 1'b0;  addr_rom[ 6646]='h00001458;  wr_data_rom[ 6646]='h00000000;
    rd_cycle[ 6647] = 1'b1;  wr_cycle[ 6647] = 1'b0;  addr_rom[ 6647]='h00001954;  wr_data_rom[ 6647]='h00000000;
    rd_cycle[ 6648] = 1'b1;  wr_cycle[ 6648] = 1'b0;  addr_rom[ 6648]='h000004ac;  wr_data_rom[ 6648]='h00000000;
    rd_cycle[ 6649] = 1'b1;  wr_cycle[ 6649] = 1'b0;  addr_rom[ 6649]='h00001918;  wr_data_rom[ 6649]='h00000000;
    rd_cycle[ 6650] = 1'b1;  wr_cycle[ 6650] = 1'b0;  addr_rom[ 6650]='h00000bf4;  wr_data_rom[ 6650]='h00000000;
    rd_cycle[ 6651] = 1'b0;  wr_cycle[ 6651] = 1'b1;  addr_rom[ 6651]='h000007f4;  wr_data_rom[ 6651]='h0000095d;
    rd_cycle[ 6652] = 1'b0;  wr_cycle[ 6652] = 1'b1;  addr_rom[ 6652]='h00000d18;  wr_data_rom[ 6652]='h00000baf;
    rd_cycle[ 6653] = 1'b0;  wr_cycle[ 6653] = 1'b1;  addr_rom[ 6653]='h00001330;  wr_data_rom[ 6653]='h00000754;
    rd_cycle[ 6654] = 1'b1;  wr_cycle[ 6654] = 1'b0;  addr_rom[ 6654]='h00000194;  wr_data_rom[ 6654]='h00000000;
    rd_cycle[ 6655] = 1'b1;  wr_cycle[ 6655] = 1'b0;  addr_rom[ 6655]='h00001688;  wr_data_rom[ 6655]='h00000000;
    rd_cycle[ 6656] = 1'b1;  wr_cycle[ 6656] = 1'b0;  addr_rom[ 6656]='h000001f4;  wr_data_rom[ 6656]='h00000000;
    rd_cycle[ 6657] = 1'b1;  wr_cycle[ 6657] = 1'b0;  addr_rom[ 6657]='h0000165c;  wr_data_rom[ 6657]='h00000000;
    rd_cycle[ 6658] = 1'b1;  wr_cycle[ 6658] = 1'b0;  addr_rom[ 6658]='h00001160;  wr_data_rom[ 6658]='h00000000;
    rd_cycle[ 6659] = 1'b0;  wr_cycle[ 6659] = 1'b1;  addr_rom[ 6659]='h00000efc;  wr_data_rom[ 6659]='h000001b5;
    rd_cycle[ 6660] = 1'b0;  wr_cycle[ 6660] = 1'b1;  addr_rom[ 6660]='h00000b90;  wr_data_rom[ 6660]='h0000127e;
    rd_cycle[ 6661] = 1'b0;  wr_cycle[ 6661] = 1'b1;  addr_rom[ 6661]='h000005f0;  wr_data_rom[ 6661]='h00000c73;
    rd_cycle[ 6662] = 1'b1;  wr_cycle[ 6662] = 1'b0;  addr_rom[ 6662]='h00000cd0;  wr_data_rom[ 6662]='h00000000;
    rd_cycle[ 6663] = 1'b0;  wr_cycle[ 6663] = 1'b1;  addr_rom[ 6663]='h00001474;  wr_data_rom[ 6663]='h00001f1e;
    rd_cycle[ 6664] = 1'b1;  wr_cycle[ 6664] = 1'b0;  addr_rom[ 6664]='h00000ae0;  wr_data_rom[ 6664]='h00000000;
    rd_cycle[ 6665] = 1'b0;  wr_cycle[ 6665] = 1'b1;  addr_rom[ 6665]='h00000a3c;  wr_data_rom[ 6665]='h00001cda;
    rd_cycle[ 6666] = 1'b1;  wr_cycle[ 6666] = 1'b0;  addr_rom[ 6666]='h00000854;  wr_data_rom[ 6666]='h00000000;
    rd_cycle[ 6667] = 1'b0;  wr_cycle[ 6667] = 1'b1;  addr_rom[ 6667]='h00001e6c;  wr_data_rom[ 6667]='h00001386;
    rd_cycle[ 6668] = 1'b0;  wr_cycle[ 6668] = 1'b1;  addr_rom[ 6668]='h000013b0;  wr_data_rom[ 6668]='h00001579;
    rd_cycle[ 6669] = 1'b0;  wr_cycle[ 6669] = 1'b1;  addr_rom[ 6669]='h00000b38;  wr_data_rom[ 6669]='h00000336;
    rd_cycle[ 6670] = 1'b1;  wr_cycle[ 6670] = 1'b0;  addr_rom[ 6670]='h00000984;  wr_data_rom[ 6670]='h00000000;
    rd_cycle[ 6671] = 1'b0;  wr_cycle[ 6671] = 1'b1;  addr_rom[ 6671]='h00001434;  wr_data_rom[ 6671]='h00000260;
    rd_cycle[ 6672] = 1'b1;  wr_cycle[ 6672] = 1'b0;  addr_rom[ 6672]='h000007e8;  wr_data_rom[ 6672]='h00000000;
    rd_cycle[ 6673] = 1'b1;  wr_cycle[ 6673] = 1'b0;  addr_rom[ 6673]='h00000b4c;  wr_data_rom[ 6673]='h00000000;
    rd_cycle[ 6674] = 1'b1;  wr_cycle[ 6674] = 1'b0;  addr_rom[ 6674]='h0000014c;  wr_data_rom[ 6674]='h00000000;
    rd_cycle[ 6675] = 1'b0;  wr_cycle[ 6675] = 1'b1;  addr_rom[ 6675]='h00001628;  wr_data_rom[ 6675]='h00000506;
    rd_cycle[ 6676] = 1'b1;  wr_cycle[ 6676] = 1'b0;  addr_rom[ 6676]='h00001878;  wr_data_rom[ 6676]='h00000000;
    rd_cycle[ 6677] = 1'b1;  wr_cycle[ 6677] = 1'b0;  addr_rom[ 6677]='h00001e5c;  wr_data_rom[ 6677]='h00000000;
    rd_cycle[ 6678] = 1'b0;  wr_cycle[ 6678] = 1'b1;  addr_rom[ 6678]='h00001554;  wr_data_rom[ 6678]='h00000d72;
    rd_cycle[ 6679] = 1'b1;  wr_cycle[ 6679] = 1'b0;  addr_rom[ 6679]='h0000122c;  wr_data_rom[ 6679]='h00000000;
    rd_cycle[ 6680] = 1'b1;  wr_cycle[ 6680] = 1'b0;  addr_rom[ 6680]='h00001444;  wr_data_rom[ 6680]='h00000000;
    rd_cycle[ 6681] = 1'b0;  wr_cycle[ 6681] = 1'b1;  addr_rom[ 6681]='h000014a8;  wr_data_rom[ 6681]='h00000993;
    rd_cycle[ 6682] = 1'b0;  wr_cycle[ 6682] = 1'b1;  addr_rom[ 6682]='h00000a5c;  wr_data_rom[ 6682]='h000001f9;
    rd_cycle[ 6683] = 1'b1;  wr_cycle[ 6683] = 1'b0;  addr_rom[ 6683]='h00001d3c;  wr_data_rom[ 6683]='h00000000;
    rd_cycle[ 6684] = 1'b0;  wr_cycle[ 6684] = 1'b1;  addr_rom[ 6684]='h00001c84;  wr_data_rom[ 6684]='h00001994;
    rd_cycle[ 6685] = 1'b0;  wr_cycle[ 6685] = 1'b1;  addr_rom[ 6685]='h00001134;  wr_data_rom[ 6685]='h000003db;
    rd_cycle[ 6686] = 1'b1;  wr_cycle[ 6686] = 1'b0;  addr_rom[ 6686]='h0000049c;  wr_data_rom[ 6686]='h00000000;
    rd_cycle[ 6687] = 1'b0;  wr_cycle[ 6687] = 1'b1;  addr_rom[ 6687]='h00000abc;  wr_data_rom[ 6687]='h000003f7;
    rd_cycle[ 6688] = 1'b0;  wr_cycle[ 6688] = 1'b1;  addr_rom[ 6688]='h00000ba0;  wr_data_rom[ 6688]='h00000c9c;
    rd_cycle[ 6689] = 1'b0;  wr_cycle[ 6689] = 1'b1;  addr_rom[ 6689]='h000000f4;  wr_data_rom[ 6689]='h00001e74;
    rd_cycle[ 6690] = 1'b1;  wr_cycle[ 6690] = 1'b0;  addr_rom[ 6690]='h00000064;  wr_data_rom[ 6690]='h00000000;
    rd_cycle[ 6691] = 1'b1;  wr_cycle[ 6691] = 1'b0;  addr_rom[ 6691]='h00001960;  wr_data_rom[ 6691]='h00000000;
    rd_cycle[ 6692] = 1'b0;  wr_cycle[ 6692] = 1'b1;  addr_rom[ 6692]='h0000048c;  wr_data_rom[ 6692]='h00000259;
    rd_cycle[ 6693] = 1'b1;  wr_cycle[ 6693] = 1'b0;  addr_rom[ 6693]='h00001754;  wr_data_rom[ 6693]='h00000000;
    rd_cycle[ 6694] = 1'b0;  wr_cycle[ 6694] = 1'b1;  addr_rom[ 6694]='h00000288;  wr_data_rom[ 6694]='h00000de2;
    rd_cycle[ 6695] = 1'b1;  wr_cycle[ 6695] = 1'b0;  addr_rom[ 6695]='h00000ad0;  wr_data_rom[ 6695]='h00000000;
    rd_cycle[ 6696] = 1'b0;  wr_cycle[ 6696] = 1'b1;  addr_rom[ 6696]='h00000f10;  wr_data_rom[ 6696]='h00001763;
    rd_cycle[ 6697] = 1'b0;  wr_cycle[ 6697] = 1'b1;  addr_rom[ 6697]='h00001108;  wr_data_rom[ 6697]='h00000476;
    rd_cycle[ 6698] = 1'b0;  wr_cycle[ 6698] = 1'b1;  addr_rom[ 6698]='h00000908;  wr_data_rom[ 6698]='h00001729;
    rd_cycle[ 6699] = 1'b0;  wr_cycle[ 6699] = 1'b1;  addr_rom[ 6699]='h00000304;  wr_data_rom[ 6699]='h0000188e;
    rd_cycle[ 6700] = 1'b1;  wr_cycle[ 6700] = 1'b0;  addr_rom[ 6700]='h00000ab0;  wr_data_rom[ 6700]='h00000000;
    rd_cycle[ 6701] = 1'b1;  wr_cycle[ 6701] = 1'b0;  addr_rom[ 6701]='h00001134;  wr_data_rom[ 6701]='h00000000;
    rd_cycle[ 6702] = 1'b1;  wr_cycle[ 6702] = 1'b0;  addr_rom[ 6702]='h00001bc4;  wr_data_rom[ 6702]='h00000000;
    rd_cycle[ 6703] = 1'b1;  wr_cycle[ 6703] = 1'b0;  addr_rom[ 6703]='h000002d4;  wr_data_rom[ 6703]='h00000000;
    rd_cycle[ 6704] = 1'b0;  wr_cycle[ 6704] = 1'b1;  addr_rom[ 6704]='h000000cc;  wr_data_rom[ 6704]='h00000f15;
    rd_cycle[ 6705] = 1'b0;  wr_cycle[ 6705] = 1'b1;  addr_rom[ 6705]='h00000600;  wr_data_rom[ 6705]='h0000009c;
    rd_cycle[ 6706] = 1'b1;  wr_cycle[ 6706] = 1'b0;  addr_rom[ 6706]='h0000048c;  wr_data_rom[ 6706]='h00000000;
    rd_cycle[ 6707] = 1'b1;  wr_cycle[ 6707] = 1'b0;  addr_rom[ 6707]='h00001104;  wr_data_rom[ 6707]='h00000000;
    rd_cycle[ 6708] = 1'b1;  wr_cycle[ 6708] = 1'b0;  addr_rom[ 6708]='h00001b80;  wr_data_rom[ 6708]='h00000000;
    rd_cycle[ 6709] = 1'b1;  wr_cycle[ 6709] = 1'b0;  addr_rom[ 6709]='h00000350;  wr_data_rom[ 6709]='h00000000;
    rd_cycle[ 6710] = 1'b1;  wr_cycle[ 6710] = 1'b0;  addr_rom[ 6710]='h000004fc;  wr_data_rom[ 6710]='h00000000;
    rd_cycle[ 6711] = 1'b1;  wr_cycle[ 6711] = 1'b0;  addr_rom[ 6711]='h00001748;  wr_data_rom[ 6711]='h00000000;
    rd_cycle[ 6712] = 1'b1;  wr_cycle[ 6712] = 1'b0;  addr_rom[ 6712]='h00000528;  wr_data_rom[ 6712]='h00000000;
    rd_cycle[ 6713] = 1'b0;  wr_cycle[ 6713] = 1'b1;  addr_rom[ 6713]='h00000214;  wr_data_rom[ 6713]='h00000551;
    rd_cycle[ 6714] = 1'b1;  wr_cycle[ 6714] = 1'b0;  addr_rom[ 6714]='h000010f4;  wr_data_rom[ 6714]='h00000000;
    rd_cycle[ 6715] = 1'b0;  wr_cycle[ 6715] = 1'b1;  addr_rom[ 6715]='h000016a4;  wr_data_rom[ 6715]='h00001d8f;
    rd_cycle[ 6716] = 1'b0;  wr_cycle[ 6716] = 1'b1;  addr_rom[ 6716]='h00001558;  wr_data_rom[ 6716]='h00000fad;
    rd_cycle[ 6717] = 1'b1;  wr_cycle[ 6717] = 1'b0;  addr_rom[ 6717]='h00001e30;  wr_data_rom[ 6717]='h00000000;
    rd_cycle[ 6718] = 1'b1;  wr_cycle[ 6718] = 1'b0;  addr_rom[ 6718]='h00000bc0;  wr_data_rom[ 6718]='h00000000;
    rd_cycle[ 6719] = 1'b0;  wr_cycle[ 6719] = 1'b1;  addr_rom[ 6719]='h000019c4;  wr_data_rom[ 6719]='h0000105f;
    rd_cycle[ 6720] = 1'b0;  wr_cycle[ 6720] = 1'b1;  addr_rom[ 6720]='h000006bc;  wr_data_rom[ 6720]='h000016fe;
    rd_cycle[ 6721] = 1'b1;  wr_cycle[ 6721] = 1'b0;  addr_rom[ 6721]='h00000670;  wr_data_rom[ 6721]='h00000000;
    rd_cycle[ 6722] = 1'b1;  wr_cycle[ 6722] = 1'b0;  addr_rom[ 6722]='h00000ee4;  wr_data_rom[ 6722]='h00000000;
    rd_cycle[ 6723] = 1'b1;  wr_cycle[ 6723] = 1'b0;  addr_rom[ 6723]='h000009cc;  wr_data_rom[ 6723]='h00000000;
    rd_cycle[ 6724] = 1'b1;  wr_cycle[ 6724] = 1'b0;  addr_rom[ 6724]='h00001b20;  wr_data_rom[ 6724]='h00000000;
    rd_cycle[ 6725] = 1'b1;  wr_cycle[ 6725] = 1'b0;  addr_rom[ 6725]='h0000015c;  wr_data_rom[ 6725]='h00000000;
    rd_cycle[ 6726] = 1'b0;  wr_cycle[ 6726] = 1'b1;  addr_rom[ 6726]='h000005e8;  wr_data_rom[ 6726]='h00000115;
    rd_cycle[ 6727] = 1'b1;  wr_cycle[ 6727] = 1'b0;  addr_rom[ 6727]='h00001a34;  wr_data_rom[ 6727]='h00000000;
    rd_cycle[ 6728] = 1'b1;  wr_cycle[ 6728] = 1'b0;  addr_rom[ 6728]='h000006d0;  wr_data_rom[ 6728]='h00000000;
    rd_cycle[ 6729] = 1'b1;  wr_cycle[ 6729] = 1'b0;  addr_rom[ 6729]='h000006cc;  wr_data_rom[ 6729]='h00000000;
    rd_cycle[ 6730] = 1'b0;  wr_cycle[ 6730] = 1'b1;  addr_rom[ 6730]='h000006a4;  wr_data_rom[ 6730]='h00000d29;
    rd_cycle[ 6731] = 1'b1;  wr_cycle[ 6731] = 1'b0;  addr_rom[ 6731]='h00001cd0;  wr_data_rom[ 6731]='h00000000;
    rd_cycle[ 6732] = 1'b1;  wr_cycle[ 6732] = 1'b0;  addr_rom[ 6732]='h00001318;  wr_data_rom[ 6732]='h00000000;
    rd_cycle[ 6733] = 1'b1;  wr_cycle[ 6733] = 1'b0;  addr_rom[ 6733]='h00001334;  wr_data_rom[ 6733]='h00000000;
    rd_cycle[ 6734] = 1'b1;  wr_cycle[ 6734] = 1'b0;  addr_rom[ 6734]='h00001094;  wr_data_rom[ 6734]='h00000000;
    rd_cycle[ 6735] = 1'b0;  wr_cycle[ 6735] = 1'b1;  addr_rom[ 6735]='h00000670;  wr_data_rom[ 6735]='h000004a8;
    rd_cycle[ 6736] = 1'b1;  wr_cycle[ 6736] = 1'b0;  addr_rom[ 6736]='h000002b8;  wr_data_rom[ 6736]='h00000000;
    rd_cycle[ 6737] = 1'b1;  wr_cycle[ 6737] = 1'b0;  addr_rom[ 6737]='h0000148c;  wr_data_rom[ 6737]='h00000000;
    rd_cycle[ 6738] = 1'b1;  wr_cycle[ 6738] = 1'b0;  addr_rom[ 6738]='h000015d8;  wr_data_rom[ 6738]='h00000000;
    rd_cycle[ 6739] = 1'b0;  wr_cycle[ 6739] = 1'b1;  addr_rom[ 6739]='h00001744;  wr_data_rom[ 6739]='h00001559;
    rd_cycle[ 6740] = 1'b1;  wr_cycle[ 6740] = 1'b0;  addr_rom[ 6740]='h0000069c;  wr_data_rom[ 6740]='h00000000;
    rd_cycle[ 6741] = 1'b0;  wr_cycle[ 6741] = 1'b1;  addr_rom[ 6741]='h00001e68;  wr_data_rom[ 6741]='h00000f45;
    rd_cycle[ 6742] = 1'b1;  wr_cycle[ 6742] = 1'b0;  addr_rom[ 6742]='h00001c30;  wr_data_rom[ 6742]='h00000000;
    rd_cycle[ 6743] = 1'b0;  wr_cycle[ 6743] = 1'b1;  addr_rom[ 6743]='h00000240;  wr_data_rom[ 6743]='h00001458;
    rd_cycle[ 6744] = 1'b0;  wr_cycle[ 6744] = 1'b1;  addr_rom[ 6744]='h000004f8;  wr_data_rom[ 6744]='h00000662;
    rd_cycle[ 6745] = 1'b1;  wr_cycle[ 6745] = 1'b0;  addr_rom[ 6745]='h00000798;  wr_data_rom[ 6745]='h00000000;
    rd_cycle[ 6746] = 1'b1;  wr_cycle[ 6746] = 1'b0;  addr_rom[ 6746]='h000017f8;  wr_data_rom[ 6746]='h00000000;
    rd_cycle[ 6747] = 1'b1;  wr_cycle[ 6747] = 1'b0;  addr_rom[ 6747]='h000006a8;  wr_data_rom[ 6747]='h00000000;
    rd_cycle[ 6748] = 1'b1;  wr_cycle[ 6748] = 1'b0;  addr_rom[ 6748]='h0000111c;  wr_data_rom[ 6748]='h00000000;
    rd_cycle[ 6749] = 1'b0;  wr_cycle[ 6749] = 1'b1;  addr_rom[ 6749]='h00000648;  wr_data_rom[ 6749]='h00000d4b;
    rd_cycle[ 6750] = 1'b1;  wr_cycle[ 6750] = 1'b0;  addr_rom[ 6750]='h000006c0;  wr_data_rom[ 6750]='h00000000;
    rd_cycle[ 6751] = 1'b1;  wr_cycle[ 6751] = 1'b0;  addr_rom[ 6751]='h0000112c;  wr_data_rom[ 6751]='h00000000;
    rd_cycle[ 6752] = 1'b1;  wr_cycle[ 6752] = 1'b0;  addr_rom[ 6752]='h00001a28;  wr_data_rom[ 6752]='h00000000;
    rd_cycle[ 6753] = 1'b1;  wr_cycle[ 6753] = 1'b0;  addr_rom[ 6753]='h000008f0;  wr_data_rom[ 6753]='h00000000;
    rd_cycle[ 6754] = 1'b0;  wr_cycle[ 6754] = 1'b1;  addr_rom[ 6754]='h00001200;  wr_data_rom[ 6754]='h000013ed;
    rd_cycle[ 6755] = 1'b0;  wr_cycle[ 6755] = 1'b1;  addr_rom[ 6755]='h00000924;  wr_data_rom[ 6755]='h00000491;
    rd_cycle[ 6756] = 1'b0;  wr_cycle[ 6756] = 1'b1;  addr_rom[ 6756]='h000005b4;  wr_data_rom[ 6756]='h000016c6;
    rd_cycle[ 6757] = 1'b0;  wr_cycle[ 6757] = 1'b1;  addr_rom[ 6757]='h00001e24;  wr_data_rom[ 6757]='h00000cbf;
    rd_cycle[ 6758] = 1'b0;  wr_cycle[ 6758] = 1'b1;  addr_rom[ 6758]='h00001934;  wr_data_rom[ 6758]='h00000095;
    rd_cycle[ 6759] = 1'b0;  wr_cycle[ 6759] = 1'b1;  addr_rom[ 6759]='h00001914;  wr_data_rom[ 6759]='h000010dc;
    rd_cycle[ 6760] = 1'b1;  wr_cycle[ 6760] = 1'b0;  addr_rom[ 6760]='h00000480;  wr_data_rom[ 6760]='h00000000;
    rd_cycle[ 6761] = 1'b1;  wr_cycle[ 6761] = 1'b0;  addr_rom[ 6761]='h00000e0c;  wr_data_rom[ 6761]='h00000000;
    rd_cycle[ 6762] = 1'b0;  wr_cycle[ 6762] = 1'b1;  addr_rom[ 6762]='h000008fc;  wr_data_rom[ 6762]='h00000fa4;
    rd_cycle[ 6763] = 1'b1;  wr_cycle[ 6763] = 1'b0;  addr_rom[ 6763]='h00000a38;  wr_data_rom[ 6763]='h00000000;
    rd_cycle[ 6764] = 1'b1;  wr_cycle[ 6764] = 1'b0;  addr_rom[ 6764]='h000007b4;  wr_data_rom[ 6764]='h00000000;
    rd_cycle[ 6765] = 1'b0;  wr_cycle[ 6765] = 1'b1;  addr_rom[ 6765]='h00001c50;  wr_data_rom[ 6765]='h00000024;
    rd_cycle[ 6766] = 1'b0;  wr_cycle[ 6766] = 1'b1;  addr_rom[ 6766]='h00000bac;  wr_data_rom[ 6766]='h000017b5;
    rd_cycle[ 6767] = 1'b0;  wr_cycle[ 6767] = 1'b1;  addr_rom[ 6767]='h00000a20;  wr_data_rom[ 6767]='h00000497;
    rd_cycle[ 6768] = 1'b1;  wr_cycle[ 6768] = 1'b0;  addr_rom[ 6768]='h00000fcc;  wr_data_rom[ 6768]='h00000000;
    rd_cycle[ 6769] = 1'b0;  wr_cycle[ 6769] = 1'b1;  addr_rom[ 6769]='h0000157c;  wr_data_rom[ 6769]='h00001631;
    rd_cycle[ 6770] = 1'b1;  wr_cycle[ 6770] = 1'b0;  addr_rom[ 6770]='h00001d64;  wr_data_rom[ 6770]='h00000000;
    rd_cycle[ 6771] = 1'b0;  wr_cycle[ 6771] = 1'b1;  addr_rom[ 6771]='h00000924;  wr_data_rom[ 6771]='h0000070a;
    rd_cycle[ 6772] = 1'b0;  wr_cycle[ 6772] = 1'b1;  addr_rom[ 6772]='h00000970;  wr_data_rom[ 6772]='h00000f0a;
    rd_cycle[ 6773] = 1'b0;  wr_cycle[ 6773] = 1'b1;  addr_rom[ 6773]='h00001450;  wr_data_rom[ 6773]='h00001398;
    rd_cycle[ 6774] = 1'b1;  wr_cycle[ 6774] = 1'b0;  addr_rom[ 6774]='h000017b4;  wr_data_rom[ 6774]='h00000000;
    rd_cycle[ 6775] = 1'b0;  wr_cycle[ 6775] = 1'b1;  addr_rom[ 6775]='h00000a14;  wr_data_rom[ 6775]='h0000113f;
    rd_cycle[ 6776] = 1'b0;  wr_cycle[ 6776] = 1'b1;  addr_rom[ 6776]='h0000123c;  wr_data_rom[ 6776]='h0000084a;
    rd_cycle[ 6777] = 1'b1;  wr_cycle[ 6777] = 1'b0;  addr_rom[ 6777]='h00001ecc;  wr_data_rom[ 6777]='h00000000;
    rd_cycle[ 6778] = 1'b0;  wr_cycle[ 6778] = 1'b1;  addr_rom[ 6778]='h00001530;  wr_data_rom[ 6778]='h00001f3b;
    rd_cycle[ 6779] = 1'b1;  wr_cycle[ 6779] = 1'b0;  addr_rom[ 6779]='h00001c8c;  wr_data_rom[ 6779]='h00000000;
    rd_cycle[ 6780] = 1'b0;  wr_cycle[ 6780] = 1'b1;  addr_rom[ 6780]='h000018d8;  wr_data_rom[ 6780]='h000014eb;
    rd_cycle[ 6781] = 1'b1;  wr_cycle[ 6781] = 1'b0;  addr_rom[ 6781]='h00001434;  wr_data_rom[ 6781]='h00000000;
    rd_cycle[ 6782] = 1'b0;  wr_cycle[ 6782] = 1'b1;  addr_rom[ 6782]='h00001270;  wr_data_rom[ 6782]='h0000192e;
    rd_cycle[ 6783] = 1'b1;  wr_cycle[ 6783] = 1'b0;  addr_rom[ 6783]='h00000a48;  wr_data_rom[ 6783]='h00000000;
    rd_cycle[ 6784] = 1'b1;  wr_cycle[ 6784] = 1'b0;  addr_rom[ 6784]='h00001a78;  wr_data_rom[ 6784]='h00000000;
    rd_cycle[ 6785] = 1'b1;  wr_cycle[ 6785] = 1'b0;  addr_rom[ 6785]='h00001284;  wr_data_rom[ 6785]='h00000000;
    rd_cycle[ 6786] = 1'b1;  wr_cycle[ 6786] = 1'b0;  addr_rom[ 6786]='h00000e24;  wr_data_rom[ 6786]='h00000000;
    rd_cycle[ 6787] = 1'b1;  wr_cycle[ 6787] = 1'b0;  addr_rom[ 6787]='h00001d04;  wr_data_rom[ 6787]='h00000000;
    rd_cycle[ 6788] = 1'b0;  wr_cycle[ 6788] = 1'b1;  addr_rom[ 6788]='h00000258;  wr_data_rom[ 6788]='h00000c51;
    rd_cycle[ 6789] = 1'b1;  wr_cycle[ 6789] = 1'b0;  addr_rom[ 6789]='h000006d4;  wr_data_rom[ 6789]='h00000000;
    rd_cycle[ 6790] = 1'b0;  wr_cycle[ 6790] = 1'b1;  addr_rom[ 6790]='h00000c30;  wr_data_rom[ 6790]='h000015dc;
    rd_cycle[ 6791] = 1'b1;  wr_cycle[ 6791] = 1'b0;  addr_rom[ 6791]='h00000610;  wr_data_rom[ 6791]='h00000000;
    rd_cycle[ 6792] = 1'b0;  wr_cycle[ 6792] = 1'b1;  addr_rom[ 6792]='h00000a90;  wr_data_rom[ 6792]='h00000aa7;
    rd_cycle[ 6793] = 1'b0;  wr_cycle[ 6793] = 1'b1;  addr_rom[ 6793]='h00000074;  wr_data_rom[ 6793]='h00000967;
    rd_cycle[ 6794] = 1'b1;  wr_cycle[ 6794] = 1'b0;  addr_rom[ 6794]='h00000eb0;  wr_data_rom[ 6794]='h00000000;
    rd_cycle[ 6795] = 1'b0;  wr_cycle[ 6795] = 1'b1;  addr_rom[ 6795]='h00000a24;  wr_data_rom[ 6795]='h000009b5;
    rd_cycle[ 6796] = 1'b1;  wr_cycle[ 6796] = 1'b0;  addr_rom[ 6796]='h000013e4;  wr_data_rom[ 6796]='h00000000;
    rd_cycle[ 6797] = 1'b0;  wr_cycle[ 6797] = 1'b1;  addr_rom[ 6797]='h00000188;  wr_data_rom[ 6797]='h00000902;
    rd_cycle[ 6798] = 1'b0;  wr_cycle[ 6798] = 1'b1;  addr_rom[ 6798]='h00001e1c;  wr_data_rom[ 6798]='h00000b01;
    rd_cycle[ 6799] = 1'b0;  wr_cycle[ 6799] = 1'b1;  addr_rom[ 6799]='h00001778;  wr_data_rom[ 6799]='h00000e9f;
    rd_cycle[ 6800] = 1'b1;  wr_cycle[ 6800] = 1'b0;  addr_rom[ 6800]='h00000768;  wr_data_rom[ 6800]='h00000000;
    rd_cycle[ 6801] = 1'b1;  wr_cycle[ 6801] = 1'b0;  addr_rom[ 6801]='h00001d18;  wr_data_rom[ 6801]='h00000000;
    rd_cycle[ 6802] = 1'b0;  wr_cycle[ 6802] = 1'b1;  addr_rom[ 6802]='h00001ebc;  wr_data_rom[ 6802]='h00001ed8;
    rd_cycle[ 6803] = 1'b1;  wr_cycle[ 6803] = 1'b0;  addr_rom[ 6803]='h00001500;  wr_data_rom[ 6803]='h00000000;
    rd_cycle[ 6804] = 1'b0;  wr_cycle[ 6804] = 1'b1;  addr_rom[ 6804]='h0000042c;  wr_data_rom[ 6804]='h000014f8;
    rd_cycle[ 6805] = 1'b0;  wr_cycle[ 6805] = 1'b1;  addr_rom[ 6805]='h00001164;  wr_data_rom[ 6805]='h00000fc6;
    rd_cycle[ 6806] = 1'b1;  wr_cycle[ 6806] = 1'b0;  addr_rom[ 6806]='h00001f08;  wr_data_rom[ 6806]='h00000000;
    rd_cycle[ 6807] = 1'b0;  wr_cycle[ 6807] = 1'b1;  addr_rom[ 6807]='h000004f0;  wr_data_rom[ 6807]='h000015b0;
    rd_cycle[ 6808] = 1'b0;  wr_cycle[ 6808] = 1'b1;  addr_rom[ 6808]='h00001af8;  wr_data_rom[ 6808]='h00001c84;
    rd_cycle[ 6809] = 1'b1;  wr_cycle[ 6809] = 1'b0;  addr_rom[ 6809]='h00000950;  wr_data_rom[ 6809]='h00000000;
    rd_cycle[ 6810] = 1'b1;  wr_cycle[ 6810] = 1'b0;  addr_rom[ 6810]='h00001034;  wr_data_rom[ 6810]='h00000000;
    rd_cycle[ 6811] = 1'b1;  wr_cycle[ 6811] = 1'b0;  addr_rom[ 6811]='h000015a8;  wr_data_rom[ 6811]='h00000000;
    rd_cycle[ 6812] = 1'b1;  wr_cycle[ 6812] = 1'b0;  addr_rom[ 6812]='h00000728;  wr_data_rom[ 6812]='h00000000;
    rd_cycle[ 6813] = 1'b1;  wr_cycle[ 6813] = 1'b0;  addr_rom[ 6813]='h000002e8;  wr_data_rom[ 6813]='h00000000;
    rd_cycle[ 6814] = 1'b0;  wr_cycle[ 6814] = 1'b1;  addr_rom[ 6814]='h000009f8;  wr_data_rom[ 6814]='h00001ca3;
    rd_cycle[ 6815] = 1'b0;  wr_cycle[ 6815] = 1'b1;  addr_rom[ 6815]='h00001320;  wr_data_rom[ 6815]='h00000b35;
    rd_cycle[ 6816] = 1'b0;  wr_cycle[ 6816] = 1'b1;  addr_rom[ 6816]='h00001b38;  wr_data_rom[ 6816]='h00001076;
    rd_cycle[ 6817] = 1'b1;  wr_cycle[ 6817] = 1'b0;  addr_rom[ 6817]='h00001554;  wr_data_rom[ 6817]='h00000000;
    rd_cycle[ 6818] = 1'b1;  wr_cycle[ 6818] = 1'b0;  addr_rom[ 6818]='h00001130;  wr_data_rom[ 6818]='h00000000;
    rd_cycle[ 6819] = 1'b1;  wr_cycle[ 6819] = 1'b0;  addr_rom[ 6819]='h00000980;  wr_data_rom[ 6819]='h00000000;
    rd_cycle[ 6820] = 1'b0;  wr_cycle[ 6820] = 1'b1;  addr_rom[ 6820]='h00001198;  wr_data_rom[ 6820]='h00001a7b;
    rd_cycle[ 6821] = 1'b0;  wr_cycle[ 6821] = 1'b1;  addr_rom[ 6821]='h00001554;  wr_data_rom[ 6821]='h000004bc;
    rd_cycle[ 6822] = 1'b1;  wr_cycle[ 6822] = 1'b0;  addr_rom[ 6822]='h0000072c;  wr_data_rom[ 6822]='h00000000;
    rd_cycle[ 6823] = 1'b0;  wr_cycle[ 6823] = 1'b1;  addr_rom[ 6823]='h00001560;  wr_data_rom[ 6823]='h00000358;
    rd_cycle[ 6824] = 1'b0;  wr_cycle[ 6824] = 1'b1;  addr_rom[ 6824]='h00000f8c;  wr_data_rom[ 6824]='h0000132a;
    rd_cycle[ 6825] = 1'b1;  wr_cycle[ 6825] = 1'b0;  addr_rom[ 6825]='h00000f2c;  wr_data_rom[ 6825]='h00000000;
    rd_cycle[ 6826] = 1'b0;  wr_cycle[ 6826] = 1'b1;  addr_rom[ 6826]='h00000fec;  wr_data_rom[ 6826]='h00001a75;
    rd_cycle[ 6827] = 1'b1;  wr_cycle[ 6827] = 1'b0;  addr_rom[ 6827]='h00001804;  wr_data_rom[ 6827]='h00000000;
    rd_cycle[ 6828] = 1'b1;  wr_cycle[ 6828] = 1'b0;  addr_rom[ 6828]='h00000fc0;  wr_data_rom[ 6828]='h00000000;
    rd_cycle[ 6829] = 1'b0;  wr_cycle[ 6829] = 1'b1;  addr_rom[ 6829]='h00000268;  wr_data_rom[ 6829]='h000002b3;
    rd_cycle[ 6830] = 1'b0;  wr_cycle[ 6830] = 1'b1;  addr_rom[ 6830]='h00000f58;  wr_data_rom[ 6830]='h00000491;
    rd_cycle[ 6831] = 1'b0;  wr_cycle[ 6831] = 1'b1;  addr_rom[ 6831]='h000002f0;  wr_data_rom[ 6831]='h000009c0;
    rd_cycle[ 6832] = 1'b1;  wr_cycle[ 6832] = 1'b0;  addr_rom[ 6832]='h000014c8;  wr_data_rom[ 6832]='h00000000;
    rd_cycle[ 6833] = 1'b0;  wr_cycle[ 6833] = 1'b1;  addr_rom[ 6833]='h00001838;  wr_data_rom[ 6833]='h00000446;
    rd_cycle[ 6834] = 1'b0;  wr_cycle[ 6834] = 1'b1;  addr_rom[ 6834]='h000018f8;  wr_data_rom[ 6834]='h000008cd;
    rd_cycle[ 6835] = 1'b0;  wr_cycle[ 6835] = 1'b1;  addr_rom[ 6835]='h0000048c;  wr_data_rom[ 6835]='h0000055d;
    rd_cycle[ 6836] = 1'b0;  wr_cycle[ 6836] = 1'b1;  addr_rom[ 6836]='h0000070c;  wr_data_rom[ 6836]='h000011e9;
    rd_cycle[ 6837] = 1'b1;  wr_cycle[ 6837] = 1'b0;  addr_rom[ 6837]='h00000a6c;  wr_data_rom[ 6837]='h00000000;
    rd_cycle[ 6838] = 1'b0;  wr_cycle[ 6838] = 1'b1;  addr_rom[ 6838]='h00001360;  wr_data_rom[ 6838]='h00001748;
    rd_cycle[ 6839] = 1'b1;  wr_cycle[ 6839] = 1'b0;  addr_rom[ 6839]='h00000668;  wr_data_rom[ 6839]='h00000000;
    rd_cycle[ 6840] = 1'b1;  wr_cycle[ 6840] = 1'b0;  addr_rom[ 6840]='h00001064;  wr_data_rom[ 6840]='h00000000;
    rd_cycle[ 6841] = 1'b0;  wr_cycle[ 6841] = 1'b1;  addr_rom[ 6841]='h00000c6c;  wr_data_rom[ 6841]='h0000132b;
    rd_cycle[ 6842] = 1'b0;  wr_cycle[ 6842] = 1'b1;  addr_rom[ 6842]='h00000d28;  wr_data_rom[ 6842]='h00000206;
    rd_cycle[ 6843] = 1'b1;  wr_cycle[ 6843] = 1'b0;  addr_rom[ 6843]='h0000196c;  wr_data_rom[ 6843]='h00000000;
    rd_cycle[ 6844] = 1'b0;  wr_cycle[ 6844] = 1'b1;  addr_rom[ 6844]='h00000518;  wr_data_rom[ 6844]='h000000e4;
    rd_cycle[ 6845] = 1'b0;  wr_cycle[ 6845] = 1'b1;  addr_rom[ 6845]='h000013fc;  wr_data_rom[ 6845]='h0000133f;
    rd_cycle[ 6846] = 1'b0;  wr_cycle[ 6846] = 1'b1;  addr_rom[ 6846]='h00001b48;  wr_data_rom[ 6846]='h0000151c;
    rd_cycle[ 6847] = 1'b0;  wr_cycle[ 6847] = 1'b1;  addr_rom[ 6847]='h0000121c;  wr_data_rom[ 6847]='h00001eef;
    rd_cycle[ 6848] = 1'b1;  wr_cycle[ 6848] = 1'b0;  addr_rom[ 6848]='h00001898;  wr_data_rom[ 6848]='h00000000;
    rd_cycle[ 6849] = 1'b1;  wr_cycle[ 6849] = 1'b0;  addr_rom[ 6849]='h00000c64;  wr_data_rom[ 6849]='h00000000;
    rd_cycle[ 6850] = 1'b0;  wr_cycle[ 6850] = 1'b1;  addr_rom[ 6850]='h00000b34;  wr_data_rom[ 6850]='h00000d88;
    rd_cycle[ 6851] = 1'b0;  wr_cycle[ 6851] = 1'b1;  addr_rom[ 6851]='h00001378;  wr_data_rom[ 6851]='h0000166f;
    rd_cycle[ 6852] = 1'b0;  wr_cycle[ 6852] = 1'b1;  addr_rom[ 6852]='h00001cc0;  wr_data_rom[ 6852]='h000009e7;
    rd_cycle[ 6853] = 1'b1;  wr_cycle[ 6853] = 1'b0;  addr_rom[ 6853]='h000017f4;  wr_data_rom[ 6853]='h00000000;
    rd_cycle[ 6854] = 1'b0;  wr_cycle[ 6854] = 1'b1;  addr_rom[ 6854]='h0000015c;  wr_data_rom[ 6854]='h00001516;
    rd_cycle[ 6855] = 1'b0;  wr_cycle[ 6855] = 1'b1;  addr_rom[ 6855]='h00001e6c;  wr_data_rom[ 6855]='h0000008c;
    rd_cycle[ 6856] = 1'b0;  wr_cycle[ 6856] = 1'b1;  addr_rom[ 6856]='h00000fd0;  wr_data_rom[ 6856]='h0000105c;
    rd_cycle[ 6857] = 1'b0;  wr_cycle[ 6857] = 1'b1;  addr_rom[ 6857]='h00001bd8;  wr_data_rom[ 6857]='h0000159c;
    rd_cycle[ 6858] = 1'b0;  wr_cycle[ 6858] = 1'b1;  addr_rom[ 6858]='h00001610;  wr_data_rom[ 6858]='h000002ee;
    rd_cycle[ 6859] = 1'b1;  wr_cycle[ 6859] = 1'b0;  addr_rom[ 6859]='h00001d10;  wr_data_rom[ 6859]='h00000000;
    rd_cycle[ 6860] = 1'b0;  wr_cycle[ 6860] = 1'b1;  addr_rom[ 6860]='h00000638;  wr_data_rom[ 6860]='h0000057b;
    rd_cycle[ 6861] = 1'b0;  wr_cycle[ 6861] = 1'b1;  addr_rom[ 6861]='h0000022c;  wr_data_rom[ 6861]='h00001632;
    rd_cycle[ 6862] = 1'b0;  wr_cycle[ 6862] = 1'b1;  addr_rom[ 6862]='h00000f80;  wr_data_rom[ 6862]='h00000187;
    rd_cycle[ 6863] = 1'b0;  wr_cycle[ 6863] = 1'b1;  addr_rom[ 6863]='h00001288;  wr_data_rom[ 6863]='h000004a5;
    rd_cycle[ 6864] = 1'b1;  wr_cycle[ 6864] = 1'b0;  addr_rom[ 6864]='h00001d74;  wr_data_rom[ 6864]='h00000000;
    rd_cycle[ 6865] = 1'b0;  wr_cycle[ 6865] = 1'b1;  addr_rom[ 6865]='h000012f8;  wr_data_rom[ 6865]='h00000581;
    rd_cycle[ 6866] = 1'b0;  wr_cycle[ 6866] = 1'b1;  addr_rom[ 6866]='h00001b0c;  wr_data_rom[ 6866]='h00001a0c;
    rd_cycle[ 6867] = 1'b1;  wr_cycle[ 6867] = 1'b0;  addr_rom[ 6867]='h00001c5c;  wr_data_rom[ 6867]='h00000000;
    rd_cycle[ 6868] = 1'b1;  wr_cycle[ 6868] = 1'b0;  addr_rom[ 6868]='h0000014c;  wr_data_rom[ 6868]='h00000000;
    rd_cycle[ 6869] = 1'b1;  wr_cycle[ 6869] = 1'b0;  addr_rom[ 6869]='h00001144;  wr_data_rom[ 6869]='h00000000;
    rd_cycle[ 6870] = 1'b0;  wr_cycle[ 6870] = 1'b1;  addr_rom[ 6870]='h000010f4;  wr_data_rom[ 6870]='h000006ba;
    rd_cycle[ 6871] = 1'b0;  wr_cycle[ 6871] = 1'b1;  addr_rom[ 6871]='h00000508;  wr_data_rom[ 6871]='h000004dd;
    rd_cycle[ 6872] = 1'b0;  wr_cycle[ 6872] = 1'b1;  addr_rom[ 6872]='h00001148;  wr_data_rom[ 6872]='h00000e61;
    rd_cycle[ 6873] = 1'b0;  wr_cycle[ 6873] = 1'b1;  addr_rom[ 6873]='h000015bc;  wr_data_rom[ 6873]='h0000175e;
    rd_cycle[ 6874] = 1'b1;  wr_cycle[ 6874] = 1'b0;  addr_rom[ 6874]='h00000c08;  wr_data_rom[ 6874]='h00000000;
    rd_cycle[ 6875] = 1'b1;  wr_cycle[ 6875] = 1'b0;  addr_rom[ 6875]='h00001040;  wr_data_rom[ 6875]='h00000000;
    rd_cycle[ 6876] = 1'b1;  wr_cycle[ 6876] = 1'b0;  addr_rom[ 6876]='h00000d9c;  wr_data_rom[ 6876]='h00000000;
    rd_cycle[ 6877] = 1'b0;  wr_cycle[ 6877] = 1'b1;  addr_rom[ 6877]='h0000066c;  wr_data_rom[ 6877]='h0000125e;
    rd_cycle[ 6878] = 1'b0;  wr_cycle[ 6878] = 1'b1;  addr_rom[ 6878]='h00001034;  wr_data_rom[ 6878]='h0000099f;
    rd_cycle[ 6879] = 1'b0;  wr_cycle[ 6879] = 1'b1;  addr_rom[ 6879]='h0000119c;  wr_data_rom[ 6879]='h00001269;
    rd_cycle[ 6880] = 1'b0;  wr_cycle[ 6880] = 1'b1;  addr_rom[ 6880]='h00001bfc;  wr_data_rom[ 6880]='h0000093f;
    rd_cycle[ 6881] = 1'b0;  wr_cycle[ 6881] = 1'b1;  addr_rom[ 6881]='h0000147c;  wr_data_rom[ 6881]='h00000d53;
    rd_cycle[ 6882] = 1'b0;  wr_cycle[ 6882] = 1'b1;  addr_rom[ 6882]='h000016b4;  wr_data_rom[ 6882]='h00001918;
    rd_cycle[ 6883] = 1'b1;  wr_cycle[ 6883] = 1'b0;  addr_rom[ 6883]='h000012b8;  wr_data_rom[ 6883]='h00000000;
    rd_cycle[ 6884] = 1'b0;  wr_cycle[ 6884] = 1'b1;  addr_rom[ 6884]='h00000b3c;  wr_data_rom[ 6884]='h0000141b;
    rd_cycle[ 6885] = 1'b0;  wr_cycle[ 6885] = 1'b1;  addr_rom[ 6885]='h000015e8;  wr_data_rom[ 6885]='h0000188e;
    rd_cycle[ 6886] = 1'b0;  wr_cycle[ 6886] = 1'b1;  addr_rom[ 6886]='h00001ab0;  wr_data_rom[ 6886]='h00001223;
    rd_cycle[ 6887] = 1'b0;  wr_cycle[ 6887] = 1'b1;  addr_rom[ 6887]='h000005d8;  wr_data_rom[ 6887]='h00000009;
    rd_cycle[ 6888] = 1'b1;  wr_cycle[ 6888] = 1'b0;  addr_rom[ 6888]='h00001968;  wr_data_rom[ 6888]='h00000000;
    rd_cycle[ 6889] = 1'b1;  wr_cycle[ 6889] = 1'b0;  addr_rom[ 6889]='h000004fc;  wr_data_rom[ 6889]='h00000000;
    rd_cycle[ 6890] = 1'b1;  wr_cycle[ 6890] = 1'b0;  addr_rom[ 6890]='h00000808;  wr_data_rom[ 6890]='h00000000;
    rd_cycle[ 6891] = 1'b0;  wr_cycle[ 6891] = 1'b1;  addr_rom[ 6891]='h00000414;  wr_data_rom[ 6891]='h00000c48;
    rd_cycle[ 6892] = 1'b1;  wr_cycle[ 6892] = 1'b0;  addr_rom[ 6892]='h00000dd4;  wr_data_rom[ 6892]='h00000000;
    rd_cycle[ 6893] = 1'b1;  wr_cycle[ 6893] = 1'b0;  addr_rom[ 6893]='h00000698;  wr_data_rom[ 6893]='h00000000;
    rd_cycle[ 6894] = 1'b0;  wr_cycle[ 6894] = 1'b1;  addr_rom[ 6894]='h00001118;  wr_data_rom[ 6894]='h000015fb;
    rd_cycle[ 6895] = 1'b0;  wr_cycle[ 6895] = 1'b1;  addr_rom[ 6895]='h000017ac;  wr_data_rom[ 6895]='h000018c0;
    rd_cycle[ 6896] = 1'b1;  wr_cycle[ 6896] = 1'b0;  addr_rom[ 6896]='h00001db8;  wr_data_rom[ 6896]='h00000000;
    rd_cycle[ 6897] = 1'b1;  wr_cycle[ 6897] = 1'b0;  addr_rom[ 6897]='h00001b74;  wr_data_rom[ 6897]='h00000000;
    rd_cycle[ 6898] = 1'b1;  wr_cycle[ 6898] = 1'b0;  addr_rom[ 6898]='h00000b8c;  wr_data_rom[ 6898]='h00000000;
    rd_cycle[ 6899] = 1'b1;  wr_cycle[ 6899] = 1'b0;  addr_rom[ 6899]='h0000109c;  wr_data_rom[ 6899]='h00000000;
    rd_cycle[ 6900] = 1'b1;  wr_cycle[ 6900] = 1'b0;  addr_rom[ 6900]='h00001030;  wr_data_rom[ 6900]='h00000000;
    rd_cycle[ 6901] = 1'b1;  wr_cycle[ 6901] = 1'b0;  addr_rom[ 6901]='h00001b08;  wr_data_rom[ 6901]='h00000000;
    rd_cycle[ 6902] = 1'b0;  wr_cycle[ 6902] = 1'b1;  addr_rom[ 6902]='h00001108;  wr_data_rom[ 6902]='h000000dd;
    rd_cycle[ 6903] = 1'b1;  wr_cycle[ 6903] = 1'b0;  addr_rom[ 6903]='h00001624;  wr_data_rom[ 6903]='h00000000;
    rd_cycle[ 6904] = 1'b1;  wr_cycle[ 6904] = 1'b0;  addr_rom[ 6904]='h0000068c;  wr_data_rom[ 6904]='h00000000;
    rd_cycle[ 6905] = 1'b0;  wr_cycle[ 6905] = 1'b1;  addr_rom[ 6905]='h000017f4;  wr_data_rom[ 6905]='h000001b3;
    rd_cycle[ 6906] = 1'b0;  wr_cycle[ 6906] = 1'b1;  addr_rom[ 6906]='h00000e04;  wr_data_rom[ 6906]='h00001ae3;
    rd_cycle[ 6907] = 1'b1;  wr_cycle[ 6907] = 1'b0;  addr_rom[ 6907]='h00001e2c;  wr_data_rom[ 6907]='h00000000;
    rd_cycle[ 6908] = 1'b0;  wr_cycle[ 6908] = 1'b1;  addr_rom[ 6908]='h00000600;  wr_data_rom[ 6908]='h00000251;
    rd_cycle[ 6909] = 1'b0;  wr_cycle[ 6909] = 1'b1;  addr_rom[ 6909]='h0000146c;  wr_data_rom[ 6909]='h000002c4;
    rd_cycle[ 6910] = 1'b0;  wr_cycle[ 6910] = 1'b1;  addr_rom[ 6910]='h00000c38;  wr_data_rom[ 6910]='h0000195d;
    rd_cycle[ 6911] = 1'b0;  wr_cycle[ 6911] = 1'b1;  addr_rom[ 6911]='h000019f4;  wr_data_rom[ 6911]='h0000006c;
    rd_cycle[ 6912] = 1'b1;  wr_cycle[ 6912] = 1'b0;  addr_rom[ 6912]='h00001670;  wr_data_rom[ 6912]='h00000000;
    rd_cycle[ 6913] = 1'b1;  wr_cycle[ 6913] = 1'b0;  addr_rom[ 6913]='h00000a40;  wr_data_rom[ 6913]='h00000000;
    rd_cycle[ 6914] = 1'b1;  wr_cycle[ 6914] = 1'b0;  addr_rom[ 6914]='h000004fc;  wr_data_rom[ 6914]='h00000000;
    rd_cycle[ 6915] = 1'b0;  wr_cycle[ 6915] = 1'b1;  addr_rom[ 6915]='h00000644;  wr_data_rom[ 6915]='h00001278;
    rd_cycle[ 6916] = 1'b1;  wr_cycle[ 6916] = 1'b0;  addr_rom[ 6916]='h00001044;  wr_data_rom[ 6916]='h00000000;
    rd_cycle[ 6917] = 1'b1;  wr_cycle[ 6917] = 1'b0;  addr_rom[ 6917]='h00000494;  wr_data_rom[ 6917]='h00000000;
    rd_cycle[ 6918] = 1'b1;  wr_cycle[ 6918] = 1'b0;  addr_rom[ 6918]='h000007f4;  wr_data_rom[ 6918]='h00000000;
    rd_cycle[ 6919] = 1'b1;  wr_cycle[ 6919] = 1'b0;  addr_rom[ 6919]='h000012ac;  wr_data_rom[ 6919]='h00000000;
    rd_cycle[ 6920] = 1'b0;  wr_cycle[ 6920] = 1'b1;  addr_rom[ 6920]='h00000958;  wr_data_rom[ 6920]='h000019b5;
    rd_cycle[ 6921] = 1'b1;  wr_cycle[ 6921] = 1'b0;  addr_rom[ 6921]='h00000234;  wr_data_rom[ 6921]='h00000000;
    rd_cycle[ 6922] = 1'b1;  wr_cycle[ 6922] = 1'b0;  addr_rom[ 6922]='h00000874;  wr_data_rom[ 6922]='h00000000;
    rd_cycle[ 6923] = 1'b1;  wr_cycle[ 6923] = 1'b0;  addr_rom[ 6923]='h00000600;  wr_data_rom[ 6923]='h00000000;
    rd_cycle[ 6924] = 1'b1;  wr_cycle[ 6924] = 1'b0;  addr_rom[ 6924]='h00000918;  wr_data_rom[ 6924]='h00000000;
    rd_cycle[ 6925] = 1'b1;  wr_cycle[ 6925] = 1'b0;  addr_rom[ 6925]='h00001540;  wr_data_rom[ 6925]='h00000000;
    rd_cycle[ 6926] = 1'b0;  wr_cycle[ 6926] = 1'b1;  addr_rom[ 6926]='h00000d08;  wr_data_rom[ 6926]='h00000dd8;
    rd_cycle[ 6927] = 1'b0;  wr_cycle[ 6927] = 1'b1;  addr_rom[ 6927]='h00000718;  wr_data_rom[ 6927]='h0000022c;
    rd_cycle[ 6928] = 1'b1;  wr_cycle[ 6928] = 1'b0;  addr_rom[ 6928]='h00001b28;  wr_data_rom[ 6928]='h00000000;
    rd_cycle[ 6929] = 1'b1;  wr_cycle[ 6929] = 1'b0;  addr_rom[ 6929]='h000014e0;  wr_data_rom[ 6929]='h00000000;
    rd_cycle[ 6930] = 1'b0;  wr_cycle[ 6930] = 1'b1;  addr_rom[ 6930]='h0000035c;  wr_data_rom[ 6930]='h000013d4;
    rd_cycle[ 6931] = 1'b1;  wr_cycle[ 6931] = 1'b0;  addr_rom[ 6931]='h000011b8;  wr_data_rom[ 6931]='h00000000;
    rd_cycle[ 6932] = 1'b1;  wr_cycle[ 6932] = 1'b0;  addr_rom[ 6932]='h000008f8;  wr_data_rom[ 6932]='h00000000;
    rd_cycle[ 6933] = 1'b1;  wr_cycle[ 6933] = 1'b0;  addr_rom[ 6933]='h00001c6c;  wr_data_rom[ 6933]='h00000000;
    rd_cycle[ 6934] = 1'b0;  wr_cycle[ 6934] = 1'b1;  addr_rom[ 6934]='h00000f60;  wr_data_rom[ 6934]='h00001358;
    rd_cycle[ 6935] = 1'b1;  wr_cycle[ 6935] = 1'b0;  addr_rom[ 6935]='h000016d0;  wr_data_rom[ 6935]='h00000000;
    rd_cycle[ 6936] = 1'b0;  wr_cycle[ 6936] = 1'b1;  addr_rom[ 6936]='h000011ec;  wr_data_rom[ 6936]='h00001e87;
    rd_cycle[ 6937] = 1'b0;  wr_cycle[ 6937] = 1'b1;  addr_rom[ 6937]='h00000008;  wr_data_rom[ 6937]='h00001650;
    rd_cycle[ 6938] = 1'b1;  wr_cycle[ 6938] = 1'b0;  addr_rom[ 6938]='h0000190c;  wr_data_rom[ 6938]='h00000000;
    rd_cycle[ 6939] = 1'b1;  wr_cycle[ 6939] = 1'b0;  addr_rom[ 6939]='h000007d0;  wr_data_rom[ 6939]='h00000000;
    rd_cycle[ 6940] = 1'b0;  wr_cycle[ 6940] = 1'b1;  addr_rom[ 6940]='h00001638;  wr_data_rom[ 6940]='h0000080b;
    rd_cycle[ 6941] = 1'b1;  wr_cycle[ 6941] = 1'b0;  addr_rom[ 6941]='h0000044c;  wr_data_rom[ 6941]='h00000000;
    rd_cycle[ 6942] = 1'b0;  wr_cycle[ 6942] = 1'b1;  addr_rom[ 6942]='h0000079c;  wr_data_rom[ 6942]='h000012a9;
    rd_cycle[ 6943] = 1'b0;  wr_cycle[ 6943] = 1'b1;  addr_rom[ 6943]='h00000ef4;  wr_data_rom[ 6943]='h000009dd;
    rd_cycle[ 6944] = 1'b1;  wr_cycle[ 6944] = 1'b0;  addr_rom[ 6944]='h000014a0;  wr_data_rom[ 6944]='h00000000;
    rd_cycle[ 6945] = 1'b1;  wr_cycle[ 6945] = 1'b0;  addr_rom[ 6945]='h000004c8;  wr_data_rom[ 6945]='h00000000;
    rd_cycle[ 6946] = 1'b0;  wr_cycle[ 6946] = 1'b1;  addr_rom[ 6946]='h0000109c;  wr_data_rom[ 6946]='h00001d67;
    rd_cycle[ 6947] = 1'b0;  wr_cycle[ 6947] = 1'b1;  addr_rom[ 6947]='h00000620;  wr_data_rom[ 6947]='h000011b1;
    rd_cycle[ 6948] = 1'b0;  wr_cycle[ 6948] = 1'b1;  addr_rom[ 6948]='h00001b68;  wr_data_rom[ 6948]='h00000cab;
    rd_cycle[ 6949] = 1'b1;  wr_cycle[ 6949] = 1'b0;  addr_rom[ 6949]='h00000d78;  wr_data_rom[ 6949]='h00000000;
    rd_cycle[ 6950] = 1'b1;  wr_cycle[ 6950] = 1'b0;  addr_rom[ 6950]='h000019c0;  wr_data_rom[ 6950]='h00000000;
    rd_cycle[ 6951] = 1'b0;  wr_cycle[ 6951] = 1'b1;  addr_rom[ 6951]='h0000078c;  wr_data_rom[ 6951]='h00000ac5;
    rd_cycle[ 6952] = 1'b1;  wr_cycle[ 6952] = 1'b0;  addr_rom[ 6952]='h000019b4;  wr_data_rom[ 6952]='h00000000;
    rd_cycle[ 6953] = 1'b1;  wr_cycle[ 6953] = 1'b0;  addr_rom[ 6953]='h000016a4;  wr_data_rom[ 6953]='h00000000;
    rd_cycle[ 6954] = 1'b1;  wr_cycle[ 6954] = 1'b0;  addr_rom[ 6954]='h00001050;  wr_data_rom[ 6954]='h00000000;
    rd_cycle[ 6955] = 1'b1;  wr_cycle[ 6955] = 1'b0;  addr_rom[ 6955]='h00001b20;  wr_data_rom[ 6955]='h00000000;
    rd_cycle[ 6956] = 1'b0;  wr_cycle[ 6956] = 1'b1;  addr_rom[ 6956]='h00001014;  wr_data_rom[ 6956]='h00001a5a;
    rd_cycle[ 6957] = 1'b1;  wr_cycle[ 6957] = 1'b0;  addr_rom[ 6957]='h00000e04;  wr_data_rom[ 6957]='h00000000;
    rd_cycle[ 6958] = 1'b1;  wr_cycle[ 6958] = 1'b0;  addr_rom[ 6958]='h00001864;  wr_data_rom[ 6958]='h00000000;
    rd_cycle[ 6959] = 1'b1;  wr_cycle[ 6959] = 1'b0;  addr_rom[ 6959]='h00000f20;  wr_data_rom[ 6959]='h00000000;
    rd_cycle[ 6960] = 1'b1;  wr_cycle[ 6960] = 1'b0;  addr_rom[ 6960]='h00000b28;  wr_data_rom[ 6960]='h00000000;
    rd_cycle[ 6961] = 1'b0;  wr_cycle[ 6961] = 1'b1;  addr_rom[ 6961]='h00000698;  wr_data_rom[ 6961]='h000005ce;
    rd_cycle[ 6962] = 1'b1;  wr_cycle[ 6962] = 1'b0;  addr_rom[ 6962]='h00001538;  wr_data_rom[ 6962]='h00000000;
    rd_cycle[ 6963] = 1'b1;  wr_cycle[ 6963] = 1'b0;  addr_rom[ 6963]='h000003ec;  wr_data_rom[ 6963]='h00000000;
    rd_cycle[ 6964] = 1'b1;  wr_cycle[ 6964] = 1'b0;  addr_rom[ 6964]='h0000009c;  wr_data_rom[ 6964]='h00000000;
    rd_cycle[ 6965] = 1'b1;  wr_cycle[ 6965] = 1'b0;  addr_rom[ 6965]='h00000340;  wr_data_rom[ 6965]='h00000000;
    rd_cycle[ 6966] = 1'b0;  wr_cycle[ 6966] = 1'b1;  addr_rom[ 6966]='h00001218;  wr_data_rom[ 6966]='h00000acc;
    rd_cycle[ 6967] = 1'b1;  wr_cycle[ 6967] = 1'b0;  addr_rom[ 6967]='h00000d20;  wr_data_rom[ 6967]='h00000000;
    rd_cycle[ 6968] = 1'b1;  wr_cycle[ 6968] = 1'b0;  addr_rom[ 6968]='h00000754;  wr_data_rom[ 6968]='h00000000;
    rd_cycle[ 6969] = 1'b0;  wr_cycle[ 6969] = 1'b1;  addr_rom[ 6969]='h000014c4;  wr_data_rom[ 6969]='h000004ad;
    rd_cycle[ 6970] = 1'b1;  wr_cycle[ 6970] = 1'b0;  addr_rom[ 6970]='h0000051c;  wr_data_rom[ 6970]='h00000000;
    rd_cycle[ 6971] = 1'b0;  wr_cycle[ 6971] = 1'b1;  addr_rom[ 6971]='h00000960;  wr_data_rom[ 6971]='h00001c64;
    rd_cycle[ 6972] = 1'b1;  wr_cycle[ 6972] = 1'b0;  addr_rom[ 6972]='h00000fd8;  wr_data_rom[ 6972]='h00000000;
    rd_cycle[ 6973] = 1'b0;  wr_cycle[ 6973] = 1'b1;  addr_rom[ 6973]='h000010b8;  wr_data_rom[ 6973]='h00001783;
    rd_cycle[ 6974] = 1'b1;  wr_cycle[ 6974] = 1'b0;  addr_rom[ 6974]='h00001980;  wr_data_rom[ 6974]='h00000000;
    rd_cycle[ 6975] = 1'b0;  wr_cycle[ 6975] = 1'b1;  addr_rom[ 6975]='h00000654;  wr_data_rom[ 6975]='h000001ec;
    rd_cycle[ 6976] = 1'b1;  wr_cycle[ 6976] = 1'b0;  addr_rom[ 6976]='h0000187c;  wr_data_rom[ 6976]='h00000000;
    rd_cycle[ 6977] = 1'b0;  wr_cycle[ 6977] = 1'b1;  addr_rom[ 6977]='h0000189c;  wr_data_rom[ 6977]='h00000578;
    rd_cycle[ 6978] = 1'b0;  wr_cycle[ 6978] = 1'b1;  addr_rom[ 6978]='h00001828;  wr_data_rom[ 6978]='h0000048c;
    rd_cycle[ 6979] = 1'b0;  wr_cycle[ 6979] = 1'b1;  addr_rom[ 6979]='h000008e8;  wr_data_rom[ 6979]='h0000056e;
    rd_cycle[ 6980] = 1'b0;  wr_cycle[ 6980] = 1'b1;  addr_rom[ 6980]='h00001788;  wr_data_rom[ 6980]='h00001871;
    rd_cycle[ 6981] = 1'b0;  wr_cycle[ 6981] = 1'b1;  addr_rom[ 6981]='h000015c0;  wr_data_rom[ 6981]='h00001890;
    rd_cycle[ 6982] = 1'b1;  wr_cycle[ 6982] = 1'b0;  addr_rom[ 6982]='h000003a0;  wr_data_rom[ 6982]='h00000000;
    rd_cycle[ 6983] = 1'b1;  wr_cycle[ 6983] = 1'b0;  addr_rom[ 6983]='h00001bf8;  wr_data_rom[ 6983]='h00000000;
    rd_cycle[ 6984] = 1'b1;  wr_cycle[ 6984] = 1'b0;  addr_rom[ 6984]='h00001a80;  wr_data_rom[ 6984]='h00000000;
    rd_cycle[ 6985] = 1'b0;  wr_cycle[ 6985] = 1'b1;  addr_rom[ 6985]='h00000820;  wr_data_rom[ 6985]='h000011ae;
    rd_cycle[ 6986] = 1'b1;  wr_cycle[ 6986] = 1'b0;  addr_rom[ 6986]='h00001a28;  wr_data_rom[ 6986]='h00000000;
    rd_cycle[ 6987] = 1'b0;  wr_cycle[ 6987] = 1'b1;  addr_rom[ 6987]='h00001530;  wr_data_rom[ 6987]='h00000d7a;
    rd_cycle[ 6988] = 1'b0;  wr_cycle[ 6988] = 1'b1;  addr_rom[ 6988]='h00000208;  wr_data_rom[ 6988]='h0000185e;
    rd_cycle[ 6989] = 1'b0;  wr_cycle[ 6989] = 1'b1;  addr_rom[ 6989]='h00000894;  wr_data_rom[ 6989]='h00000226;
    rd_cycle[ 6990] = 1'b1;  wr_cycle[ 6990] = 1'b0;  addr_rom[ 6990]='h000015a0;  wr_data_rom[ 6990]='h00000000;
    rd_cycle[ 6991] = 1'b1;  wr_cycle[ 6991] = 1'b0;  addr_rom[ 6991]='h00000a44;  wr_data_rom[ 6991]='h00000000;
    rd_cycle[ 6992] = 1'b0;  wr_cycle[ 6992] = 1'b1;  addr_rom[ 6992]='h00001018;  wr_data_rom[ 6992]='h00000537;
    rd_cycle[ 6993] = 1'b0;  wr_cycle[ 6993] = 1'b1;  addr_rom[ 6993]='h00000eb8;  wr_data_rom[ 6993]='h0000138e;
    rd_cycle[ 6994] = 1'b0;  wr_cycle[ 6994] = 1'b1;  addr_rom[ 6994]='h0000155c;  wr_data_rom[ 6994]='h000015d0;
    rd_cycle[ 6995] = 1'b0;  wr_cycle[ 6995] = 1'b1;  addr_rom[ 6995]='h00001af4;  wr_data_rom[ 6995]='h000013fd;
    rd_cycle[ 6996] = 1'b1;  wr_cycle[ 6996] = 1'b0;  addr_rom[ 6996]='h00000ac0;  wr_data_rom[ 6996]='h00000000;
    rd_cycle[ 6997] = 1'b0;  wr_cycle[ 6997] = 1'b1;  addr_rom[ 6997]='h00000e14;  wr_data_rom[ 6997]='h0000029a;
    rd_cycle[ 6998] = 1'b1;  wr_cycle[ 6998] = 1'b0;  addr_rom[ 6998]='h00001b54;  wr_data_rom[ 6998]='h00000000;
    rd_cycle[ 6999] = 1'b0;  wr_cycle[ 6999] = 1'b1;  addr_rom[ 6999]='h00000794;  wr_data_rom[ 6999]='h00000532;
    rd_cycle[ 7000] = 1'b1;  wr_cycle[ 7000] = 1'b0;  addr_rom[ 7000]='h0000174c;  wr_data_rom[ 7000]='h00000000;
    rd_cycle[ 7001] = 1'b1;  wr_cycle[ 7001] = 1'b0;  addr_rom[ 7001]='h00001020;  wr_data_rom[ 7001]='h00000000;
    rd_cycle[ 7002] = 1'b0;  wr_cycle[ 7002] = 1'b1;  addr_rom[ 7002]='h0000138c;  wr_data_rom[ 7002]='h0000071c;
    rd_cycle[ 7003] = 1'b0;  wr_cycle[ 7003] = 1'b1;  addr_rom[ 7003]='h00001758;  wr_data_rom[ 7003]='h00000f62;
    rd_cycle[ 7004] = 1'b0;  wr_cycle[ 7004] = 1'b1;  addr_rom[ 7004]='h00001bd4;  wr_data_rom[ 7004]='h00001928;
    rd_cycle[ 7005] = 1'b1;  wr_cycle[ 7005] = 1'b0;  addr_rom[ 7005]='h00000d98;  wr_data_rom[ 7005]='h00000000;
    rd_cycle[ 7006] = 1'b0;  wr_cycle[ 7006] = 1'b1;  addr_rom[ 7006]='h00000fa8;  wr_data_rom[ 7006]='h00000f42;
    rd_cycle[ 7007] = 1'b0;  wr_cycle[ 7007] = 1'b1;  addr_rom[ 7007]='h0000158c;  wr_data_rom[ 7007]='h00000ae8;
    rd_cycle[ 7008] = 1'b1;  wr_cycle[ 7008] = 1'b0;  addr_rom[ 7008]='h00000604;  wr_data_rom[ 7008]='h00000000;
    rd_cycle[ 7009] = 1'b0;  wr_cycle[ 7009] = 1'b1;  addr_rom[ 7009]='h000002dc;  wr_data_rom[ 7009]='h000004d5;
    rd_cycle[ 7010] = 1'b1;  wr_cycle[ 7010] = 1'b0;  addr_rom[ 7010]='h00000b30;  wr_data_rom[ 7010]='h00000000;
    rd_cycle[ 7011] = 1'b1;  wr_cycle[ 7011] = 1'b0;  addr_rom[ 7011]='h00000688;  wr_data_rom[ 7011]='h00000000;
    rd_cycle[ 7012] = 1'b0;  wr_cycle[ 7012] = 1'b1;  addr_rom[ 7012]='h00000d88;  wr_data_rom[ 7012]='h00000f1b;
    rd_cycle[ 7013] = 1'b1;  wr_cycle[ 7013] = 1'b0;  addr_rom[ 7013]='h00000d38;  wr_data_rom[ 7013]='h00000000;
    rd_cycle[ 7014] = 1'b0;  wr_cycle[ 7014] = 1'b1;  addr_rom[ 7014]='h00000e24;  wr_data_rom[ 7014]='h00001e76;
    rd_cycle[ 7015] = 1'b0;  wr_cycle[ 7015] = 1'b1;  addr_rom[ 7015]='h00000c38;  wr_data_rom[ 7015]='h00001a2f;
    rd_cycle[ 7016] = 1'b1;  wr_cycle[ 7016] = 1'b0;  addr_rom[ 7016]='h0000087c;  wr_data_rom[ 7016]='h00000000;
    rd_cycle[ 7017] = 1'b0;  wr_cycle[ 7017] = 1'b1;  addr_rom[ 7017]='h000010ec;  wr_data_rom[ 7017]='h000007cc;
    rd_cycle[ 7018] = 1'b1;  wr_cycle[ 7018] = 1'b0;  addr_rom[ 7018]='h00001288;  wr_data_rom[ 7018]='h00000000;
    rd_cycle[ 7019] = 1'b0;  wr_cycle[ 7019] = 1'b1;  addr_rom[ 7019]='h00000420;  wr_data_rom[ 7019]='h00001ebf;
    rd_cycle[ 7020] = 1'b1;  wr_cycle[ 7020] = 1'b0;  addr_rom[ 7020]='h00000b78;  wr_data_rom[ 7020]='h00000000;
    rd_cycle[ 7021] = 1'b1;  wr_cycle[ 7021] = 1'b0;  addr_rom[ 7021]='h00000f44;  wr_data_rom[ 7021]='h00000000;
    rd_cycle[ 7022] = 1'b0;  wr_cycle[ 7022] = 1'b1;  addr_rom[ 7022]='h00001774;  wr_data_rom[ 7022]='h00000f15;
    rd_cycle[ 7023] = 1'b0;  wr_cycle[ 7023] = 1'b1;  addr_rom[ 7023]='h00000e74;  wr_data_rom[ 7023]='h00001359;
    rd_cycle[ 7024] = 1'b0;  wr_cycle[ 7024] = 1'b1;  addr_rom[ 7024]='h00000ad8;  wr_data_rom[ 7024]='h000010a7;
    rd_cycle[ 7025] = 1'b1;  wr_cycle[ 7025] = 1'b0;  addr_rom[ 7025]='h0000025c;  wr_data_rom[ 7025]='h00000000;
    rd_cycle[ 7026] = 1'b0;  wr_cycle[ 7026] = 1'b1;  addr_rom[ 7026]='h00000724;  wr_data_rom[ 7026]='h00000db4;
    rd_cycle[ 7027] = 1'b0;  wr_cycle[ 7027] = 1'b1;  addr_rom[ 7027]='h00000c48;  wr_data_rom[ 7027]='h000004b9;
    rd_cycle[ 7028] = 1'b0;  wr_cycle[ 7028] = 1'b1;  addr_rom[ 7028]='h0000039c;  wr_data_rom[ 7028]='h00000238;
    rd_cycle[ 7029] = 1'b1;  wr_cycle[ 7029] = 1'b0;  addr_rom[ 7029]='h00001590;  wr_data_rom[ 7029]='h00000000;
    rd_cycle[ 7030] = 1'b1;  wr_cycle[ 7030] = 1'b0;  addr_rom[ 7030]='h000005e4;  wr_data_rom[ 7030]='h00000000;
    rd_cycle[ 7031] = 1'b1;  wr_cycle[ 7031] = 1'b0;  addr_rom[ 7031]='h000012a0;  wr_data_rom[ 7031]='h00000000;
    rd_cycle[ 7032] = 1'b1;  wr_cycle[ 7032] = 1'b0;  addr_rom[ 7032]='h0000087c;  wr_data_rom[ 7032]='h00000000;
    rd_cycle[ 7033] = 1'b1;  wr_cycle[ 7033] = 1'b0;  addr_rom[ 7033]='h000003cc;  wr_data_rom[ 7033]='h00000000;
    rd_cycle[ 7034] = 1'b0;  wr_cycle[ 7034] = 1'b1;  addr_rom[ 7034]='h000009d8;  wr_data_rom[ 7034]='h00000cf2;
    rd_cycle[ 7035] = 1'b1;  wr_cycle[ 7035] = 1'b0;  addr_rom[ 7035]='h000000d0;  wr_data_rom[ 7035]='h00000000;
    rd_cycle[ 7036] = 1'b0;  wr_cycle[ 7036] = 1'b1;  addr_rom[ 7036]='h0000091c;  wr_data_rom[ 7036]='h00000ce2;
    rd_cycle[ 7037] = 1'b0;  wr_cycle[ 7037] = 1'b1;  addr_rom[ 7037]='h00001554;  wr_data_rom[ 7037]='h00000245;
    rd_cycle[ 7038] = 1'b0;  wr_cycle[ 7038] = 1'b1;  addr_rom[ 7038]='h00001e24;  wr_data_rom[ 7038]='h00001a53;
    rd_cycle[ 7039] = 1'b1;  wr_cycle[ 7039] = 1'b0;  addr_rom[ 7039]='h0000004c;  wr_data_rom[ 7039]='h00000000;
    rd_cycle[ 7040] = 1'b1;  wr_cycle[ 7040] = 1'b0;  addr_rom[ 7040]='h00000c04;  wr_data_rom[ 7040]='h00000000;
    rd_cycle[ 7041] = 1'b1;  wr_cycle[ 7041] = 1'b0;  addr_rom[ 7041]='h00000bc4;  wr_data_rom[ 7041]='h00000000;
    rd_cycle[ 7042] = 1'b1;  wr_cycle[ 7042] = 1'b0;  addr_rom[ 7042]='h00001174;  wr_data_rom[ 7042]='h00000000;
    rd_cycle[ 7043] = 1'b1;  wr_cycle[ 7043] = 1'b0;  addr_rom[ 7043]='h00001eac;  wr_data_rom[ 7043]='h00000000;
    rd_cycle[ 7044] = 1'b0;  wr_cycle[ 7044] = 1'b1;  addr_rom[ 7044]='h00001708;  wr_data_rom[ 7044]='h000011cd;
    rd_cycle[ 7045] = 1'b0;  wr_cycle[ 7045] = 1'b1;  addr_rom[ 7045]='h0000101c;  wr_data_rom[ 7045]='h00001bfc;
    rd_cycle[ 7046] = 1'b1;  wr_cycle[ 7046] = 1'b0;  addr_rom[ 7046]='h00001798;  wr_data_rom[ 7046]='h00000000;
    rd_cycle[ 7047] = 1'b0;  wr_cycle[ 7047] = 1'b1;  addr_rom[ 7047]='h00000aac;  wr_data_rom[ 7047]='h00000ddc;
    rd_cycle[ 7048] = 1'b1;  wr_cycle[ 7048] = 1'b0;  addr_rom[ 7048]='h00000c60;  wr_data_rom[ 7048]='h00000000;
    rd_cycle[ 7049] = 1'b0;  wr_cycle[ 7049] = 1'b1;  addr_rom[ 7049]='h000002b8;  wr_data_rom[ 7049]='h00000261;
    rd_cycle[ 7050] = 1'b0;  wr_cycle[ 7050] = 1'b1;  addr_rom[ 7050]='h00001900;  wr_data_rom[ 7050]='h0000076d;
    rd_cycle[ 7051] = 1'b0;  wr_cycle[ 7051] = 1'b1;  addr_rom[ 7051]='h000008d8;  wr_data_rom[ 7051]='h00001df3;
    rd_cycle[ 7052] = 1'b1;  wr_cycle[ 7052] = 1'b0;  addr_rom[ 7052]='h00000584;  wr_data_rom[ 7052]='h00000000;
    rd_cycle[ 7053] = 1'b1;  wr_cycle[ 7053] = 1'b0;  addr_rom[ 7053]='h00000c60;  wr_data_rom[ 7053]='h00000000;
    rd_cycle[ 7054] = 1'b1;  wr_cycle[ 7054] = 1'b0;  addr_rom[ 7054]='h00001e8c;  wr_data_rom[ 7054]='h00000000;
    rd_cycle[ 7055] = 1'b1;  wr_cycle[ 7055] = 1'b0;  addr_rom[ 7055]='h00000014;  wr_data_rom[ 7055]='h00000000;
    rd_cycle[ 7056] = 1'b1;  wr_cycle[ 7056] = 1'b0;  addr_rom[ 7056]='h000014a0;  wr_data_rom[ 7056]='h00000000;
    rd_cycle[ 7057] = 1'b1;  wr_cycle[ 7057] = 1'b0;  addr_rom[ 7057]='h00001944;  wr_data_rom[ 7057]='h00000000;
    rd_cycle[ 7058] = 1'b0;  wr_cycle[ 7058] = 1'b1;  addr_rom[ 7058]='h00001278;  wr_data_rom[ 7058]='h000005b6;
    rd_cycle[ 7059] = 1'b0;  wr_cycle[ 7059] = 1'b1;  addr_rom[ 7059]='h00000c7c;  wr_data_rom[ 7059]='h00000817;
    rd_cycle[ 7060] = 1'b1;  wr_cycle[ 7060] = 1'b0;  addr_rom[ 7060]='h0000176c;  wr_data_rom[ 7060]='h00000000;
    rd_cycle[ 7061] = 1'b1;  wr_cycle[ 7061] = 1'b0;  addr_rom[ 7061]='h00001844;  wr_data_rom[ 7061]='h00000000;
    rd_cycle[ 7062] = 1'b1;  wr_cycle[ 7062] = 1'b0;  addr_rom[ 7062]='h00001d28;  wr_data_rom[ 7062]='h00000000;
    rd_cycle[ 7063] = 1'b1;  wr_cycle[ 7063] = 1'b0;  addr_rom[ 7063]='h000005b8;  wr_data_rom[ 7063]='h00000000;
    rd_cycle[ 7064] = 1'b1;  wr_cycle[ 7064] = 1'b0;  addr_rom[ 7064]='h00001164;  wr_data_rom[ 7064]='h00000000;
    rd_cycle[ 7065] = 1'b0;  wr_cycle[ 7065] = 1'b1;  addr_rom[ 7065]='h0000177c;  wr_data_rom[ 7065]='h00001d3a;
    rd_cycle[ 7066] = 1'b1;  wr_cycle[ 7066] = 1'b0;  addr_rom[ 7066]='h00000874;  wr_data_rom[ 7066]='h00000000;
    rd_cycle[ 7067] = 1'b1;  wr_cycle[ 7067] = 1'b0;  addr_rom[ 7067]='h0000024c;  wr_data_rom[ 7067]='h00000000;
    rd_cycle[ 7068] = 1'b1;  wr_cycle[ 7068] = 1'b0;  addr_rom[ 7068]='h000013e0;  wr_data_rom[ 7068]='h00000000;
    rd_cycle[ 7069] = 1'b0;  wr_cycle[ 7069] = 1'b1;  addr_rom[ 7069]='h00001c68;  wr_data_rom[ 7069]='h000008e4;
    rd_cycle[ 7070] = 1'b1;  wr_cycle[ 7070] = 1'b0;  addr_rom[ 7070]='h00001898;  wr_data_rom[ 7070]='h00000000;
    rd_cycle[ 7071] = 1'b0;  wr_cycle[ 7071] = 1'b1;  addr_rom[ 7071]='h000001b8;  wr_data_rom[ 7071]='h00000ae3;
    rd_cycle[ 7072] = 1'b1;  wr_cycle[ 7072] = 1'b0;  addr_rom[ 7072]='h00000070;  wr_data_rom[ 7072]='h00000000;
    rd_cycle[ 7073] = 1'b1;  wr_cycle[ 7073] = 1'b0;  addr_rom[ 7073]='h00000678;  wr_data_rom[ 7073]='h00000000;
    rd_cycle[ 7074] = 1'b0;  wr_cycle[ 7074] = 1'b1;  addr_rom[ 7074]='h000018f8;  wr_data_rom[ 7074]='h00000d99;
    rd_cycle[ 7075] = 1'b1;  wr_cycle[ 7075] = 1'b0;  addr_rom[ 7075]='h0000103c;  wr_data_rom[ 7075]='h00000000;
    rd_cycle[ 7076] = 1'b1;  wr_cycle[ 7076] = 1'b0;  addr_rom[ 7076]='h000014c0;  wr_data_rom[ 7076]='h00000000;
    rd_cycle[ 7077] = 1'b0;  wr_cycle[ 7077] = 1'b1;  addr_rom[ 7077]='h00000c70;  wr_data_rom[ 7077]='h0000015d;
    rd_cycle[ 7078] = 1'b0;  wr_cycle[ 7078] = 1'b1;  addr_rom[ 7078]='h00001134;  wr_data_rom[ 7078]='h00000834;
    rd_cycle[ 7079] = 1'b0;  wr_cycle[ 7079] = 1'b1;  addr_rom[ 7079]='h000000b4;  wr_data_rom[ 7079]='h00000ede;
    rd_cycle[ 7080] = 1'b1;  wr_cycle[ 7080] = 1'b0;  addr_rom[ 7080]='h000011f8;  wr_data_rom[ 7080]='h00000000;
    rd_cycle[ 7081] = 1'b1;  wr_cycle[ 7081] = 1'b0;  addr_rom[ 7081]='h00001338;  wr_data_rom[ 7081]='h00000000;
    rd_cycle[ 7082] = 1'b1;  wr_cycle[ 7082] = 1'b0;  addr_rom[ 7082]='h00001528;  wr_data_rom[ 7082]='h00000000;
    rd_cycle[ 7083] = 1'b0;  wr_cycle[ 7083] = 1'b1;  addr_rom[ 7083]='h000003c4;  wr_data_rom[ 7083]='h000005fd;
    rd_cycle[ 7084] = 1'b0;  wr_cycle[ 7084] = 1'b1;  addr_rom[ 7084]='h00000a60;  wr_data_rom[ 7084]='h000003e1;
    rd_cycle[ 7085] = 1'b1;  wr_cycle[ 7085] = 1'b0;  addr_rom[ 7085]='h000013b0;  wr_data_rom[ 7085]='h00000000;
    rd_cycle[ 7086] = 1'b1;  wr_cycle[ 7086] = 1'b0;  addr_rom[ 7086]='h00000b20;  wr_data_rom[ 7086]='h00000000;
    rd_cycle[ 7087] = 1'b1;  wr_cycle[ 7087] = 1'b0;  addr_rom[ 7087]='h00001450;  wr_data_rom[ 7087]='h00000000;
    rd_cycle[ 7088] = 1'b1;  wr_cycle[ 7088] = 1'b0;  addr_rom[ 7088]='h00001ae0;  wr_data_rom[ 7088]='h00000000;
    rd_cycle[ 7089] = 1'b0;  wr_cycle[ 7089] = 1'b1;  addr_rom[ 7089]='h00000f2c;  wr_data_rom[ 7089]='h00001dc2;
    rd_cycle[ 7090] = 1'b1;  wr_cycle[ 7090] = 1'b0;  addr_rom[ 7090]='h000004ec;  wr_data_rom[ 7090]='h00000000;
    rd_cycle[ 7091] = 1'b0;  wr_cycle[ 7091] = 1'b1;  addr_rom[ 7091]='h000006f4;  wr_data_rom[ 7091]='h0000154e;
    rd_cycle[ 7092] = 1'b0;  wr_cycle[ 7092] = 1'b1;  addr_rom[ 7092]='h0000018c;  wr_data_rom[ 7092]='h0000141e;
    rd_cycle[ 7093] = 1'b0;  wr_cycle[ 7093] = 1'b1;  addr_rom[ 7093]='h00000788;  wr_data_rom[ 7093]='h000006a9;
    rd_cycle[ 7094] = 1'b0;  wr_cycle[ 7094] = 1'b1;  addr_rom[ 7094]='h000017ac;  wr_data_rom[ 7094]='h000000f7;
    rd_cycle[ 7095] = 1'b1;  wr_cycle[ 7095] = 1'b0;  addr_rom[ 7095]='h000008cc;  wr_data_rom[ 7095]='h00000000;
    rd_cycle[ 7096] = 1'b1;  wr_cycle[ 7096] = 1'b0;  addr_rom[ 7096]='h00000c1c;  wr_data_rom[ 7096]='h00000000;
    rd_cycle[ 7097] = 1'b0;  wr_cycle[ 7097] = 1'b1;  addr_rom[ 7097]='h0000051c;  wr_data_rom[ 7097]='h00001a7a;
    rd_cycle[ 7098] = 1'b1;  wr_cycle[ 7098] = 1'b0;  addr_rom[ 7098]='h00000504;  wr_data_rom[ 7098]='h00000000;
    rd_cycle[ 7099] = 1'b1;  wr_cycle[ 7099] = 1'b0;  addr_rom[ 7099]='h00001088;  wr_data_rom[ 7099]='h00000000;
    rd_cycle[ 7100] = 1'b1;  wr_cycle[ 7100] = 1'b0;  addr_rom[ 7100]='h000009cc;  wr_data_rom[ 7100]='h00000000;
    rd_cycle[ 7101] = 1'b1;  wr_cycle[ 7101] = 1'b0;  addr_rom[ 7101]='h000013bc;  wr_data_rom[ 7101]='h00000000;
    rd_cycle[ 7102] = 1'b0;  wr_cycle[ 7102] = 1'b1;  addr_rom[ 7102]='h000006a0;  wr_data_rom[ 7102]='h00001d8c;
    rd_cycle[ 7103] = 1'b1;  wr_cycle[ 7103] = 1'b0;  addr_rom[ 7103]='h00000328;  wr_data_rom[ 7103]='h00000000;
    rd_cycle[ 7104] = 1'b0;  wr_cycle[ 7104] = 1'b1;  addr_rom[ 7104]='h00000ec0;  wr_data_rom[ 7104]='h00001bea;
    rd_cycle[ 7105] = 1'b0;  wr_cycle[ 7105] = 1'b1;  addr_rom[ 7105]='h00001204;  wr_data_rom[ 7105]='h00000061;
    rd_cycle[ 7106] = 1'b1;  wr_cycle[ 7106] = 1'b0;  addr_rom[ 7106]='h00001844;  wr_data_rom[ 7106]='h00000000;
    rd_cycle[ 7107] = 1'b1;  wr_cycle[ 7107] = 1'b0;  addr_rom[ 7107]='h00001158;  wr_data_rom[ 7107]='h00000000;
    rd_cycle[ 7108] = 1'b1;  wr_cycle[ 7108] = 1'b0;  addr_rom[ 7108]='h00000f08;  wr_data_rom[ 7108]='h00000000;
    rd_cycle[ 7109] = 1'b1;  wr_cycle[ 7109] = 1'b0;  addr_rom[ 7109]='h00001e80;  wr_data_rom[ 7109]='h00000000;
    rd_cycle[ 7110] = 1'b0;  wr_cycle[ 7110] = 1'b1;  addr_rom[ 7110]='h00000c20;  wr_data_rom[ 7110]='h000007e8;
    rd_cycle[ 7111] = 1'b0;  wr_cycle[ 7111] = 1'b1;  addr_rom[ 7111]='h00000b2c;  wr_data_rom[ 7111]='h000014a7;
    rd_cycle[ 7112] = 1'b0;  wr_cycle[ 7112] = 1'b1;  addr_rom[ 7112]='h00001de0;  wr_data_rom[ 7112]='h000014c2;
    rd_cycle[ 7113] = 1'b0;  wr_cycle[ 7113] = 1'b1;  addr_rom[ 7113]='h00000828;  wr_data_rom[ 7113]='h000017cd;
    rd_cycle[ 7114] = 1'b1;  wr_cycle[ 7114] = 1'b0;  addr_rom[ 7114]='h00001ea4;  wr_data_rom[ 7114]='h00000000;
    rd_cycle[ 7115] = 1'b0;  wr_cycle[ 7115] = 1'b1;  addr_rom[ 7115]='h00000920;  wr_data_rom[ 7115]='h00000ce1;
    rd_cycle[ 7116] = 1'b0;  wr_cycle[ 7116] = 1'b1;  addr_rom[ 7116]='h000005ac;  wr_data_rom[ 7116]='h00000ee6;
    rd_cycle[ 7117] = 1'b1;  wr_cycle[ 7117] = 1'b0;  addr_rom[ 7117]='h000012ec;  wr_data_rom[ 7117]='h00000000;
    rd_cycle[ 7118] = 1'b0;  wr_cycle[ 7118] = 1'b1;  addr_rom[ 7118]='h00001190;  wr_data_rom[ 7118]='h00001935;
    rd_cycle[ 7119] = 1'b0;  wr_cycle[ 7119] = 1'b1;  addr_rom[ 7119]='h00000b1c;  wr_data_rom[ 7119]='h00001c3d;
    rd_cycle[ 7120] = 1'b1;  wr_cycle[ 7120] = 1'b0;  addr_rom[ 7120]='h00001dd0;  wr_data_rom[ 7120]='h00000000;
    rd_cycle[ 7121] = 1'b1;  wr_cycle[ 7121] = 1'b0;  addr_rom[ 7121]='h00001cd0;  wr_data_rom[ 7121]='h00000000;
    rd_cycle[ 7122] = 1'b0;  wr_cycle[ 7122] = 1'b1;  addr_rom[ 7122]='h00000450;  wr_data_rom[ 7122]='h000015bc;
    rd_cycle[ 7123] = 1'b1;  wr_cycle[ 7123] = 1'b0;  addr_rom[ 7123]='h000012cc;  wr_data_rom[ 7123]='h00000000;
    rd_cycle[ 7124] = 1'b0;  wr_cycle[ 7124] = 1'b1;  addr_rom[ 7124]='h00001a78;  wr_data_rom[ 7124]='h00001043;
    rd_cycle[ 7125] = 1'b0;  wr_cycle[ 7125] = 1'b1;  addr_rom[ 7125]='h00000d5c;  wr_data_rom[ 7125]='h000012ba;
    rd_cycle[ 7126] = 1'b1;  wr_cycle[ 7126] = 1'b0;  addr_rom[ 7126]='h00000870;  wr_data_rom[ 7126]='h00000000;
    rd_cycle[ 7127] = 1'b1;  wr_cycle[ 7127] = 1'b0;  addr_rom[ 7127]='h00000924;  wr_data_rom[ 7127]='h00000000;
    rd_cycle[ 7128] = 1'b1;  wr_cycle[ 7128] = 1'b0;  addr_rom[ 7128]='h00001354;  wr_data_rom[ 7128]='h00000000;
    rd_cycle[ 7129] = 1'b0;  wr_cycle[ 7129] = 1'b1;  addr_rom[ 7129]='h00001b88;  wr_data_rom[ 7129]='h000005ed;
    rd_cycle[ 7130] = 1'b1;  wr_cycle[ 7130] = 1'b0;  addr_rom[ 7130]='h000014f8;  wr_data_rom[ 7130]='h00000000;
    rd_cycle[ 7131] = 1'b0;  wr_cycle[ 7131] = 1'b1;  addr_rom[ 7131]='h000001ac;  wr_data_rom[ 7131]='h0000050f;
    rd_cycle[ 7132] = 1'b1;  wr_cycle[ 7132] = 1'b0;  addr_rom[ 7132]='h00000ee8;  wr_data_rom[ 7132]='h00000000;
    rd_cycle[ 7133] = 1'b1;  wr_cycle[ 7133] = 1'b0;  addr_rom[ 7133]='h000012e0;  wr_data_rom[ 7133]='h00000000;
    rd_cycle[ 7134] = 1'b1;  wr_cycle[ 7134] = 1'b0;  addr_rom[ 7134]='h00000048;  wr_data_rom[ 7134]='h00000000;
    rd_cycle[ 7135] = 1'b1;  wr_cycle[ 7135] = 1'b0;  addr_rom[ 7135]='h000011a8;  wr_data_rom[ 7135]='h00000000;
    rd_cycle[ 7136] = 1'b0;  wr_cycle[ 7136] = 1'b1;  addr_rom[ 7136]='h00000ed8;  wr_data_rom[ 7136]='h00000849;
    rd_cycle[ 7137] = 1'b0;  wr_cycle[ 7137] = 1'b1;  addr_rom[ 7137]='h000015e0;  wr_data_rom[ 7137]='h000009e4;
    rd_cycle[ 7138] = 1'b1;  wr_cycle[ 7138] = 1'b0;  addr_rom[ 7138]='h00001448;  wr_data_rom[ 7138]='h00000000;
    rd_cycle[ 7139] = 1'b1;  wr_cycle[ 7139] = 1'b0;  addr_rom[ 7139]='h00001310;  wr_data_rom[ 7139]='h00000000;
    rd_cycle[ 7140] = 1'b0;  wr_cycle[ 7140] = 1'b1;  addr_rom[ 7140]='h000011a4;  wr_data_rom[ 7140]='h000009b3;
    rd_cycle[ 7141] = 1'b1;  wr_cycle[ 7141] = 1'b0;  addr_rom[ 7141]='h00001240;  wr_data_rom[ 7141]='h00000000;
    rd_cycle[ 7142] = 1'b1;  wr_cycle[ 7142] = 1'b0;  addr_rom[ 7142]='h00000d10;  wr_data_rom[ 7142]='h00000000;
    rd_cycle[ 7143] = 1'b1;  wr_cycle[ 7143] = 1'b0;  addr_rom[ 7143]='h00001e90;  wr_data_rom[ 7143]='h00000000;
    rd_cycle[ 7144] = 1'b0;  wr_cycle[ 7144] = 1'b1;  addr_rom[ 7144]='h00001948;  wr_data_rom[ 7144]='h0000137c;
    rd_cycle[ 7145] = 1'b1;  wr_cycle[ 7145] = 1'b0;  addr_rom[ 7145]='h00001e24;  wr_data_rom[ 7145]='h00000000;
    rd_cycle[ 7146] = 1'b0;  wr_cycle[ 7146] = 1'b1;  addr_rom[ 7146]='h0000120c;  wr_data_rom[ 7146]='h000010e1;
    rd_cycle[ 7147] = 1'b0;  wr_cycle[ 7147] = 1'b1;  addr_rom[ 7147]='h000006ec;  wr_data_rom[ 7147]='h00001c28;
    rd_cycle[ 7148] = 1'b0;  wr_cycle[ 7148] = 1'b1;  addr_rom[ 7148]='h0000106c;  wr_data_rom[ 7148]='h0000036f;
    rd_cycle[ 7149] = 1'b1;  wr_cycle[ 7149] = 1'b0;  addr_rom[ 7149]='h00000304;  wr_data_rom[ 7149]='h00000000;
    rd_cycle[ 7150] = 1'b1;  wr_cycle[ 7150] = 1'b0;  addr_rom[ 7150]='h00001908;  wr_data_rom[ 7150]='h00000000;
    rd_cycle[ 7151] = 1'b0;  wr_cycle[ 7151] = 1'b1;  addr_rom[ 7151]='h000006e4;  wr_data_rom[ 7151]='h000018e0;
    rd_cycle[ 7152] = 1'b1;  wr_cycle[ 7152] = 1'b0;  addr_rom[ 7152]='h00000edc;  wr_data_rom[ 7152]='h00000000;
    rd_cycle[ 7153] = 1'b1;  wr_cycle[ 7153] = 1'b0;  addr_rom[ 7153]='h00000e74;  wr_data_rom[ 7153]='h00000000;
    rd_cycle[ 7154] = 1'b1;  wr_cycle[ 7154] = 1'b0;  addr_rom[ 7154]='h00000d74;  wr_data_rom[ 7154]='h00000000;
    rd_cycle[ 7155] = 1'b1;  wr_cycle[ 7155] = 1'b0;  addr_rom[ 7155]='h000018e8;  wr_data_rom[ 7155]='h00000000;
    rd_cycle[ 7156] = 1'b1;  wr_cycle[ 7156] = 1'b0;  addr_rom[ 7156]='h000009cc;  wr_data_rom[ 7156]='h00000000;
    rd_cycle[ 7157] = 1'b0;  wr_cycle[ 7157] = 1'b1;  addr_rom[ 7157]='h00001778;  wr_data_rom[ 7157]='h00001da8;
    rd_cycle[ 7158] = 1'b1;  wr_cycle[ 7158] = 1'b0;  addr_rom[ 7158]='h00001814;  wr_data_rom[ 7158]='h00000000;
    rd_cycle[ 7159] = 1'b0;  wr_cycle[ 7159] = 1'b1;  addr_rom[ 7159]='h00000408;  wr_data_rom[ 7159]='h000017d3;
    rd_cycle[ 7160] = 1'b1;  wr_cycle[ 7160] = 1'b0;  addr_rom[ 7160]='h000008fc;  wr_data_rom[ 7160]='h00000000;
    rd_cycle[ 7161] = 1'b1;  wr_cycle[ 7161] = 1'b0;  addr_rom[ 7161]='h000019c8;  wr_data_rom[ 7161]='h00000000;
    rd_cycle[ 7162] = 1'b1;  wr_cycle[ 7162] = 1'b0;  addr_rom[ 7162]='h000001fc;  wr_data_rom[ 7162]='h00000000;
    rd_cycle[ 7163] = 1'b0;  wr_cycle[ 7163] = 1'b1;  addr_rom[ 7163]='h000012b0;  wr_data_rom[ 7163]='h00000941;
    rd_cycle[ 7164] = 1'b1;  wr_cycle[ 7164] = 1'b0;  addr_rom[ 7164]='h00000488;  wr_data_rom[ 7164]='h00000000;
    rd_cycle[ 7165] = 1'b0;  wr_cycle[ 7165] = 1'b1;  addr_rom[ 7165]='h00001004;  wr_data_rom[ 7165]='h00000268;
    rd_cycle[ 7166] = 1'b1;  wr_cycle[ 7166] = 1'b0;  addr_rom[ 7166]='h00001490;  wr_data_rom[ 7166]='h00000000;
    rd_cycle[ 7167] = 1'b0;  wr_cycle[ 7167] = 1'b1;  addr_rom[ 7167]='h00001cec;  wr_data_rom[ 7167]='h00000406;
    rd_cycle[ 7168] = 1'b0;  wr_cycle[ 7168] = 1'b1;  addr_rom[ 7168]='h00001ce8;  wr_data_rom[ 7168]='h00000433;
    rd_cycle[ 7169] = 1'b1;  wr_cycle[ 7169] = 1'b0;  addr_rom[ 7169]='h0000145c;  wr_data_rom[ 7169]='h00000000;
    rd_cycle[ 7170] = 1'b1;  wr_cycle[ 7170] = 1'b0;  addr_rom[ 7170]='h00001378;  wr_data_rom[ 7170]='h00000000;
    rd_cycle[ 7171] = 1'b0;  wr_cycle[ 7171] = 1'b1;  addr_rom[ 7171]='h00000da8;  wr_data_rom[ 7171]='h00000979;
    rd_cycle[ 7172] = 1'b1;  wr_cycle[ 7172] = 1'b0;  addr_rom[ 7172]='h00000484;  wr_data_rom[ 7172]='h00000000;
    rd_cycle[ 7173] = 1'b1;  wr_cycle[ 7173] = 1'b0;  addr_rom[ 7173]='h000019ec;  wr_data_rom[ 7173]='h00000000;
    rd_cycle[ 7174] = 1'b1;  wr_cycle[ 7174] = 1'b0;  addr_rom[ 7174]='h000011f0;  wr_data_rom[ 7174]='h00000000;
    rd_cycle[ 7175] = 1'b0;  wr_cycle[ 7175] = 1'b1;  addr_rom[ 7175]='h00000c88;  wr_data_rom[ 7175]='h0000137b;
    rd_cycle[ 7176] = 1'b0;  wr_cycle[ 7176] = 1'b1;  addr_rom[ 7176]='h0000108c;  wr_data_rom[ 7176]='h0000012f;
    rd_cycle[ 7177] = 1'b0;  wr_cycle[ 7177] = 1'b1;  addr_rom[ 7177]='h0000018c;  wr_data_rom[ 7177]='h0000143d;
    rd_cycle[ 7178] = 1'b0;  wr_cycle[ 7178] = 1'b1;  addr_rom[ 7178]='h00001044;  wr_data_rom[ 7178]='h00000620;
    rd_cycle[ 7179] = 1'b1;  wr_cycle[ 7179] = 1'b0;  addr_rom[ 7179]='h000001d0;  wr_data_rom[ 7179]='h00000000;
    rd_cycle[ 7180] = 1'b0;  wr_cycle[ 7180] = 1'b1;  addr_rom[ 7180]='h000001f0;  wr_data_rom[ 7180]='h00000dd4;
    rd_cycle[ 7181] = 1'b0;  wr_cycle[ 7181] = 1'b1;  addr_rom[ 7181]='h00000070;  wr_data_rom[ 7181]='h000019d3;
    rd_cycle[ 7182] = 1'b1;  wr_cycle[ 7182] = 1'b0;  addr_rom[ 7182]='h0000167c;  wr_data_rom[ 7182]='h00000000;
    rd_cycle[ 7183] = 1'b1;  wr_cycle[ 7183] = 1'b0;  addr_rom[ 7183]='h0000197c;  wr_data_rom[ 7183]='h00000000;
    rd_cycle[ 7184] = 1'b0;  wr_cycle[ 7184] = 1'b1;  addr_rom[ 7184]='h0000005c;  wr_data_rom[ 7184]='h000004d1;
    rd_cycle[ 7185] = 1'b1;  wr_cycle[ 7185] = 1'b0;  addr_rom[ 7185]='h000017e4;  wr_data_rom[ 7185]='h00000000;
    rd_cycle[ 7186] = 1'b0;  wr_cycle[ 7186] = 1'b1;  addr_rom[ 7186]='h00000374;  wr_data_rom[ 7186]='h000019a4;
    rd_cycle[ 7187] = 1'b0;  wr_cycle[ 7187] = 1'b1;  addr_rom[ 7187]='h00001150;  wr_data_rom[ 7187]='h00001635;
    rd_cycle[ 7188] = 1'b0;  wr_cycle[ 7188] = 1'b1;  addr_rom[ 7188]='h00001760;  wr_data_rom[ 7188]='h000000b2;
    rd_cycle[ 7189] = 1'b0;  wr_cycle[ 7189] = 1'b1;  addr_rom[ 7189]='h00000a00;  wr_data_rom[ 7189]='h000001d6;
    rd_cycle[ 7190] = 1'b0;  wr_cycle[ 7190] = 1'b1;  addr_rom[ 7190]='h0000108c;  wr_data_rom[ 7190]='h000019f9;
    rd_cycle[ 7191] = 1'b0;  wr_cycle[ 7191] = 1'b1;  addr_rom[ 7191]='h000006cc;  wr_data_rom[ 7191]='h00001507;
    rd_cycle[ 7192] = 1'b1;  wr_cycle[ 7192] = 1'b0;  addr_rom[ 7192]='h00001e98;  wr_data_rom[ 7192]='h00000000;
    rd_cycle[ 7193] = 1'b0;  wr_cycle[ 7193] = 1'b1;  addr_rom[ 7193]='h0000050c;  wr_data_rom[ 7193]='h00001173;
    rd_cycle[ 7194] = 1'b1;  wr_cycle[ 7194] = 1'b0;  addr_rom[ 7194]='h00001ae0;  wr_data_rom[ 7194]='h00000000;
    rd_cycle[ 7195] = 1'b1;  wr_cycle[ 7195] = 1'b0;  addr_rom[ 7195]='h00000654;  wr_data_rom[ 7195]='h00000000;
    rd_cycle[ 7196] = 1'b0;  wr_cycle[ 7196] = 1'b1;  addr_rom[ 7196]='h00001704;  wr_data_rom[ 7196]='h00001a1d;
    rd_cycle[ 7197] = 1'b0;  wr_cycle[ 7197] = 1'b1;  addr_rom[ 7197]='h00000f4c;  wr_data_rom[ 7197]='h00001cae;
    rd_cycle[ 7198] = 1'b0;  wr_cycle[ 7198] = 1'b1;  addr_rom[ 7198]='h00001c00;  wr_data_rom[ 7198]='h000006db;
    rd_cycle[ 7199] = 1'b1;  wr_cycle[ 7199] = 1'b0;  addr_rom[ 7199]='h00001dec;  wr_data_rom[ 7199]='h00000000;
    rd_cycle[ 7200] = 1'b1;  wr_cycle[ 7200] = 1'b0;  addr_rom[ 7200]='h00001f1c;  wr_data_rom[ 7200]='h00000000;
    rd_cycle[ 7201] = 1'b0;  wr_cycle[ 7201] = 1'b1;  addr_rom[ 7201]='h00001a0c;  wr_data_rom[ 7201]='h00001b72;
    rd_cycle[ 7202] = 1'b1;  wr_cycle[ 7202] = 1'b0;  addr_rom[ 7202]='h000004d0;  wr_data_rom[ 7202]='h00000000;
    rd_cycle[ 7203] = 1'b0;  wr_cycle[ 7203] = 1'b1;  addr_rom[ 7203]='h00000cfc;  wr_data_rom[ 7203]='h00000075;
    rd_cycle[ 7204] = 1'b1;  wr_cycle[ 7204] = 1'b0;  addr_rom[ 7204]='h00001450;  wr_data_rom[ 7204]='h00000000;
    rd_cycle[ 7205] = 1'b0;  wr_cycle[ 7205] = 1'b1;  addr_rom[ 7205]='h00001bbc;  wr_data_rom[ 7205]='h00001c6f;
    rd_cycle[ 7206] = 1'b0;  wr_cycle[ 7206] = 1'b1;  addr_rom[ 7206]='h000015c4;  wr_data_rom[ 7206]='h0000139c;
    rd_cycle[ 7207] = 1'b0;  wr_cycle[ 7207] = 1'b1;  addr_rom[ 7207]='h000019dc;  wr_data_rom[ 7207]='h00000456;
    rd_cycle[ 7208] = 1'b0;  wr_cycle[ 7208] = 1'b1;  addr_rom[ 7208]='h000014b0;  wr_data_rom[ 7208]='h00001bab;
    rd_cycle[ 7209] = 1'b1;  wr_cycle[ 7209] = 1'b0;  addr_rom[ 7209]='h00000668;  wr_data_rom[ 7209]='h00000000;
    rd_cycle[ 7210] = 1'b0;  wr_cycle[ 7210] = 1'b1;  addr_rom[ 7210]='h000003a8;  wr_data_rom[ 7210]='h00001bfb;
    rd_cycle[ 7211] = 1'b1;  wr_cycle[ 7211] = 1'b0;  addr_rom[ 7211]='h00000fbc;  wr_data_rom[ 7211]='h00000000;
    rd_cycle[ 7212] = 1'b0;  wr_cycle[ 7212] = 1'b1;  addr_rom[ 7212]='h00001b44;  wr_data_rom[ 7212]='h00000027;
    rd_cycle[ 7213] = 1'b1;  wr_cycle[ 7213] = 1'b0;  addr_rom[ 7213]='h000013d4;  wr_data_rom[ 7213]='h00000000;
    rd_cycle[ 7214] = 1'b1;  wr_cycle[ 7214] = 1'b0;  addr_rom[ 7214]='h000009c4;  wr_data_rom[ 7214]='h00000000;
    rd_cycle[ 7215] = 1'b0;  wr_cycle[ 7215] = 1'b1;  addr_rom[ 7215]='h000014a8;  wr_data_rom[ 7215]='h00001323;
    rd_cycle[ 7216] = 1'b1;  wr_cycle[ 7216] = 1'b0;  addr_rom[ 7216]='h00000628;  wr_data_rom[ 7216]='h00000000;
    rd_cycle[ 7217] = 1'b0;  wr_cycle[ 7217] = 1'b1;  addr_rom[ 7217]='h00000350;  wr_data_rom[ 7217]='h00001b42;
    rd_cycle[ 7218] = 1'b0;  wr_cycle[ 7218] = 1'b1;  addr_rom[ 7218]='h00000800;  wr_data_rom[ 7218]='h00000d56;
    rd_cycle[ 7219] = 1'b0;  wr_cycle[ 7219] = 1'b1;  addr_rom[ 7219]='h00000f84;  wr_data_rom[ 7219]='h000016ea;
    rd_cycle[ 7220] = 1'b0;  wr_cycle[ 7220] = 1'b1;  addr_rom[ 7220]='h00000890;  wr_data_rom[ 7220]='h000005c2;
    rd_cycle[ 7221] = 1'b1;  wr_cycle[ 7221] = 1'b0;  addr_rom[ 7221]='h00001024;  wr_data_rom[ 7221]='h00000000;
    rd_cycle[ 7222] = 1'b1;  wr_cycle[ 7222] = 1'b0;  addr_rom[ 7222]='h000018f4;  wr_data_rom[ 7222]='h00000000;
    rd_cycle[ 7223] = 1'b0;  wr_cycle[ 7223] = 1'b1;  addr_rom[ 7223]='h000002d0;  wr_data_rom[ 7223]='h00000b0f;
    rd_cycle[ 7224] = 1'b1;  wr_cycle[ 7224] = 1'b0;  addr_rom[ 7224]='h00001a34;  wr_data_rom[ 7224]='h00000000;
    rd_cycle[ 7225] = 1'b1;  wr_cycle[ 7225] = 1'b0;  addr_rom[ 7225]='h00001a8c;  wr_data_rom[ 7225]='h00000000;
    rd_cycle[ 7226] = 1'b1;  wr_cycle[ 7226] = 1'b0;  addr_rom[ 7226]='h000006c4;  wr_data_rom[ 7226]='h00000000;
    rd_cycle[ 7227] = 1'b0;  wr_cycle[ 7227] = 1'b1;  addr_rom[ 7227]='h0000097c;  wr_data_rom[ 7227]='h00000e3d;
    rd_cycle[ 7228] = 1'b1;  wr_cycle[ 7228] = 1'b0;  addr_rom[ 7228]='h00000ed8;  wr_data_rom[ 7228]='h00000000;
    rd_cycle[ 7229] = 1'b1;  wr_cycle[ 7229] = 1'b0;  addr_rom[ 7229]='h000006dc;  wr_data_rom[ 7229]='h00000000;
    rd_cycle[ 7230] = 1'b0;  wr_cycle[ 7230] = 1'b1;  addr_rom[ 7230]='h000016c8;  wr_data_rom[ 7230]='h00001aa3;
    rd_cycle[ 7231] = 1'b0;  wr_cycle[ 7231] = 1'b1;  addr_rom[ 7231]='h000009ec;  wr_data_rom[ 7231]='h000008c6;
    rd_cycle[ 7232] = 1'b0;  wr_cycle[ 7232] = 1'b1;  addr_rom[ 7232]='h00000c68;  wr_data_rom[ 7232]='h0000173e;
    rd_cycle[ 7233] = 1'b1;  wr_cycle[ 7233] = 1'b0;  addr_rom[ 7233]='h00000490;  wr_data_rom[ 7233]='h00000000;
    rd_cycle[ 7234] = 1'b1;  wr_cycle[ 7234] = 1'b0;  addr_rom[ 7234]='h0000150c;  wr_data_rom[ 7234]='h00000000;
    rd_cycle[ 7235] = 1'b1;  wr_cycle[ 7235] = 1'b0;  addr_rom[ 7235]='h000006e8;  wr_data_rom[ 7235]='h00000000;
    rd_cycle[ 7236] = 1'b1;  wr_cycle[ 7236] = 1'b0;  addr_rom[ 7236]='h00001ab0;  wr_data_rom[ 7236]='h00000000;
    rd_cycle[ 7237] = 1'b0;  wr_cycle[ 7237] = 1'b1;  addr_rom[ 7237]='h0000194c;  wr_data_rom[ 7237]='h00001abe;
    rd_cycle[ 7238] = 1'b1;  wr_cycle[ 7238] = 1'b0;  addr_rom[ 7238]='h00000e1c;  wr_data_rom[ 7238]='h00000000;
    rd_cycle[ 7239] = 1'b0;  wr_cycle[ 7239] = 1'b1;  addr_rom[ 7239]='h000004ec;  wr_data_rom[ 7239]='h00001c24;
    rd_cycle[ 7240] = 1'b0;  wr_cycle[ 7240] = 1'b1;  addr_rom[ 7240]='h00000034;  wr_data_rom[ 7240]='h0000057a;
    rd_cycle[ 7241] = 1'b0;  wr_cycle[ 7241] = 1'b1;  addr_rom[ 7241]='h00001560;  wr_data_rom[ 7241]='h00001548;
    rd_cycle[ 7242] = 1'b1;  wr_cycle[ 7242] = 1'b0;  addr_rom[ 7242]='h00001d08;  wr_data_rom[ 7242]='h00000000;
    rd_cycle[ 7243] = 1'b1;  wr_cycle[ 7243] = 1'b0;  addr_rom[ 7243]='h00001154;  wr_data_rom[ 7243]='h00000000;
    rd_cycle[ 7244] = 1'b1;  wr_cycle[ 7244] = 1'b0;  addr_rom[ 7244]='h000014c8;  wr_data_rom[ 7244]='h00000000;
    rd_cycle[ 7245] = 1'b0;  wr_cycle[ 7245] = 1'b1;  addr_rom[ 7245]='h000003c4;  wr_data_rom[ 7245]='h00000279;
    rd_cycle[ 7246] = 1'b1;  wr_cycle[ 7246] = 1'b0;  addr_rom[ 7246]='h00001c6c;  wr_data_rom[ 7246]='h00000000;
    rd_cycle[ 7247] = 1'b0;  wr_cycle[ 7247] = 1'b1;  addr_rom[ 7247]='h00001840;  wr_data_rom[ 7247]='h00000873;
    rd_cycle[ 7248] = 1'b0;  wr_cycle[ 7248] = 1'b1;  addr_rom[ 7248]='h00000260;  wr_data_rom[ 7248]='h0000118f;
    rd_cycle[ 7249] = 1'b0;  wr_cycle[ 7249] = 1'b1;  addr_rom[ 7249]='h00001968;  wr_data_rom[ 7249]='h0000057b;
    rd_cycle[ 7250] = 1'b0;  wr_cycle[ 7250] = 1'b1;  addr_rom[ 7250]='h00000498;  wr_data_rom[ 7250]='h00000e25;
    rd_cycle[ 7251] = 1'b1;  wr_cycle[ 7251] = 1'b0;  addr_rom[ 7251]='h00001d8c;  wr_data_rom[ 7251]='h00000000;
    rd_cycle[ 7252] = 1'b0;  wr_cycle[ 7252] = 1'b1;  addr_rom[ 7252]='h00000ed0;  wr_data_rom[ 7252]='h000012e3;
    rd_cycle[ 7253] = 1'b0;  wr_cycle[ 7253] = 1'b1;  addr_rom[ 7253]='h000017f0;  wr_data_rom[ 7253]='h00001952;
    rd_cycle[ 7254] = 1'b0;  wr_cycle[ 7254] = 1'b1;  addr_rom[ 7254]='h00001370;  wr_data_rom[ 7254]='h00001838;
    rd_cycle[ 7255] = 1'b1;  wr_cycle[ 7255] = 1'b0;  addr_rom[ 7255]='h00001180;  wr_data_rom[ 7255]='h00000000;
    rd_cycle[ 7256] = 1'b1;  wr_cycle[ 7256] = 1'b0;  addr_rom[ 7256]='h00000468;  wr_data_rom[ 7256]='h00000000;
    rd_cycle[ 7257] = 1'b0;  wr_cycle[ 7257] = 1'b1;  addr_rom[ 7257]='h000009dc;  wr_data_rom[ 7257]='h00001284;
    rd_cycle[ 7258] = 1'b1;  wr_cycle[ 7258] = 1'b0;  addr_rom[ 7258]='h00001c44;  wr_data_rom[ 7258]='h00000000;
    rd_cycle[ 7259] = 1'b0;  wr_cycle[ 7259] = 1'b1;  addr_rom[ 7259]='h00000ac8;  wr_data_rom[ 7259]='h00001640;
    rd_cycle[ 7260] = 1'b0;  wr_cycle[ 7260] = 1'b1;  addr_rom[ 7260]='h00001b64;  wr_data_rom[ 7260]='h00001996;
    rd_cycle[ 7261] = 1'b1;  wr_cycle[ 7261] = 1'b0;  addr_rom[ 7261]='h0000076c;  wr_data_rom[ 7261]='h00000000;
    rd_cycle[ 7262] = 1'b1;  wr_cycle[ 7262] = 1'b0;  addr_rom[ 7262]='h0000056c;  wr_data_rom[ 7262]='h00000000;
    rd_cycle[ 7263] = 1'b1;  wr_cycle[ 7263] = 1'b0;  addr_rom[ 7263]='h00000ae0;  wr_data_rom[ 7263]='h00000000;
    rd_cycle[ 7264] = 1'b0;  wr_cycle[ 7264] = 1'b1;  addr_rom[ 7264]='h00000cf4;  wr_data_rom[ 7264]='h00000e58;
    rd_cycle[ 7265] = 1'b1;  wr_cycle[ 7265] = 1'b0;  addr_rom[ 7265]='h00001444;  wr_data_rom[ 7265]='h00000000;
    rd_cycle[ 7266] = 1'b1;  wr_cycle[ 7266] = 1'b0;  addr_rom[ 7266]='h00000f28;  wr_data_rom[ 7266]='h00000000;
    rd_cycle[ 7267] = 1'b1;  wr_cycle[ 7267] = 1'b0;  addr_rom[ 7267]='h000009c4;  wr_data_rom[ 7267]='h00000000;
    rd_cycle[ 7268] = 1'b1;  wr_cycle[ 7268] = 1'b0;  addr_rom[ 7268]='h00001650;  wr_data_rom[ 7268]='h00000000;
    rd_cycle[ 7269] = 1'b1;  wr_cycle[ 7269] = 1'b0;  addr_rom[ 7269]='h000012ac;  wr_data_rom[ 7269]='h00000000;
    rd_cycle[ 7270] = 1'b1;  wr_cycle[ 7270] = 1'b0;  addr_rom[ 7270]='h00000600;  wr_data_rom[ 7270]='h00000000;
    rd_cycle[ 7271] = 1'b0;  wr_cycle[ 7271] = 1'b1;  addr_rom[ 7271]='h00000e10;  wr_data_rom[ 7271]='h000011f4;
    rd_cycle[ 7272] = 1'b1;  wr_cycle[ 7272] = 1'b0;  addr_rom[ 7272]='h00000764;  wr_data_rom[ 7272]='h00000000;
    rd_cycle[ 7273] = 1'b1;  wr_cycle[ 7273] = 1'b0;  addr_rom[ 7273]='h00001318;  wr_data_rom[ 7273]='h00000000;
    rd_cycle[ 7274] = 1'b1;  wr_cycle[ 7274] = 1'b0;  addr_rom[ 7274]='h00000274;  wr_data_rom[ 7274]='h00000000;
    rd_cycle[ 7275] = 1'b1;  wr_cycle[ 7275] = 1'b0;  addr_rom[ 7275]='h00000278;  wr_data_rom[ 7275]='h00000000;
    rd_cycle[ 7276] = 1'b0;  wr_cycle[ 7276] = 1'b1;  addr_rom[ 7276]='h00001224;  wr_data_rom[ 7276]='h000009c0;
    rd_cycle[ 7277] = 1'b0;  wr_cycle[ 7277] = 1'b1;  addr_rom[ 7277]='h000007d0;  wr_data_rom[ 7277]='h000003bf;
    rd_cycle[ 7278] = 1'b0;  wr_cycle[ 7278] = 1'b1;  addr_rom[ 7278]='h00000984;  wr_data_rom[ 7278]='h00001872;
    rd_cycle[ 7279] = 1'b1;  wr_cycle[ 7279] = 1'b0;  addr_rom[ 7279]='h00000088;  wr_data_rom[ 7279]='h00000000;
    rd_cycle[ 7280] = 1'b1;  wr_cycle[ 7280] = 1'b0;  addr_rom[ 7280]='h000017e0;  wr_data_rom[ 7280]='h00000000;
    rd_cycle[ 7281] = 1'b1;  wr_cycle[ 7281] = 1'b0;  addr_rom[ 7281]='h00001d0c;  wr_data_rom[ 7281]='h00000000;
    rd_cycle[ 7282] = 1'b1;  wr_cycle[ 7282] = 1'b0;  addr_rom[ 7282]='h0000096c;  wr_data_rom[ 7282]='h00000000;
    rd_cycle[ 7283] = 1'b1;  wr_cycle[ 7283] = 1'b0;  addr_rom[ 7283]='h00001afc;  wr_data_rom[ 7283]='h00000000;
    rd_cycle[ 7284] = 1'b1;  wr_cycle[ 7284] = 1'b0;  addr_rom[ 7284]='h00000748;  wr_data_rom[ 7284]='h00000000;
    rd_cycle[ 7285] = 1'b1;  wr_cycle[ 7285] = 1'b0;  addr_rom[ 7285]='h000015a0;  wr_data_rom[ 7285]='h00000000;
    rd_cycle[ 7286] = 1'b0;  wr_cycle[ 7286] = 1'b1;  addr_rom[ 7286]='h000012a4;  wr_data_rom[ 7286]='h00000639;
    rd_cycle[ 7287] = 1'b0;  wr_cycle[ 7287] = 1'b1;  addr_rom[ 7287]='h000002b4;  wr_data_rom[ 7287]='h00001884;
    rd_cycle[ 7288] = 1'b0;  wr_cycle[ 7288] = 1'b1;  addr_rom[ 7288]='h00001ab8;  wr_data_rom[ 7288]='h000018a5;
    rd_cycle[ 7289] = 1'b0;  wr_cycle[ 7289] = 1'b1;  addr_rom[ 7289]='h00001a34;  wr_data_rom[ 7289]='h00000da6;
    rd_cycle[ 7290] = 1'b1;  wr_cycle[ 7290] = 1'b0;  addr_rom[ 7290]='h000004ec;  wr_data_rom[ 7290]='h00000000;
    rd_cycle[ 7291] = 1'b1;  wr_cycle[ 7291] = 1'b0;  addr_rom[ 7291]='h00000648;  wr_data_rom[ 7291]='h00000000;
    rd_cycle[ 7292] = 1'b1;  wr_cycle[ 7292] = 1'b0;  addr_rom[ 7292]='h00001528;  wr_data_rom[ 7292]='h00000000;
    rd_cycle[ 7293] = 1'b0;  wr_cycle[ 7293] = 1'b1;  addr_rom[ 7293]='h00001c90;  wr_data_rom[ 7293]='h00000f5d;
    rd_cycle[ 7294] = 1'b1;  wr_cycle[ 7294] = 1'b0;  addr_rom[ 7294]='h0000102c;  wr_data_rom[ 7294]='h00000000;
    rd_cycle[ 7295] = 1'b1;  wr_cycle[ 7295] = 1'b0;  addr_rom[ 7295]='h00000614;  wr_data_rom[ 7295]='h00000000;
    rd_cycle[ 7296] = 1'b0;  wr_cycle[ 7296] = 1'b1;  addr_rom[ 7296]='h00000ebc;  wr_data_rom[ 7296]='h0000047a;
    rd_cycle[ 7297] = 1'b1;  wr_cycle[ 7297] = 1'b0;  addr_rom[ 7297]='h00000798;  wr_data_rom[ 7297]='h00000000;
    rd_cycle[ 7298] = 1'b0;  wr_cycle[ 7298] = 1'b1;  addr_rom[ 7298]='h00000fb0;  wr_data_rom[ 7298]='h00000f91;
    rd_cycle[ 7299] = 1'b0;  wr_cycle[ 7299] = 1'b1;  addr_rom[ 7299]='h000004bc;  wr_data_rom[ 7299]='h0000063c;
    rd_cycle[ 7300] = 1'b1;  wr_cycle[ 7300] = 1'b0;  addr_rom[ 7300]='h00000808;  wr_data_rom[ 7300]='h00000000;
    rd_cycle[ 7301] = 1'b1;  wr_cycle[ 7301] = 1'b0;  addr_rom[ 7301]='h00000720;  wr_data_rom[ 7301]='h00000000;
    rd_cycle[ 7302] = 1'b0;  wr_cycle[ 7302] = 1'b1;  addr_rom[ 7302]='h0000145c;  wr_data_rom[ 7302]='h000000af;
    rd_cycle[ 7303] = 1'b0;  wr_cycle[ 7303] = 1'b1;  addr_rom[ 7303]='h00000f94;  wr_data_rom[ 7303]='h0000157f;
    rd_cycle[ 7304] = 1'b0;  wr_cycle[ 7304] = 1'b1;  addr_rom[ 7304]='h00000f00;  wr_data_rom[ 7304]='h000002df;
    rd_cycle[ 7305] = 1'b1;  wr_cycle[ 7305] = 1'b0;  addr_rom[ 7305]='h00001d8c;  wr_data_rom[ 7305]='h00000000;
    rd_cycle[ 7306] = 1'b1;  wr_cycle[ 7306] = 1'b0;  addr_rom[ 7306]='h00001200;  wr_data_rom[ 7306]='h00000000;
    rd_cycle[ 7307] = 1'b0;  wr_cycle[ 7307] = 1'b1;  addr_rom[ 7307]='h00000e58;  wr_data_rom[ 7307]='h00001677;
    rd_cycle[ 7308] = 1'b0;  wr_cycle[ 7308] = 1'b1;  addr_rom[ 7308]='h000007cc;  wr_data_rom[ 7308]='h00001f27;
    rd_cycle[ 7309] = 1'b0;  wr_cycle[ 7309] = 1'b1;  addr_rom[ 7309]='h000000e8;  wr_data_rom[ 7309]='h00000997;
    rd_cycle[ 7310] = 1'b0;  wr_cycle[ 7310] = 1'b1;  addr_rom[ 7310]='h000018d0;  wr_data_rom[ 7310]='h0000141e;
    rd_cycle[ 7311] = 1'b0;  wr_cycle[ 7311] = 1'b1;  addr_rom[ 7311]='h00001be0;  wr_data_rom[ 7311]='h00000b12;
    rd_cycle[ 7312] = 1'b1;  wr_cycle[ 7312] = 1'b0;  addr_rom[ 7312]='h000011dc;  wr_data_rom[ 7312]='h00000000;
    rd_cycle[ 7313] = 1'b1;  wr_cycle[ 7313] = 1'b0;  addr_rom[ 7313]='h0000169c;  wr_data_rom[ 7313]='h00000000;
    rd_cycle[ 7314] = 1'b0;  wr_cycle[ 7314] = 1'b1;  addr_rom[ 7314]='h00000b74;  wr_data_rom[ 7314]='h00001ae9;
    rd_cycle[ 7315] = 1'b1;  wr_cycle[ 7315] = 1'b0;  addr_rom[ 7315]='h00000d00;  wr_data_rom[ 7315]='h00000000;
    rd_cycle[ 7316] = 1'b1;  wr_cycle[ 7316] = 1'b0;  addr_rom[ 7316]='h00000124;  wr_data_rom[ 7316]='h00000000;
    rd_cycle[ 7317] = 1'b1;  wr_cycle[ 7317] = 1'b0;  addr_rom[ 7317]='h00001954;  wr_data_rom[ 7317]='h00000000;
    rd_cycle[ 7318] = 1'b1;  wr_cycle[ 7318] = 1'b0;  addr_rom[ 7318]='h0000052c;  wr_data_rom[ 7318]='h00000000;
    rd_cycle[ 7319] = 1'b0;  wr_cycle[ 7319] = 1'b1;  addr_rom[ 7319]='h000007dc;  wr_data_rom[ 7319]='h00000f80;
    rd_cycle[ 7320] = 1'b0;  wr_cycle[ 7320] = 1'b1;  addr_rom[ 7320]='h00001004;  wr_data_rom[ 7320]='h000009f3;
    rd_cycle[ 7321] = 1'b1;  wr_cycle[ 7321] = 1'b0;  addr_rom[ 7321]='h000013e4;  wr_data_rom[ 7321]='h00000000;
    rd_cycle[ 7322] = 1'b0;  wr_cycle[ 7322] = 1'b1;  addr_rom[ 7322]='h00000b84;  wr_data_rom[ 7322]='h00000092;
    rd_cycle[ 7323] = 1'b1;  wr_cycle[ 7323] = 1'b0;  addr_rom[ 7323]='h00001090;  wr_data_rom[ 7323]='h00000000;
    rd_cycle[ 7324] = 1'b1;  wr_cycle[ 7324] = 1'b0;  addr_rom[ 7324]='h000003fc;  wr_data_rom[ 7324]='h00000000;
    rd_cycle[ 7325] = 1'b1;  wr_cycle[ 7325] = 1'b0;  addr_rom[ 7325]='h00000f88;  wr_data_rom[ 7325]='h00000000;
    rd_cycle[ 7326] = 1'b1;  wr_cycle[ 7326] = 1'b0;  addr_rom[ 7326]='h00001950;  wr_data_rom[ 7326]='h00000000;
    rd_cycle[ 7327] = 1'b0;  wr_cycle[ 7327] = 1'b1;  addr_rom[ 7327]='h00001284;  wr_data_rom[ 7327]='h000015fd;
    rd_cycle[ 7328] = 1'b0;  wr_cycle[ 7328] = 1'b1;  addr_rom[ 7328]='h0000099c;  wr_data_rom[ 7328]='h00000fc0;
    rd_cycle[ 7329] = 1'b0;  wr_cycle[ 7329] = 1'b1;  addr_rom[ 7329]='h00000680;  wr_data_rom[ 7329]='h0000111d;
    rd_cycle[ 7330] = 1'b1;  wr_cycle[ 7330] = 1'b0;  addr_rom[ 7330]='h00000a64;  wr_data_rom[ 7330]='h00000000;
    rd_cycle[ 7331] = 1'b1;  wr_cycle[ 7331] = 1'b0;  addr_rom[ 7331]='h00001338;  wr_data_rom[ 7331]='h00000000;
    rd_cycle[ 7332] = 1'b1;  wr_cycle[ 7332] = 1'b0;  addr_rom[ 7332]='h00001ac4;  wr_data_rom[ 7332]='h00000000;
    rd_cycle[ 7333] = 1'b1;  wr_cycle[ 7333] = 1'b0;  addr_rom[ 7333]='h00000228;  wr_data_rom[ 7333]='h00000000;
    rd_cycle[ 7334] = 1'b0;  wr_cycle[ 7334] = 1'b1;  addr_rom[ 7334]='h00001d38;  wr_data_rom[ 7334]='h00001d2e;
    rd_cycle[ 7335] = 1'b0;  wr_cycle[ 7335] = 1'b1;  addr_rom[ 7335]='h00000e44;  wr_data_rom[ 7335]='h00001974;
    rd_cycle[ 7336] = 1'b0;  wr_cycle[ 7336] = 1'b1;  addr_rom[ 7336]='h0000008c;  wr_data_rom[ 7336]='h000010f4;
    rd_cycle[ 7337] = 1'b1;  wr_cycle[ 7337] = 1'b0;  addr_rom[ 7337]='h000016b4;  wr_data_rom[ 7337]='h00000000;
    rd_cycle[ 7338] = 1'b1;  wr_cycle[ 7338] = 1'b0;  addr_rom[ 7338]='h00000478;  wr_data_rom[ 7338]='h00000000;
    rd_cycle[ 7339] = 1'b1;  wr_cycle[ 7339] = 1'b0;  addr_rom[ 7339]='h00001000;  wr_data_rom[ 7339]='h00000000;
    rd_cycle[ 7340] = 1'b0;  wr_cycle[ 7340] = 1'b1;  addr_rom[ 7340]='h00000ae0;  wr_data_rom[ 7340]='h00001932;
    rd_cycle[ 7341] = 1'b1;  wr_cycle[ 7341] = 1'b0;  addr_rom[ 7341]='h000006f4;  wr_data_rom[ 7341]='h00000000;
    rd_cycle[ 7342] = 1'b0;  wr_cycle[ 7342] = 1'b1;  addr_rom[ 7342]='h00001628;  wr_data_rom[ 7342]='h00001a47;
    rd_cycle[ 7343] = 1'b0;  wr_cycle[ 7343] = 1'b1;  addr_rom[ 7343]='h00000a70;  wr_data_rom[ 7343]='h00001619;
    rd_cycle[ 7344] = 1'b1;  wr_cycle[ 7344] = 1'b0;  addr_rom[ 7344]='h00001f3c;  wr_data_rom[ 7344]='h00000000;
    rd_cycle[ 7345] = 1'b1;  wr_cycle[ 7345] = 1'b0;  addr_rom[ 7345]='h00001070;  wr_data_rom[ 7345]='h00000000;
    rd_cycle[ 7346] = 1'b0;  wr_cycle[ 7346] = 1'b1;  addr_rom[ 7346]='h000003bc;  wr_data_rom[ 7346]='h0000137d;
    rd_cycle[ 7347] = 1'b0;  wr_cycle[ 7347] = 1'b1;  addr_rom[ 7347]='h00000eb0;  wr_data_rom[ 7347]='h00000f2d;
    rd_cycle[ 7348] = 1'b1;  wr_cycle[ 7348] = 1'b0;  addr_rom[ 7348]='h00000be8;  wr_data_rom[ 7348]='h00000000;
    rd_cycle[ 7349] = 1'b0;  wr_cycle[ 7349] = 1'b1;  addr_rom[ 7349]='h00000b4c;  wr_data_rom[ 7349]='h00000631;
    rd_cycle[ 7350] = 1'b0;  wr_cycle[ 7350] = 1'b1;  addr_rom[ 7350]='h00000fe8;  wr_data_rom[ 7350]='h00001df1;
    rd_cycle[ 7351] = 1'b1;  wr_cycle[ 7351] = 1'b0;  addr_rom[ 7351]='h000003a4;  wr_data_rom[ 7351]='h00000000;
    rd_cycle[ 7352] = 1'b1;  wr_cycle[ 7352] = 1'b0;  addr_rom[ 7352]='h00001468;  wr_data_rom[ 7352]='h00000000;
    rd_cycle[ 7353] = 1'b1;  wr_cycle[ 7353] = 1'b0;  addr_rom[ 7353]='h00001588;  wr_data_rom[ 7353]='h00000000;
    rd_cycle[ 7354] = 1'b0;  wr_cycle[ 7354] = 1'b1;  addr_rom[ 7354]='h00001dd8;  wr_data_rom[ 7354]='h0000037d;
    rd_cycle[ 7355] = 1'b0;  wr_cycle[ 7355] = 1'b1;  addr_rom[ 7355]='h00000e54;  wr_data_rom[ 7355]='h00000c47;
    rd_cycle[ 7356] = 1'b0;  wr_cycle[ 7356] = 1'b1;  addr_rom[ 7356]='h00001920;  wr_data_rom[ 7356]='h00000871;
    rd_cycle[ 7357] = 1'b0;  wr_cycle[ 7357] = 1'b1;  addr_rom[ 7357]='h00001a5c;  wr_data_rom[ 7357]='h00000d4c;
    rd_cycle[ 7358] = 1'b1;  wr_cycle[ 7358] = 1'b0;  addr_rom[ 7358]='h000011b8;  wr_data_rom[ 7358]='h00000000;
    rd_cycle[ 7359] = 1'b0;  wr_cycle[ 7359] = 1'b1;  addr_rom[ 7359]='h00000c20;  wr_data_rom[ 7359]='h00000663;
    rd_cycle[ 7360] = 1'b0;  wr_cycle[ 7360] = 1'b1;  addr_rom[ 7360]='h000018e4;  wr_data_rom[ 7360]='h0000087d;
    rd_cycle[ 7361] = 1'b0;  wr_cycle[ 7361] = 1'b1;  addr_rom[ 7361]='h00001dd4;  wr_data_rom[ 7361]='h0000084f;
    rd_cycle[ 7362] = 1'b1;  wr_cycle[ 7362] = 1'b0;  addr_rom[ 7362]='h00000294;  wr_data_rom[ 7362]='h00000000;
    rd_cycle[ 7363] = 1'b0;  wr_cycle[ 7363] = 1'b1;  addr_rom[ 7363]='h000016c4;  wr_data_rom[ 7363]='h0000009e;
    rd_cycle[ 7364] = 1'b0;  wr_cycle[ 7364] = 1'b1;  addr_rom[ 7364]='h00001800;  wr_data_rom[ 7364]='h000007eb;
    rd_cycle[ 7365] = 1'b0;  wr_cycle[ 7365] = 1'b1;  addr_rom[ 7365]='h0000129c;  wr_data_rom[ 7365]='h00001ac9;
    rd_cycle[ 7366] = 1'b0;  wr_cycle[ 7366] = 1'b1;  addr_rom[ 7366]='h00001330;  wr_data_rom[ 7366]='h000001b1;
    rd_cycle[ 7367] = 1'b0;  wr_cycle[ 7367] = 1'b1;  addr_rom[ 7367]='h000009c4;  wr_data_rom[ 7367]='h00000444;
    rd_cycle[ 7368] = 1'b0;  wr_cycle[ 7368] = 1'b1;  addr_rom[ 7368]='h00000340;  wr_data_rom[ 7368]='h000010d0;
    rd_cycle[ 7369] = 1'b1;  wr_cycle[ 7369] = 1'b0;  addr_rom[ 7369]='h00001794;  wr_data_rom[ 7369]='h00000000;
    rd_cycle[ 7370] = 1'b1;  wr_cycle[ 7370] = 1'b0;  addr_rom[ 7370]='h00001dec;  wr_data_rom[ 7370]='h00000000;
    rd_cycle[ 7371] = 1'b0;  wr_cycle[ 7371] = 1'b1;  addr_rom[ 7371]='h00001db0;  wr_data_rom[ 7371]='h00001574;
    rd_cycle[ 7372] = 1'b0;  wr_cycle[ 7372] = 1'b1;  addr_rom[ 7372]='h00000b3c;  wr_data_rom[ 7372]='h000000ff;
    rd_cycle[ 7373] = 1'b0;  wr_cycle[ 7373] = 1'b1;  addr_rom[ 7373]='h00001dc4;  wr_data_rom[ 7373]='h00000b7c;
    rd_cycle[ 7374] = 1'b0;  wr_cycle[ 7374] = 1'b1;  addr_rom[ 7374]='h00001dfc;  wr_data_rom[ 7374]='h0000012c;
    rd_cycle[ 7375] = 1'b1;  wr_cycle[ 7375] = 1'b0;  addr_rom[ 7375]='h00000630;  wr_data_rom[ 7375]='h00000000;
    rd_cycle[ 7376] = 1'b0;  wr_cycle[ 7376] = 1'b1;  addr_rom[ 7376]='h00000324;  wr_data_rom[ 7376]='h00001cf3;
    rd_cycle[ 7377] = 1'b1;  wr_cycle[ 7377] = 1'b0;  addr_rom[ 7377]='h000011c8;  wr_data_rom[ 7377]='h00000000;
    rd_cycle[ 7378] = 1'b1;  wr_cycle[ 7378] = 1'b0;  addr_rom[ 7378]='h00000fa8;  wr_data_rom[ 7378]='h00000000;
    rd_cycle[ 7379] = 1'b0;  wr_cycle[ 7379] = 1'b1;  addr_rom[ 7379]='h000000b0;  wr_data_rom[ 7379]='h00001219;
    rd_cycle[ 7380] = 1'b1;  wr_cycle[ 7380] = 1'b0;  addr_rom[ 7380]='h00001b74;  wr_data_rom[ 7380]='h00000000;
    rd_cycle[ 7381] = 1'b0;  wr_cycle[ 7381] = 1'b1;  addr_rom[ 7381]='h0000118c;  wr_data_rom[ 7381]='h00001e77;
    rd_cycle[ 7382] = 1'b1;  wr_cycle[ 7382] = 1'b0;  addr_rom[ 7382]='h00001b80;  wr_data_rom[ 7382]='h00000000;
    rd_cycle[ 7383] = 1'b0;  wr_cycle[ 7383] = 1'b1;  addr_rom[ 7383]='h00000180;  wr_data_rom[ 7383]='h00001967;
    rd_cycle[ 7384] = 1'b0;  wr_cycle[ 7384] = 1'b1;  addr_rom[ 7384]='h00001de4;  wr_data_rom[ 7384]='h000000e5;
    rd_cycle[ 7385] = 1'b1;  wr_cycle[ 7385] = 1'b0;  addr_rom[ 7385]='h00000240;  wr_data_rom[ 7385]='h00000000;
    rd_cycle[ 7386] = 1'b0;  wr_cycle[ 7386] = 1'b1;  addr_rom[ 7386]='h00000458;  wr_data_rom[ 7386]='h000015ff;
    rd_cycle[ 7387] = 1'b1;  wr_cycle[ 7387] = 1'b0;  addr_rom[ 7387]='h00000c10;  wr_data_rom[ 7387]='h00000000;
    rd_cycle[ 7388] = 1'b1;  wr_cycle[ 7388] = 1'b0;  addr_rom[ 7388]='h000016a4;  wr_data_rom[ 7388]='h00000000;
    rd_cycle[ 7389] = 1'b1;  wr_cycle[ 7389] = 1'b0;  addr_rom[ 7389]='h00000168;  wr_data_rom[ 7389]='h00000000;
    rd_cycle[ 7390] = 1'b0;  wr_cycle[ 7390] = 1'b1;  addr_rom[ 7390]='h00000104;  wr_data_rom[ 7390]='h00000d73;
    rd_cycle[ 7391] = 1'b1;  wr_cycle[ 7391] = 1'b0;  addr_rom[ 7391]='h00001ae0;  wr_data_rom[ 7391]='h00000000;
    rd_cycle[ 7392] = 1'b1;  wr_cycle[ 7392] = 1'b0;  addr_rom[ 7392]='h00001ec0;  wr_data_rom[ 7392]='h00000000;
    rd_cycle[ 7393] = 1'b1;  wr_cycle[ 7393] = 1'b0;  addr_rom[ 7393]='h00001118;  wr_data_rom[ 7393]='h00000000;
    rd_cycle[ 7394] = 1'b0;  wr_cycle[ 7394] = 1'b1;  addr_rom[ 7394]='h000013f4;  wr_data_rom[ 7394]='h000012e2;
    rd_cycle[ 7395] = 1'b0;  wr_cycle[ 7395] = 1'b1;  addr_rom[ 7395]='h00001d6c;  wr_data_rom[ 7395]='h0000072c;
    rd_cycle[ 7396] = 1'b0;  wr_cycle[ 7396] = 1'b1;  addr_rom[ 7396]='h000012e0;  wr_data_rom[ 7396]='h0000162d;
    rd_cycle[ 7397] = 1'b1;  wr_cycle[ 7397] = 1'b0;  addr_rom[ 7397]='h00001b68;  wr_data_rom[ 7397]='h00000000;
    rd_cycle[ 7398] = 1'b0;  wr_cycle[ 7398] = 1'b1;  addr_rom[ 7398]='h00001e44;  wr_data_rom[ 7398]='h00000665;
    rd_cycle[ 7399] = 1'b0;  wr_cycle[ 7399] = 1'b1;  addr_rom[ 7399]='h00000fb8;  wr_data_rom[ 7399]='h00001ad7;
    rd_cycle[ 7400] = 1'b1;  wr_cycle[ 7400] = 1'b0;  addr_rom[ 7400]='h00000790;  wr_data_rom[ 7400]='h00000000;
    rd_cycle[ 7401] = 1'b1;  wr_cycle[ 7401] = 1'b0;  addr_rom[ 7401]='h00001a78;  wr_data_rom[ 7401]='h00000000;
    rd_cycle[ 7402] = 1'b0;  wr_cycle[ 7402] = 1'b1;  addr_rom[ 7402]='h00001b64;  wr_data_rom[ 7402]='h00000843;
    rd_cycle[ 7403] = 1'b0;  wr_cycle[ 7403] = 1'b1;  addr_rom[ 7403]='h000010c8;  wr_data_rom[ 7403]='h000001e7;
    rd_cycle[ 7404] = 1'b1;  wr_cycle[ 7404] = 1'b0;  addr_rom[ 7404]='h00000aa0;  wr_data_rom[ 7404]='h00000000;
    rd_cycle[ 7405] = 1'b0;  wr_cycle[ 7405] = 1'b1;  addr_rom[ 7405]='h00000928;  wr_data_rom[ 7405]='h00001b3d;
    rd_cycle[ 7406] = 1'b0;  wr_cycle[ 7406] = 1'b1;  addr_rom[ 7406]='h00001684;  wr_data_rom[ 7406]='h00001515;
    rd_cycle[ 7407] = 1'b0;  wr_cycle[ 7407] = 1'b1;  addr_rom[ 7407]='h000011bc;  wr_data_rom[ 7407]='h00000a95;
    rd_cycle[ 7408] = 1'b0;  wr_cycle[ 7408] = 1'b1;  addr_rom[ 7408]='h000006e0;  wr_data_rom[ 7408]='h00000324;
    rd_cycle[ 7409] = 1'b0;  wr_cycle[ 7409] = 1'b1;  addr_rom[ 7409]='h00000240;  wr_data_rom[ 7409]='h00000243;
    rd_cycle[ 7410] = 1'b1;  wr_cycle[ 7410] = 1'b0;  addr_rom[ 7410]='h00000ac4;  wr_data_rom[ 7410]='h00000000;
    rd_cycle[ 7411] = 1'b0;  wr_cycle[ 7411] = 1'b1;  addr_rom[ 7411]='h00001730;  wr_data_rom[ 7411]='h0000188b;
    rd_cycle[ 7412] = 1'b1;  wr_cycle[ 7412] = 1'b0;  addr_rom[ 7412]='h00000244;  wr_data_rom[ 7412]='h00000000;
    rd_cycle[ 7413] = 1'b1;  wr_cycle[ 7413] = 1'b0;  addr_rom[ 7413]='h0000172c;  wr_data_rom[ 7413]='h00000000;
    rd_cycle[ 7414] = 1'b0;  wr_cycle[ 7414] = 1'b1;  addr_rom[ 7414]='h00001ad0;  wr_data_rom[ 7414]='h0000013f;
    rd_cycle[ 7415] = 1'b1;  wr_cycle[ 7415] = 1'b0;  addr_rom[ 7415]='h000012d0;  wr_data_rom[ 7415]='h00000000;
    rd_cycle[ 7416] = 1'b0;  wr_cycle[ 7416] = 1'b1;  addr_rom[ 7416]='h00000cc4;  wr_data_rom[ 7416]='h0000088c;
    rd_cycle[ 7417] = 1'b1;  wr_cycle[ 7417] = 1'b0;  addr_rom[ 7417]='h000007d0;  wr_data_rom[ 7417]='h00000000;
    rd_cycle[ 7418] = 1'b1;  wr_cycle[ 7418] = 1'b0;  addr_rom[ 7418]='h00000fdc;  wr_data_rom[ 7418]='h00000000;
    rd_cycle[ 7419] = 1'b0;  wr_cycle[ 7419] = 1'b1;  addr_rom[ 7419]='h00000f04;  wr_data_rom[ 7419]='h00000d0f;
    rd_cycle[ 7420] = 1'b1;  wr_cycle[ 7420] = 1'b0;  addr_rom[ 7420]='h000008ac;  wr_data_rom[ 7420]='h00000000;
    rd_cycle[ 7421] = 1'b0;  wr_cycle[ 7421] = 1'b1;  addr_rom[ 7421]='h000014d8;  wr_data_rom[ 7421]='h00000a3e;
    rd_cycle[ 7422] = 1'b0;  wr_cycle[ 7422] = 1'b1;  addr_rom[ 7422]='h00000c0c;  wr_data_rom[ 7422]='h00001cec;
    rd_cycle[ 7423] = 1'b1;  wr_cycle[ 7423] = 1'b0;  addr_rom[ 7423]='h00001ed0;  wr_data_rom[ 7423]='h00000000;
    rd_cycle[ 7424] = 1'b1;  wr_cycle[ 7424] = 1'b0;  addr_rom[ 7424]='h00000a00;  wr_data_rom[ 7424]='h00000000;
    rd_cycle[ 7425] = 1'b0;  wr_cycle[ 7425] = 1'b1;  addr_rom[ 7425]='h00001ae0;  wr_data_rom[ 7425]='h0000157c;
    rd_cycle[ 7426] = 1'b1;  wr_cycle[ 7426] = 1'b0;  addr_rom[ 7426]='h00001768;  wr_data_rom[ 7426]='h00000000;
    rd_cycle[ 7427] = 1'b0;  wr_cycle[ 7427] = 1'b1;  addr_rom[ 7427]='h00000e68;  wr_data_rom[ 7427]='h00001864;
    rd_cycle[ 7428] = 1'b1;  wr_cycle[ 7428] = 1'b0;  addr_rom[ 7428]='h00001d10;  wr_data_rom[ 7428]='h00000000;
    rd_cycle[ 7429] = 1'b1;  wr_cycle[ 7429] = 1'b0;  addr_rom[ 7429]='h00001b78;  wr_data_rom[ 7429]='h00000000;
    rd_cycle[ 7430] = 1'b1;  wr_cycle[ 7430] = 1'b0;  addr_rom[ 7430]='h00001e80;  wr_data_rom[ 7430]='h00000000;
    rd_cycle[ 7431] = 1'b0;  wr_cycle[ 7431] = 1'b1;  addr_rom[ 7431]='h000004b8;  wr_data_rom[ 7431]='h00000f3f;
    rd_cycle[ 7432] = 1'b1;  wr_cycle[ 7432] = 1'b0;  addr_rom[ 7432]='h00000ef8;  wr_data_rom[ 7432]='h00000000;
    rd_cycle[ 7433] = 1'b0;  wr_cycle[ 7433] = 1'b1;  addr_rom[ 7433]='h000015f0;  wr_data_rom[ 7433]='h0000178d;
    rd_cycle[ 7434] = 1'b1;  wr_cycle[ 7434] = 1'b0;  addr_rom[ 7434]='h000009c4;  wr_data_rom[ 7434]='h00000000;
    rd_cycle[ 7435] = 1'b0;  wr_cycle[ 7435] = 1'b1;  addr_rom[ 7435]='h00001138;  wr_data_rom[ 7435]='h00001457;
    rd_cycle[ 7436] = 1'b0;  wr_cycle[ 7436] = 1'b1;  addr_rom[ 7436]='h00000734;  wr_data_rom[ 7436]='h00001cf5;
    rd_cycle[ 7437] = 1'b0;  wr_cycle[ 7437] = 1'b1;  addr_rom[ 7437]='h00001180;  wr_data_rom[ 7437]='h000000a2;
    rd_cycle[ 7438] = 1'b0;  wr_cycle[ 7438] = 1'b1;  addr_rom[ 7438]='h0000059c;  wr_data_rom[ 7438]='h00000ab0;
    rd_cycle[ 7439] = 1'b0;  wr_cycle[ 7439] = 1'b1;  addr_rom[ 7439]='h00001b4c;  wr_data_rom[ 7439]='h000016fa;
    rd_cycle[ 7440] = 1'b0;  wr_cycle[ 7440] = 1'b1;  addr_rom[ 7440]='h00001450;  wr_data_rom[ 7440]='h00001def;
    rd_cycle[ 7441] = 1'b0;  wr_cycle[ 7441] = 1'b1;  addr_rom[ 7441]='h00001bc0;  wr_data_rom[ 7441]='h00000eb5;
    rd_cycle[ 7442] = 1'b1;  wr_cycle[ 7442] = 1'b0;  addr_rom[ 7442]='h00000ef8;  wr_data_rom[ 7442]='h00000000;
    rd_cycle[ 7443] = 1'b1;  wr_cycle[ 7443] = 1'b0;  addr_rom[ 7443]='h00000f14;  wr_data_rom[ 7443]='h00000000;
    rd_cycle[ 7444] = 1'b0;  wr_cycle[ 7444] = 1'b1;  addr_rom[ 7444]='h00000318;  wr_data_rom[ 7444]='h00001aa0;
    rd_cycle[ 7445] = 1'b0;  wr_cycle[ 7445] = 1'b1;  addr_rom[ 7445]='h000018dc;  wr_data_rom[ 7445]='h0000093a;
    rd_cycle[ 7446] = 1'b1;  wr_cycle[ 7446] = 1'b0;  addr_rom[ 7446]='h00000f00;  wr_data_rom[ 7446]='h00000000;
    rd_cycle[ 7447] = 1'b1;  wr_cycle[ 7447] = 1'b0;  addr_rom[ 7447]='h0000120c;  wr_data_rom[ 7447]='h00000000;
    rd_cycle[ 7448] = 1'b1;  wr_cycle[ 7448] = 1'b0;  addr_rom[ 7448]='h000019e0;  wr_data_rom[ 7448]='h00000000;
    rd_cycle[ 7449] = 1'b1;  wr_cycle[ 7449] = 1'b0;  addr_rom[ 7449]='h000004f4;  wr_data_rom[ 7449]='h00000000;
    rd_cycle[ 7450] = 1'b0;  wr_cycle[ 7450] = 1'b1;  addr_rom[ 7450]='h00001614;  wr_data_rom[ 7450]='h00001db6;
    rd_cycle[ 7451] = 1'b0;  wr_cycle[ 7451] = 1'b1;  addr_rom[ 7451]='h00001cd0;  wr_data_rom[ 7451]='h00001734;
    rd_cycle[ 7452] = 1'b1;  wr_cycle[ 7452] = 1'b0;  addr_rom[ 7452]='h00001bb8;  wr_data_rom[ 7452]='h00000000;
    rd_cycle[ 7453] = 1'b1;  wr_cycle[ 7453] = 1'b0;  addr_rom[ 7453]='h000010dc;  wr_data_rom[ 7453]='h00000000;
    rd_cycle[ 7454] = 1'b0;  wr_cycle[ 7454] = 1'b1;  addr_rom[ 7454]='h00000d64;  wr_data_rom[ 7454]='h00001ecf;
    rd_cycle[ 7455] = 1'b1;  wr_cycle[ 7455] = 1'b0;  addr_rom[ 7455]='h000016fc;  wr_data_rom[ 7455]='h00000000;
    rd_cycle[ 7456] = 1'b0;  wr_cycle[ 7456] = 1'b1;  addr_rom[ 7456]='h00000500;  wr_data_rom[ 7456]='h0000042a;
    rd_cycle[ 7457] = 1'b1;  wr_cycle[ 7457] = 1'b0;  addr_rom[ 7457]='h00000b9c;  wr_data_rom[ 7457]='h00000000;
    rd_cycle[ 7458] = 1'b1;  wr_cycle[ 7458] = 1'b0;  addr_rom[ 7458]='h000009fc;  wr_data_rom[ 7458]='h00000000;
    rd_cycle[ 7459] = 1'b1;  wr_cycle[ 7459] = 1'b0;  addr_rom[ 7459]='h000008d0;  wr_data_rom[ 7459]='h00000000;
    rd_cycle[ 7460] = 1'b1;  wr_cycle[ 7460] = 1'b0;  addr_rom[ 7460]='h00001714;  wr_data_rom[ 7460]='h00000000;
    rd_cycle[ 7461] = 1'b0;  wr_cycle[ 7461] = 1'b1;  addr_rom[ 7461]='h00001ebc;  wr_data_rom[ 7461]='h00000a2a;
    rd_cycle[ 7462] = 1'b1;  wr_cycle[ 7462] = 1'b0;  addr_rom[ 7462]='h00001c80;  wr_data_rom[ 7462]='h00000000;
    rd_cycle[ 7463] = 1'b0;  wr_cycle[ 7463] = 1'b1;  addr_rom[ 7463]='h00000180;  wr_data_rom[ 7463]='h00000a68;
    rd_cycle[ 7464] = 1'b1;  wr_cycle[ 7464] = 1'b0;  addr_rom[ 7464]='h00001ca4;  wr_data_rom[ 7464]='h00000000;
    rd_cycle[ 7465] = 1'b0;  wr_cycle[ 7465] = 1'b1;  addr_rom[ 7465]='h00001b7c;  wr_data_rom[ 7465]='h00001c92;
    rd_cycle[ 7466] = 1'b1;  wr_cycle[ 7466] = 1'b0;  addr_rom[ 7466]='h00000670;  wr_data_rom[ 7466]='h00000000;
    rd_cycle[ 7467] = 1'b0;  wr_cycle[ 7467] = 1'b1;  addr_rom[ 7467]='h00000d30;  wr_data_rom[ 7467]='h0000126a;
    rd_cycle[ 7468] = 1'b0;  wr_cycle[ 7468] = 1'b1;  addr_rom[ 7468]='h00000090;  wr_data_rom[ 7468]='h0000078a;
    rd_cycle[ 7469] = 1'b0;  wr_cycle[ 7469] = 1'b1;  addr_rom[ 7469]='h000004dc;  wr_data_rom[ 7469]='h00001aa7;
    rd_cycle[ 7470] = 1'b0;  wr_cycle[ 7470] = 1'b1;  addr_rom[ 7470]='h00001340;  wr_data_rom[ 7470]='h00001b61;
    rd_cycle[ 7471] = 1'b1;  wr_cycle[ 7471] = 1'b0;  addr_rom[ 7471]='h00001a7c;  wr_data_rom[ 7471]='h00000000;
    rd_cycle[ 7472] = 1'b0;  wr_cycle[ 7472] = 1'b1;  addr_rom[ 7472]='h00000450;  wr_data_rom[ 7472]='h00000096;
    rd_cycle[ 7473] = 1'b0;  wr_cycle[ 7473] = 1'b1;  addr_rom[ 7473]='h000012b0;  wr_data_rom[ 7473]='h000002f6;
    rd_cycle[ 7474] = 1'b1;  wr_cycle[ 7474] = 1'b0;  addr_rom[ 7474]='h00000c64;  wr_data_rom[ 7474]='h00000000;
    rd_cycle[ 7475] = 1'b1;  wr_cycle[ 7475] = 1'b0;  addr_rom[ 7475]='h0000163c;  wr_data_rom[ 7475]='h00000000;
    rd_cycle[ 7476] = 1'b0;  wr_cycle[ 7476] = 1'b1;  addr_rom[ 7476]='h000010f4;  wr_data_rom[ 7476]='h000015c9;
    rd_cycle[ 7477] = 1'b0;  wr_cycle[ 7477] = 1'b1;  addr_rom[ 7477]='h0000032c;  wr_data_rom[ 7477]='h00001e03;
    rd_cycle[ 7478] = 1'b0;  wr_cycle[ 7478] = 1'b1;  addr_rom[ 7478]='h000019f8;  wr_data_rom[ 7478]='h00000a4a;
    rd_cycle[ 7479] = 1'b0;  wr_cycle[ 7479] = 1'b1;  addr_rom[ 7479]='h00001440;  wr_data_rom[ 7479]='h00001698;
    rd_cycle[ 7480] = 1'b1;  wr_cycle[ 7480] = 1'b0;  addr_rom[ 7480]='h00000e98;  wr_data_rom[ 7480]='h00000000;
    rd_cycle[ 7481] = 1'b1;  wr_cycle[ 7481] = 1'b0;  addr_rom[ 7481]='h00000818;  wr_data_rom[ 7481]='h00000000;
    rd_cycle[ 7482] = 1'b1;  wr_cycle[ 7482] = 1'b0;  addr_rom[ 7482]='h00000ba4;  wr_data_rom[ 7482]='h00000000;
    rd_cycle[ 7483] = 1'b1;  wr_cycle[ 7483] = 1'b0;  addr_rom[ 7483]='h00001720;  wr_data_rom[ 7483]='h00000000;
    rd_cycle[ 7484] = 1'b1;  wr_cycle[ 7484] = 1'b0;  addr_rom[ 7484]='h00000374;  wr_data_rom[ 7484]='h00000000;
    rd_cycle[ 7485] = 1'b1;  wr_cycle[ 7485] = 1'b0;  addr_rom[ 7485]='h0000075c;  wr_data_rom[ 7485]='h00000000;
    rd_cycle[ 7486] = 1'b1;  wr_cycle[ 7486] = 1'b0;  addr_rom[ 7486]='h000002e4;  wr_data_rom[ 7486]='h00000000;
    rd_cycle[ 7487] = 1'b0;  wr_cycle[ 7487] = 1'b1;  addr_rom[ 7487]='h00000fc4;  wr_data_rom[ 7487]='h00001af7;
    rd_cycle[ 7488] = 1'b1;  wr_cycle[ 7488] = 1'b0;  addr_rom[ 7488]='h0000053c;  wr_data_rom[ 7488]='h00000000;
    rd_cycle[ 7489] = 1'b1;  wr_cycle[ 7489] = 1'b0;  addr_rom[ 7489]='h000014c0;  wr_data_rom[ 7489]='h00000000;
    rd_cycle[ 7490] = 1'b0;  wr_cycle[ 7490] = 1'b1;  addr_rom[ 7490]='h00001620;  wr_data_rom[ 7490]='h00001c7c;
    rd_cycle[ 7491] = 1'b0;  wr_cycle[ 7491] = 1'b1;  addr_rom[ 7491]='h00000d3c;  wr_data_rom[ 7491]='h00001b4d;
    rd_cycle[ 7492] = 1'b0;  wr_cycle[ 7492] = 1'b1;  addr_rom[ 7492]='h000002d4;  wr_data_rom[ 7492]='h00001f2c;
    rd_cycle[ 7493] = 1'b1;  wr_cycle[ 7493] = 1'b0;  addr_rom[ 7493]='h0000029c;  wr_data_rom[ 7493]='h00000000;
    rd_cycle[ 7494] = 1'b1;  wr_cycle[ 7494] = 1'b0;  addr_rom[ 7494]='h00000540;  wr_data_rom[ 7494]='h00000000;
    rd_cycle[ 7495] = 1'b1;  wr_cycle[ 7495] = 1'b0;  addr_rom[ 7495]='h0000032c;  wr_data_rom[ 7495]='h00000000;
    rd_cycle[ 7496] = 1'b1;  wr_cycle[ 7496] = 1'b0;  addr_rom[ 7496]='h0000120c;  wr_data_rom[ 7496]='h00000000;
    rd_cycle[ 7497] = 1'b0;  wr_cycle[ 7497] = 1'b1;  addr_rom[ 7497]='h000015b8;  wr_data_rom[ 7497]='h000008d5;
    rd_cycle[ 7498] = 1'b1;  wr_cycle[ 7498] = 1'b0;  addr_rom[ 7498]='h000016bc;  wr_data_rom[ 7498]='h00000000;
    rd_cycle[ 7499] = 1'b0;  wr_cycle[ 7499] = 1'b1;  addr_rom[ 7499]='h0000093c;  wr_data_rom[ 7499]='h000003af;
    rd_cycle[ 7500] = 1'b0;  wr_cycle[ 7500] = 1'b1;  addr_rom[ 7500]='h00001cb8;  wr_data_rom[ 7500]='h00000ea1;
    rd_cycle[ 7501] = 1'b1;  wr_cycle[ 7501] = 1'b0;  addr_rom[ 7501]='h00000fdc;  wr_data_rom[ 7501]='h00000000;
    rd_cycle[ 7502] = 1'b1;  wr_cycle[ 7502] = 1'b0;  addr_rom[ 7502]='h000003b4;  wr_data_rom[ 7502]='h00000000;
    rd_cycle[ 7503] = 1'b1;  wr_cycle[ 7503] = 1'b0;  addr_rom[ 7503]='h00001a68;  wr_data_rom[ 7503]='h00000000;
    rd_cycle[ 7504] = 1'b1;  wr_cycle[ 7504] = 1'b0;  addr_rom[ 7504]='h00001134;  wr_data_rom[ 7504]='h00000000;
    rd_cycle[ 7505] = 1'b0;  wr_cycle[ 7505] = 1'b1;  addr_rom[ 7505]='h00000078;  wr_data_rom[ 7505]='h0000127b;
    rd_cycle[ 7506] = 1'b0;  wr_cycle[ 7506] = 1'b1;  addr_rom[ 7506]='h00001528;  wr_data_rom[ 7506]='h000007a8;
    rd_cycle[ 7507] = 1'b1;  wr_cycle[ 7507] = 1'b0;  addr_rom[ 7507]='h00001ea0;  wr_data_rom[ 7507]='h00000000;
    rd_cycle[ 7508] = 1'b1;  wr_cycle[ 7508] = 1'b0;  addr_rom[ 7508]='h00000ae4;  wr_data_rom[ 7508]='h00000000;
    rd_cycle[ 7509] = 1'b0;  wr_cycle[ 7509] = 1'b1;  addr_rom[ 7509]='h000000ec;  wr_data_rom[ 7509]='h00000008;
    rd_cycle[ 7510] = 1'b1;  wr_cycle[ 7510] = 1'b0;  addr_rom[ 7510]='h00001370;  wr_data_rom[ 7510]='h00000000;
    rd_cycle[ 7511] = 1'b1;  wr_cycle[ 7511] = 1'b0;  addr_rom[ 7511]='h00001f04;  wr_data_rom[ 7511]='h00000000;
    rd_cycle[ 7512] = 1'b0;  wr_cycle[ 7512] = 1'b1;  addr_rom[ 7512]='h000001d0;  wr_data_rom[ 7512]='h00001eac;
    rd_cycle[ 7513] = 1'b0;  wr_cycle[ 7513] = 1'b1;  addr_rom[ 7513]='h00000d5c;  wr_data_rom[ 7513]='h00001c5a;
    rd_cycle[ 7514] = 1'b0;  wr_cycle[ 7514] = 1'b1;  addr_rom[ 7514]='h00000320;  wr_data_rom[ 7514]='h00000996;
    rd_cycle[ 7515] = 1'b0;  wr_cycle[ 7515] = 1'b1;  addr_rom[ 7515]='h00001058;  wr_data_rom[ 7515]='h0000188b;
    rd_cycle[ 7516] = 1'b0;  wr_cycle[ 7516] = 1'b1;  addr_rom[ 7516]='h00000634;  wr_data_rom[ 7516]='h00000cce;
    rd_cycle[ 7517] = 1'b1;  wr_cycle[ 7517] = 1'b0;  addr_rom[ 7517]='h00001dc0;  wr_data_rom[ 7517]='h00000000;
    rd_cycle[ 7518] = 1'b1;  wr_cycle[ 7518] = 1'b0;  addr_rom[ 7518]='h00001258;  wr_data_rom[ 7518]='h00000000;
    rd_cycle[ 7519] = 1'b0;  wr_cycle[ 7519] = 1'b1;  addr_rom[ 7519]='h000009a0;  wr_data_rom[ 7519]='h00000293;
    rd_cycle[ 7520] = 1'b1;  wr_cycle[ 7520] = 1'b0;  addr_rom[ 7520]='h00000240;  wr_data_rom[ 7520]='h00000000;
    rd_cycle[ 7521] = 1'b1;  wr_cycle[ 7521] = 1'b0;  addr_rom[ 7521]='h000011d8;  wr_data_rom[ 7521]='h00000000;
    rd_cycle[ 7522] = 1'b0;  wr_cycle[ 7522] = 1'b1;  addr_rom[ 7522]='h00000b20;  wr_data_rom[ 7522]='h00001ae8;
    rd_cycle[ 7523] = 1'b1;  wr_cycle[ 7523] = 1'b0;  addr_rom[ 7523]='h00001410;  wr_data_rom[ 7523]='h00000000;
    rd_cycle[ 7524] = 1'b1;  wr_cycle[ 7524] = 1'b0;  addr_rom[ 7524]='h00001758;  wr_data_rom[ 7524]='h00000000;
    rd_cycle[ 7525] = 1'b1;  wr_cycle[ 7525] = 1'b0;  addr_rom[ 7525]='h00000a80;  wr_data_rom[ 7525]='h00000000;
    rd_cycle[ 7526] = 1'b1;  wr_cycle[ 7526] = 1'b0;  addr_rom[ 7526]='h00000270;  wr_data_rom[ 7526]='h00000000;
    rd_cycle[ 7527] = 1'b0;  wr_cycle[ 7527] = 1'b1;  addr_rom[ 7527]='h00001ed4;  wr_data_rom[ 7527]='h00001661;
    rd_cycle[ 7528] = 1'b0;  wr_cycle[ 7528] = 1'b1;  addr_rom[ 7528]='h000002d0;  wr_data_rom[ 7528]='h00000fde;
    rd_cycle[ 7529] = 1'b1;  wr_cycle[ 7529] = 1'b0;  addr_rom[ 7529]='h00001014;  wr_data_rom[ 7529]='h00000000;
    rd_cycle[ 7530] = 1'b0;  wr_cycle[ 7530] = 1'b1;  addr_rom[ 7530]='h0000031c;  wr_data_rom[ 7530]='h00000fd7;
    rd_cycle[ 7531] = 1'b0;  wr_cycle[ 7531] = 1'b1;  addr_rom[ 7531]='h00001c80;  wr_data_rom[ 7531]='h00001d44;
    rd_cycle[ 7532] = 1'b0;  wr_cycle[ 7532] = 1'b1;  addr_rom[ 7532]='h00000b94;  wr_data_rom[ 7532]='h00000dde;
    rd_cycle[ 7533] = 1'b0;  wr_cycle[ 7533] = 1'b1;  addr_rom[ 7533]='h000004d0;  wr_data_rom[ 7533]='h00001ce1;
    rd_cycle[ 7534] = 1'b1;  wr_cycle[ 7534] = 1'b0;  addr_rom[ 7534]='h00001290;  wr_data_rom[ 7534]='h00000000;
    rd_cycle[ 7535] = 1'b0;  wr_cycle[ 7535] = 1'b1;  addr_rom[ 7535]='h00001874;  wr_data_rom[ 7535]='h00000bdb;
    rd_cycle[ 7536] = 1'b1;  wr_cycle[ 7536] = 1'b0;  addr_rom[ 7536]='h00001194;  wr_data_rom[ 7536]='h00000000;
    rd_cycle[ 7537] = 1'b0;  wr_cycle[ 7537] = 1'b1;  addr_rom[ 7537]='h0000103c;  wr_data_rom[ 7537]='h0000166e;
    rd_cycle[ 7538] = 1'b1;  wr_cycle[ 7538] = 1'b0;  addr_rom[ 7538]='h00001124;  wr_data_rom[ 7538]='h00000000;
    rd_cycle[ 7539] = 1'b0;  wr_cycle[ 7539] = 1'b1;  addr_rom[ 7539]='h0000010c;  wr_data_rom[ 7539]='h00001002;
    rd_cycle[ 7540] = 1'b1;  wr_cycle[ 7540] = 1'b0;  addr_rom[ 7540]='h00001454;  wr_data_rom[ 7540]='h00000000;
    rd_cycle[ 7541] = 1'b1;  wr_cycle[ 7541] = 1'b0;  addr_rom[ 7541]='h00000650;  wr_data_rom[ 7541]='h00000000;
    rd_cycle[ 7542] = 1'b0;  wr_cycle[ 7542] = 1'b1;  addr_rom[ 7542]='h00000448;  wr_data_rom[ 7542]='h00001095;
    rd_cycle[ 7543] = 1'b1;  wr_cycle[ 7543] = 1'b0;  addr_rom[ 7543]='h00001150;  wr_data_rom[ 7543]='h00000000;
    rd_cycle[ 7544] = 1'b1;  wr_cycle[ 7544] = 1'b0;  addr_rom[ 7544]='h00000aac;  wr_data_rom[ 7544]='h00000000;
    rd_cycle[ 7545] = 1'b0;  wr_cycle[ 7545] = 1'b1;  addr_rom[ 7545]='h00001b14;  wr_data_rom[ 7545]='h00000777;
    rd_cycle[ 7546] = 1'b1;  wr_cycle[ 7546] = 1'b0;  addr_rom[ 7546]='h000007d4;  wr_data_rom[ 7546]='h00000000;
    rd_cycle[ 7547] = 1'b1;  wr_cycle[ 7547] = 1'b0;  addr_rom[ 7547]='h00000ac8;  wr_data_rom[ 7547]='h00000000;
    rd_cycle[ 7548] = 1'b1;  wr_cycle[ 7548] = 1'b0;  addr_rom[ 7548]='h000001d8;  wr_data_rom[ 7548]='h00000000;
    rd_cycle[ 7549] = 1'b1;  wr_cycle[ 7549] = 1'b0;  addr_rom[ 7549]='h00001c58;  wr_data_rom[ 7549]='h00000000;
    rd_cycle[ 7550] = 1'b1;  wr_cycle[ 7550] = 1'b0;  addr_rom[ 7550]='h00000994;  wr_data_rom[ 7550]='h00000000;
    rd_cycle[ 7551] = 1'b0;  wr_cycle[ 7551] = 1'b1;  addr_rom[ 7551]='h00001344;  wr_data_rom[ 7551]='h000019a2;
    rd_cycle[ 7552] = 1'b1;  wr_cycle[ 7552] = 1'b0;  addr_rom[ 7552]='h00000238;  wr_data_rom[ 7552]='h00000000;
    rd_cycle[ 7553] = 1'b0;  wr_cycle[ 7553] = 1'b1;  addr_rom[ 7553]='h00000bf4;  wr_data_rom[ 7553]='h0000044b;
    rd_cycle[ 7554] = 1'b0;  wr_cycle[ 7554] = 1'b1;  addr_rom[ 7554]='h00000df4;  wr_data_rom[ 7554]='h00000b73;
    rd_cycle[ 7555] = 1'b0;  wr_cycle[ 7555] = 1'b1;  addr_rom[ 7555]='h0000033c;  wr_data_rom[ 7555]='h000000fe;
    rd_cycle[ 7556] = 1'b1;  wr_cycle[ 7556] = 1'b0;  addr_rom[ 7556]='h00000e90;  wr_data_rom[ 7556]='h00000000;
    rd_cycle[ 7557] = 1'b0;  wr_cycle[ 7557] = 1'b1;  addr_rom[ 7557]='h00001ed0;  wr_data_rom[ 7557]='h0000108e;
    rd_cycle[ 7558] = 1'b0;  wr_cycle[ 7558] = 1'b1;  addr_rom[ 7558]='h000003a8;  wr_data_rom[ 7558]='h000009ef;
    rd_cycle[ 7559] = 1'b1;  wr_cycle[ 7559] = 1'b0;  addr_rom[ 7559]='h00001d40;  wr_data_rom[ 7559]='h00000000;
    rd_cycle[ 7560] = 1'b0;  wr_cycle[ 7560] = 1'b1;  addr_rom[ 7560]='h000012b8;  wr_data_rom[ 7560]='h00001f0d;
    rd_cycle[ 7561] = 1'b1;  wr_cycle[ 7561] = 1'b0;  addr_rom[ 7561]='h00001aa4;  wr_data_rom[ 7561]='h00000000;
    rd_cycle[ 7562] = 1'b0;  wr_cycle[ 7562] = 1'b1;  addr_rom[ 7562]='h00000b98;  wr_data_rom[ 7562]='h0000011d;
    rd_cycle[ 7563] = 1'b0;  wr_cycle[ 7563] = 1'b1;  addr_rom[ 7563]='h000009f4;  wr_data_rom[ 7563]='h000019c0;
    rd_cycle[ 7564] = 1'b0;  wr_cycle[ 7564] = 1'b1;  addr_rom[ 7564]='h00000e00;  wr_data_rom[ 7564]='h000009b6;
    rd_cycle[ 7565] = 1'b0;  wr_cycle[ 7565] = 1'b1;  addr_rom[ 7565]='h000003d4;  wr_data_rom[ 7565]='h00001247;
    rd_cycle[ 7566] = 1'b0;  wr_cycle[ 7566] = 1'b1;  addr_rom[ 7566]='h000001f8;  wr_data_rom[ 7566]='h00001f2e;
    rd_cycle[ 7567] = 1'b0;  wr_cycle[ 7567] = 1'b1;  addr_rom[ 7567]='h00001dc0;  wr_data_rom[ 7567]='h00000654;
    rd_cycle[ 7568] = 1'b1;  wr_cycle[ 7568] = 1'b0;  addr_rom[ 7568]='h000006b8;  wr_data_rom[ 7568]='h00000000;
    rd_cycle[ 7569] = 1'b1;  wr_cycle[ 7569] = 1'b0;  addr_rom[ 7569]='h000013e8;  wr_data_rom[ 7569]='h00000000;
    rd_cycle[ 7570] = 1'b0;  wr_cycle[ 7570] = 1'b1;  addr_rom[ 7570]='h00001034;  wr_data_rom[ 7570]='h00001c38;
    rd_cycle[ 7571] = 1'b1;  wr_cycle[ 7571] = 1'b0;  addr_rom[ 7571]='h00001c54;  wr_data_rom[ 7571]='h00000000;
    rd_cycle[ 7572] = 1'b1;  wr_cycle[ 7572] = 1'b0;  addr_rom[ 7572]='h00000ec4;  wr_data_rom[ 7572]='h00000000;
    rd_cycle[ 7573] = 1'b1;  wr_cycle[ 7573] = 1'b0;  addr_rom[ 7573]='h00001854;  wr_data_rom[ 7573]='h00000000;
    rd_cycle[ 7574] = 1'b0;  wr_cycle[ 7574] = 1'b1;  addr_rom[ 7574]='h000000c8;  wr_data_rom[ 7574]='h0000197f;
    rd_cycle[ 7575] = 1'b0;  wr_cycle[ 7575] = 1'b1;  addr_rom[ 7575]='h00001e6c;  wr_data_rom[ 7575]='h0000091c;
    rd_cycle[ 7576] = 1'b1;  wr_cycle[ 7576] = 1'b0;  addr_rom[ 7576]='h000019b4;  wr_data_rom[ 7576]='h00000000;
    rd_cycle[ 7577] = 1'b0;  wr_cycle[ 7577] = 1'b1;  addr_rom[ 7577]='h000010a8;  wr_data_rom[ 7577]='h00001edd;
    rd_cycle[ 7578] = 1'b0;  wr_cycle[ 7578] = 1'b1;  addr_rom[ 7578]='h000016ac;  wr_data_rom[ 7578]='h00001eaf;
    rd_cycle[ 7579] = 1'b1;  wr_cycle[ 7579] = 1'b0;  addr_rom[ 7579]='h0000073c;  wr_data_rom[ 7579]='h00000000;
    rd_cycle[ 7580] = 1'b0;  wr_cycle[ 7580] = 1'b1;  addr_rom[ 7580]='h00000b00;  wr_data_rom[ 7580]='h0000140c;
    rd_cycle[ 7581] = 1'b1;  wr_cycle[ 7581] = 1'b0;  addr_rom[ 7581]='h0000093c;  wr_data_rom[ 7581]='h00000000;
    rd_cycle[ 7582] = 1'b1;  wr_cycle[ 7582] = 1'b0;  addr_rom[ 7582]='h0000156c;  wr_data_rom[ 7582]='h00000000;
    rd_cycle[ 7583] = 1'b0;  wr_cycle[ 7583] = 1'b1;  addr_rom[ 7583]='h00001314;  wr_data_rom[ 7583]='h00000f82;
    rd_cycle[ 7584] = 1'b1;  wr_cycle[ 7584] = 1'b0;  addr_rom[ 7584]='h00001b1c;  wr_data_rom[ 7584]='h00000000;
    rd_cycle[ 7585] = 1'b0;  wr_cycle[ 7585] = 1'b1;  addr_rom[ 7585]='h0000156c;  wr_data_rom[ 7585]='h00001b72;
    rd_cycle[ 7586] = 1'b0;  wr_cycle[ 7586] = 1'b1;  addr_rom[ 7586]='h00000034;  wr_data_rom[ 7586]='h00001b9b;
    rd_cycle[ 7587] = 1'b0;  wr_cycle[ 7587] = 1'b1;  addr_rom[ 7587]='h00000360;  wr_data_rom[ 7587]='h00000462;
    rd_cycle[ 7588] = 1'b1;  wr_cycle[ 7588] = 1'b0;  addr_rom[ 7588]='h000006cc;  wr_data_rom[ 7588]='h00000000;
    rd_cycle[ 7589] = 1'b0;  wr_cycle[ 7589] = 1'b1;  addr_rom[ 7589]='h00000454;  wr_data_rom[ 7589]='h00000eb3;
    rd_cycle[ 7590] = 1'b0;  wr_cycle[ 7590] = 1'b1;  addr_rom[ 7590]='h00001364;  wr_data_rom[ 7590]='h000017f6;
    rd_cycle[ 7591] = 1'b1;  wr_cycle[ 7591] = 1'b0;  addr_rom[ 7591]='h00000bf0;  wr_data_rom[ 7591]='h00000000;
    rd_cycle[ 7592] = 1'b1;  wr_cycle[ 7592] = 1'b0;  addr_rom[ 7592]='h00001c10;  wr_data_rom[ 7592]='h00000000;
    rd_cycle[ 7593] = 1'b0;  wr_cycle[ 7593] = 1'b1;  addr_rom[ 7593]='h000014b0;  wr_data_rom[ 7593]='h00001036;
    rd_cycle[ 7594] = 1'b0;  wr_cycle[ 7594] = 1'b1;  addr_rom[ 7594]='h0000064c;  wr_data_rom[ 7594]='h000007c8;
    rd_cycle[ 7595] = 1'b0;  wr_cycle[ 7595] = 1'b1;  addr_rom[ 7595]='h000019cc;  wr_data_rom[ 7595]='h00000681;
    rd_cycle[ 7596] = 1'b0;  wr_cycle[ 7596] = 1'b1;  addr_rom[ 7596]='h00000190;  wr_data_rom[ 7596]='h00001590;
    rd_cycle[ 7597] = 1'b0;  wr_cycle[ 7597] = 1'b1;  addr_rom[ 7597]='h00001c0c;  wr_data_rom[ 7597]='h00000efb;
    rd_cycle[ 7598] = 1'b1;  wr_cycle[ 7598] = 1'b0;  addr_rom[ 7598]='h000001e8;  wr_data_rom[ 7598]='h00000000;
    rd_cycle[ 7599] = 1'b0;  wr_cycle[ 7599] = 1'b1;  addr_rom[ 7599]='h00000268;  wr_data_rom[ 7599]='h00000070;
    rd_cycle[ 7600] = 1'b0;  wr_cycle[ 7600] = 1'b1;  addr_rom[ 7600]='h0000137c;  wr_data_rom[ 7600]='h000010ed;
    rd_cycle[ 7601] = 1'b0;  wr_cycle[ 7601] = 1'b1;  addr_rom[ 7601]='h000001e8;  wr_data_rom[ 7601]='h000004eb;
    rd_cycle[ 7602] = 1'b1;  wr_cycle[ 7602] = 1'b0;  addr_rom[ 7602]='h00001da4;  wr_data_rom[ 7602]='h00000000;
    rd_cycle[ 7603] = 1'b0;  wr_cycle[ 7603] = 1'b1;  addr_rom[ 7603]='h00000bf0;  wr_data_rom[ 7603]='h00000a6a;
    rd_cycle[ 7604] = 1'b0;  wr_cycle[ 7604] = 1'b1;  addr_rom[ 7604]='h000019c4;  wr_data_rom[ 7604]='h000016c3;
    rd_cycle[ 7605] = 1'b0;  wr_cycle[ 7605] = 1'b1;  addr_rom[ 7605]='h00000170;  wr_data_rom[ 7605]='h0000062f;
    rd_cycle[ 7606] = 1'b1;  wr_cycle[ 7606] = 1'b0;  addr_rom[ 7606]='h00000920;  wr_data_rom[ 7606]='h00000000;
    rd_cycle[ 7607] = 1'b1;  wr_cycle[ 7607] = 1'b0;  addr_rom[ 7607]='h0000080c;  wr_data_rom[ 7607]='h00000000;
    rd_cycle[ 7608] = 1'b1;  wr_cycle[ 7608] = 1'b0;  addr_rom[ 7608]='h00001074;  wr_data_rom[ 7608]='h00000000;
    rd_cycle[ 7609] = 1'b1;  wr_cycle[ 7609] = 1'b0;  addr_rom[ 7609]='h000009cc;  wr_data_rom[ 7609]='h00000000;
    rd_cycle[ 7610] = 1'b1;  wr_cycle[ 7610] = 1'b0;  addr_rom[ 7610]='h00001a18;  wr_data_rom[ 7610]='h00000000;
    rd_cycle[ 7611] = 1'b1;  wr_cycle[ 7611] = 1'b0;  addr_rom[ 7611]='h000019b4;  wr_data_rom[ 7611]='h00000000;
    rd_cycle[ 7612] = 1'b1;  wr_cycle[ 7612] = 1'b0;  addr_rom[ 7612]='h0000135c;  wr_data_rom[ 7612]='h00000000;
    rd_cycle[ 7613] = 1'b1;  wr_cycle[ 7613] = 1'b0;  addr_rom[ 7613]='h000016d8;  wr_data_rom[ 7613]='h00000000;
    rd_cycle[ 7614] = 1'b1;  wr_cycle[ 7614] = 1'b0;  addr_rom[ 7614]='h00001d64;  wr_data_rom[ 7614]='h00000000;
    rd_cycle[ 7615] = 1'b0;  wr_cycle[ 7615] = 1'b1;  addr_rom[ 7615]='h000019e8;  wr_data_rom[ 7615]='h0000123e;
    rd_cycle[ 7616] = 1'b0;  wr_cycle[ 7616] = 1'b1;  addr_rom[ 7616]='h00001e6c;  wr_data_rom[ 7616]='h00001cb8;
    rd_cycle[ 7617] = 1'b1;  wr_cycle[ 7617] = 1'b0;  addr_rom[ 7617]='h0000121c;  wr_data_rom[ 7617]='h00000000;
    rd_cycle[ 7618] = 1'b0;  wr_cycle[ 7618] = 1'b1;  addr_rom[ 7618]='h00000e20;  wr_data_rom[ 7618]='h00000f95;
    rd_cycle[ 7619] = 1'b1;  wr_cycle[ 7619] = 1'b0;  addr_rom[ 7619]='h000010e0;  wr_data_rom[ 7619]='h00000000;
    rd_cycle[ 7620] = 1'b0;  wr_cycle[ 7620] = 1'b1;  addr_rom[ 7620]='h00000158;  wr_data_rom[ 7620]='h00000cd9;
    rd_cycle[ 7621] = 1'b1;  wr_cycle[ 7621] = 1'b0;  addr_rom[ 7621]='h000013f8;  wr_data_rom[ 7621]='h00000000;
    rd_cycle[ 7622] = 1'b1;  wr_cycle[ 7622] = 1'b0;  addr_rom[ 7622]='h00000674;  wr_data_rom[ 7622]='h00000000;
    rd_cycle[ 7623] = 1'b1;  wr_cycle[ 7623] = 1'b0;  addr_rom[ 7623]='h000019b4;  wr_data_rom[ 7623]='h00000000;
    rd_cycle[ 7624] = 1'b1;  wr_cycle[ 7624] = 1'b0;  addr_rom[ 7624]='h00001620;  wr_data_rom[ 7624]='h00000000;
    rd_cycle[ 7625] = 1'b0;  wr_cycle[ 7625] = 1'b1;  addr_rom[ 7625]='h000005b8;  wr_data_rom[ 7625]='h00001979;
    rd_cycle[ 7626] = 1'b0;  wr_cycle[ 7626] = 1'b1;  addr_rom[ 7626]='h00001ea8;  wr_data_rom[ 7626]='h0000171c;
    rd_cycle[ 7627] = 1'b0;  wr_cycle[ 7627] = 1'b1;  addr_rom[ 7627]='h000008b4;  wr_data_rom[ 7627]='h0000046b;
    rd_cycle[ 7628] = 1'b0;  wr_cycle[ 7628] = 1'b1;  addr_rom[ 7628]='h00001c90;  wr_data_rom[ 7628]='h00000916;
    rd_cycle[ 7629] = 1'b0;  wr_cycle[ 7629] = 1'b1;  addr_rom[ 7629]='h000003b4;  wr_data_rom[ 7629]='h00001216;
    rd_cycle[ 7630] = 1'b0;  wr_cycle[ 7630] = 1'b1;  addr_rom[ 7630]='h00000f2c;  wr_data_rom[ 7630]='h000015a3;
    rd_cycle[ 7631] = 1'b1;  wr_cycle[ 7631] = 1'b0;  addr_rom[ 7631]='h00001b3c;  wr_data_rom[ 7631]='h00000000;
    rd_cycle[ 7632] = 1'b0;  wr_cycle[ 7632] = 1'b1;  addr_rom[ 7632]='h00000600;  wr_data_rom[ 7632]='h000005e8;
    rd_cycle[ 7633] = 1'b0;  wr_cycle[ 7633] = 1'b1;  addr_rom[ 7633]='h000010b0;  wr_data_rom[ 7633]='h00001d69;
    rd_cycle[ 7634] = 1'b1;  wr_cycle[ 7634] = 1'b0;  addr_rom[ 7634]='h00000498;  wr_data_rom[ 7634]='h00000000;
    rd_cycle[ 7635] = 1'b1;  wr_cycle[ 7635] = 1'b0;  addr_rom[ 7635]='h00000228;  wr_data_rom[ 7635]='h00000000;
    rd_cycle[ 7636] = 1'b1;  wr_cycle[ 7636] = 1'b0;  addr_rom[ 7636]='h00000a4c;  wr_data_rom[ 7636]='h00000000;
    rd_cycle[ 7637] = 1'b1;  wr_cycle[ 7637] = 1'b0;  addr_rom[ 7637]='h00000860;  wr_data_rom[ 7637]='h00000000;
    rd_cycle[ 7638] = 1'b0;  wr_cycle[ 7638] = 1'b1;  addr_rom[ 7638]='h0000098c;  wr_data_rom[ 7638]='h00001171;
    rd_cycle[ 7639] = 1'b1;  wr_cycle[ 7639] = 1'b0;  addr_rom[ 7639]='h00001a2c;  wr_data_rom[ 7639]='h00000000;
    rd_cycle[ 7640] = 1'b0;  wr_cycle[ 7640] = 1'b1;  addr_rom[ 7640]='h00001198;  wr_data_rom[ 7640]='h00001d78;
    rd_cycle[ 7641] = 1'b0;  wr_cycle[ 7641] = 1'b1;  addr_rom[ 7641]='h00001794;  wr_data_rom[ 7641]='h00001e89;
    rd_cycle[ 7642] = 1'b1;  wr_cycle[ 7642] = 1'b0;  addr_rom[ 7642]='h000015bc;  wr_data_rom[ 7642]='h00000000;
    rd_cycle[ 7643] = 1'b0;  wr_cycle[ 7643] = 1'b1;  addr_rom[ 7643]='h00000ff0;  wr_data_rom[ 7643]='h00000bfc;
    rd_cycle[ 7644] = 1'b0;  wr_cycle[ 7644] = 1'b1;  addr_rom[ 7644]='h00001e6c;  wr_data_rom[ 7644]='h000000eb;
    rd_cycle[ 7645] = 1'b1;  wr_cycle[ 7645] = 1'b0;  addr_rom[ 7645]='h000016f8;  wr_data_rom[ 7645]='h00000000;
    rd_cycle[ 7646] = 1'b0;  wr_cycle[ 7646] = 1'b1;  addr_rom[ 7646]='h00000620;  wr_data_rom[ 7646]='h00000dda;
    rd_cycle[ 7647] = 1'b1;  wr_cycle[ 7647] = 1'b0;  addr_rom[ 7647]='h0000035c;  wr_data_rom[ 7647]='h00000000;
    rd_cycle[ 7648] = 1'b0;  wr_cycle[ 7648] = 1'b1;  addr_rom[ 7648]='h00000f74;  wr_data_rom[ 7648]='h00000bc1;
    rd_cycle[ 7649] = 1'b0;  wr_cycle[ 7649] = 1'b1;  addr_rom[ 7649]='h00001978;  wr_data_rom[ 7649]='h000019cb;
    rd_cycle[ 7650] = 1'b1;  wr_cycle[ 7650] = 1'b0;  addr_rom[ 7650]='h00001a44;  wr_data_rom[ 7650]='h00000000;
    rd_cycle[ 7651] = 1'b1;  wr_cycle[ 7651] = 1'b0;  addr_rom[ 7651]='h00000bf8;  wr_data_rom[ 7651]='h00000000;
    rd_cycle[ 7652] = 1'b0;  wr_cycle[ 7652] = 1'b1;  addr_rom[ 7652]='h00000ba8;  wr_data_rom[ 7652]='h00001df2;
    rd_cycle[ 7653] = 1'b1;  wr_cycle[ 7653] = 1'b0;  addr_rom[ 7653]='h000012d0;  wr_data_rom[ 7653]='h00000000;
    rd_cycle[ 7654] = 1'b1;  wr_cycle[ 7654] = 1'b0;  addr_rom[ 7654]='h00001bc8;  wr_data_rom[ 7654]='h00000000;
    rd_cycle[ 7655] = 1'b0;  wr_cycle[ 7655] = 1'b1;  addr_rom[ 7655]='h00001c1c;  wr_data_rom[ 7655]='h00000168;
    rd_cycle[ 7656] = 1'b1;  wr_cycle[ 7656] = 1'b0;  addr_rom[ 7656]='h00001568;  wr_data_rom[ 7656]='h00000000;
    rd_cycle[ 7657] = 1'b0;  wr_cycle[ 7657] = 1'b1;  addr_rom[ 7657]='h0000087c;  wr_data_rom[ 7657]='h00000e2b;
    rd_cycle[ 7658] = 1'b1;  wr_cycle[ 7658] = 1'b0;  addr_rom[ 7658]='h00000670;  wr_data_rom[ 7658]='h00000000;
    rd_cycle[ 7659] = 1'b1;  wr_cycle[ 7659] = 1'b0;  addr_rom[ 7659]='h00001e70;  wr_data_rom[ 7659]='h00000000;
    rd_cycle[ 7660] = 1'b1;  wr_cycle[ 7660] = 1'b0;  addr_rom[ 7660]='h00000990;  wr_data_rom[ 7660]='h00000000;
    rd_cycle[ 7661] = 1'b0;  wr_cycle[ 7661] = 1'b1;  addr_rom[ 7661]='h00001a3c;  wr_data_rom[ 7661]='h0000011d;
    rd_cycle[ 7662] = 1'b0;  wr_cycle[ 7662] = 1'b1;  addr_rom[ 7662]='h00001188;  wr_data_rom[ 7662]='h00001ad4;
    rd_cycle[ 7663] = 1'b0;  wr_cycle[ 7663] = 1'b1;  addr_rom[ 7663]='h000010cc;  wr_data_rom[ 7663]='h0000186b;
    rd_cycle[ 7664] = 1'b0;  wr_cycle[ 7664] = 1'b1;  addr_rom[ 7664]='h00001a6c;  wr_data_rom[ 7664]='h00001705;
    rd_cycle[ 7665] = 1'b1;  wr_cycle[ 7665] = 1'b0;  addr_rom[ 7665]='h00000f98;  wr_data_rom[ 7665]='h00000000;
    rd_cycle[ 7666] = 1'b1;  wr_cycle[ 7666] = 1'b0;  addr_rom[ 7666]='h00000988;  wr_data_rom[ 7666]='h00000000;
    rd_cycle[ 7667] = 1'b1;  wr_cycle[ 7667] = 1'b0;  addr_rom[ 7667]='h00001830;  wr_data_rom[ 7667]='h00000000;
    rd_cycle[ 7668] = 1'b1;  wr_cycle[ 7668] = 1'b0;  addr_rom[ 7668]='h000004f0;  wr_data_rom[ 7668]='h00000000;
    rd_cycle[ 7669] = 1'b1;  wr_cycle[ 7669] = 1'b0;  addr_rom[ 7669]='h00000eb0;  wr_data_rom[ 7669]='h00000000;
    rd_cycle[ 7670] = 1'b0;  wr_cycle[ 7670] = 1'b1;  addr_rom[ 7670]='h00001790;  wr_data_rom[ 7670]='h0000139d;
    rd_cycle[ 7671] = 1'b1;  wr_cycle[ 7671] = 1'b0;  addr_rom[ 7671]='h000008fc;  wr_data_rom[ 7671]='h00000000;
    rd_cycle[ 7672] = 1'b1;  wr_cycle[ 7672] = 1'b0;  addr_rom[ 7672]='h00000bc4;  wr_data_rom[ 7672]='h00000000;
    rd_cycle[ 7673] = 1'b0;  wr_cycle[ 7673] = 1'b1;  addr_rom[ 7673]='h00001278;  wr_data_rom[ 7673]='h00000b20;
    rd_cycle[ 7674] = 1'b0;  wr_cycle[ 7674] = 1'b1;  addr_rom[ 7674]='h000010a4;  wr_data_rom[ 7674]='h00001139;
    rd_cycle[ 7675] = 1'b1;  wr_cycle[ 7675] = 1'b0;  addr_rom[ 7675]='h00000378;  wr_data_rom[ 7675]='h00000000;
    rd_cycle[ 7676] = 1'b0;  wr_cycle[ 7676] = 1'b1;  addr_rom[ 7676]='h00001058;  wr_data_rom[ 7676]='h000011f3;
    rd_cycle[ 7677] = 1'b0;  wr_cycle[ 7677] = 1'b1;  addr_rom[ 7677]='h0000111c;  wr_data_rom[ 7677]='h000008d2;
    rd_cycle[ 7678] = 1'b1;  wr_cycle[ 7678] = 1'b0;  addr_rom[ 7678]='h00000efc;  wr_data_rom[ 7678]='h00000000;
    rd_cycle[ 7679] = 1'b1;  wr_cycle[ 7679] = 1'b0;  addr_rom[ 7679]='h000002f0;  wr_data_rom[ 7679]='h00000000;
    rd_cycle[ 7680] = 1'b1;  wr_cycle[ 7680] = 1'b0;  addr_rom[ 7680]='h000006a4;  wr_data_rom[ 7680]='h00000000;
    rd_cycle[ 7681] = 1'b0;  wr_cycle[ 7681] = 1'b1;  addr_rom[ 7681]='h00000ef8;  wr_data_rom[ 7681]='h000006df;
    rd_cycle[ 7682] = 1'b1;  wr_cycle[ 7682] = 1'b0;  addr_rom[ 7682]='h000018fc;  wr_data_rom[ 7682]='h00000000;
    rd_cycle[ 7683] = 1'b0;  wr_cycle[ 7683] = 1'b1;  addr_rom[ 7683]='h00000f00;  wr_data_rom[ 7683]='h0000113e;
    rd_cycle[ 7684] = 1'b1;  wr_cycle[ 7684] = 1'b0;  addr_rom[ 7684]='h00001920;  wr_data_rom[ 7684]='h00000000;
    rd_cycle[ 7685] = 1'b1;  wr_cycle[ 7685] = 1'b0;  addr_rom[ 7685]='h00001de0;  wr_data_rom[ 7685]='h00000000;
    rd_cycle[ 7686] = 1'b0;  wr_cycle[ 7686] = 1'b1;  addr_rom[ 7686]='h00000774;  wr_data_rom[ 7686]='h000006c5;
    rd_cycle[ 7687] = 1'b1;  wr_cycle[ 7687] = 1'b0;  addr_rom[ 7687]='h000016dc;  wr_data_rom[ 7687]='h00000000;
    rd_cycle[ 7688] = 1'b1;  wr_cycle[ 7688] = 1'b0;  addr_rom[ 7688]='h00000ba4;  wr_data_rom[ 7688]='h00000000;
    rd_cycle[ 7689] = 1'b1;  wr_cycle[ 7689] = 1'b0;  addr_rom[ 7689]='h00001c3c;  wr_data_rom[ 7689]='h00000000;
    rd_cycle[ 7690] = 1'b1;  wr_cycle[ 7690] = 1'b0;  addr_rom[ 7690]='h00001950;  wr_data_rom[ 7690]='h00000000;
    rd_cycle[ 7691] = 1'b1;  wr_cycle[ 7691] = 1'b0;  addr_rom[ 7691]='h00000288;  wr_data_rom[ 7691]='h00000000;
    rd_cycle[ 7692] = 1'b0;  wr_cycle[ 7692] = 1'b1;  addr_rom[ 7692]='h00000c48;  wr_data_rom[ 7692]='h00001813;
    rd_cycle[ 7693] = 1'b0;  wr_cycle[ 7693] = 1'b1;  addr_rom[ 7693]='h000003b8;  wr_data_rom[ 7693]='h00001924;
    rd_cycle[ 7694] = 1'b0;  wr_cycle[ 7694] = 1'b1;  addr_rom[ 7694]='h000002ac;  wr_data_rom[ 7694]='h00000e39;
    rd_cycle[ 7695] = 1'b1;  wr_cycle[ 7695] = 1'b0;  addr_rom[ 7695]='h00001c0c;  wr_data_rom[ 7695]='h00000000;
    rd_cycle[ 7696] = 1'b1;  wr_cycle[ 7696] = 1'b0;  addr_rom[ 7696]='h00000640;  wr_data_rom[ 7696]='h00000000;
    rd_cycle[ 7697] = 1'b0;  wr_cycle[ 7697] = 1'b1;  addr_rom[ 7697]='h00001e64;  wr_data_rom[ 7697]='h00001a36;
    rd_cycle[ 7698] = 1'b0;  wr_cycle[ 7698] = 1'b1;  addr_rom[ 7698]='h00001df0;  wr_data_rom[ 7698]='h00001934;
    rd_cycle[ 7699] = 1'b0;  wr_cycle[ 7699] = 1'b1;  addr_rom[ 7699]='h00001868;  wr_data_rom[ 7699]='h00000df9;
    rd_cycle[ 7700] = 1'b0;  wr_cycle[ 7700] = 1'b1;  addr_rom[ 7700]='h00000c50;  wr_data_rom[ 7700]='h00001eb3;
    rd_cycle[ 7701] = 1'b0;  wr_cycle[ 7701] = 1'b1;  addr_rom[ 7701]='h00001590;  wr_data_rom[ 7701]='h000014cd;
    rd_cycle[ 7702] = 1'b0;  wr_cycle[ 7702] = 1'b1;  addr_rom[ 7702]='h00001608;  wr_data_rom[ 7702]='h00000dbc;
    rd_cycle[ 7703] = 1'b0;  wr_cycle[ 7703] = 1'b1;  addr_rom[ 7703]='h00001810;  wr_data_rom[ 7703]='h0000012a;
    rd_cycle[ 7704] = 1'b0;  wr_cycle[ 7704] = 1'b1;  addr_rom[ 7704]='h000013c8;  wr_data_rom[ 7704]='h000013d6;
    rd_cycle[ 7705] = 1'b1;  wr_cycle[ 7705] = 1'b0;  addr_rom[ 7705]='h00001300;  wr_data_rom[ 7705]='h00000000;
    rd_cycle[ 7706] = 1'b1;  wr_cycle[ 7706] = 1'b0;  addr_rom[ 7706]='h0000030c;  wr_data_rom[ 7706]='h00000000;
    rd_cycle[ 7707] = 1'b0;  wr_cycle[ 7707] = 1'b1;  addr_rom[ 7707]='h00000544;  wr_data_rom[ 7707]='h00000a68;
    rd_cycle[ 7708] = 1'b1;  wr_cycle[ 7708] = 1'b0;  addr_rom[ 7708]='h00000d3c;  wr_data_rom[ 7708]='h00000000;
    rd_cycle[ 7709] = 1'b1;  wr_cycle[ 7709] = 1'b0;  addr_rom[ 7709]='h00001d94;  wr_data_rom[ 7709]='h00000000;
    rd_cycle[ 7710] = 1'b1;  wr_cycle[ 7710] = 1'b0;  addr_rom[ 7710]='h00001220;  wr_data_rom[ 7710]='h00000000;
    rd_cycle[ 7711] = 1'b0;  wr_cycle[ 7711] = 1'b1;  addr_rom[ 7711]='h0000171c;  wr_data_rom[ 7711]='h00000a23;
    rd_cycle[ 7712] = 1'b1;  wr_cycle[ 7712] = 1'b0;  addr_rom[ 7712]='h000018c0;  wr_data_rom[ 7712]='h00000000;
    rd_cycle[ 7713] = 1'b0;  wr_cycle[ 7713] = 1'b1;  addr_rom[ 7713]='h00000274;  wr_data_rom[ 7713]='h000002bc;
    rd_cycle[ 7714] = 1'b1;  wr_cycle[ 7714] = 1'b0;  addr_rom[ 7714]='h00000844;  wr_data_rom[ 7714]='h00000000;
    rd_cycle[ 7715] = 1'b0;  wr_cycle[ 7715] = 1'b1;  addr_rom[ 7715]='h00000944;  wr_data_rom[ 7715]='h000015d0;
    rd_cycle[ 7716] = 1'b1;  wr_cycle[ 7716] = 1'b0;  addr_rom[ 7716]='h00000e08;  wr_data_rom[ 7716]='h00000000;
    rd_cycle[ 7717] = 1'b0;  wr_cycle[ 7717] = 1'b1;  addr_rom[ 7717]='h00000914;  wr_data_rom[ 7717]='h00000418;
    rd_cycle[ 7718] = 1'b1;  wr_cycle[ 7718] = 1'b0;  addr_rom[ 7718]='h00000be8;  wr_data_rom[ 7718]='h00000000;
    rd_cycle[ 7719] = 1'b1;  wr_cycle[ 7719] = 1'b0;  addr_rom[ 7719]='h000016dc;  wr_data_rom[ 7719]='h00000000;
    rd_cycle[ 7720] = 1'b0;  wr_cycle[ 7720] = 1'b1;  addr_rom[ 7720]='h00001d34;  wr_data_rom[ 7720]='h0000191a;
    rd_cycle[ 7721] = 1'b0;  wr_cycle[ 7721] = 1'b1;  addr_rom[ 7721]='h000019ac;  wr_data_rom[ 7721]='h00001c5d;
    rd_cycle[ 7722] = 1'b1;  wr_cycle[ 7722] = 1'b0;  addr_rom[ 7722]='h0000178c;  wr_data_rom[ 7722]='h00000000;
    rd_cycle[ 7723] = 1'b0;  wr_cycle[ 7723] = 1'b1;  addr_rom[ 7723]='h00000f2c;  wr_data_rom[ 7723]='h00001725;
    rd_cycle[ 7724] = 1'b0;  wr_cycle[ 7724] = 1'b1;  addr_rom[ 7724]='h000017cc;  wr_data_rom[ 7724]='h000012c5;
    rd_cycle[ 7725] = 1'b0;  wr_cycle[ 7725] = 1'b1;  addr_rom[ 7725]='h00001e94;  wr_data_rom[ 7725]='h0000050c;
    rd_cycle[ 7726] = 1'b0;  wr_cycle[ 7726] = 1'b1;  addr_rom[ 7726]='h0000086c;  wr_data_rom[ 7726]='h0000038a;
    rd_cycle[ 7727] = 1'b1;  wr_cycle[ 7727] = 1'b0;  addr_rom[ 7727]='h00001e1c;  wr_data_rom[ 7727]='h00000000;
    rd_cycle[ 7728] = 1'b1;  wr_cycle[ 7728] = 1'b0;  addr_rom[ 7728]='h000002e8;  wr_data_rom[ 7728]='h00000000;
    rd_cycle[ 7729] = 1'b0;  wr_cycle[ 7729] = 1'b1;  addr_rom[ 7729]='h0000063c;  wr_data_rom[ 7729]='h0000110e;
    rd_cycle[ 7730] = 1'b0;  wr_cycle[ 7730] = 1'b1;  addr_rom[ 7730]='h00001524;  wr_data_rom[ 7730]='h000006ea;
    rd_cycle[ 7731] = 1'b0;  wr_cycle[ 7731] = 1'b1;  addr_rom[ 7731]='h00000008;  wr_data_rom[ 7731]='h0000142c;
    rd_cycle[ 7732] = 1'b1;  wr_cycle[ 7732] = 1'b0;  addr_rom[ 7732]='h00000e8c;  wr_data_rom[ 7732]='h00000000;
    rd_cycle[ 7733] = 1'b0;  wr_cycle[ 7733] = 1'b1;  addr_rom[ 7733]='h00001730;  wr_data_rom[ 7733]='h00000b79;
    rd_cycle[ 7734] = 1'b0;  wr_cycle[ 7734] = 1'b1;  addr_rom[ 7734]='h00001ef4;  wr_data_rom[ 7734]='h00001110;
    rd_cycle[ 7735] = 1'b0;  wr_cycle[ 7735] = 1'b1;  addr_rom[ 7735]='h00000ce4;  wr_data_rom[ 7735]='h000012c9;
    rd_cycle[ 7736] = 1'b1;  wr_cycle[ 7736] = 1'b0;  addr_rom[ 7736]='h000016f8;  wr_data_rom[ 7736]='h00000000;
    rd_cycle[ 7737] = 1'b0;  wr_cycle[ 7737] = 1'b1;  addr_rom[ 7737]='h00000ba0;  wr_data_rom[ 7737]='h00000887;
    rd_cycle[ 7738] = 1'b1;  wr_cycle[ 7738] = 1'b0;  addr_rom[ 7738]='h000005bc;  wr_data_rom[ 7738]='h00000000;
    rd_cycle[ 7739] = 1'b0;  wr_cycle[ 7739] = 1'b1;  addr_rom[ 7739]='h000007b0;  wr_data_rom[ 7739]='h000003fc;
    rd_cycle[ 7740] = 1'b0;  wr_cycle[ 7740] = 1'b1;  addr_rom[ 7740]='h00000bf4;  wr_data_rom[ 7740]='h000007dc;
    rd_cycle[ 7741] = 1'b0;  wr_cycle[ 7741] = 1'b1;  addr_rom[ 7741]='h000012bc;  wr_data_rom[ 7741]='h00000ceb;
    rd_cycle[ 7742] = 1'b0;  wr_cycle[ 7742] = 1'b1;  addr_rom[ 7742]='h00000578;  wr_data_rom[ 7742]='h00000e41;
    rd_cycle[ 7743] = 1'b1;  wr_cycle[ 7743] = 1'b0;  addr_rom[ 7743]='h0000021c;  wr_data_rom[ 7743]='h00000000;
    rd_cycle[ 7744] = 1'b0;  wr_cycle[ 7744] = 1'b1;  addr_rom[ 7744]='h0000134c;  wr_data_rom[ 7744]='h00000a2c;
    rd_cycle[ 7745] = 1'b0;  wr_cycle[ 7745] = 1'b1;  addr_rom[ 7745]='h00000724;  wr_data_rom[ 7745]='h00000509;
    rd_cycle[ 7746] = 1'b1;  wr_cycle[ 7746] = 1'b0;  addr_rom[ 7746]='h00001b68;  wr_data_rom[ 7746]='h00000000;
    rd_cycle[ 7747] = 1'b1;  wr_cycle[ 7747] = 1'b0;  addr_rom[ 7747]='h00001c48;  wr_data_rom[ 7747]='h00000000;
    rd_cycle[ 7748] = 1'b1;  wr_cycle[ 7748] = 1'b0;  addr_rom[ 7748]='h00001d34;  wr_data_rom[ 7748]='h00000000;
    rd_cycle[ 7749] = 1'b0;  wr_cycle[ 7749] = 1'b1;  addr_rom[ 7749]='h000002c4;  wr_data_rom[ 7749]='h00000ef3;
    rd_cycle[ 7750] = 1'b1;  wr_cycle[ 7750] = 1'b0;  addr_rom[ 7750]='h00000a04;  wr_data_rom[ 7750]='h00000000;
    rd_cycle[ 7751] = 1'b1;  wr_cycle[ 7751] = 1'b0;  addr_rom[ 7751]='h000016b8;  wr_data_rom[ 7751]='h00000000;
    rd_cycle[ 7752] = 1'b0;  wr_cycle[ 7752] = 1'b1;  addr_rom[ 7752]='h00001738;  wr_data_rom[ 7752]='h000000ab;
    rd_cycle[ 7753] = 1'b0;  wr_cycle[ 7753] = 1'b1;  addr_rom[ 7753]='h00001980;  wr_data_rom[ 7753]='h00000694;
    rd_cycle[ 7754] = 1'b1;  wr_cycle[ 7754] = 1'b0;  addr_rom[ 7754]='h00001db8;  wr_data_rom[ 7754]='h00000000;
    rd_cycle[ 7755] = 1'b1;  wr_cycle[ 7755] = 1'b0;  addr_rom[ 7755]='h0000158c;  wr_data_rom[ 7755]='h00000000;
    rd_cycle[ 7756] = 1'b1;  wr_cycle[ 7756] = 1'b0;  addr_rom[ 7756]='h00000414;  wr_data_rom[ 7756]='h00000000;
    rd_cycle[ 7757] = 1'b0;  wr_cycle[ 7757] = 1'b1;  addr_rom[ 7757]='h000013a8;  wr_data_rom[ 7757]='h00001b39;
    rd_cycle[ 7758] = 1'b0;  wr_cycle[ 7758] = 1'b1;  addr_rom[ 7758]='h00000b38;  wr_data_rom[ 7758]='h00001946;
    rd_cycle[ 7759] = 1'b0;  wr_cycle[ 7759] = 1'b1;  addr_rom[ 7759]='h0000188c;  wr_data_rom[ 7759]='h00000501;
    rd_cycle[ 7760] = 1'b0;  wr_cycle[ 7760] = 1'b1;  addr_rom[ 7760]='h00000320;  wr_data_rom[ 7760]='h00000e37;
    rd_cycle[ 7761] = 1'b1;  wr_cycle[ 7761] = 1'b0;  addr_rom[ 7761]='h000010dc;  wr_data_rom[ 7761]='h00000000;
    rd_cycle[ 7762] = 1'b1;  wr_cycle[ 7762] = 1'b0;  addr_rom[ 7762]='h00000b7c;  wr_data_rom[ 7762]='h00000000;
    rd_cycle[ 7763] = 1'b0;  wr_cycle[ 7763] = 1'b1;  addr_rom[ 7763]='h000005a4;  wr_data_rom[ 7763]='h00000c53;
    rd_cycle[ 7764] = 1'b1;  wr_cycle[ 7764] = 1'b0;  addr_rom[ 7764]='h00001c30;  wr_data_rom[ 7764]='h00000000;
    rd_cycle[ 7765] = 1'b1;  wr_cycle[ 7765] = 1'b0;  addr_rom[ 7765]='h00000fd0;  wr_data_rom[ 7765]='h00000000;
    rd_cycle[ 7766] = 1'b1;  wr_cycle[ 7766] = 1'b0;  addr_rom[ 7766]='h0000027c;  wr_data_rom[ 7766]='h00000000;
    rd_cycle[ 7767] = 1'b1;  wr_cycle[ 7767] = 1'b0;  addr_rom[ 7767]='h00001bac;  wr_data_rom[ 7767]='h00000000;
    rd_cycle[ 7768] = 1'b0;  wr_cycle[ 7768] = 1'b1;  addr_rom[ 7768]='h00000934;  wr_data_rom[ 7768]='h00001ef0;
    rd_cycle[ 7769] = 1'b1;  wr_cycle[ 7769] = 1'b0;  addr_rom[ 7769]='h00000388;  wr_data_rom[ 7769]='h00000000;
    rd_cycle[ 7770] = 1'b0;  wr_cycle[ 7770] = 1'b1;  addr_rom[ 7770]='h00001364;  wr_data_rom[ 7770]='h00000b94;
    rd_cycle[ 7771] = 1'b0;  wr_cycle[ 7771] = 1'b1;  addr_rom[ 7771]='h000004b8;  wr_data_rom[ 7771]='h00000dfc;
    rd_cycle[ 7772] = 1'b1;  wr_cycle[ 7772] = 1'b0;  addr_rom[ 7772]='h0000106c;  wr_data_rom[ 7772]='h00000000;
    rd_cycle[ 7773] = 1'b1;  wr_cycle[ 7773] = 1'b0;  addr_rom[ 7773]='h000017ac;  wr_data_rom[ 7773]='h00000000;
    rd_cycle[ 7774] = 1'b1;  wr_cycle[ 7774] = 1'b0;  addr_rom[ 7774]='h000008bc;  wr_data_rom[ 7774]='h00000000;
    rd_cycle[ 7775] = 1'b1;  wr_cycle[ 7775] = 1'b0;  addr_rom[ 7775]='h0000097c;  wr_data_rom[ 7775]='h00000000;
    rd_cycle[ 7776] = 1'b0;  wr_cycle[ 7776] = 1'b1;  addr_rom[ 7776]='h00001250;  wr_data_rom[ 7776]='h00001b1c;
    rd_cycle[ 7777] = 1'b0;  wr_cycle[ 7777] = 1'b1;  addr_rom[ 7777]='h00001bcc;  wr_data_rom[ 7777]='h00000c83;
    rd_cycle[ 7778] = 1'b0;  wr_cycle[ 7778] = 1'b1;  addr_rom[ 7778]='h0000126c;  wr_data_rom[ 7778]='h00000a7b;
    rd_cycle[ 7779] = 1'b0;  wr_cycle[ 7779] = 1'b1;  addr_rom[ 7779]='h000017fc;  wr_data_rom[ 7779]='h0000046e;
    rd_cycle[ 7780] = 1'b1;  wr_cycle[ 7780] = 1'b0;  addr_rom[ 7780]='h0000123c;  wr_data_rom[ 7780]='h00000000;
    rd_cycle[ 7781] = 1'b1;  wr_cycle[ 7781] = 1'b0;  addr_rom[ 7781]='h00001724;  wr_data_rom[ 7781]='h00000000;
    rd_cycle[ 7782] = 1'b0;  wr_cycle[ 7782] = 1'b1;  addr_rom[ 7782]='h00000ae4;  wr_data_rom[ 7782]='h000007f7;
    rd_cycle[ 7783] = 1'b1;  wr_cycle[ 7783] = 1'b0;  addr_rom[ 7783]='h00000098;  wr_data_rom[ 7783]='h00000000;
    rd_cycle[ 7784] = 1'b1;  wr_cycle[ 7784] = 1'b0;  addr_rom[ 7784]='h00001b50;  wr_data_rom[ 7784]='h00000000;
    rd_cycle[ 7785] = 1'b1;  wr_cycle[ 7785] = 1'b0;  addr_rom[ 7785]='h00001c6c;  wr_data_rom[ 7785]='h00000000;
    rd_cycle[ 7786] = 1'b1;  wr_cycle[ 7786] = 1'b0;  addr_rom[ 7786]='h00000338;  wr_data_rom[ 7786]='h00000000;
    rd_cycle[ 7787] = 1'b1;  wr_cycle[ 7787] = 1'b0;  addr_rom[ 7787]='h0000145c;  wr_data_rom[ 7787]='h00000000;
    rd_cycle[ 7788] = 1'b0;  wr_cycle[ 7788] = 1'b1;  addr_rom[ 7788]='h000012c4;  wr_data_rom[ 7788]='h00000466;
    rd_cycle[ 7789] = 1'b1;  wr_cycle[ 7789] = 1'b0;  addr_rom[ 7789]='h00000988;  wr_data_rom[ 7789]='h00000000;
    rd_cycle[ 7790] = 1'b0;  wr_cycle[ 7790] = 1'b1;  addr_rom[ 7790]='h000011a0;  wr_data_rom[ 7790]='h0000131e;
    rd_cycle[ 7791] = 1'b0;  wr_cycle[ 7791] = 1'b1;  addr_rom[ 7791]='h00001094;  wr_data_rom[ 7791]='h00000675;
    rd_cycle[ 7792] = 1'b1;  wr_cycle[ 7792] = 1'b0;  addr_rom[ 7792]='h00000674;  wr_data_rom[ 7792]='h00000000;
    rd_cycle[ 7793] = 1'b1;  wr_cycle[ 7793] = 1'b0;  addr_rom[ 7793]='h000016a0;  wr_data_rom[ 7793]='h00000000;
    rd_cycle[ 7794] = 1'b1;  wr_cycle[ 7794] = 1'b0;  addr_rom[ 7794]='h00001810;  wr_data_rom[ 7794]='h00000000;
    rd_cycle[ 7795] = 1'b1;  wr_cycle[ 7795] = 1'b0;  addr_rom[ 7795]='h0000154c;  wr_data_rom[ 7795]='h00000000;
    rd_cycle[ 7796] = 1'b1;  wr_cycle[ 7796] = 1'b0;  addr_rom[ 7796]='h00000480;  wr_data_rom[ 7796]='h00000000;
    rd_cycle[ 7797] = 1'b0;  wr_cycle[ 7797] = 1'b1;  addr_rom[ 7797]='h00001514;  wr_data_rom[ 7797]='h0000053d;
    rd_cycle[ 7798] = 1'b0;  wr_cycle[ 7798] = 1'b1;  addr_rom[ 7798]='h0000155c;  wr_data_rom[ 7798]='h00000a30;
    rd_cycle[ 7799] = 1'b1;  wr_cycle[ 7799] = 1'b0;  addr_rom[ 7799]='h00000690;  wr_data_rom[ 7799]='h00000000;
    rd_cycle[ 7800] = 1'b1;  wr_cycle[ 7800] = 1'b0;  addr_rom[ 7800]='h0000022c;  wr_data_rom[ 7800]='h00000000;
    rd_cycle[ 7801] = 1'b0;  wr_cycle[ 7801] = 1'b1;  addr_rom[ 7801]='h000004f0;  wr_data_rom[ 7801]='h000017d3;
    rd_cycle[ 7802] = 1'b0;  wr_cycle[ 7802] = 1'b1;  addr_rom[ 7802]='h00000e80;  wr_data_rom[ 7802]='h000010a6;
    rd_cycle[ 7803] = 1'b0;  wr_cycle[ 7803] = 1'b1;  addr_rom[ 7803]='h00001678;  wr_data_rom[ 7803]='h000017ed;
    rd_cycle[ 7804] = 1'b0;  wr_cycle[ 7804] = 1'b1;  addr_rom[ 7804]='h00000098;  wr_data_rom[ 7804]='h000016db;
    rd_cycle[ 7805] = 1'b1;  wr_cycle[ 7805] = 1'b0;  addr_rom[ 7805]='h00000bcc;  wr_data_rom[ 7805]='h00000000;
    rd_cycle[ 7806] = 1'b1;  wr_cycle[ 7806] = 1'b0;  addr_rom[ 7806]='h0000123c;  wr_data_rom[ 7806]='h00000000;
    rd_cycle[ 7807] = 1'b0;  wr_cycle[ 7807] = 1'b1;  addr_rom[ 7807]='h00000084;  wr_data_rom[ 7807]='h00001766;
    rd_cycle[ 7808] = 1'b1;  wr_cycle[ 7808] = 1'b0;  addr_rom[ 7808]='h00001024;  wr_data_rom[ 7808]='h00000000;
    rd_cycle[ 7809] = 1'b0;  wr_cycle[ 7809] = 1'b1;  addr_rom[ 7809]='h000005f0;  wr_data_rom[ 7809]='h00001b14;
    rd_cycle[ 7810] = 1'b1;  wr_cycle[ 7810] = 1'b0;  addr_rom[ 7810]='h00000284;  wr_data_rom[ 7810]='h00000000;
    rd_cycle[ 7811] = 1'b1;  wr_cycle[ 7811] = 1'b0;  addr_rom[ 7811]='h000013f0;  wr_data_rom[ 7811]='h00000000;
    rd_cycle[ 7812] = 1'b1;  wr_cycle[ 7812] = 1'b0;  addr_rom[ 7812]='h000015cc;  wr_data_rom[ 7812]='h00000000;
    rd_cycle[ 7813] = 1'b1;  wr_cycle[ 7813] = 1'b0;  addr_rom[ 7813]='h00001570;  wr_data_rom[ 7813]='h00000000;
    rd_cycle[ 7814] = 1'b1;  wr_cycle[ 7814] = 1'b0;  addr_rom[ 7814]='h00000704;  wr_data_rom[ 7814]='h00000000;
    rd_cycle[ 7815] = 1'b0;  wr_cycle[ 7815] = 1'b1;  addr_rom[ 7815]='h000001b4;  wr_data_rom[ 7815]='h00000f69;
    rd_cycle[ 7816] = 1'b0;  wr_cycle[ 7816] = 1'b1;  addr_rom[ 7816]='h00001d30;  wr_data_rom[ 7816]='h00000932;
    rd_cycle[ 7817] = 1'b0;  wr_cycle[ 7817] = 1'b1;  addr_rom[ 7817]='h00001d2c;  wr_data_rom[ 7817]='h000011e2;
    rd_cycle[ 7818] = 1'b1;  wr_cycle[ 7818] = 1'b0;  addr_rom[ 7818]='h000002c8;  wr_data_rom[ 7818]='h00000000;
    rd_cycle[ 7819] = 1'b0;  wr_cycle[ 7819] = 1'b1;  addr_rom[ 7819]='h00000eb0;  wr_data_rom[ 7819]='h00000bda;
    rd_cycle[ 7820] = 1'b1;  wr_cycle[ 7820] = 1'b0;  addr_rom[ 7820]='h000000f8;  wr_data_rom[ 7820]='h00000000;
    rd_cycle[ 7821] = 1'b0;  wr_cycle[ 7821] = 1'b1;  addr_rom[ 7821]='h00001af0;  wr_data_rom[ 7821]='h000012a5;
    rd_cycle[ 7822] = 1'b0;  wr_cycle[ 7822] = 1'b1;  addr_rom[ 7822]='h000010e0;  wr_data_rom[ 7822]='h00001380;
    rd_cycle[ 7823] = 1'b1;  wr_cycle[ 7823] = 1'b0;  addr_rom[ 7823]='h000011d0;  wr_data_rom[ 7823]='h00000000;
    rd_cycle[ 7824] = 1'b0;  wr_cycle[ 7824] = 1'b1;  addr_rom[ 7824]='h00001320;  wr_data_rom[ 7824]='h00001e10;
    rd_cycle[ 7825] = 1'b0;  wr_cycle[ 7825] = 1'b1;  addr_rom[ 7825]='h00001554;  wr_data_rom[ 7825]='h00001ec1;
    rd_cycle[ 7826] = 1'b1;  wr_cycle[ 7826] = 1'b0;  addr_rom[ 7826]='h000018f0;  wr_data_rom[ 7826]='h00000000;
    rd_cycle[ 7827] = 1'b1;  wr_cycle[ 7827] = 1'b0;  addr_rom[ 7827]='h0000087c;  wr_data_rom[ 7827]='h00000000;
    rd_cycle[ 7828] = 1'b1;  wr_cycle[ 7828] = 1'b0;  addr_rom[ 7828]='h00001748;  wr_data_rom[ 7828]='h00000000;
    rd_cycle[ 7829] = 1'b0;  wr_cycle[ 7829] = 1'b1;  addr_rom[ 7829]='h000001dc;  wr_data_rom[ 7829]='h00001aca;
    rd_cycle[ 7830] = 1'b0;  wr_cycle[ 7830] = 1'b1;  addr_rom[ 7830]='h00000d58;  wr_data_rom[ 7830]='h00001abe;
    rd_cycle[ 7831] = 1'b0;  wr_cycle[ 7831] = 1'b1;  addr_rom[ 7831]='h00001e3c;  wr_data_rom[ 7831]='h00000eea;
    rd_cycle[ 7832] = 1'b1;  wr_cycle[ 7832] = 1'b0;  addr_rom[ 7832]='h00000c68;  wr_data_rom[ 7832]='h00000000;
    rd_cycle[ 7833] = 1'b0;  wr_cycle[ 7833] = 1'b1;  addr_rom[ 7833]='h0000191c;  wr_data_rom[ 7833]='h00001d26;
    rd_cycle[ 7834] = 1'b1;  wr_cycle[ 7834] = 1'b0;  addr_rom[ 7834]='h00000530;  wr_data_rom[ 7834]='h00000000;
    rd_cycle[ 7835] = 1'b0;  wr_cycle[ 7835] = 1'b1;  addr_rom[ 7835]='h00001a98;  wr_data_rom[ 7835]='h00001d2c;
    rd_cycle[ 7836] = 1'b0;  wr_cycle[ 7836] = 1'b1;  addr_rom[ 7836]='h00001284;  wr_data_rom[ 7836]='h00000d05;
    rd_cycle[ 7837] = 1'b1;  wr_cycle[ 7837] = 1'b0;  addr_rom[ 7837]='h00001294;  wr_data_rom[ 7837]='h00000000;
    rd_cycle[ 7838] = 1'b1;  wr_cycle[ 7838] = 1'b0;  addr_rom[ 7838]='h00001158;  wr_data_rom[ 7838]='h00000000;
    rd_cycle[ 7839] = 1'b1;  wr_cycle[ 7839] = 1'b0;  addr_rom[ 7839]='h00001958;  wr_data_rom[ 7839]='h00000000;
    rd_cycle[ 7840] = 1'b1;  wr_cycle[ 7840] = 1'b0;  addr_rom[ 7840]='h000008a4;  wr_data_rom[ 7840]='h00000000;
    rd_cycle[ 7841] = 1'b0;  wr_cycle[ 7841] = 1'b1;  addr_rom[ 7841]='h000003ac;  wr_data_rom[ 7841]='h0000023d;
    rd_cycle[ 7842] = 1'b1;  wr_cycle[ 7842] = 1'b0;  addr_rom[ 7842]='h0000171c;  wr_data_rom[ 7842]='h00000000;
    rd_cycle[ 7843] = 1'b1;  wr_cycle[ 7843] = 1'b0;  addr_rom[ 7843]='h000008d4;  wr_data_rom[ 7843]='h00000000;
    rd_cycle[ 7844] = 1'b1;  wr_cycle[ 7844] = 1'b0;  addr_rom[ 7844]='h0000020c;  wr_data_rom[ 7844]='h00000000;
    rd_cycle[ 7845] = 1'b0;  wr_cycle[ 7845] = 1'b1;  addr_rom[ 7845]='h00001b40;  wr_data_rom[ 7845]='h000003bd;
    rd_cycle[ 7846] = 1'b1;  wr_cycle[ 7846] = 1'b0;  addr_rom[ 7846]='h000017a4;  wr_data_rom[ 7846]='h00000000;
    rd_cycle[ 7847] = 1'b1;  wr_cycle[ 7847] = 1'b0;  addr_rom[ 7847]='h00001d48;  wr_data_rom[ 7847]='h00000000;
    rd_cycle[ 7848] = 1'b0;  wr_cycle[ 7848] = 1'b1;  addr_rom[ 7848]='h00001080;  wr_data_rom[ 7848]='h00000616;
    rd_cycle[ 7849] = 1'b0;  wr_cycle[ 7849] = 1'b1;  addr_rom[ 7849]='h000009e4;  wr_data_rom[ 7849]='h0000148f;
    rd_cycle[ 7850] = 1'b0;  wr_cycle[ 7850] = 1'b1;  addr_rom[ 7850]='h00000ed8;  wr_data_rom[ 7850]='h000001d5;
    rd_cycle[ 7851] = 1'b0;  wr_cycle[ 7851] = 1'b1;  addr_rom[ 7851]='h00000c90;  wr_data_rom[ 7851]='h00000dab;
    rd_cycle[ 7852] = 1'b1;  wr_cycle[ 7852] = 1'b0;  addr_rom[ 7852]='h00000f60;  wr_data_rom[ 7852]='h00000000;
    rd_cycle[ 7853] = 1'b1;  wr_cycle[ 7853] = 1'b0;  addr_rom[ 7853]='h000018f8;  wr_data_rom[ 7853]='h00000000;
    rd_cycle[ 7854] = 1'b0;  wr_cycle[ 7854] = 1'b1;  addr_rom[ 7854]='h000003cc;  wr_data_rom[ 7854]='h00001b38;
    rd_cycle[ 7855] = 1'b1;  wr_cycle[ 7855] = 1'b0;  addr_rom[ 7855]='h00000990;  wr_data_rom[ 7855]='h00000000;
    rd_cycle[ 7856] = 1'b0;  wr_cycle[ 7856] = 1'b1;  addr_rom[ 7856]='h00001a2c;  wr_data_rom[ 7856]='h000007e2;
    rd_cycle[ 7857] = 1'b1;  wr_cycle[ 7857] = 1'b0;  addr_rom[ 7857]='h000019b0;  wr_data_rom[ 7857]='h00000000;
    rd_cycle[ 7858] = 1'b1;  wr_cycle[ 7858] = 1'b0;  addr_rom[ 7858]='h00000590;  wr_data_rom[ 7858]='h00000000;
    rd_cycle[ 7859] = 1'b0;  wr_cycle[ 7859] = 1'b1;  addr_rom[ 7859]='h000003dc;  wr_data_rom[ 7859]='h00001689;
    rd_cycle[ 7860] = 1'b1;  wr_cycle[ 7860] = 1'b0;  addr_rom[ 7860]='h00001074;  wr_data_rom[ 7860]='h00000000;
    rd_cycle[ 7861] = 1'b1;  wr_cycle[ 7861] = 1'b0;  addr_rom[ 7861]='h00000b80;  wr_data_rom[ 7861]='h00000000;
    rd_cycle[ 7862] = 1'b0;  wr_cycle[ 7862] = 1'b1;  addr_rom[ 7862]='h00000f10;  wr_data_rom[ 7862]='h000003e3;
    rd_cycle[ 7863] = 1'b1;  wr_cycle[ 7863] = 1'b0;  addr_rom[ 7863]='h000013b4;  wr_data_rom[ 7863]='h00000000;
    rd_cycle[ 7864] = 1'b1;  wr_cycle[ 7864] = 1'b0;  addr_rom[ 7864]='h00001530;  wr_data_rom[ 7864]='h00000000;
    rd_cycle[ 7865] = 1'b0;  wr_cycle[ 7865] = 1'b1;  addr_rom[ 7865]='h00000520;  wr_data_rom[ 7865]='h000015ef;
    rd_cycle[ 7866] = 1'b0;  wr_cycle[ 7866] = 1'b1;  addr_rom[ 7866]='h00001cf8;  wr_data_rom[ 7866]='h00001380;
    rd_cycle[ 7867] = 1'b0;  wr_cycle[ 7867] = 1'b1;  addr_rom[ 7867]='h00001124;  wr_data_rom[ 7867]='h00000193;
    rd_cycle[ 7868] = 1'b1;  wr_cycle[ 7868] = 1'b0;  addr_rom[ 7868]='h0000003c;  wr_data_rom[ 7868]='h00000000;
    rd_cycle[ 7869] = 1'b0;  wr_cycle[ 7869] = 1'b1;  addr_rom[ 7869]='h000005c0;  wr_data_rom[ 7869]='h000011f5;
    rd_cycle[ 7870] = 1'b1;  wr_cycle[ 7870] = 1'b0;  addr_rom[ 7870]='h000018c8;  wr_data_rom[ 7870]='h00000000;
    rd_cycle[ 7871] = 1'b0;  wr_cycle[ 7871] = 1'b1;  addr_rom[ 7871]='h00001a78;  wr_data_rom[ 7871]='h00001dcd;
    rd_cycle[ 7872] = 1'b0;  wr_cycle[ 7872] = 1'b1;  addr_rom[ 7872]='h00000dfc;  wr_data_rom[ 7872]='h00001245;
    rd_cycle[ 7873] = 1'b1;  wr_cycle[ 7873] = 1'b0;  addr_rom[ 7873]='h00001a54;  wr_data_rom[ 7873]='h00000000;
    rd_cycle[ 7874] = 1'b0;  wr_cycle[ 7874] = 1'b1;  addr_rom[ 7874]='h00000cdc;  wr_data_rom[ 7874]='h0000078f;
    rd_cycle[ 7875] = 1'b0;  wr_cycle[ 7875] = 1'b1;  addr_rom[ 7875]='h00000eac;  wr_data_rom[ 7875]='h0000128a;
    rd_cycle[ 7876] = 1'b1;  wr_cycle[ 7876] = 1'b0;  addr_rom[ 7876]='h00000fb4;  wr_data_rom[ 7876]='h00000000;
    rd_cycle[ 7877] = 1'b0;  wr_cycle[ 7877] = 1'b1;  addr_rom[ 7877]='h00000d48;  wr_data_rom[ 7877]='h00000851;
    rd_cycle[ 7878] = 1'b0;  wr_cycle[ 7878] = 1'b1;  addr_rom[ 7878]='h00000f78;  wr_data_rom[ 7878]='h00000b08;
    rd_cycle[ 7879] = 1'b0;  wr_cycle[ 7879] = 1'b1;  addr_rom[ 7879]='h00000908;  wr_data_rom[ 7879]='h000011e1;
    rd_cycle[ 7880] = 1'b1;  wr_cycle[ 7880] = 1'b0;  addr_rom[ 7880]='h00000ffc;  wr_data_rom[ 7880]='h00000000;
    rd_cycle[ 7881] = 1'b0;  wr_cycle[ 7881] = 1'b1;  addr_rom[ 7881]='h00000550;  wr_data_rom[ 7881]='h000013f7;
    rd_cycle[ 7882] = 1'b1;  wr_cycle[ 7882] = 1'b0;  addr_rom[ 7882]='h00000d88;  wr_data_rom[ 7882]='h00000000;
    rd_cycle[ 7883] = 1'b0;  wr_cycle[ 7883] = 1'b1;  addr_rom[ 7883]='h00000184;  wr_data_rom[ 7883]='h00000802;
    rd_cycle[ 7884] = 1'b1;  wr_cycle[ 7884] = 1'b0;  addr_rom[ 7884]='h00000318;  wr_data_rom[ 7884]='h00000000;
    rd_cycle[ 7885] = 1'b0;  wr_cycle[ 7885] = 1'b1;  addr_rom[ 7885]='h00000520;  wr_data_rom[ 7885]='h00000d53;
    rd_cycle[ 7886] = 1'b0;  wr_cycle[ 7886] = 1'b1;  addr_rom[ 7886]='h00000b04;  wr_data_rom[ 7886]='h0000177b;
    rd_cycle[ 7887] = 1'b0;  wr_cycle[ 7887] = 1'b1;  addr_rom[ 7887]='h00001e64;  wr_data_rom[ 7887]='h00001a9d;
    rd_cycle[ 7888] = 1'b1;  wr_cycle[ 7888] = 1'b0;  addr_rom[ 7888]='h0000124c;  wr_data_rom[ 7888]='h00000000;
    rd_cycle[ 7889] = 1'b1;  wr_cycle[ 7889] = 1'b0;  addr_rom[ 7889]='h00000b8c;  wr_data_rom[ 7889]='h00000000;
    rd_cycle[ 7890] = 1'b0;  wr_cycle[ 7890] = 1'b1;  addr_rom[ 7890]='h000004c4;  wr_data_rom[ 7890]='h00000416;
    rd_cycle[ 7891] = 1'b0;  wr_cycle[ 7891] = 1'b1;  addr_rom[ 7891]='h00000840;  wr_data_rom[ 7891]='h00001693;
    rd_cycle[ 7892] = 1'b0;  wr_cycle[ 7892] = 1'b1;  addr_rom[ 7892]='h000013f8;  wr_data_rom[ 7892]='h00001c23;
    rd_cycle[ 7893] = 1'b1;  wr_cycle[ 7893] = 1'b0;  addr_rom[ 7893]='h00000fec;  wr_data_rom[ 7893]='h00000000;
    rd_cycle[ 7894] = 1'b0;  wr_cycle[ 7894] = 1'b1;  addr_rom[ 7894]='h00000958;  wr_data_rom[ 7894]='h00000217;
    rd_cycle[ 7895] = 1'b1;  wr_cycle[ 7895] = 1'b0;  addr_rom[ 7895]='h00001774;  wr_data_rom[ 7895]='h00000000;
    rd_cycle[ 7896] = 1'b0;  wr_cycle[ 7896] = 1'b1;  addr_rom[ 7896]='h00001124;  wr_data_rom[ 7896]='h00000a00;
    rd_cycle[ 7897] = 1'b0;  wr_cycle[ 7897] = 1'b1;  addr_rom[ 7897]='h000014f0;  wr_data_rom[ 7897]='h0000132b;
    rd_cycle[ 7898] = 1'b1;  wr_cycle[ 7898] = 1'b0;  addr_rom[ 7898]='h00001544;  wr_data_rom[ 7898]='h00000000;
    rd_cycle[ 7899] = 1'b0;  wr_cycle[ 7899] = 1'b1;  addr_rom[ 7899]='h000006a0;  wr_data_rom[ 7899]='h00001595;
    rd_cycle[ 7900] = 1'b0;  wr_cycle[ 7900] = 1'b1;  addr_rom[ 7900]='h00001518;  wr_data_rom[ 7900]='h00000fca;
    rd_cycle[ 7901] = 1'b1;  wr_cycle[ 7901] = 1'b0;  addr_rom[ 7901]='h00000e00;  wr_data_rom[ 7901]='h00000000;
    rd_cycle[ 7902] = 1'b1;  wr_cycle[ 7902] = 1'b0;  addr_rom[ 7902]='h00000044;  wr_data_rom[ 7902]='h00000000;
    rd_cycle[ 7903] = 1'b0;  wr_cycle[ 7903] = 1'b1;  addr_rom[ 7903]='h00000200;  wr_data_rom[ 7903]='h00000176;
    rd_cycle[ 7904] = 1'b0;  wr_cycle[ 7904] = 1'b1;  addr_rom[ 7904]='h0000053c;  wr_data_rom[ 7904]='h00001169;
    rd_cycle[ 7905] = 1'b1;  wr_cycle[ 7905] = 1'b0;  addr_rom[ 7905]='h00000f3c;  wr_data_rom[ 7905]='h00000000;
    rd_cycle[ 7906] = 1'b0;  wr_cycle[ 7906] = 1'b1;  addr_rom[ 7906]='h00001300;  wr_data_rom[ 7906]='h000010c2;
    rd_cycle[ 7907] = 1'b1;  wr_cycle[ 7907] = 1'b0;  addr_rom[ 7907]='h00001308;  wr_data_rom[ 7907]='h00000000;
    rd_cycle[ 7908] = 1'b1;  wr_cycle[ 7908] = 1'b0;  addr_rom[ 7908]='h00000d2c;  wr_data_rom[ 7908]='h00000000;
    rd_cycle[ 7909] = 1'b1;  wr_cycle[ 7909] = 1'b0;  addr_rom[ 7909]='h00001234;  wr_data_rom[ 7909]='h00000000;
    rd_cycle[ 7910] = 1'b0;  wr_cycle[ 7910] = 1'b1;  addr_rom[ 7910]='h000018a0;  wr_data_rom[ 7910]='h000000ec;
    rd_cycle[ 7911] = 1'b1;  wr_cycle[ 7911] = 1'b0;  addr_rom[ 7911]='h00001b94;  wr_data_rom[ 7911]='h00000000;
    rd_cycle[ 7912] = 1'b0;  wr_cycle[ 7912] = 1'b1;  addr_rom[ 7912]='h00001248;  wr_data_rom[ 7912]='h00000ce3;
    rd_cycle[ 7913] = 1'b1;  wr_cycle[ 7913] = 1'b0;  addr_rom[ 7913]='h00001b88;  wr_data_rom[ 7913]='h00000000;
    rd_cycle[ 7914] = 1'b1;  wr_cycle[ 7914] = 1'b0;  addr_rom[ 7914]='h00000f7c;  wr_data_rom[ 7914]='h00000000;
    rd_cycle[ 7915] = 1'b1;  wr_cycle[ 7915] = 1'b0;  addr_rom[ 7915]='h00001c04;  wr_data_rom[ 7915]='h00000000;
    rd_cycle[ 7916] = 1'b0;  wr_cycle[ 7916] = 1'b1;  addr_rom[ 7916]='h00000464;  wr_data_rom[ 7916]='h000015e8;
    rd_cycle[ 7917] = 1'b1;  wr_cycle[ 7917] = 1'b0;  addr_rom[ 7917]='h000010ec;  wr_data_rom[ 7917]='h00000000;
    rd_cycle[ 7918] = 1'b0;  wr_cycle[ 7918] = 1'b1;  addr_rom[ 7918]='h000009f4;  wr_data_rom[ 7918]='h00001e50;
    rd_cycle[ 7919] = 1'b0;  wr_cycle[ 7919] = 1'b1;  addr_rom[ 7919]='h00001d98;  wr_data_rom[ 7919]='h00001c11;
    rd_cycle[ 7920] = 1'b0;  wr_cycle[ 7920] = 1'b1;  addr_rom[ 7920]='h000013d4;  wr_data_rom[ 7920]='h00001549;
    rd_cycle[ 7921] = 1'b1;  wr_cycle[ 7921] = 1'b0;  addr_rom[ 7921]='h00001d8c;  wr_data_rom[ 7921]='h00000000;
    rd_cycle[ 7922] = 1'b0;  wr_cycle[ 7922] = 1'b1;  addr_rom[ 7922]='h0000129c;  wr_data_rom[ 7922]='h00001dd3;
    rd_cycle[ 7923] = 1'b0;  wr_cycle[ 7923] = 1'b1;  addr_rom[ 7923]='h0000178c;  wr_data_rom[ 7923]='h00000a68;
    rd_cycle[ 7924] = 1'b0;  wr_cycle[ 7924] = 1'b1;  addr_rom[ 7924]='h000016e8;  wr_data_rom[ 7924]='h000005be;
    rd_cycle[ 7925] = 1'b1;  wr_cycle[ 7925] = 1'b0;  addr_rom[ 7925]='h0000000c;  wr_data_rom[ 7925]='h00000000;
    rd_cycle[ 7926] = 1'b0;  wr_cycle[ 7926] = 1'b1;  addr_rom[ 7926]='h000013e0;  wr_data_rom[ 7926]='h000004c7;
    rd_cycle[ 7927] = 1'b1;  wr_cycle[ 7927] = 1'b0;  addr_rom[ 7927]='h00000c30;  wr_data_rom[ 7927]='h00000000;
    rd_cycle[ 7928] = 1'b0;  wr_cycle[ 7928] = 1'b1;  addr_rom[ 7928]='h00001f00;  wr_data_rom[ 7928]='h00001a0e;
    rd_cycle[ 7929] = 1'b1;  wr_cycle[ 7929] = 1'b0;  addr_rom[ 7929]='h000005c4;  wr_data_rom[ 7929]='h00000000;
    rd_cycle[ 7930] = 1'b0;  wr_cycle[ 7930] = 1'b1;  addr_rom[ 7930]='h00000284;  wr_data_rom[ 7930]='h00001326;
    rd_cycle[ 7931] = 1'b1;  wr_cycle[ 7931] = 1'b0;  addr_rom[ 7931]='h00000884;  wr_data_rom[ 7931]='h00000000;
    rd_cycle[ 7932] = 1'b0;  wr_cycle[ 7932] = 1'b1;  addr_rom[ 7932]='h000006e0;  wr_data_rom[ 7932]='h00000e5c;
    rd_cycle[ 7933] = 1'b0;  wr_cycle[ 7933] = 1'b1;  addr_rom[ 7933]='h000019c0;  wr_data_rom[ 7933]='h00000ba9;
    rd_cycle[ 7934] = 1'b1;  wr_cycle[ 7934] = 1'b0;  addr_rom[ 7934]='h00001730;  wr_data_rom[ 7934]='h00000000;
    rd_cycle[ 7935] = 1'b1;  wr_cycle[ 7935] = 1'b0;  addr_rom[ 7935]='h00001c2c;  wr_data_rom[ 7935]='h00000000;
    rd_cycle[ 7936] = 1'b1;  wr_cycle[ 7936] = 1'b0;  addr_rom[ 7936]='h000010ac;  wr_data_rom[ 7936]='h00000000;
    rd_cycle[ 7937] = 1'b0;  wr_cycle[ 7937] = 1'b1;  addr_rom[ 7937]='h00000ed0;  wr_data_rom[ 7937]='h00000f8e;
    rd_cycle[ 7938] = 1'b1;  wr_cycle[ 7938] = 1'b0;  addr_rom[ 7938]='h00000c60;  wr_data_rom[ 7938]='h00000000;
    rd_cycle[ 7939] = 1'b1;  wr_cycle[ 7939] = 1'b0;  addr_rom[ 7939]='h00000cc4;  wr_data_rom[ 7939]='h00000000;
    rd_cycle[ 7940] = 1'b1;  wr_cycle[ 7940] = 1'b0;  addr_rom[ 7940]='h00001aa0;  wr_data_rom[ 7940]='h00000000;
    rd_cycle[ 7941] = 1'b1;  wr_cycle[ 7941] = 1'b0;  addr_rom[ 7941]='h000002e8;  wr_data_rom[ 7941]='h00000000;
    rd_cycle[ 7942] = 1'b1;  wr_cycle[ 7942] = 1'b0;  addr_rom[ 7942]='h00000df4;  wr_data_rom[ 7942]='h00000000;
    rd_cycle[ 7943] = 1'b0;  wr_cycle[ 7943] = 1'b1;  addr_rom[ 7943]='h000016e0;  wr_data_rom[ 7943]='h00001d57;
    rd_cycle[ 7944] = 1'b0;  wr_cycle[ 7944] = 1'b1;  addr_rom[ 7944]='h00001048;  wr_data_rom[ 7944]='h00000839;
    rd_cycle[ 7945] = 1'b0;  wr_cycle[ 7945] = 1'b1;  addr_rom[ 7945]='h000015cc;  wr_data_rom[ 7945]='h00000008;
    rd_cycle[ 7946] = 1'b0;  wr_cycle[ 7946] = 1'b1;  addr_rom[ 7946]='h00001100;  wr_data_rom[ 7946]='h0000003c;
    rd_cycle[ 7947] = 1'b1;  wr_cycle[ 7947] = 1'b0;  addr_rom[ 7947]='h00000fa0;  wr_data_rom[ 7947]='h00000000;
    rd_cycle[ 7948] = 1'b1;  wr_cycle[ 7948] = 1'b0;  addr_rom[ 7948]='h00000a00;  wr_data_rom[ 7948]='h00000000;
    rd_cycle[ 7949] = 1'b1;  wr_cycle[ 7949] = 1'b0;  addr_rom[ 7949]='h0000026c;  wr_data_rom[ 7949]='h00000000;
    rd_cycle[ 7950] = 1'b0;  wr_cycle[ 7950] = 1'b1;  addr_rom[ 7950]='h000007bc;  wr_data_rom[ 7950]='h00001c9a;
    rd_cycle[ 7951] = 1'b0;  wr_cycle[ 7951] = 1'b1;  addr_rom[ 7951]='h00000808;  wr_data_rom[ 7951]='h000015f5;
    rd_cycle[ 7952] = 1'b0;  wr_cycle[ 7952] = 1'b1;  addr_rom[ 7952]='h00001238;  wr_data_rom[ 7952]='h000005c8;
    rd_cycle[ 7953] = 1'b0;  wr_cycle[ 7953] = 1'b1;  addr_rom[ 7953]='h000011d0;  wr_data_rom[ 7953]='h000010d1;
    rd_cycle[ 7954] = 1'b1;  wr_cycle[ 7954] = 1'b0;  addr_rom[ 7954]='h000014fc;  wr_data_rom[ 7954]='h00000000;
    rd_cycle[ 7955] = 1'b1;  wr_cycle[ 7955] = 1'b0;  addr_rom[ 7955]='h00001de0;  wr_data_rom[ 7955]='h00000000;
    rd_cycle[ 7956] = 1'b0;  wr_cycle[ 7956] = 1'b1;  addr_rom[ 7956]='h00000920;  wr_data_rom[ 7956]='h00000d21;
    rd_cycle[ 7957] = 1'b0;  wr_cycle[ 7957] = 1'b1;  addr_rom[ 7957]='h00001d70;  wr_data_rom[ 7957]='h000016c6;
    rd_cycle[ 7958] = 1'b0;  wr_cycle[ 7958] = 1'b1;  addr_rom[ 7958]='h00000184;  wr_data_rom[ 7958]='h0000187f;
    rd_cycle[ 7959] = 1'b0;  wr_cycle[ 7959] = 1'b1;  addr_rom[ 7959]='h00000cb4;  wr_data_rom[ 7959]='h00000405;
    rd_cycle[ 7960] = 1'b1;  wr_cycle[ 7960] = 1'b0;  addr_rom[ 7960]='h00000ee0;  wr_data_rom[ 7960]='h00000000;
    rd_cycle[ 7961] = 1'b0;  wr_cycle[ 7961] = 1'b1;  addr_rom[ 7961]='h00000694;  wr_data_rom[ 7961]='h000012cf;
    rd_cycle[ 7962] = 1'b0;  wr_cycle[ 7962] = 1'b1;  addr_rom[ 7962]='h0000149c;  wr_data_rom[ 7962]='h00000310;
    rd_cycle[ 7963] = 1'b1;  wr_cycle[ 7963] = 1'b0;  addr_rom[ 7963]='h0000183c;  wr_data_rom[ 7963]='h00000000;
    rd_cycle[ 7964] = 1'b0;  wr_cycle[ 7964] = 1'b1;  addr_rom[ 7964]='h00000320;  wr_data_rom[ 7964]='h00000327;
    rd_cycle[ 7965] = 1'b1;  wr_cycle[ 7965] = 1'b0;  addr_rom[ 7965]='h00001d90;  wr_data_rom[ 7965]='h00000000;
    rd_cycle[ 7966] = 1'b0;  wr_cycle[ 7966] = 1'b1;  addr_rom[ 7966]='h0000061c;  wr_data_rom[ 7966]='h00000765;
    rd_cycle[ 7967] = 1'b0;  wr_cycle[ 7967] = 1'b1;  addr_rom[ 7967]='h0000192c;  wr_data_rom[ 7967]='h00001406;
    rd_cycle[ 7968] = 1'b0;  wr_cycle[ 7968] = 1'b1;  addr_rom[ 7968]='h00000cac;  wr_data_rom[ 7968]='h00000e9b;
    rd_cycle[ 7969] = 1'b1;  wr_cycle[ 7969] = 1'b0;  addr_rom[ 7969]='h00001a80;  wr_data_rom[ 7969]='h00000000;
    rd_cycle[ 7970] = 1'b1;  wr_cycle[ 7970] = 1'b0;  addr_rom[ 7970]='h00000720;  wr_data_rom[ 7970]='h00000000;
    rd_cycle[ 7971] = 1'b0;  wr_cycle[ 7971] = 1'b1;  addr_rom[ 7971]='h00000254;  wr_data_rom[ 7971]='h00001352;
    rd_cycle[ 7972] = 1'b0;  wr_cycle[ 7972] = 1'b1;  addr_rom[ 7972]='h00000ab4;  wr_data_rom[ 7972]='h00000513;
    rd_cycle[ 7973] = 1'b1;  wr_cycle[ 7973] = 1'b0;  addr_rom[ 7973]='h00000d40;  wr_data_rom[ 7973]='h00000000;
    rd_cycle[ 7974] = 1'b1;  wr_cycle[ 7974] = 1'b0;  addr_rom[ 7974]='h00000d4c;  wr_data_rom[ 7974]='h00000000;
    rd_cycle[ 7975] = 1'b0;  wr_cycle[ 7975] = 1'b1;  addr_rom[ 7975]='h00001590;  wr_data_rom[ 7975]='h000005c7;
    rd_cycle[ 7976] = 1'b0;  wr_cycle[ 7976] = 1'b1;  addr_rom[ 7976]='h00001620;  wr_data_rom[ 7976]='h00000acb;
    rd_cycle[ 7977] = 1'b0;  wr_cycle[ 7977] = 1'b1;  addr_rom[ 7977]='h0000127c;  wr_data_rom[ 7977]='h00001ee5;
    rd_cycle[ 7978] = 1'b0;  wr_cycle[ 7978] = 1'b1;  addr_rom[ 7978]='h00000c34;  wr_data_rom[ 7978]='h00001a24;
    rd_cycle[ 7979] = 1'b0;  wr_cycle[ 7979] = 1'b1;  addr_rom[ 7979]='h00000698;  wr_data_rom[ 7979]='h000007ac;
    rd_cycle[ 7980] = 1'b0;  wr_cycle[ 7980] = 1'b1;  addr_rom[ 7980]='h00001280;  wr_data_rom[ 7980]='h000001de;
    rd_cycle[ 7981] = 1'b0;  wr_cycle[ 7981] = 1'b1;  addr_rom[ 7981]='h00001dac;  wr_data_rom[ 7981]='h00000790;
    rd_cycle[ 7982] = 1'b0;  wr_cycle[ 7982] = 1'b1;  addr_rom[ 7982]='h000000d4;  wr_data_rom[ 7982]='h00001e4e;
    rd_cycle[ 7983] = 1'b0;  wr_cycle[ 7983] = 1'b1;  addr_rom[ 7983]='h00001388;  wr_data_rom[ 7983]='h000012c5;
    rd_cycle[ 7984] = 1'b0;  wr_cycle[ 7984] = 1'b1;  addr_rom[ 7984]='h000012dc;  wr_data_rom[ 7984]='h00001d7c;
    rd_cycle[ 7985] = 1'b1;  wr_cycle[ 7985] = 1'b0;  addr_rom[ 7985]='h0000015c;  wr_data_rom[ 7985]='h00000000;
    rd_cycle[ 7986] = 1'b0;  wr_cycle[ 7986] = 1'b1;  addr_rom[ 7986]='h00001ac8;  wr_data_rom[ 7986]='h00001e3b;
    rd_cycle[ 7987] = 1'b1;  wr_cycle[ 7987] = 1'b0;  addr_rom[ 7987]='h00000d0c;  wr_data_rom[ 7987]='h00000000;
    rd_cycle[ 7988] = 1'b1;  wr_cycle[ 7988] = 1'b0;  addr_rom[ 7988]='h00000408;  wr_data_rom[ 7988]='h00000000;
    rd_cycle[ 7989] = 1'b0;  wr_cycle[ 7989] = 1'b1;  addr_rom[ 7989]='h000010ac;  wr_data_rom[ 7989]='h0000006a;
    rd_cycle[ 7990] = 1'b1;  wr_cycle[ 7990] = 1'b0;  addr_rom[ 7990]='h00001db0;  wr_data_rom[ 7990]='h00000000;
    rd_cycle[ 7991] = 1'b0;  wr_cycle[ 7991] = 1'b1;  addr_rom[ 7991]='h00000388;  wr_data_rom[ 7991]='h000010aa;
    rd_cycle[ 7992] = 1'b0;  wr_cycle[ 7992] = 1'b1;  addr_rom[ 7992]='h00001cb8;  wr_data_rom[ 7992]='h00000951;
    rd_cycle[ 7993] = 1'b1;  wr_cycle[ 7993] = 1'b0;  addr_rom[ 7993]='h00000b94;  wr_data_rom[ 7993]='h00000000;
    rd_cycle[ 7994] = 1'b1;  wr_cycle[ 7994] = 1'b0;  addr_rom[ 7994]='h00001ba8;  wr_data_rom[ 7994]='h00000000;
    rd_cycle[ 7995] = 1'b0;  wr_cycle[ 7995] = 1'b1;  addr_rom[ 7995]='h00000938;  wr_data_rom[ 7995]='h00001c11;
    rd_cycle[ 7996] = 1'b1;  wr_cycle[ 7996] = 1'b0;  addr_rom[ 7996]='h0000018c;  wr_data_rom[ 7996]='h00000000;
    rd_cycle[ 7997] = 1'b0;  wr_cycle[ 7997] = 1'b1;  addr_rom[ 7997]='h000011d0;  wr_data_rom[ 7997]='h00000ccf;
    rd_cycle[ 7998] = 1'b1;  wr_cycle[ 7998] = 1'b0;  addr_rom[ 7998]='h0000063c;  wr_data_rom[ 7998]='h00000000;
    rd_cycle[ 7999] = 1'b1;  wr_cycle[ 7999] = 1'b0;  addr_rom[ 7999]='h00001d30;  wr_data_rom[ 7999]='h00000000;
    // 2000 silence cycles
    rd_cycle[ 8000] = 1'b0;  wr_cycle[ 8000] = 1'b0;  addr_rom[ 8000]='h00000000;  wr_data_rom[ 8000]='h00000000;
    rd_cycle[ 8001] = 1'b0;  wr_cycle[ 8001] = 1'b0;  addr_rom[ 8001]='h00000000;  wr_data_rom[ 8001]='h00000000;
    rd_cycle[ 8002] = 1'b0;  wr_cycle[ 8002] = 1'b0;  addr_rom[ 8002]='h00000000;  wr_data_rom[ 8002]='h00000000;
    rd_cycle[ 8003] = 1'b0;  wr_cycle[ 8003] = 1'b0;  addr_rom[ 8003]='h00000000;  wr_data_rom[ 8003]='h00000000;
    rd_cycle[ 8004] = 1'b0;  wr_cycle[ 8004] = 1'b0;  addr_rom[ 8004]='h00000000;  wr_data_rom[ 8004]='h00000000;
    rd_cycle[ 8005] = 1'b0;  wr_cycle[ 8005] = 1'b0;  addr_rom[ 8005]='h00000000;  wr_data_rom[ 8005]='h00000000;
    rd_cycle[ 8006] = 1'b0;  wr_cycle[ 8006] = 1'b0;  addr_rom[ 8006]='h00000000;  wr_data_rom[ 8006]='h00000000;
    rd_cycle[ 8007] = 1'b0;  wr_cycle[ 8007] = 1'b0;  addr_rom[ 8007]='h00000000;  wr_data_rom[ 8007]='h00000000;
    rd_cycle[ 8008] = 1'b0;  wr_cycle[ 8008] = 1'b0;  addr_rom[ 8008]='h00000000;  wr_data_rom[ 8008]='h00000000;
    rd_cycle[ 8009] = 1'b0;  wr_cycle[ 8009] = 1'b0;  addr_rom[ 8009]='h00000000;  wr_data_rom[ 8009]='h00000000;
    rd_cycle[ 8010] = 1'b0;  wr_cycle[ 8010] = 1'b0;  addr_rom[ 8010]='h00000000;  wr_data_rom[ 8010]='h00000000;
    rd_cycle[ 8011] = 1'b0;  wr_cycle[ 8011] = 1'b0;  addr_rom[ 8011]='h00000000;  wr_data_rom[ 8011]='h00000000;
    rd_cycle[ 8012] = 1'b0;  wr_cycle[ 8012] = 1'b0;  addr_rom[ 8012]='h00000000;  wr_data_rom[ 8012]='h00000000;
    rd_cycle[ 8013] = 1'b0;  wr_cycle[ 8013] = 1'b0;  addr_rom[ 8013]='h00000000;  wr_data_rom[ 8013]='h00000000;
    rd_cycle[ 8014] = 1'b0;  wr_cycle[ 8014] = 1'b0;  addr_rom[ 8014]='h00000000;  wr_data_rom[ 8014]='h00000000;
    rd_cycle[ 8015] = 1'b0;  wr_cycle[ 8015] = 1'b0;  addr_rom[ 8015]='h00000000;  wr_data_rom[ 8015]='h00000000;
    rd_cycle[ 8016] = 1'b0;  wr_cycle[ 8016] = 1'b0;  addr_rom[ 8016]='h00000000;  wr_data_rom[ 8016]='h00000000;
    rd_cycle[ 8017] = 1'b0;  wr_cycle[ 8017] = 1'b0;  addr_rom[ 8017]='h00000000;  wr_data_rom[ 8017]='h00000000;
    rd_cycle[ 8018] = 1'b0;  wr_cycle[ 8018] = 1'b0;  addr_rom[ 8018]='h00000000;  wr_data_rom[ 8018]='h00000000;
    rd_cycle[ 8019] = 1'b0;  wr_cycle[ 8019] = 1'b0;  addr_rom[ 8019]='h00000000;  wr_data_rom[ 8019]='h00000000;
    rd_cycle[ 8020] = 1'b0;  wr_cycle[ 8020] = 1'b0;  addr_rom[ 8020]='h00000000;  wr_data_rom[ 8020]='h00000000;
    rd_cycle[ 8021] = 1'b0;  wr_cycle[ 8021] = 1'b0;  addr_rom[ 8021]='h00000000;  wr_data_rom[ 8021]='h00000000;
    rd_cycle[ 8022] = 1'b0;  wr_cycle[ 8022] = 1'b0;  addr_rom[ 8022]='h00000000;  wr_data_rom[ 8022]='h00000000;
    rd_cycle[ 8023] = 1'b0;  wr_cycle[ 8023] = 1'b0;  addr_rom[ 8023]='h00000000;  wr_data_rom[ 8023]='h00000000;
    rd_cycle[ 8024] = 1'b0;  wr_cycle[ 8024] = 1'b0;  addr_rom[ 8024]='h00000000;  wr_data_rom[ 8024]='h00000000;
    rd_cycle[ 8025] = 1'b0;  wr_cycle[ 8025] = 1'b0;  addr_rom[ 8025]='h00000000;  wr_data_rom[ 8025]='h00000000;
    rd_cycle[ 8026] = 1'b0;  wr_cycle[ 8026] = 1'b0;  addr_rom[ 8026]='h00000000;  wr_data_rom[ 8026]='h00000000;
    rd_cycle[ 8027] = 1'b0;  wr_cycle[ 8027] = 1'b0;  addr_rom[ 8027]='h00000000;  wr_data_rom[ 8027]='h00000000;
    rd_cycle[ 8028] = 1'b0;  wr_cycle[ 8028] = 1'b0;  addr_rom[ 8028]='h00000000;  wr_data_rom[ 8028]='h00000000;
    rd_cycle[ 8029] = 1'b0;  wr_cycle[ 8029] = 1'b0;  addr_rom[ 8029]='h00000000;  wr_data_rom[ 8029]='h00000000;
    rd_cycle[ 8030] = 1'b0;  wr_cycle[ 8030] = 1'b0;  addr_rom[ 8030]='h00000000;  wr_data_rom[ 8030]='h00000000;
    rd_cycle[ 8031] = 1'b0;  wr_cycle[ 8031] = 1'b0;  addr_rom[ 8031]='h00000000;  wr_data_rom[ 8031]='h00000000;
    rd_cycle[ 8032] = 1'b0;  wr_cycle[ 8032] = 1'b0;  addr_rom[ 8032]='h00000000;  wr_data_rom[ 8032]='h00000000;
    rd_cycle[ 8033] = 1'b0;  wr_cycle[ 8033] = 1'b0;  addr_rom[ 8033]='h00000000;  wr_data_rom[ 8033]='h00000000;
    rd_cycle[ 8034] = 1'b0;  wr_cycle[ 8034] = 1'b0;  addr_rom[ 8034]='h00000000;  wr_data_rom[ 8034]='h00000000;
    rd_cycle[ 8035] = 1'b0;  wr_cycle[ 8035] = 1'b0;  addr_rom[ 8035]='h00000000;  wr_data_rom[ 8035]='h00000000;
    rd_cycle[ 8036] = 1'b0;  wr_cycle[ 8036] = 1'b0;  addr_rom[ 8036]='h00000000;  wr_data_rom[ 8036]='h00000000;
    rd_cycle[ 8037] = 1'b0;  wr_cycle[ 8037] = 1'b0;  addr_rom[ 8037]='h00000000;  wr_data_rom[ 8037]='h00000000;
    rd_cycle[ 8038] = 1'b0;  wr_cycle[ 8038] = 1'b0;  addr_rom[ 8038]='h00000000;  wr_data_rom[ 8038]='h00000000;
    rd_cycle[ 8039] = 1'b0;  wr_cycle[ 8039] = 1'b0;  addr_rom[ 8039]='h00000000;  wr_data_rom[ 8039]='h00000000;
    rd_cycle[ 8040] = 1'b0;  wr_cycle[ 8040] = 1'b0;  addr_rom[ 8040]='h00000000;  wr_data_rom[ 8040]='h00000000;
    rd_cycle[ 8041] = 1'b0;  wr_cycle[ 8041] = 1'b0;  addr_rom[ 8041]='h00000000;  wr_data_rom[ 8041]='h00000000;
    rd_cycle[ 8042] = 1'b0;  wr_cycle[ 8042] = 1'b0;  addr_rom[ 8042]='h00000000;  wr_data_rom[ 8042]='h00000000;
    rd_cycle[ 8043] = 1'b0;  wr_cycle[ 8043] = 1'b0;  addr_rom[ 8043]='h00000000;  wr_data_rom[ 8043]='h00000000;
    rd_cycle[ 8044] = 1'b0;  wr_cycle[ 8044] = 1'b0;  addr_rom[ 8044]='h00000000;  wr_data_rom[ 8044]='h00000000;
    rd_cycle[ 8045] = 1'b0;  wr_cycle[ 8045] = 1'b0;  addr_rom[ 8045]='h00000000;  wr_data_rom[ 8045]='h00000000;
    rd_cycle[ 8046] = 1'b0;  wr_cycle[ 8046] = 1'b0;  addr_rom[ 8046]='h00000000;  wr_data_rom[ 8046]='h00000000;
    rd_cycle[ 8047] = 1'b0;  wr_cycle[ 8047] = 1'b0;  addr_rom[ 8047]='h00000000;  wr_data_rom[ 8047]='h00000000;
    rd_cycle[ 8048] = 1'b0;  wr_cycle[ 8048] = 1'b0;  addr_rom[ 8048]='h00000000;  wr_data_rom[ 8048]='h00000000;
    rd_cycle[ 8049] = 1'b0;  wr_cycle[ 8049] = 1'b0;  addr_rom[ 8049]='h00000000;  wr_data_rom[ 8049]='h00000000;
    rd_cycle[ 8050] = 1'b0;  wr_cycle[ 8050] = 1'b0;  addr_rom[ 8050]='h00000000;  wr_data_rom[ 8050]='h00000000;
    rd_cycle[ 8051] = 1'b0;  wr_cycle[ 8051] = 1'b0;  addr_rom[ 8051]='h00000000;  wr_data_rom[ 8051]='h00000000;
    rd_cycle[ 8052] = 1'b0;  wr_cycle[ 8052] = 1'b0;  addr_rom[ 8052]='h00000000;  wr_data_rom[ 8052]='h00000000;
    rd_cycle[ 8053] = 1'b0;  wr_cycle[ 8053] = 1'b0;  addr_rom[ 8053]='h00000000;  wr_data_rom[ 8053]='h00000000;
    rd_cycle[ 8054] = 1'b0;  wr_cycle[ 8054] = 1'b0;  addr_rom[ 8054]='h00000000;  wr_data_rom[ 8054]='h00000000;
    rd_cycle[ 8055] = 1'b0;  wr_cycle[ 8055] = 1'b0;  addr_rom[ 8055]='h00000000;  wr_data_rom[ 8055]='h00000000;
    rd_cycle[ 8056] = 1'b0;  wr_cycle[ 8056] = 1'b0;  addr_rom[ 8056]='h00000000;  wr_data_rom[ 8056]='h00000000;
    rd_cycle[ 8057] = 1'b0;  wr_cycle[ 8057] = 1'b0;  addr_rom[ 8057]='h00000000;  wr_data_rom[ 8057]='h00000000;
    rd_cycle[ 8058] = 1'b0;  wr_cycle[ 8058] = 1'b0;  addr_rom[ 8058]='h00000000;  wr_data_rom[ 8058]='h00000000;
    rd_cycle[ 8059] = 1'b0;  wr_cycle[ 8059] = 1'b0;  addr_rom[ 8059]='h00000000;  wr_data_rom[ 8059]='h00000000;
    rd_cycle[ 8060] = 1'b0;  wr_cycle[ 8060] = 1'b0;  addr_rom[ 8060]='h00000000;  wr_data_rom[ 8060]='h00000000;
    rd_cycle[ 8061] = 1'b0;  wr_cycle[ 8061] = 1'b0;  addr_rom[ 8061]='h00000000;  wr_data_rom[ 8061]='h00000000;
    rd_cycle[ 8062] = 1'b0;  wr_cycle[ 8062] = 1'b0;  addr_rom[ 8062]='h00000000;  wr_data_rom[ 8062]='h00000000;
    rd_cycle[ 8063] = 1'b0;  wr_cycle[ 8063] = 1'b0;  addr_rom[ 8063]='h00000000;  wr_data_rom[ 8063]='h00000000;
    rd_cycle[ 8064] = 1'b0;  wr_cycle[ 8064] = 1'b0;  addr_rom[ 8064]='h00000000;  wr_data_rom[ 8064]='h00000000;
    rd_cycle[ 8065] = 1'b0;  wr_cycle[ 8065] = 1'b0;  addr_rom[ 8065]='h00000000;  wr_data_rom[ 8065]='h00000000;
    rd_cycle[ 8066] = 1'b0;  wr_cycle[ 8066] = 1'b0;  addr_rom[ 8066]='h00000000;  wr_data_rom[ 8066]='h00000000;
    rd_cycle[ 8067] = 1'b0;  wr_cycle[ 8067] = 1'b0;  addr_rom[ 8067]='h00000000;  wr_data_rom[ 8067]='h00000000;
    rd_cycle[ 8068] = 1'b0;  wr_cycle[ 8068] = 1'b0;  addr_rom[ 8068]='h00000000;  wr_data_rom[ 8068]='h00000000;
    rd_cycle[ 8069] = 1'b0;  wr_cycle[ 8069] = 1'b0;  addr_rom[ 8069]='h00000000;  wr_data_rom[ 8069]='h00000000;
    rd_cycle[ 8070] = 1'b0;  wr_cycle[ 8070] = 1'b0;  addr_rom[ 8070]='h00000000;  wr_data_rom[ 8070]='h00000000;
    rd_cycle[ 8071] = 1'b0;  wr_cycle[ 8071] = 1'b0;  addr_rom[ 8071]='h00000000;  wr_data_rom[ 8071]='h00000000;
    rd_cycle[ 8072] = 1'b0;  wr_cycle[ 8072] = 1'b0;  addr_rom[ 8072]='h00000000;  wr_data_rom[ 8072]='h00000000;
    rd_cycle[ 8073] = 1'b0;  wr_cycle[ 8073] = 1'b0;  addr_rom[ 8073]='h00000000;  wr_data_rom[ 8073]='h00000000;
    rd_cycle[ 8074] = 1'b0;  wr_cycle[ 8074] = 1'b0;  addr_rom[ 8074]='h00000000;  wr_data_rom[ 8074]='h00000000;
    rd_cycle[ 8075] = 1'b0;  wr_cycle[ 8075] = 1'b0;  addr_rom[ 8075]='h00000000;  wr_data_rom[ 8075]='h00000000;
    rd_cycle[ 8076] = 1'b0;  wr_cycle[ 8076] = 1'b0;  addr_rom[ 8076]='h00000000;  wr_data_rom[ 8076]='h00000000;
    rd_cycle[ 8077] = 1'b0;  wr_cycle[ 8077] = 1'b0;  addr_rom[ 8077]='h00000000;  wr_data_rom[ 8077]='h00000000;
    rd_cycle[ 8078] = 1'b0;  wr_cycle[ 8078] = 1'b0;  addr_rom[ 8078]='h00000000;  wr_data_rom[ 8078]='h00000000;
    rd_cycle[ 8079] = 1'b0;  wr_cycle[ 8079] = 1'b0;  addr_rom[ 8079]='h00000000;  wr_data_rom[ 8079]='h00000000;
    rd_cycle[ 8080] = 1'b0;  wr_cycle[ 8080] = 1'b0;  addr_rom[ 8080]='h00000000;  wr_data_rom[ 8080]='h00000000;
    rd_cycle[ 8081] = 1'b0;  wr_cycle[ 8081] = 1'b0;  addr_rom[ 8081]='h00000000;  wr_data_rom[ 8081]='h00000000;
    rd_cycle[ 8082] = 1'b0;  wr_cycle[ 8082] = 1'b0;  addr_rom[ 8082]='h00000000;  wr_data_rom[ 8082]='h00000000;
    rd_cycle[ 8083] = 1'b0;  wr_cycle[ 8083] = 1'b0;  addr_rom[ 8083]='h00000000;  wr_data_rom[ 8083]='h00000000;
    rd_cycle[ 8084] = 1'b0;  wr_cycle[ 8084] = 1'b0;  addr_rom[ 8084]='h00000000;  wr_data_rom[ 8084]='h00000000;
    rd_cycle[ 8085] = 1'b0;  wr_cycle[ 8085] = 1'b0;  addr_rom[ 8085]='h00000000;  wr_data_rom[ 8085]='h00000000;
    rd_cycle[ 8086] = 1'b0;  wr_cycle[ 8086] = 1'b0;  addr_rom[ 8086]='h00000000;  wr_data_rom[ 8086]='h00000000;
    rd_cycle[ 8087] = 1'b0;  wr_cycle[ 8087] = 1'b0;  addr_rom[ 8087]='h00000000;  wr_data_rom[ 8087]='h00000000;
    rd_cycle[ 8088] = 1'b0;  wr_cycle[ 8088] = 1'b0;  addr_rom[ 8088]='h00000000;  wr_data_rom[ 8088]='h00000000;
    rd_cycle[ 8089] = 1'b0;  wr_cycle[ 8089] = 1'b0;  addr_rom[ 8089]='h00000000;  wr_data_rom[ 8089]='h00000000;
    rd_cycle[ 8090] = 1'b0;  wr_cycle[ 8090] = 1'b0;  addr_rom[ 8090]='h00000000;  wr_data_rom[ 8090]='h00000000;
    rd_cycle[ 8091] = 1'b0;  wr_cycle[ 8091] = 1'b0;  addr_rom[ 8091]='h00000000;  wr_data_rom[ 8091]='h00000000;
    rd_cycle[ 8092] = 1'b0;  wr_cycle[ 8092] = 1'b0;  addr_rom[ 8092]='h00000000;  wr_data_rom[ 8092]='h00000000;
    rd_cycle[ 8093] = 1'b0;  wr_cycle[ 8093] = 1'b0;  addr_rom[ 8093]='h00000000;  wr_data_rom[ 8093]='h00000000;
    rd_cycle[ 8094] = 1'b0;  wr_cycle[ 8094] = 1'b0;  addr_rom[ 8094]='h00000000;  wr_data_rom[ 8094]='h00000000;
    rd_cycle[ 8095] = 1'b0;  wr_cycle[ 8095] = 1'b0;  addr_rom[ 8095]='h00000000;  wr_data_rom[ 8095]='h00000000;
    rd_cycle[ 8096] = 1'b0;  wr_cycle[ 8096] = 1'b0;  addr_rom[ 8096]='h00000000;  wr_data_rom[ 8096]='h00000000;
    rd_cycle[ 8097] = 1'b0;  wr_cycle[ 8097] = 1'b0;  addr_rom[ 8097]='h00000000;  wr_data_rom[ 8097]='h00000000;
    rd_cycle[ 8098] = 1'b0;  wr_cycle[ 8098] = 1'b0;  addr_rom[ 8098]='h00000000;  wr_data_rom[ 8098]='h00000000;
    rd_cycle[ 8099] = 1'b0;  wr_cycle[ 8099] = 1'b0;  addr_rom[ 8099]='h00000000;  wr_data_rom[ 8099]='h00000000;
    rd_cycle[ 8100] = 1'b0;  wr_cycle[ 8100] = 1'b0;  addr_rom[ 8100]='h00000000;  wr_data_rom[ 8100]='h00000000;
    rd_cycle[ 8101] = 1'b0;  wr_cycle[ 8101] = 1'b0;  addr_rom[ 8101]='h00000000;  wr_data_rom[ 8101]='h00000000;
    rd_cycle[ 8102] = 1'b0;  wr_cycle[ 8102] = 1'b0;  addr_rom[ 8102]='h00000000;  wr_data_rom[ 8102]='h00000000;
    rd_cycle[ 8103] = 1'b0;  wr_cycle[ 8103] = 1'b0;  addr_rom[ 8103]='h00000000;  wr_data_rom[ 8103]='h00000000;
    rd_cycle[ 8104] = 1'b0;  wr_cycle[ 8104] = 1'b0;  addr_rom[ 8104]='h00000000;  wr_data_rom[ 8104]='h00000000;
    rd_cycle[ 8105] = 1'b0;  wr_cycle[ 8105] = 1'b0;  addr_rom[ 8105]='h00000000;  wr_data_rom[ 8105]='h00000000;
    rd_cycle[ 8106] = 1'b0;  wr_cycle[ 8106] = 1'b0;  addr_rom[ 8106]='h00000000;  wr_data_rom[ 8106]='h00000000;
    rd_cycle[ 8107] = 1'b0;  wr_cycle[ 8107] = 1'b0;  addr_rom[ 8107]='h00000000;  wr_data_rom[ 8107]='h00000000;
    rd_cycle[ 8108] = 1'b0;  wr_cycle[ 8108] = 1'b0;  addr_rom[ 8108]='h00000000;  wr_data_rom[ 8108]='h00000000;
    rd_cycle[ 8109] = 1'b0;  wr_cycle[ 8109] = 1'b0;  addr_rom[ 8109]='h00000000;  wr_data_rom[ 8109]='h00000000;
    rd_cycle[ 8110] = 1'b0;  wr_cycle[ 8110] = 1'b0;  addr_rom[ 8110]='h00000000;  wr_data_rom[ 8110]='h00000000;
    rd_cycle[ 8111] = 1'b0;  wr_cycle[ 8111] = 1'b0;  addr_rom[ 8111]='h00000000;  wr_data_rom[ 8111]='h00000000;
    rd_cycle[ 8112] = 1'b0;  wr_cycle[ 8112] = 1'b0;  addr_rom[ 8112]='h00000000;  wr_data_rom[ 8112]='h00000000;
    rd_cycle[ 8113] = 1'b0;  wr_cycle[ 8113] = 1'b0;  addr_rom[ 8113]='h00000000;  wr_data_rom[ 8113]='h00000000;
    rd_cycle[ 8114] = 1'b0;  wr_cycle[ 8114] = 1'b0;  addr_rom[ 8114]='h00000000;  wr_data_rom[ 8114]='h00000000;
    rd_cycle[ 8115] = 1'b0;  wr_cycle[ 8115] = 1'b0;  addr_rom[ 8115]='h00000000;  wr_data_rom[ 8115]='h00000000;
    rd_cycle[ 8116] = 1'b0;  wr_cycle[ 8116] = 1'b0;  addr_rom[ 8116]='h00000000;  wr_data_rom[ 8116]='h00000000;
    rd_cycle[ 8117] = 1'b0;  wr_cycle[ 8117] = 1'b0;  addr_rom[ 8117]='h00000000;  wr_data_rom[ 8117]='h00000000;
    rd_cycle[ 8118] = 1'b0;  wr_cycle[ 8118] = 1'b0;  addr_rom[ 8118]='h00000000;  wr_data_rom[ 8118]='h00000000;
    rd_cycle[ 8119] = 1'b0;  wr_cycle[ 8119] = 1'b0;  addr_rom[ 8119]='h00000000;  wr_data_rom[ 8119]='h00000000;
    rd_cycle[ 8120] = 1'b0;  wr_cycle[ 8120] = 1'b0;  addr_rom[ 8120]='h00000000;  wr_data_rom[ 8120]='h00000000;
    rd_cycle[ 8121] = 1'b0;  wr_cycle[ 8121] = 1'b0;  addr_rom[ 8121]='h00000000;  wr_data_rom[ 8121]='h00000000;
    rd_cycle[ 8122] = 1'b0;  wr_cycle[ 8122] = 1'b0;  addr_rom[ 8122]='h00000000;  wr_data_rom[ 8122]='h00000000;
    rd_cycle[ 8123] = 1'b0;  wr_cycle[ 8123] = 1'b0;  addr_rom[ 8123]='h00000000;  wr_data_rom[ 8123]='h00000000;
    rd_cycle[ 8124] = 1'b0;  wr_cycle[ 8124] = 1'b0;  addr_rom[ 8124]='h00000000;  wr_data_rom[ 8124]='h00000000;
    rd_cycle[ 8125] = 1'b0;  wr_cycle[ 8125] = 1'b0;  addr_rom[ 8125]='h00000000;  wr_data_rom[ 8125]='h00000000;
    rd_cycle[ 8126] = 1'b0;  wr_cycle[ 8126] = 1'b0;  addr_rom[ 8126]='h00000000;  wr_data_rom[ 8126]='h00000000;
    rd_cycle[ 8127] = 1'b0;  wr_cycle[ 8127] = 1'b0;  addr_rom[ 8127]='h00000000;  wr_data_rom[ 8127]='h00000000;
    rd_cycle[ 8128] = 1'b0;  wr_cycle[ 8128] = 1'b0;  addr_rom[ 8128]='h00000000;  wr_data_rom[ 8128]='h00000000;
    rd_cycle[ 8129] = 1'b0;  wr_cycle[ 8129] = 1'b0;  addr_rom[ 8129]='h00000000;  wr_data_rom[ 8129]='h00000000;
    rd_cycle[ 8130] = 1'b0;  wr_cycle[ 8130] = 1'b0;  addr_rom[ 8130]='h00000000;  wr_data_rom[ 8130]='h00000000;
    rd_cycle[ 8131] = 1'b0;  wr_cycle[ 8131] = 1'b0;  addr_rom[ 8131]='h00000000;  wr_data_rom[ 8131]='h00000000;
    rd_cycle[ 8132] = 1'b0;  wr_cycle[ 8132] = 1'b0;  addr_rom[ 8132]='h00000000;  wr_data_rom[ 8132]='h00000000;
    rd_cycle[ 8133] = 1'b0;  wr_cycle[ 8133] = 1'b0;  addr_rom[ 8133]='h00000000;  wr_data_rom[ 8133]='h00000000;
    rd_cycle[ 8134] = 1'b0;  wr_cycle[ 8134] = 1'b0;  addr_rom[ 8134]='h00000000;  wr_data_rom[ 8134]='h00000000;
    rd_cycle[ 8135] = 1'b0;  wr_cycle[ 8135] = 1'b0;  addr_rom[ 8135]='h00000000;  wr_data_rom[ 8135]='h00000000;
    rd_cycle[ 8136] = 1'b0;  wr_cycle[ 8136] = 1'b0;  addr_rom[ 8136]='h00000000;  wr_data_rom[ 8136]='h00000000;
    rd_cycle[ 8137] = 1'b0;  wr_cycle[ 8137] = 1'b0;  addr_rom[ 8137]='h00000000;  wr_data_rom[ 8137]='h00000000;
    rd_cycle[ 8138] = 1'b0;  wr_cycle[ 8138] = 1'b0;  addr_rom[ 8138]='h00000000;  wr_data_rom[ 8138]='h00000000;
    rd_cycle[ 8139] = 1'b0;  wr_cycle[ 8139] = 1'b0;  addr_rom[ 8139]='h00000000;  wr_data_rom[ 8139]='h00000000;
    rd_cycle[ 8140] = 1'b0;  wr_cycle[ 8140] = 1'b0;  addr_rom[ 8140]='h00000000;  wr_data_rom[ 8140]='h00000000;
    rd_cycle[ 8141] = 1'b0;  wr_cycle[ 8141] = 1'b0;  addr_rom[ 8141]='h00000000;  wr_data_rom[ 8141]='h00000000;
    rd_cycle[ 8142] = 1'b0;  wr_cycle[ 8142] = 1'b0;  addr_rom[ 8142]='h00000000;  wr_data_rom[ 8142]='h00000000;
    rd_cycle[ 8143] = 1'b0;  wr_cycle[ 8143] = 1'b0;  addr_rom[ 8143]='h00000000;  wr_data_rom[ 8143]='h00000000;
    rd_cycle[ 8144] = 1'b0;  wr_cycle[ 8144] = 1'b0;  addr_rom[ 8144]='h00000000;  wr_data_rom[ 8144]='h00000000;
    rd_cycle[ 8145] = 1'b0;  wr_cycle[ 8145] = 1'b0;  addr_rom[ 8145]='h00000000;  wr_data_rom[ 8145]='h00000000;
    rd_cycle[ 8146] = 1'b0;  wr_cycle[ 8146] = 1'b0;  addr_rom[ 8146]='h00000000;  wr_data_rom[ 8146]='h00000000;
    rd_cycle[ 8147] = 1'b0;  wr_cycle[ 8147] = 1'b0;  addr_rom[ 8147]='h00000000;  wr_data_rom[ 8147]='h00000000;
    rd_cycle[ 8148] = 1'b0;  wr_cycle[ 8148] = 1'b0;  addr_rom[ 8148]='h00000000;  wr_data_rom[ 8148]='h00000000;
    rd_cycle[ 8149] = 1'b0;  wr_cycle[ 8149] = 1'b0;  addr_rom[ 8149]='h00000000;  wr_data_rom[ 8149]='h00000000;
    rd_cycle[ 8150] = 1'b0;  wr_cycle[ 8150] = 1'b0;  addr_rom[ 8150]='h00000000;  wr_data_rom[ 8150]='h00000000;
    rd_cycle[ 8151] = 1'b0;  wr_cycle[ 8151] = 1'b0;  addr_rom[ 8151]='h00000000;  wr_data_rom[ 8151]='h00000000;
    rd_cycle[ 8152] = 1'b0;  wr_cycle[ 8152] = 1'b0;  addr_rom[ 8152]='h00000000;  wr_data_rom[ 8152]='h00000000;
    rd_cycle[ 8153] = 1'b0;  wr_cycle[ 8153] = 1'b0;  addr_rom[ 8153]='h00000000;  wr_data_rom[ 8153]='h00000000;
    rd_cycle[ 8154] = 1'b0;  wr_cycle[ 8154] = 1'b0;  addr_rom[ 8154]='h00000000;  wr_data_rom[ 8154]='h00000000;
    rd_cycle[ 8155] = 1'b0;  wr_cycle[ 8155] = 1'b0;  addr_rom[ 8155]='h00000000;  wr_data_rom[ 8155]='h00000000;
    rd_cycle[ 8156] = 1'b0;  wr_cycle[ 8156] = 1'b0;  addr_rom[ 8156]='h00000000;  wr_data_rom[ 8156]='h00000000;
    rd_cycle[ 8157] = 1'b0;  wr_cycle[ 8157] = 1'b0;  addr_rom[ 8157]='h00000000;  wr_data_rom[ 8157]='h00000000;
    rd_cycle[ 8158] = 1'b0;  wr_cycle[ 8158] = 1'b0;  addr_rom[ 8158]='h00000000;  wr_data_rom[ 8158]='h00000000;
    rd_cycle[ 8159] = 1'b0;  wr_cycle[ 8159] = 1'b0;  addr_rom[ 8159]='h00000000;  wr_data_rom[ 8159]='h00000000;
    rd_cycle[ 8160] = 1'b0;  wr_cycle[ 8160] = 1'b0;  addr_rom[ 8160]='h00000000;  wr_data_rom[ 8160]='h00000000;
    rd_cycle[ 8161] = 1'b0;  wr_cycle[ 8161] = 1'b0;  addr_rom[ 8161]='h00000000;  wr_data_rom[ 8161]='h00000000;
    rd_cycle[ 8162] = 1'b0;  wr_cycle[ 8162] = 1'b0;  addr_rom[ 8162]='h00000000;  wr_data_rom[ 8162]='h00000000;
    rd_cycle[ 8163] = 1'b0;  wr_cycle[ 8163] = 1'b0;  addr_rom[ 8163]='h00000000;  wr_data_rom[ 8163]='h00000000;
    rd_cycle[ 8164] = 1'b0;  wr_cycle[ 8164] = 1'b0;  addr_rom[ 8164]='h00000000;  wr_data_rom[ 8164]='h00000000;
    rd_cycle[ 8165] = 1'b0;  wr_cycle[ 8165] = 1'b0;  addr_rom[ 8165]='h00000000;  wr_data_rom[ 8165]='h00000000;
    rd_cycle[ 8166] = 1'b0;  wr_cycle[ 8166] = 1'b0;  addr_rom[ 8166]='h00000000;  wr_data_rom[ 8166]='h00000000;
    rd_cycle[ 8167] = 1'b0;  wr_cycle[ 8167] = 1'b0;  addr_rom[ 8167]='h00000000;  wr_data_rom[ 8167]='h00000000;
    rd_cycle[ 8168] = 1'b0;  wr_cycle[ 8168] = 1'b0;  addr_rom[ 8168]='h00000000;  wr_data_rom[ 8168]='h00000000;
    rd_cycle[ 8169] = 1'b0;  wr_cycle[ 8169] = 1'b0;  addr_rom[ 8169]='h00000000;  wr_data_rom[ 8169]='h00000000;
    rd_cycle[ 8170] = 1'b0;  wr_cycle[ 8170] = 1'b0;  addr_rom[ 8170]='h00000000;  wr_data_rom[ 8170]='h00000000;
    rd_cycle[ 8171] = 1'b0;  wr_cycle[ 8171] = 1'b0;  addr_rom[ 8171]='h00000000;  wr_data_rom[ 8171]='h00000000;
    rd_cycle[ 8172] = 1'b0;  wr_cycle[ 8172] = 1'b0;  addr_rom[ 8172]='h00000000;  wr_data_rom[ 8172]='h00000000;
    rd_cycle[ 8173] = 1'b0;  wr_cycle[ 8173] = 1'b0;  addr_rom[ 8173]='h00000000;  wr_data_rom[ 8173]='h00000000;
    rd_cycle[ 8174] = 1'b0;  wr_cycle[ 8174] = 1'b0;  addr_rom[ 8174]='h00000000;  wr_data_rom[ 8174]='h00000000;
    rd_cycle[ 8175] = 1'b0;  wr_cycle[ 8175] = 1'b0;  addr_rom[ 8175]='h00000000;  wr_data_rom[ 8175]='h00000000;
    rd_cycle[ 8176] = 1'b0;  wr_cycle[ 8176] = 1'b0;  addr_rom[ 8176]='h00000000;  wr_data_rom[ 8176]='h00000000;
    rd_cycle[ 8177] = 1'b0;  wr_cycle[ 8177] = 1'b0;  addr_rom[ 8177]='h00000000;  wr_data_rom[ 8177]='h00000000;
    rd_cycle[ 8178] = 1'b0;  wr_cycle[ 8178] = 1'b0;  addr_rom[ 8178]='h00000000;  wr_data_rom[ 8178]='h00000000;
    rd_cycle[ 8179] = 1'b0;  wr_cycle[ 8179] = 1'b0;  addr_rom[ 8179]='h00000000;  wr_data_rom[ 8179]='h00000000;
    rd_cycle[ 8180] = 1'b0;  wr_cycle[ 8180] = 1'b0;  addr_rom[ 8180]='h00000000;  wr_data_rom[ 8180]='h00000000;
    rd_cycle[ 8181] = 1'b0;  wr_cycle[ 8181] = 1'b0;  addr_rom[ 8181]='h00000000;  wr_data_rom[ 8181]='h00000000;
    rd_cycle[ 8182] = 1'b0;  wr_cycle[ 8182] = 1'b0;  addr_rom[ 8182]='h00000000;  wr_data_rom[ 8182]='h00000000;
    rd_cycle[ 8183] = 1'b0;  wr_cycle[ 8183] = 1'b0;  addr_rom[ 8183]='h00000000;  wr_data_rom[ 8183]='h00000000;
    rd_cycle[ 8184] = 1'b0;  wr_cycle[ 8184] = 1'b0;  addr_rom[ 8184]='h00000000;  wr_data_rom[ 8184]='h00000000;
    rd_cycle[ 8185] = 1'b0;  wr_cycle[ 8185] = 1'b0;  addr_rom[ 8185]='h00000000;  wr_data_rom[ 8185]='h00000000;
    rd_cycle[ 8186] = 1'b0;  wr_cycle[ 8186] = 1'b0;  addr_rom[ 8186]='h00000000;  wr_data_rom[ 8186]='h00000000;
    rd_cycle[ 8187] = 1'b0;  wr_cycle[ 8187] = 1'b0;  addr_rom[ 8187]='h00000000;  wr_data_rom[ 8187]='h00000000;
    rd_cycle[ 8188] = 1'b0;  wr_cycle[ 8188] = 1'b0;  addr_rom[ 8188]='h00000000;  wr_data_rom[ 8188]='h00000000;
    rd_cycle[ 8189] = 1'b0;  wr_cycle[ 8189] = 1'b0;  addr_rom[ 8189]='h00000000;  wr_data_rom[ 8189]='h00000000;
    rd_cycle[ 8190] = 1'b0;  wr_cycle[ 8190] = 1'b0;  addr_rom[ 8190]='h00000000;  wr_data_rom[ 8190]='h00000000;
    rd_cycle[ 8191] = 1'b0;  wr_cycle[ 8191] = 1'b0;  addr_rom[ 8191]='h00000000;  wr_data_rom[ 8191]='h00000000;
    rd_cycle[ 8192] = 1'b0;  wr_cycle[ 8192] = 1'b0;  addr_rom[ 8192]='h00000000;  wr_data_rom[ 8192]='h00000000;
    rd_cycle[ 8193] = 1'b0;  wr_cycle[ 8193] = 1'b0;  addr_rom[ 8193]='h00000000;  wr_data_rom[ 8193]='h00000000;
    rd_cycle[ 8194] = 1'b0;  wr_cycle[ 8194] = 1'b0;  addr_rom[ 8194]='h00000000;  wr_data_rom[ 8194]='h00000000;
    rd_cycle[ 8195] = 1'b0;  wr_cycle[ 8195] = 1'b0;  addr_rom[ 8195]='h00000000;  wr_data_rom[ 8195]='h00000000;
    rd_cycle[ 8196] = 1'b0;  wr_cycle[ 8196] = 1'b0;  addr_rom[ 8196]='h00000000;  wr_data_rom[ 8196]='h00000000;
    rd_cycle[ 8197] = 1'b0;  wr_cycle[ 8197] = 1'b0;  addr_rom[ 8197]='h00000000;  wr_data_rom[ 8197]='h00000000;
    rd_cycle[ 8198] = 1'b0;  wr_cycle[ 8198] = 1'b0;  addr_rom[ 8198]='h00000000;  wr_data_rom[ 8198]='h00000000;
    rd_cycle[ 8199] = 1'b0;  wr_cycle[ 8199] = 1'b0;  addr_rom[ 8199]='h00000000;  wr_data_rom[ 8199]='h00000000;
    rd_cycle[ 8200] = 1'b0;  wr_cycle[ 8200] = 1'b0;  addr_rom[ 8200]='h00000000;  wr_data_rom[ 8200]='h00000000;
    rd_cycle[ 8201] = 1'b0;  wr_cycle[ 8201] = 1'b0;  addr_rom[ 8201]='h00000000;  wr_data_rom[ 8201]='h00000000;
    rd_cycle[ 8202] = 1'b0;  wr_cycle[ 8202] = 1'b0;  addr_rom[ 8202]='h00000000;  wr_data_rom[ 8202]='h00000000;
    rd_cycle[ 8203] = 1'b0;  wr_cycle[ 8203] = 1'b0;  addr_rom[ 8203]='h00000000;  wr_data_rom[ 8203]='h00000000;
    rd_cycle[ 8204] = 1'b0;  wr_cycle[ 8204] = 1'b0;  addr_rom[ 8204]='h00000000;  wr_data_rom[ 8204]='h00000000;
    rd_cycle[ 8205] = 1'b0;  wr_cycle[ 8205] = 1'b0;  addr_rom[ 8205]='h00000000;  wr_data_rom[ 8205]='h00000000;
    rd_cycle[ 8206] = 1'b0;  wr_cycle[ 8206] = 1'b0;  addr_rom[ 8206]='h00000000;  wr_data_rom[ 8206]='h00000000;
    rd_cycle[ 8207] = 1'b0;  wr_cycle[ 8207] = 1'b0;  addr_rom[ 8207]='h00000000;  wr_data_rom[ 8207]='h00000000;
    rd_cycle[ 8208] = 1'b0;  wr_cycle[ 8208] = 1'b0;  addr_rom[ 8208]='h00000000;  wr_data_rom[ 8208]='h00000000;
    rd_cycle[ 8209] = 1'b0;  wr_cycle[ 8209] = 1'b0;  addr_rom[ 8209]='h00000000;  wr_data_rom[ 8209]='h00000000;
    rd_cycle[ 8210] = 1'b0;  wr_cycle[ 8210] = 1'b0;  addr_rom[ 8210]='h00000000;  wr_data_rom[ 8210]='h00000000;
    rd_cycle[ 8211] = 1'b0;  wr_cycle[ 8211] = 1'b0;  addr_rom[ 8211]='h00000000;  wr_data_rom[ 8211]='h00000000;
    rd_cycle[ 8212] = 1'b0;  wr_cycle[ 8212] = 1'b0;  addr_rom[ 8212]='h00000000;  wr_data_rom[ 8212]='h00000000;
    rd_cycle[ 8213] = 1'b0;  wr_cycle[ 8213] = 1'b0;  addr_rom[ 8213]='h00000000;  wr_data_rom[ 8213]='h00000000;
    rd_cycle[ 8214] = 1'b0;  wr_cycle[ 8214] = 1'b0;  addr_rom[ 8214]='h00000000;  wr_data_rom[ 8214]='h00000000;
    rd_cycle[ 8215] = 1'b0;  wr_cycle[ 8215] = 1'b0;  addr_rom[ 8215]='h00000000;  wr_data_rom[ 8215]='h00000000;
    rd_cycle[ 8216] = 1'b0;  wr_cycle[ 8216] = 1'b0;  addr_rom[ 8216]='h00000000;  wr_data_rom[ 8216]='h00000000;
    rd_cycle[ 8217] = 1'b0;  wr_cycle[ 8217] = 1'b0;  addr_rom[ 8217]='h00000000;  wr_data_rom[ 8217]='h00000000;
    rd_cycle[ 8218] = 1'b0;  wr_cycle[ 8218] = 1'b0;  addr_rom[ 8218]='h00000000;  wr_data_rom[ 8218]='h00000000;
    rd_cycle[ 8219] = 1'b0;  wr_cycle[ 8219] = 1'b0;  addr_rom[ 8219]='h00000000;  wr_data_rom[ 8219]='h00000000;
    rd_cycle[ 8220] = 1'b0;  wr_cycle[ 8220] = 1'b0;  addr_rom[ 8220]='h00000000;  wr_data_rom[ 8220]='h00000000;
    rd_cycle[ 8221] = 1'b0;  wr_cycle[ 8221] = 1'b0;  addr_rom[ 8221]='h00000000;  wr_data_rom[ 8221]='h00000000;
    rd_cycle[ 8222] = 1'b0;  wr_cycle[ 8222] = 1'b0;  addr_rom[ 8222]='h00000000;  wr_data_rom[ 8222]='h00000000;
    rd_cycle[ 8223] = 1'b0;  wr_cycle[ 8223] = 1'b0;  addr_rom[ 8223]='h00000000;  wr_data_rom[ 8223]='h00000000;
    rd_cycle[ 8224] = 1'b0;  wr_cycle[ 8224] = 1'b0;  addr_rom[ 8224]='h00000000;  wr_data_rom[ 8224]='h00000000;
    rd_cycle[ 8225] = 1'b0;  wr_cycle[ 8225] = 1'b0;  addr_rom[ 8225]='h00000000;  wr_data_rom[ 8225]='h00000000;
    rd_cycle[ 8226] = 1'b0;  wr_cycle[ 8226] = 1'b0;  addr_rom[ 8226]='h00000000;  wr_data_rom[ 8226]='h00000000;
    rd_cycle[ 8227] = 1'b0;  wr_cycle[ 8227] = 1'b0;  addr_rom[ 8227]='h00000000;  wr_data_rom[ 8227]='h00000000;
    rd_cycle[ 8228] = 1'b0;  wr_cycle[ 8228] = 1'b0;  addr_rom[ 8228]='h00000000;  wr_data_rom[ 8228]='h00000000;
    rd_cycle[ 8229] = 1'b0;  wr_cycle[ 8229] = 1'b0;  addr_rom[ 8229]='h00000000;  wr_data_rom[ 8229]='h00000000;
    rd_cycle[ 8230] = 1'b0;  wr_cycle[ 8230] = 1'b0;  addr_rom[ 8230]='h00000000;  wr_data_rom[ 8230]='h00000000;
    rd_cycle[ 8231] = 1'b0;  wr_cycle[ 8231] = 1'b0;  addr_rom[ 8231]='h00000000;  wr_data_rom[ 8231]='h00000000;
    rd_cycle[ 8232] = 1'b0;  wr_cycle[ 8232] = 1'b0;  addr_rom[ 8232]='h00000000;  wr_data_rom[ 8232]='h00000000;
    rd_cycle[ 8233] = 1'b0;  wr_cycle[ 8233] = 1'b0;  addr_rom[ 8233]='h00000000;  wr_data_rom[ 8233]='h00000000;
    rd_cycle[ 8234] = 1'b0;  wr_cycle[ 8234] = 1'b0;  addr_rom[ 8234]='h00000000;  wr_data_rom[ 8234]='h00000000;
    rd_cycle[ 8235] = 1'b0;  wr_cycle[ 8235] = 1'b0;  addr_rom[ 8235]='h00000000;  wr_data_rom[ 8235]='h00000000;
    rd_cycle[ 8236] = 1'b0;  wr_cycle[ 8236] = 1'b0;  addr_rom[ 8236]='h00000000;  wr_data_rom[ 8236]='h00000000;
    rd_cycle[ 8237] = 1'b0;  wr_cycle[ 8237] = 1'b0;  addr_rom[ 8237]='h00000000;  wr_data_rom[ 8237]='h00000000;
    rd_cycle[ 8238] = 1'b0;  wr_cycle[ 8238] = 1'b0;  addr_rom[ 8238]='h00000000;  wr_data_rom[ 8238]='h00000000;
    rd_cycle[ 8239] = 1'b0;  wr_cycle[ 8239] = 1'b0;  addr_rom[ 8239]='h00000000;  wr_data_rom[ 8239]='h00000000;
    rd_cycle[ 8240] = 1'b0;  wr_cycle[ 8240] = 1'b0;  addr_rom[ 8240]='h00000000;  wr_data_rom[ 8240]='h00000000;
    rd_cycle[ 8241] = 1'b0;  wr_cycle[ 8241] = 1'b0;  addr_rom[ 8241]='h00000000;  wr_data_rom[ 8241]='h00000000;
    rd_cycle[ 8242] = 1'b0;  wr_cycle[ 8242] = 1'b0;  addr_rom[ 8242]='h00000000;  wr_data_rom[ 8242]='h00000000;
    rd_cycle[ 8243] = 1'b0;  wr_cycle[ 8243] = 1'b0;  addr_rom[ 8243]='h00000000;  wr_data_rom[ 8243]='h00000000;
    rd_cycle[ 8244] = 1'b0;  wr_cycle[ 8244] = 1'b0;  addr_rom[ 8244]='h00000000;  wr_data_rom[ 8244]='h00000000;
    rd_cycle[ 8245] = 1'b0;  wr_cycle[ 8245] = 1'b0;  addr_rom[ 8245]='h00000000;  wr_data_rom[ 8245]='h00000000;
    rd_cycle[ 8246] = 1'b0;  wr_cycle[ 8246] = 1'b0;  addr_rom[ 8246]='h00000000;  wr_data_rom[ 8246]='h00000000;
    rd_cycle[ 8247] = 1'b0;  wr_cycle[ 8247] = 1'b0;  addr_rom[ 8247]='h00000000;  wr_data_rom[ 8247]='h00000000;
    rd_cycle[ 8248] = 1'b0;  wr_cycle[ 8248] = 1'b0;  addr_rom[ 8248]='h00000000;  wr_data_rom[ 8248]='h00000000;
    rd_cycle[ 8249] = 1'b0;  wr_cycle[ 8249] = 1'b0;  addr_rom[ 8249]='h00000000;  wr_data_rom[ 8249]='h00000000;
    rd_cycle[ 8250] = 1'b0;  wr_cycle[ 8250] = 1'b0;  addr_rom[ 8250]='h00000000;  wr_data_rom[ 8250]='h00000000;
    rd_cycle[ 8251] = 1'b0;  wr_cycle[ 8251] = 1'b0;  addr_rom[ 8251]='h00000000;  wr_data_rom[ 8251]='h00000000;
    rd_cycle[ 8252] = 1'b0;  wr_cycle[ 8252] = 1'b0;  addr_rom[ 8252]='h00000000;  wr_data_rom[ 8252]='h00000000;
    rd_cycle[ 8253] = 1'b0;  wr_cycle[ 8253] = 1'b0;  addr_rom[ 8253]='h00000000;  wr_data_rom[ 8253]='h00000000;
    rd_cycle[ 8254] = 1'b0;  wr_cycle[ 8254] = 1'b0;  addr_rom[ 8254]='h00000000;  wr_data_rom[ 8254]='h00000000;
    rd_cycle[ 8255] = 1'b0;  wr_cycle[ 8255] = 1'b0;  addr_rom[ 8255]='h00000000;  wr_data_rom[ 8255]='h00000000;
    rd_cycle[ 8256] = 1'b0;  wr_cycle[ 8256] = 1'b0;  addr_rom[ 8256]='h00000000;  wr_data_rom[ 8256]='h00000000;
    rd_cycle[ 8257] = 1'b0;  wr_cycle[ 8257] = 1'b0;  addr_rom[ 8257]='h00000000;  wr_data_rom[ 8257]='h00000000;
    rd_cycle[ 8258] = 1'b0;  wr_cycle[ 8258] = 1'b0;  addr_rom[ 8258]='h00000000;  wr_data_rom[ 8258]='h00000000;
    rd_cycle[ 8259] = 1'b0;  wr_cycle[ 8259] = 1'b0;  addr_rom[ 8259]='h00000000;  wr_data_rom[ 8259]='h00000000;
    rd_cycle[ 8260] = 1'b0;  wr_cycle[ 8260] = 1'b0;  addr_rom[ 8260]='h00000000;  wr_data_rom[ 8260]='h00000000;
    rd_cycle[ 8261] = 1'b0;  wr_cycle[ 8261] = 1'b0;  addr_rom[ 8261]='h00000000;  wr_data_rom[ 8261]='h00000000;
    rd_cycle[ 8262] = 1'b0;  wr_cycle[ 8262] = 1'b0;  addr_rom[ 8262]='h00000000;  wr_data_rom[ 8262]='h00000000;
    rd_cycle[ 8263] = 1'b0;  wr_cycle[ 8263] = 1'b0;  addr_rom[ 8263]='h00000000;  wr_data_rom[ 8263]='h00000000;
    rd_cycle[ 8264] = 1'b0;  wr_cycle[ 8264] = 1'b0;  addr_rom[ 8264]='h00000000;  wr_data_rom[ 8264]='h00000000;
    rd_cycle[ 8265] = 1'b0;  wr_cycle[ 8265] = 1'b0;  addr_rom[ 8265]='h00000000;  wr_data_rom[ 8265]='h00000000;
    rd_cycle[ 8266] = 1'b0;  wr_cycle[ 8266] = 1'b0;  addr_rom[ 8266]='h00000000;  wr_data_rom[ 8266]='h00000000;
    rd_cycle[ 8267] = 1'b0;  wr_cycle[ 8267] = 1'b0;  addr_rom[ 8267]='h00000000;  wr_data_rom[ 8267]='h00000000;
    rd_cycle[ 8268] = 1'b0;  wr_cycle[ 8268] = 1'b0;  addr_rom[ 8268]='h00000000;  wr_data_rom[ 8268]='h00000000;
    rd_cycle[ 8269] = 1'b0;  wr_cycle[ 8269] = 1'b0;  addr_rom[ 8269]='h00000000;  wr_data_rom[ 8269]='h00000000;
    rd_cycle[ 8270] = 1'b0;  wr_cycle[ 8270] = 1'b0;  addr_rom[ 8270]='h00000000;  wr_data_rom[ 8270]='h00000000;
    rd_cycle[ 8271] = 1'b0;  wr_cycle[ 8271] = 1'b0;  addr_rom[ 8271]='h00000000;  wr_data_rom[ 8271]='h00000000;
    rd_cycle[ 8272] = 1'b0;  wr_cycle[ 8272] = 1'b0;  addr_rom[ 8272]='h00000000;  wr_data_rom[ 8272]='h00000000;
    rd_cycle[ 8273] = 1'b0;  wr_cycle[ 8273] = 1'b0;  addr_rom[ 8273]='h00000000;  wr_data_rom[ 8273]='h00000000;
    rd_cycle[ 8274] = 1'b0;  wr_cycle[ 8274] = 1'b0;  addr_rom[ 8274]='h00000000;  wr_data_rom[ 8274]='h00000000;
    rd_cycle[ 8275] = 1'b0;  wr_cycle[ 8275] = 1'b0;  addr_rom[ 8275]='h00000000;  wr_data_rom[ 8275]='h00000000;
    rd_cycle[ 8276] = 1'b0;  wr_cycle[ 8276] = 1'b0;  addr_rom[ 8276]='h00000000;  wr_data_rom[ 8276]='h00000000;
    rd_cycle[ 8277] = 1'b0;  wr_cycle[ 8277] = 1'b0;  addr_rom[ 8277]='h00000000;  wr_data_rom[ 8277]='h00000000;
    rd_cycle[ 8278] = 1'b0;  wr_cycle[ 8278] = 1'b0;  addr_rom[ 8278]='h00000000;  wr_data_rom[ 8278]='h00000000;
    rd_cycle[ 8279] = 1'b0;  wr_cycle[ 8279] = 1'b0;  addr_rom[ 8279]='h00000000;  wr_data_rom[ 8279]='h00000000;
    rd_cycle[ 8280] = 1'b0;  wr_cycle[ 8280] = 1'b0;  addr_rom[ 8280]='h00000000;  wr_data_rom[ 8280]='h00000000;
    rd_cycle[ 8281] = 1'b0;  wr_cycle[ 8281] = 1'b0;  addr_rom[ 8281]='h00000000;  wr_data_rom[ 8281]='h00000000;
    rd_cycle[ 8282] = 1'b0;  wr_cycle[ 8282] = 1'b0;  addr_rom[ 8282]='h00000000;  wr_data_rom[ 8282]='h00000000;
    rd_cycle[ 8283] = 1'b0;  wr_cycle[ 8283] = 1'b0;  addr_rom[ 8283]='h00000000;  wr_data_rom[ 8283]='h00000000;
    rd_cycle[ 8284] = 1'b0;  wr_cycle[ 8284] = 1'b0;  addr_rom[ 8284]='h00000000;  wr_data_rom[ 8284]='h00000000;
    rd_cycle[ 8285] = 1'b0;  wr_cycle[ 8285] = 1'b0;  addr_rom[ 8285]='h00000000;  wr_data_rom[ 8285]='h00000000;
    rd_cycle[ 8286] = 1'b0;  wr_cycle[ 8286] = 1'b0;  addr_rom[ 8286]='h00000000;  wr_data_rom[ 8286]='h00000000;
    rd_cycle[ 8287] = 1'b0;  wr_cycle[ 8287] = 1'b0;  addr_rom[ 8287]='h00000000;  wr_data_rom[ 8287]='h00000000;
    rd_cycle[ 8288] = 1'b0;  wr_cycle[ 8288] = 1'b0;  addr_rom[ 8288]='h00000000;  wr_data_rom[ 8288]='h00000000;
    rd_cycle[ 8289] = 1'b0;  wr_cycle[ 8289] = 1'b0;  addr_rom[ 8289]='h00000000;  wr_data_rom[ 8289]='h00000000;
    rd_cycle[ 8290] = 1'b0;  wr_cycle[ 8290] = 1'b0;  addr_rom[ 8290]='h00000000;  wr_data_rom[ 8290]='h00000000;
    rd_cycle[ 8291] = 1'b0;  wr_cycle[ 8291] = 1'b0;  addr_rom[ 8291]='h00000000;  wr_data_rom[ 8291]='h00000000;
    rd_cycle[ 8292] = 1'b0;  wr_cycle[ 8292] = 1'b0;  addr_rom[ 8292]='h00000000;  wr_data_rom[ 8292]='h00000000;
    rd_cycle[ 8293] = 1'b0;  wr_cycle[ 8293] = 1'b0;  addr_rom[ 8293]='h00000000;  wr_data_rom[ 8293]='h00000000;
    rd_cycle[ 8294] = 1'b0;  wr_cycle[ 8294] = 1'b0;  addr_rom[ 8294]='h00000000;  wr_data_rom[ 8294]='h00000000;
    rd_cycle[ 8295] = 1'b0;  wr_cycle[ 8295] = 1'b0;  addr_rom[ 8295]='h00000000;  wr_data_rom[ 8295]='h00000000;
    rd_cycle[ 8296] = 1'b0;  wr_cycle[ 8296] = 1'b0;  addr_rom[ 8296]='h00000000;  wr_data_rom[ 8296]='h00000000;
    rd_cycle[ 8297] = 1'b0;  wr_cycle[ 8297] = 1'b0;  addr_rom[ 8297]='h00000000;  wr_data_rom[ 8297]='h00000000;
    rd_cycle[ 8298] = 1'b0;  wr_cycle[ 8298] = 1'b0;  addr_rom[ 8298]='h00000000;  wr_data_rom[ 8298]='h00000000;
    rd_cycle[ 8299] = 1'b0;  wr_cycle[ 8299] = 1'b0;  addr_rom[ 8299]='h00000000;  wr_data_rom[ 8299]='h00000000;
    rd_cycle[ 8300] = 1'b0;  wr_cycle[ 8300] = 1'b0;  addr_rom[ 8300]='h00000000;  wr_data_rom[ 8300]='h00000000;
    rd_cycle[ 8301] = 1'b0;  wr_cycle[ 8301] = 1'b0;  addr_rom[ 8301]='h00000000;  wr_data_rom[ 8301]='h00000000;
    rd_cycle[ 8302] = 1'b0;  wr_cycle[ 8302] = 1'b0;  addr_rom[ 8302]='h00000000;  wr_data_rom[ 8302]='h00000000;
    rd_cycle[ 8303] = 1'b0;  wr_cycle[ 8303] = 1'b0;  addr_rom[ 8303]='h00000000;  wr_data_rom[ 8303]='h00000000;
    rd_cycle[ 8304] = 1'b0;  wr_cycle[ 8304] = 1'b0;  addr_rom[ 8304]='h00000000;  wr_data_rom[ 8304]='h00000000;
    rd_cycle[ 8305] = 1'b0;  wr_cycle[ 8305] = 1'b0;  addr_rom[ 8305]='h00000000;  wr_data_rom[ 8305]='h00000000;
    rd_cycle[ 8306] = 1'b0;  wr_cycle[ 8306] = 1'b0;  addr_rom[ 8306]='h00000000;  wr_data_rom[ 8306]='h00000000;
    rd_cycle[ 8307] = 1'b0;  wr_cycle[ 8307] = 1'b0;  addr_rom[ 8307]='h00000000;  wr_data_rom[ 8307]='h00000000;
    rd_cycle[ 8308] = 1'b0;  wr_cycle[ 8308] = 1'b0;  addr_rom[ 8308]='h00000000;  wr_data_rom[ 8308]='h00000000;
    rd_cycle[ 8309] = 1'b0;  wr_cycle[ 8309] = 1'b0;  addr_rom[ 8309]='h00000000;  wr_data_rom[ 8309]='h00000000;
    rd_cycle[ 8310] = 1'b0;  wr_cycle[ 8310] = 1'b0;  addr_rom[ 8310]='h00000000;  wr_data_rom[ 8310]='h00000000;
    rd_cycle[ 8311] = 1'b0;  wr_cycle[ 8311] = 1'b0;  addr_rom[ 8311]='h00000000;  wr_data_rom[ 8311]='h00000000;
    rd_cycle[ 8312] = 1'b0;  wr_cycle[ 8312] = 1'b0;  addr_rom[ 8312]='h00000000;  wr_data_rom[ 8312]='h00000000;
    rd_cycle[ 8313] = 1'b0;  wr_cycle[ 8313] = 1'b0;  addr_rom[ 8313]='h00000000;  wr_data_rom[ 8313]='h00000000;
    rd_cycle[ 8314] = 1'b0;  wr_cycle[ 8314] = 1'b0;  addr_rom[ 8314]='h00000000;  wr_data_rom[ 8314]='h00000000;
    rd_cycle[ 8315] = 1'b0;  wr_cycle[ 8315] = 1'b0;  addr_rom[ 8315]='h00000000;  wr_data_rom[ 8315]='h00000000;
    rd_cycle[ 8316] = 1'b0;  wr_cycle[ 8316] = 1'b0;  addr_rom[ 8316]='h00000000;  wr_data_rom[ 8316]='h00000000;
    rd_cycle[ 8317] = 1'b0;  wr_cycle[ 8317] = 1'b0;  addr_rom[ 8317]='h00000000;  wr_data_rom[ 8317]='h00000000;
    rd_cycle[ 8318] = 1'b0;  wr_cycle[ 8318] = 1'b0;  addr_rom[ 8318]='h00000000;  wr_data_rom[ 8318]='h00000000;
    rd_cycle[ 8319] = 1'b0;  wr_cycle[ 8319] = 1'b0;  addr_rom[ 8319]='h00000000;  wr_data_rom[ 8319]='h00000000;
    rd_cycle[ 8320] = 1'b0;  wr_cycle[ 8320] = 1'b0;  addr_rom[ 8320]='h00000000;  wr_data_rom[ 8320]='h00000000;
    rd_cycle[ 8321] = 1'b0;  wr_cycle[ 8321] = 1'b0;  addr_rom[ 8321]='h00000000;  wr_data_rom[ 8321]='h00000000;
    rd_cycle[ 8322] = 1'b0;  wr_cycle[ 8322] = 1'b0;  addr_rom[ 8322]='h00000000;  wr_data_rom[ 8322]='h00000000;
    rd_cycle[ 8323] = 1'b0;  wr_cycle[ 8323] = 1'b0;  addr_rom[ 8323]='h00000000;  wr_data_rom[ 8323]='h00000000;
    rd_cycle[ 8324] = 1'b0;  wr_cycle[ 8324] = 1'b0;  addr_rom[ 8324]='h00000000;  wr_data_rom[ 8324]='h00000000;
    rd_cycle[ 8325] = 1'b0;  wr_cycle[ 8325] = 1'b0;  addr_rom[ 8325]='h00000000;  wr_data_rom[ 8325]='h00000000;
    rd_cycle[ 8326] = 1'b0;  wr_cycle[ 8326] = 1'b0;  addr_rom[ 8326]='h00000000;  wr_data_rom[ 8326]='h00000000;
    rd_cycle[ 8327] = 1'b0;  wr_cycle[ 8327] = 1'b0;  addr_rom[ 8327]='h00000000;  wr_data_rom[ 8327]='h00000000;
    rd_cycle[ 8328] = 1'b0;  wr_cycle[ 8328] = 1'b0;  addr_rom[ 8328]='h00000000;  wr_data_rom[ 8328]='h00000000;
    rd_cycle[ 8329] = 1'b0;  wr_cycle[ 8329] = 1'b0;  addr_rom[ 8329]='h00000000;  wr_data_rom[ 8329]='h00000000;
    rd_cycle[ 8330] = 1'b0;  wr_cycle[ 8330] = 1'b0;  addr_rom[ 8330]='h00000000;  wr_data_rom[ 8330]='h00000000;
    rd_cycle[ 8331] = 1'b0;  wr_cycle[ 8331] = 1'b0;  addr_rom[ 8331]='h00000000;  wr_data_rom[ 8331]='h00000000;
    rd_cycle[ 8332] = 1'b0;  wr_cycle[ 8332] = 1'b0;  addr_rom[ 8332]='h00000000;  wr_data_rom[ 8332]='h00000000;
    rd_cycle[ 8333] = 1'b0;  wr_cycle[ 8333] = 1'b0;  addr_rom[ 8333]='h00000000;  wr_data_rom[ 8333]='h00000000;
    rd_cycle[ 8334] = 1'b0;  wr_cycle[ 8334] = 1'b0;  addr_rom[ 8334]='h00000000;  wr_data_rom[ 8334]='h00000000;
    rd_cycle[ 8335] = 1'b0;  wr_cycle[ 8335] = 1'b0;  addr_rom[ 8335]='h00000000;  wr_data_rom[ 8335]='h00000000;
    rd_cycle[ 8336] = 1'b0;  wr_cycle[ 8336] = 1'b0;  addr_rom[ 8336]='h00000000;  wr_data_rom[ 8336]='h00000000;
    rd_cycle[ 8337] = 1'b0;  wr_cycle[ 8337] = 1'b0;  addr_rom[ 8337]='h00000000;  wr_data_rom[ 8337]='h00000000;
    rd_cycle[ 8338] = 1'b0;  wr_cycle[ 8338] = 1'b0;  addr_rom[ 8338]='h00000000;  wr_data_rom[ 8338]='h00000000;
    rd_cycle[ 8339] = 1'b0;  wr_cycle[ 8339] = 1'b0;  addr_rom[ 8339]='h00000000;  wr_data_rom[ 8339]='h00000000;
    rd_cycle[ 8340] = 1'b0;  wr_cycle[ 8340] = 1'b0;  addr_rom[ 8340]='h00000000;  wr_data_rom[ 8340]='h00000000;
    rd_cycle[ 8341] = 1'b0;  wr_cycle[ 8341] = 1'b0;  addr_rom[ 8341]='h00000000;  wr_data_rom[ 8341]='h00000000;
    rd_cycle[ 8342] = 1'b0;  wr_cycle[ 8342] = 1'b0;  addr_rom[ 8342]='h00000000;  wr_data_rom[ 8342]='h00000000;
    rd_cycle[ 8343] = 1'b0;  wr_cycle[ 8343] = 1'b0;  addr_rom[ 8343]='h00000000;  wr_data_rom[ 8343]='h00000000;
    rd_cycle[ 8344] = 1'b0;  wr_cycle[ 8344] = 1'b0;  addr_rom[ 8344]='h00000000;  wr_data_rom[ 8344]='h00000000;
    rd_cycle[ 8345] = 1'b0;  wr_cycle[ 8345] = 1'b0;  addr_rom[ 8345]='h00000000;  wr_data_rom[ 8345]='h00000000;
    rd_cycle[ 8346] = 1'b0;  wr_cycle[ 8346] = 1'b0;  addr_rom[ 8346]='h00000000;  wr_data_rom[ 8346]='h00000000;
    rd_cycle[ 8347] = 1'b0;  wr_cycle[ 8347] = 1'b0;  addr_rom[ 8347]='h00000000;  wr_data_rom[ 8347]='h00000000;
    rd_cycle[ 8348] = 1'b0;  wr_cycle[ 8348] = 1'b0;  addr_rom[ 8348]='h00000000;  wr_data_rom[ 8348]='h00000000;
    rd_cycle[ 8349] = 1'b0;  wr_cycle[ 8349] = 1'b0;  addr_rom[ 8349]='h00000000;  wr_data_rom[ 8349]='h00000000;
    rd_cycle[ 8350] = 1'b0;  wr_cycle[ 8350] = 1'b0;  addr_rom[ 8350]='h00000000;  wr_data_rom[ 8350]='h00000000;
    rd_cycle[ 8351] = 1'b0;  wr_cycle[ 8351] = 1'b0;  addr_rom[ 8351]='h00000000;  wr_data_rom[ 8351]='h00000000;
    rd_cycle[ 8352] = 1'b0;  wr_cycle[ 8352] = 1'b0;  addr_rom[ 8352]='h00000000;  wr_data_rom[ 8352]='h00000000;
    rd_cycle[ 8353] = 1'b0;  wr_cycle[ 8353] = 1'b0;  addr_rom[ 8353]='h00000000;  wr_data_rom[ 8353]='h00000000;
    rd_cycle[ 8354] = 1'b0;  wr_cycle[ 8354] = 1'b0;  addr_rom[ 8354]='h00000000;  wr_data_rom[ 8354]='h00000000;
    rd_cycle[ 8355] = 1'b0;  wr_cycle[ 8355] = 1'b0;  addr_rom[ 8355]='h00000000;  wr_data_rom[ 8355]='h00000000;
    rd_cycle[ 8356] = 1'b0;  wr_cycle[ 8356] = 1'b0;  addr_rom[ 8356]='h00000000;  wr_data_rom[ 8356]='h00000000;
    rd_cycle[ 8357] = 1'b0;  wr_cycle[ 8357] = 1'b0;  addr_rom[ 8357]='h00000000;  wr_data_rom[ 8357]='h00000000;
    rd_cycle[ 8358] = 1'b0;  wr_cycle[ 8358] = 1'b0;  addr_rom[ 8358]='h00000000;  wr_data_rom[ 8358]='h00000000;
    rd_cycle[ 8359] = 1'b0;  wr_cycle[ 8359] = 1'b0;  addr_rom[ 8359]='h00000000;  wr_data_rom[ 8359]='h00000000;
    rd_cycle[ 8360] = 1'b0;  wr_cycle[ 8360] = 1'b0;  addr_rom[ 8360]='h00000000;  wr_data_rom[ 8360]='h00000000;
    rd_cycle[ 8361] = 1'b0;  wr_cycle[ 8361] = 1'b0;  addr_rom[ 8361]='h00000000;  wr_data_rom[ 8361]='h00000000;
    rd_cycle[ 8362] = 1'b0;  wr_cycle[ 8362] = 1'b0;  addr_rom[ 8362]='h00000000;  wr_data_rom[ 8362]='h00000000;
    rd_cycle[ 8363] = 1'b0;  wr_cycle[ 8363] = 1'b0;  addr_rom[ 8363]='h00000000;  wr_data_rom[ 8363]='h00000000;
    rd_cycle[ 8364] = 1'b0;  wr_cycle[ 8364] = 1'b0;  addr_rom[ 8364]='h00000000;  wr_data_rom[ 8364]='h00000000;
    rd_cycle[ 8365] = 1'b0;  wr_cycle[ 8365] = 1'b0;  addr_rom[ 8365]='h00000000;  wr_data_rom[ 8365]='h00000000;
    rd_cycle[ 8366] = 1'b0;  wr_cycle[ 8366] = 1'b0;  addr_rom[ 8366]='h00000000;  wr_data_rom[ 8366]='h00000000;
    rd_cycle[ 8367] = 1'b0;  wr_cycle[ 8367] = 1'b0;  addr_rom[ 8367]='h00000000;  wr_data_rom[ 8367]='h00000000;
    rd_cycle[ 8368] = 1'b0;  wr_cycle[ 8368] = 1'b0;  addr_rom[ 8368]='h00000000;  wr_data_rom[ 8368]='h00000000;
    rd_cycle[ 8369] = 1'b0;  wr_cycle[ 8369] = 1'b0;  addr_rom[ 8369]='h00000000;  wr_data_rom[ 8369]='h00000000;
    rd_cycle[ 8370] = 1'b0;  wr_cycle[ 8370] = 1'b0;  addr_rom[ 8370]='h00000000;  wr_data_rom[ 8370]='h00000000;
    rd_cycle[ 8371] = 1'b0;  wr_cycle[ 8371] = 1'b0;  addr_rom[ 8371]='h00000000;  wr_data_rom[ 8371]='h00000000;
    rd_cycle[ 8372] = 1'b0;  wr_cycle[ 8372] = 1'b0;  addr_rom[ 8372]='h00000000;  wr_data_rom[ 8372]='h00000000;
    rd_cycle[ 8373] = 1'b0;  wr_cycle[ 8373] = 1'b0;  addr_rom[ 8373]='h00000000;  wr_data_rom[ 8373]='h00000000;
    rd_cycle[ 8374] = 1'b0;  wr_cycle[ 8374] = 1'b0;  addr_rom[ 8374]='h00000000;  wr_data_rom[ 8374]='h00000000;
    rd_cycle[ 8375] = 1'b0;  wr_cycle[ 8375] = 1'b0;  addr_rom[ 8375]='h00000000;  wr_data_rom[ 8375]='h00000000;
    rd_cycle[ 8376] = 1'b0;  wr_cycle[ 8376] = 1'b0;  addr_rom[ 8376]='h00000000;  wr_data_rom[ 8376]='h00000000;
    rd_cycle[ 8377] = 1'b0;  wr_cycle[ 8377] = 1'b0;  addr_rom[ 8377]='h00000000;  wr_data_rom[ 8377]='h00000000;
    rd_cycle[ 8378] = 1'b0;  wr_cycle[ 8378] = 1'b0;  addr_rom[ 8378]='h00000000;  wr_data_rom[ 8378]='h00000000;
    rd_cycle[ 8379] = 1'b0;  wr_cycle[ 8379] = 1'b0;  addr_rom[ 8379]='h00000000;  wr_data_rom[ 8379]='h00000000;
    rd_cycle[ 8380] = 1'b0;  wr_cycle[ 8380] = 1'b0;  addr_rom[ 8380]='h00000000;  wr_data_rom[ 8380]='h00000000;
    rd_cycle[ 8381] = 1'b0;  wr_cycle[ 8381] = 1'b0;  addr_rom[ 8381]='h00000000;  wr_data_rom[ 8381]='h00000000;
    rd_cycle[ 8382] = 1'b0;  wr_cycle[ 8382] = 1'b0;  addr_rom[ 8382]='h00000000;  wr_data_rom[ 8382]='h00000000;
    rd_cycle[ 8383] = 1'b0;  wr_cycle[ 8383] = 1'b0;  addr_rom[ 8383]='h00000000;  wr_data_rom[ 8383]='h00000000;
    rd_cycle[ 8384] = 1'b0;  wr_cycle[ 8384] = 1'b0;  addr_rom[ 8384]='h00000000;  wr_data_rom[ 8384]='h00000000;
    rd_cycle[ 8385] = 1'b0;  wr_cycle[ 8385] = 1'b0;  addr_rom[ 8385]='h00000000;  wr_data_rom[ 8385]='h00000000;
    rd_cycle[ 8386] = 1'b0;  wr_cycle[ 8386] = 1'b0;  addr_rom[ 8386]='h00000000;  wr_data_rom[ 8386]='h00000000;
    rd_cycle[ 8387] = 1'b0;  wr_cycle[ 8387] = 1'b0;  addr_rom[ 8387]='h00000000;  wr_data_rom[ 8387]='h00000000;
    rd_cycle[ 8388] = 1'b0;  wr_cycle[ 8388] = 1'b0;  addr_rom[ 8388]='h00000000;  wr_data_rom[ 8388]='h00000000;
    rd_cycle[ 8389] = 1'b0;  wr_cycle[ 8389] = 1'b0;  addr_rom[ 8389]='h00000000;  wr_data_rom[ 8389]='h00000000;
    rd_cycle[ 8390] = 1'b0;  wr_cycle[ 8390] = 1'b0;  addr_rom[ 8390]='h00000000;  wr_data_rom[ 8390]='h00000000;
    rd_cycle[ 8391] = 1'b0;  wr_cycle[ 8391] = 1'b0;  addr_rom[ 8391]='h00000000;  wr_data_rom[ 8391]='h00000000;
    rd_cycle[ 8392] = 1'b0;  wr_cycle[ 8392] = 1'b0;  addr_rom[ 8392]='h00000000;  wr_data_rom[ 8392]='h00000000;
    rd_cycle[ 8393] = 1'b0;  wr_cycle[ 8393] = 1'b0;  addr_rom[ 8393]='h00000000;  wr_data_rom[ 8393]='h00000000;
    rd_cycle[ 8394] = 1'b0;  wr_cycle[ 8394] = 1'b0;  addr_rom[ 8394]='h00000000;  wr_data_rom[ 8394]='h00000000;
    rd_cycle[ 8395] = 1'b0;  wr_cycle[ 8395] = 1'b0;  addr_rom[ 8395]='h00000000;  wr_data_rom[ 8395]='h00000000;
    rd_cycle[ 8396] = 1'b0;  wr_cycle[ 8396] = 1'b0;  addr_rom[ 8396]='h00000000;  wr_data_rom[ 8396]='h00000000;
    rd_cycle[ 8397] = 1'b0;  wr_cycle[ 8397] = 1'b0;  addr_rom[ 8397]='h00000000;  wr_data_rom[ 8397]='h00000000;
    rd_cycle[ 8398] = 1'b0;  wr_cycle[ 8398] = 1'b0;  addr_rom[ 8398]='h00000000;  wr_data_rom[ 8398]='h00000000;
    rd_cycle[ 8399] = 1'b0;  wr_cycle[ 8399] = 1'b0;  addr_rom[ 8399]='h00000000;  wr_data_rom[ 8399]='h00000000;
    rd_cycle[ 8400] = 1'b0;  wr_cycle[ 8400] = 1'b0;  addr_rom[ 8400]='h00000000;  wr_data_rom[ 8400]='h00000000;
    rd_cycle[ 8401] = 1'b0;  wr_cycle[ 8401] = 1'b0;  addr_rom[ 8401]='h00000000;  wr_data_rom[ 8401]='h00000000;
    rd_cycle[ 8402] = 1'b0;  wr_cycle[ 8402] = 1'b0;  addr_rom[ 8402]='h00000000;  wr_data_rom[ 8402]='h00000000;
    rd_cycle[ 8403] = 1'b0;  wr_cycle[ 8403] = 1'b0;  addr_rom[ 8403]='h00000000;  wr_data_rom[ 8403]='h00000000;
    rd_cycle[ 8404] = 1'b0;  wr_cycle[ 8404] = 1'b0;  addr_rom[ 8404]='h00000000;  wr_data_rom[ 8404]='h00000000;
    rd_cycle[ 8405] = 1'b0;  wr_cycle[ 8405] = 1'b0;  addr_rom[ 8405]='h00000000;  wr_data_rom[ 8405]='h00000000;
    rd_cycle[ 8406] = 1'b0;  wr_cycle[ 8406] = 1'b0;  addr_rom[ 8406]='h00000000;  wr_data_rom[ 8406]='h00000000;
    rd_cycle[ 8407] = 1'b0;  wr_cycle[ 8407] = 1'b0;  addr_rom[ 8407]='h00000000;  wr_data_rom[ 8407]='h00000000;
    rd_cycle[ 8408] = 1'b0;  wr_cycle[ 8408] = 1'b0;  addr_rom[ 8408]='h00000000;  wr_data_rom[ 8408]='h00000000;
    rd_cycle[ 8409] = 1'b0;  wr_cycle[ 8409] = 1'b0;  addr_rom[ 8409]='h00000000;  wr_data_rom[ 8409]='h00000000;
    rd_cycle[ 8410] = 1'b0;  wr_cycle[ 8410] = 1'b0;  addr_rom[ 8410]='h00000000;  wr_data_rom[ 8410]='h00000000;
    rd_cycle[ 8411] = 1'b0;  wr_cycle[ 8411] = 1'b0;  addr_rom[ 8411]='h00000000;  wr_data_rom[ 8411]='h00000000;
    rd_cycle[ 8412] = 1'b0;  wr_cycle[ 8412] = 1'b0;  addr_rom[ 8412]='h00000000;  wr_data_rom[ 8412]='h00000000;
    rd_cycle[ 8413] = 1'b0;  wr_cycle[ 8413] = 1'b0;  addr_rom[ 8413]='h00000000;  wr_data_rom[ 8413]='h00000000;
    rd_cycle[ 8414] = 1'b0;  wr_cycle[ 8414] = 1'b0;  addr_rom[ 8414]='h00000000;  wr_data_rom[ 8414]='h00000000;
    rd_cycle[ 8415] = 1'b0;  wr_cycle[ 8415] = 1'b0;  addr_rom[ 8415]='h00000000;  wr_data_rom[ 8415]='h00000000;
    rd_cycle[ 8416] = 1'b0;  wr_cycle[ 8416] = 1'b0;  addr_rom[ 8416]='h00000000;  wr_data_rom[ 8416]='h00000000;
    rd_cycle[ 8417] = 1'b0;  wr_cycle[ 8417] = 1'b0;  addr_rom[ 8417]='h00000000;  wr_data_rom[ 8417]='h00000000;
    rd_cycle[ 8418] = 1'b0;  wr_cycle[ 8418] = 1'b0;  addr_rom[ 8418]='h00000000;  wr_data_rom[ 8418]='h00000000;
    rd_cycle[ 8419] = 1'b0;  wr_cycle[ 8419] = 1'b0;  addr_rom[ 8419]='h00000000;  wr_data_rom[ 8419]='h00000000;
    rd_cycle[ 8420] = 1'b0;  wr_cycle[ 8420] = 1'b0;  addr_rom[ 8420]='h00000000;  wr_data_rom[ 8420]='h00000000;
    rd_cycle[ 8421] = 1'b0;  wr_cycle[ 8421] = 1'b0;  addr_rom[ 8421]='h00000000;  wr_data_rom[ 8421]='h00000000;
    rd_cycle[ 8422] = 1'b0;  wr_cycle[ 8422] = 1'b0;  addr_rom[ 8422]='h00000000;  wr_data_rom[ 8422]='h00000000;
    rd_cycle[ 8423] = 1'b0;  wr_cycle[ 8423] = 1'b0;  addr_rom[ 8423]='h00000000;  wr_data_rom[ 8423]='h00000000;
    rd_cycle[ 8424] = 1'b0;  wr_cycle[ 8424] = 1'b0;  addr_rom[ 8424]='h00000000;  wr_data_rom[ 8424]='h00000000;
    rd_cycle[ 8425] = 1'b0;  wr_cycle[ 8425] = 1'b0;  addr_rom[ 8425]='h00000000;  wr_data_rom[ 8425]='h00000000;
    rd_cycle[ 8426] = 1'b0;  wr_cycle[ 8426] = 1'b0;  addr_rom[ 8426]='h00000000;  wr_data_rom[ 8426]='h00000000;
    rd_cycle[ 8427] = 1'b0;  wr_cycle[ 8427] = 1'b0;  addr_rom[ 8427]='h00000000;  wr_data_rom[ 8427]='h00000000;
    rd_cycle[ 8428] = 1'b0;  wr_cycle[ 8428] = 1'b0;  addr_rom[ 8428]='h00000000;  wr_data_rom[ 8428]='h00000000;
    rd_cycle[ 8429] = 1'b0;  wr_cycle[ 8429] = 1'b0;  addr_rom[ 8429]='h00000000;  wr_data_rom[ 8429]='h00000000;
    rd_cycle[ 8430] = 1'b0;  wr_cycle[ 8430] = 1'b0;  addr_rom[ 8430]='h00000000;  wr_data_rom[ 8430]='h00000000;
    rd_cycle[ 8431] = 1'b0;  wr_cycle[ 8431] = 1'b0;  addr_rom[ 8431]='h00000000;  wr_data_rom[ 8431]='h00000000;
    rd_cycle[ 8432] = 1'b0;  wr_cycle[ 8432] = 1'b0;  addr_rom[ 8432]='h00000000;  wr_data_rom[ 8432]='h00000000;
    rd_cycle[ 8433] = 1'b0;  wr_cycle[ 8433] = 1'b0;  addr_rom[ 8433]='h00000000;  wr_data_rom[ 8433]='h00000000;
    rd_cycle[ 8434] = 1'b0;  wr_cycle[ 8434] = 1'b0;  addr_rom[ 8434]='h00000000;  wr_data_rom[ 8434]='h00000000;
    rd_cycle[ 8435] = 1'b0;  wr_cycle[ 8435] = 1'b0;  addr_rom[ 8435]='h00000000;  wr_data_rom[ 8435]='h00000000;
    rd_cycle[ 8436] = 1'b0;  wr_cycle[ 8436] = 1'b0;  addr_rom[ 8436]='h00000000;  wr_data_rom[ 8436]='h00000000;
    rd_cycle[ 8437] = 1'b0;  wr_cycle[ 8437] = 1'b0;  addr_rom[ 8437]='h00000000;  wr_data_rom[ 8437]='h00000000;
    rd_cycle[ 8438] = 1'b0;  wr_cycle[ 8438] = 1'b0;  addr_rom[ 8438]='h00000000;  wr_data_rom[ 8438]='h00000000;
    rd_cycle[ 8439] = 1'b0;  wr_cycle[ 8439] = 1'b0;  addr_rom[ 8439]='h00000000;  wr_data_rom[ 8439]='h00000000;
    rd_cycle[ 8440] = 1'b0;  wr_cycle[ 8440] = 1'b0;  addr_rom[ 8440]='h00000000;  wr_data_rom[ 8440]='h00000000;
    rd_cycle[ 8441] = 1'b0;  wr_cycle[ 8441] = 1'b0;  addr_rom[ 8441]='h00000000;  wr_data_rom[ 8441]='h00000000;
    rd_cycle[ 8442] = 1'b0;  wr_cycle[ 8442] = 1'b0;  addr_rom[ 8442]='h00000000;  wr_data_rom[ 8442]='h00000000;
    rd_cycle[ 8443] = 1'b0;  wr_cycle[ 8443] = 1'b0;  addr_rom[ 8443]='h00000000;  wr_data_rom[ 8443]='h00000000;
    rd_cycle[ 8444] = 1'b0;  wr_cycle[ 8444] = 1'b0;  addr_rom[ 8444]='h00000000;  wr_data_rom[ 8444]='h00000000;
    rd_cycle[ 8445] = 1'b0;  wr_cycle[ 8445] = 1'b0;  addr_rom[ 8445]='h00000000;  wr_data_rom[ 8445]='h00000000;
    rd_cycle[ 8446] = 1'b0;  wr_cycle[ 8446] = 1'b0;  addr_rom[ 8446]='h00000000;  wr_data_rom[ 8446]='h00000000;
    rd_cycle[ 8447] = 1'b0;  wr_cycle[ 8447] = 1'b0;  addr_rom[ 8447]='h00000000;  wr_data_rom[ 8447]='h00000000;
    rd_cycle[ 8448] = 1'b0;  wr_cycle[ 8448] = 1'b0;  addr_rom[ 8448]='h00000000;  wr_data_rom[ 8448]='h00000000;
    rd_cycle[ 8449] = 1'b0;  wr_cycle[ 8449] = 1'b0;  addr_rom[ 8449]='h00000000;  wr_data_rom[ 8449]='h00000000;
    rd_cycle[ 8450] = 1'b0;  wr_cycle[ 8450] = 1'b0;  addr_rom[ 8450]='h00000000;  wr_data_rom[ 8450]='h00000000;
    rd_cycle[ 8451] = 1'b0;  wr_cycle[ 8451] = 1'b0;  addr_rom[ 8451]='h00000000;  wr_data_rom[ 8451]='h00000000;
    rd_cycle[ 8452] = 1'b0;  wr_cycle[ 8452] = 1'b0;  addr_rom[ 8452]='h00000000;  wr_data_rom[ 8452]='h00000000;
    rd_cycle[ 8453] = 1'b0;  wr_cycle[ 8453] = 1'b0;  addr_rom[ 8453]='h00000000;  wr_data_rom[ 8453]='h00000000;
    rd_cycle[ 8454] = 1'b0;  wr_cycle[ 8454] = 1'b0;  addr_rom[ 8454]='h00000000;  wr_data_rom[ 8454]='h00000000;
    rd_cycle[ 8455] = 1'b0;  wr_cycle[ 8455] = 1'b0;  addr_rom[ 8455]='h00000000;  wr_data_rom[ 8455]='h00000000;
    rd_cycle[ 8456] = 1'b0;  wr_cycle[ 8456] = 1'b0;  addr_rom[ 8456]='h00000000;  wr_data_rom[ 8456]='h00000000;
    rd_cycle[ 8457] = 1'b0;  wr_cycle[ 8457] = 1'b0;  addr_rom[ 8457]='h00000000;  wr_data_rom[ 8457]='h00000000;
    rd_cycle[ 8458] = 1'b0;  wr_cycle[ 8458] = 1'b0;  addr_rom[ 8458]='h00000000;  wr_data_rom[ 8458]='h00000000;
    rd_cycle[ 8459] = 1'b0;  wr_cycle[ 8459] = 1'b0;  addr_rom[ 8459]='h00000000;  wr_data_rom[ 8459]='h00000000;
    rd_cycle[ 8460] = 1'b0;  wr_cycle[ 8460] = 1'b0;  addr_rom[ 8460]='h00000000;  wr_data_rom[ 8460]='h00000000;
    rd_cycle[ 8461] = 1'b0;  wr_cycle[ 8461] = 1'b0;  addr_rom[ 8461]='h00000000;  wr_data_rom[ 8461]='h00000000;
    rd_cycle[ 8462] = 1'b0;  wr_cycle[ 8462] = 1'b0;  addr_rom[ 8462]='h00000000;  wr_data_rom[ 8462]='h00000000;
    rd_cycle[ 8463] = 1'b0;  wr_cycle[ 8463] = 1'b0;  addr_rom[ 8463]='h00000000;  wr_data_rom[ 8463]='h00000000;
    rd_cycle[ 8464] = 1'b0;  wr_cycle[ 8464] = 1'b0;  addr_rom[ 8464]='h00000000;  wr_data_rom[ 8464]='h00000000;
    rd_cycle[ 8465] = 1'b0;  wr_cycle[ 8465] = 1'b0;  addr_rom[ 8465]='h00000000;  wr_data_rom[ 8465]='h00000000;
    rd_cycle[ 8466] = 1'b0;  wr_cycle[ 8466] = 1'b0;  addr_rom[ 8466]='h00000000;  wr_data_rom[ 8466]='h00000000;
    rd_cycle[ 8467] = 1'b0;  wr_cycle[ 8467] = 1'b0;  addr_rom[ 8467]='h00000000;  wr_data_rom[ 8467]='h00000000;
    rd_cycle[ 8468] = 1'b0;  wr_cycle[ 8468] = 1'b0;  addr_rom[ 8468]='h00000000;  wr_data_rom[ 8468]='h00000000;
    rd_cycle[ 8469] = 1'b0;  wr_cycle[ 8469] = 1'b0;  addr_rom[ 8469]='h00000000;  wr_data_rom[ 8469]='h00000000;
    rd_cycle[ 8470] = 1'b0;  wr_cycle[ 8470] = 1'b0;  addr_rom[ 8470]='h00000000;  wr_data_rom[ 8470]='h00000000;
    rd_cycle[ 8471] = 1'b0;  wr_cycle[ 8471] = 1'b0;  addr_rom[ 8471]='h00000000;  wr_data_rom[ 8471]='h00000000;
    rd_cycle[ 8472] = 1'b0;  wr_cycle[ 8472] = 1'b0;  addr_rom[ 8472]='h00000000;  wr_data_rom[ 8472]='h00000000;
    rd_cycle[ 8473] = 1'b0;  wr_cycle[ 8473] = 1'b0;  addr_rom[ 8473]='h00000000;  wr_data_rom[ 8473]='h00000000;
    rd_cycle[ 8474] = 1'b0;  wr_cycle[ 8474] = 1'b0;  addr_rom[ 8474]='h00000000;  wr_data_rom[ 8474]='h00000000;
    rd_cycle[ 8475] = 1'b0;  wr_cycle[ 8475] = 1'b0;  addr_rom[ 8475]='h00000000;  wr_data_rom[ 8475]='h00000000;
    rd_cycle[ 8476] = 1'b0;  wr_cycle[ 8476] = 1'b0;  addr_rom[ 8476]='h00000000;  wr_data_rom[ 8476]='h00000000;
    rd_cycle[ 8477] = 1'b0;  wr_cycle[ 8477] = 1'b0;  addr_rom[ 8477]='h00000000;  wr_data_rom[ 8477]='h00000000;
    rd_cycle[ 8478] = 1'b0;  wr_cycle[ 8478] = 1'b0;  addr_rom[ 8478]='h00000000;  wr_data_rom[ 8478]='h00000000;
    rd_cycle[ 8479] = 1'b0;  wr_cycle[ 8479] = 1'b0;  addr_rom[ 8479]='h00000000;  wr_data_rom[ 8479]='h00000000;
    rd_cycle[ 8480] = 1'b0;  wr_cycle[ 8480] = 1'b0;  addr_rom[ 8480]='h00000000;  wr_data_rom[ 8480]='h00000000;
    rd_cycle[ 8481] = 1'b0;  wr_cycle[ 8481] = 1'b0;  addr_rom[ 8481]='h00000000;  wr_data_rom[ 8481]='h00000000;
    rd_cycle[ 8482] = 1'b0;  wr_cycle[ 8482] = 1'b0;  addr_rom[ 8482]='h00000000;  wr_data_rom[ 8482]='h00000000;
    rd_cycle[ 8483] = 1'b0;  wr_cycle[ 8483] = 1'b0;  addr_rom[ 8483]='h00000000;  wr_data_rom[ 8483]='h00000000;
    rd_cycle[ 8484] = 1'b0;  wr_cycle[ 8484] = 1'b0;  addr_rom[ 8484]='h00000000;  wr_data_rom[ 8484]='h00000000;
    rd_cycle[ 8485] = 1'b0;  wr_cycle[ 8485] = 1'b0;  addr_rom[ 8485]='h00000000;  wr_data_rom[ 8485]='h00000000;
    rd_cycle[ 8486] = 1'b0;  wr_cycle[ 8486] = 1'b0;  addr_rom[ 8486]='h00000000;  wr_data_rom[ 8486]='h00000000;
    rd_cycle[ 8487] = 1'b0;  wr_cycle[ 8487] = 1'b0;  addr_rom[ 8487]='h00000000;  wr_data_rom[ 8487]='h00000000;
    rd_cycle[ 8488] = 1'b0;  wr_cycle[ 8488] = 1'b0;  addr_rom[ 8488]='h00000000;  wr_data_rom[ 8488]='h00000000;
    rd_cycle[ 8489] = 1'b0;  wr_cycle[ 8489] = 1'b0;  addr_rom[ 8489]='h00000000;  wr_data_rom[ 8489]='h00000000;
    rd_cycle[ 8490] = 1'b0;  wr_cycle[ 8490] = 1'b0;  addr_rom[ 8490]='h00000000;  wr_data_rom[ 8490]='h00000000;
    rd_cycle[ 8491] = 1'b0;  wr_cycle[ 8491] = 1'b0;  addr_rom[ 8491]='h00000000;  wr_data_rom[ 8491]='h00000000;
    rd_cycle[ 8492] = 1'b0;  wr_cycle[ 8492] = 1'b0;  addr_rom[ 8492]='h00000000;  wr_data_rom[ 8492]='h00000000;
    rd_cycle[ 8493] = 1'b0;  wr_cycle[ 8493] = 1'b0;  addr_rom[ 8493]='h00000000;  wr_data_rom[ 8493]='h00000000;
    rd_cycle[ 8494] = 1'b0;  wr_cycle[ 8494] = 1'b0;  addr_rom[ 8494]='h00000000;  wr_data_rom[ 8494]='h00000000;
    rd_cycle[ 8495] = 1'b0;  wr_cycle[ 8495] = 1'b0;  addr_rom[ 8495]='h00000000;  wr_data_rom[ 8495]='h00000000;
    rd_cycle[ 8496] = 1'b0;  wr_cycle[ 8496] = 1'b0;  addr_rom[ 8496]='h00000000;  wr_data_rom[ 8496]='h00000000;
    rd_cycle[ 8497] = 1'b0;  wr_cycle[ 8497] = 1'b0;  addr_rom[ 8497]='h00000000;  wr_data_rom[ 8497]='h00000000;
    rd_cycle[ 8498] = 1'b0;  wr_cycle[ 8498] = 1'b0;  addr_rom[ 8498]='h00000000;  wr_data_rom[ 8498]='h00000000;
    rd_cycle[ 8499] = 1'b0;  wr_cycle[ 8499] = 1'b0;  addr_rom[ 8499]='h00000000;  wr_data_rom[ 8499]='h00000000;
    rd_cycle[ 8500] = 1'b0;  wr_cycle[ 8500] = 1'b0;  addr_rom[ 8500]='h00000000;  wr_data_rom[ 8500]='h00000000;
    rd_cycle[ 8501] = 1'b0;  wr_cycle[ 8501] = 1'b0;  addr_rom[ 8501]='h00000000;  wr_data_rom[ 8501]='h00000000;
    rd_cycle[ 8502] = 1'b0;  wr_cycle[ 8502] = 1'b0;  addr_rom[ 8502]='h00000000;  wr_data_rom[ 8502]='h00000000;
    rd_cycle[ 8503] = 1'b0;  wr_cycle[ 8503] = 1'b0;  addr_rom[ 8503]='h00000000;  wr_data_rom[ 8503]='h00000000;
    rd_cycle[ 8504] = 1'b0;  wr_cycle[ 8504] = 1'b0;  addr_rom[ 8504]='h00000000;  wr_data_rom[ 8504]='h00000000;
    rd_cycle[ 8505] = 1'b0;  wr_cycle[ 8505] = 1'b0;  addr_rom[ 8505]='h00000000;  wr_data_rom[ 8505]='h00000000;
    rd_cycle[ 8506] = 1'b0;  wr_cycle[ 8506] = 1'b0;  addr_rom[ 8506]='h00000000;  wr_data_rom[ 8506]='h00000000;
    rd_cycle[ 8507] = 1'b0;  wr_cycle[ 8507] = 1'b0;  addr_rom[ 8507]='h00000000;  wr_data_rom[ 8507]='h00000000;
    rd_cycle[ 8508] = 1'b0;  wr_cycle[ 8508] = 1'b0;  addr_rom[ 8508]='h00000000;  wr_data_rom[ 8508]='h00000000;
    rd_cycle[ 8509] = 1'b0;  wr_cycle[ 8509] = 1'b0;  addr_rom[ 8509]='h00000000;  wr_data_rom[ 8509]='h00000000;
    rd_cycle[ 8510] = 1'b0;  wr_cycle[ 8510] = 1'b0;  addr_rom[ 8510]='h00000000;  wr_data_rom[ 8510]='h00000000;
    rd_cycle[ 8511] = 1'b0;  wr_cycle[ 8511] = 1'b0;  addr_rom[ 8511]='h00000000;  wr_data_rom[ 8511]='h00000000;
    rd_cycle[ 8512] = 1'b0;  wr_cycle[ 8512] = 1'b0;  addr_rom[ 8512]='h00000000;  wr_data_rom[ 8512]='h00000000;
    rd_cycle[ 8513] = 1'b0;  wr_cycle[ 8513] = 1'b0;  addr_rom[ 8513]='h00000000;  wr_data_rom[ 8513]='h00000000;
    rd_cycle[ 8514] = 1'b0;  wr_cycle[ 8514] = 1'b0;  addr_rom[ 8514]='h00000000;  wr_data_rom[ 8514]='h00000000;
    rd_cycle[ 8515] = 1'b0;  wr_cycle[ 8515] = 1'b0;  addr_rom[ 8515]='h00000000;  wr_data_rom[ 8515]='h00000000;
    rd_cycle[ 8516] = 1'b0;  wr_cycle[ 8516] = 1'b0;  addr_rom[ 8516]='h00000000;  wr_data_rom[ 8516]='h00000000;
    rd_cycle[ 8517] = 1'b0;  wr_cycle[ 8517] = 1'b0;  addr_rom[ 8517]='h00000000;  wr_data_rom[ 8517]='h00000000;
    rd_cycle[ 8518] = 1'b0;  wr_cycle[ 8518] = 1'b0;  addr_rom[ 8518]='h00000000;  wr_data_rom[ 8518]='h00000000;
    rd_cycle[ 8519] = 1'b0;  wr_cycle[ 8519] = 1'b0;  addr_rom[ 8519]='h00000000;  wr_data_rom[ 8519]='h00000000;
    rd_cycle[ 8520] = 1'b0;  wr_cycle[ 8520] = 1'b0;  addr_rom[ 8520]='h00000000;  wr_data_rom[ 8520]='h00000000;
    rd_cycle[ 8521] = 1'b0;  wr_cycle[ 8521] = 1'b0;  addr_rom[ 8521]='h00000000;  wr_data_rom[ 8521]='h00000000;
    rd_cycle[ 8522] = 1'b0;  wr_cycle[ 8522] = 1'b0;  addr_rom[ 8522]='h00000000;  wr_data_rom[ 8522]='h00000000;
    rd_cycle[ 8523] = 1'b0;  wr_cycle[ 8523] = 1'b0;  addr_rom[ 8523]='h00000000;  wr_data_rom[ 8523]='h00000000;
    rd_cycle[ 8524] = 1'b0;  wr_cycle[ 8524] = 1'b0;  addr_rom[ 8524]='h00000000;  wr_data_rom[ 8524]='h00000000;
    rd_cycle[ 8525] = 1'b0;  wr_cycle[ 8525] = 1'b0;  addr_rom[ 8525]='h00000000;  wr_data_rom[ 8525]='h00000000;
    rd_cycle[ 8526] = 1'b0;  wr_cycle[ 8526] = 1'b0;  addr_rom[ 8526]='h00000000;  wr_data_rom[ 8526]='h00000000;
    rd_cycle[ 8527] = 1'b0;  wr_cycle[ 8527] = 1'b0;  addr_rom[ 8527]='h00000000;  wr_data_rom[ 8527]='h00000000;
    rd_cycle[ 8528] = 1'b0;  wr_cycle[ 8528] = 1'b0;  addr_rom[ 8528]='h00000000;  wr_data_rom[ 8528]='h00000000;
    rd_cycle[ 8529] = 1'b0;  wr_cycle[ 8529] = 1'b0;  addr_rom[ 8529]='h00000000;  wr_data_rom[ 8529]='h00000000;
    rd_cycle[ 8530] = 1'b0;  wr_cycle[ 8530] = 1'b0;  addr_rom[ 8530]='h00000000;  wr_data_rom[ 8530]='h00000000;
    rd_cycle[ 8531] = 1'b0;  wr_cycle[ 8531] = 1'b0;  addr_rom[ 8531]='h00000000;  wr_data_rom[ 8531]='h00000000;
    rd_cycle[ 8532] = 1'b0;  wr_cycle[ 8532] = 1'b0;  addr_rom[ 8532]='h00000000;  wr_data_rom[ 8532]='h00000000;
    rd_cycle[ 8533] = 1'b0;  wr_cycle[ 8533] = 1'b0;  addr_rom[ 8533]='h00000000;  wr_data_rom[ 8533]='h00000000;
    rd_cycle[ 8534] = 1'b0;  wr_cycle[ 8534] = 1'b0;  addr_rom[ 8534]='h00000000;  wr_data_rom[ 8534]='h00000000;
    rd_cycle[ 8535] = 1'b0;  wr_cycle[ 8535] = 1'b0;  addr_rom[ 8535]='h00000000;  wr_data_rom[ 8535]='h00000000;
    rd_cycle[ 8536] = 1'b0;  wr_cycle[ 8536] = 1'b0;  addr_rom[ 8536]='h00000000;  wr_data_rom[ 8536]='h00000000;
    rd_cycle[ 8537] = 1'b0;  wr_cycle[ 8537] = 1'b0;  addr_rom[ 8537]='h00000000;  wr_data_rom[ 8537]='h00000000;
    rd_cycle[ 8538] = 1'b0;  wr_cycle[ 8538] = 1'b0;  addr_rom[ 8538]='h00000000;  wr_data_rom[ 8538]='h00000000;
    rd_cycle[ 8539] = 1'b0;  wr_cycle[ 8539] = 1'b0;  addr_rom[ 8539]='h00000000;  wr_data_rom[ 8539]='h00000000;
    rd_cycle[ 8540] = 1'b0;  wr_cycle[ 8540] = 1'b0;  addr_rom[ 8540]='h00000000;  wr_data_rom[ 8540]='h00000000;
    rd_cycle[ 8541] = 1'b0;  wr_cycle[ 8541] = 1'b0;  addr_rom[ 8541]='h00000000;  wr_data_rom[ 8541]='h00000000;
    rd_cycle[ 8542] = 1'b0;  wr_cycle[ 8542] = 1'b0;  addr_rom[ 8542]='h00000000;  wr_data_rom[ 8542]='h00000000;
    rd_cycle[ 8543] = 1'b0;  wr_cycle[ 8543] = 1'b0;  addr_rom[ 8543]='h00000000;  wr_data_rom[ 8543]='h00000000;
    rd_cycle[ 8544] = 1'b0;  wr_cycle[ 8544] = 1'b0;  addr_rom[ 8544]='h00000000;  wr_data_rom[ 8544]='h00000000;
    rd_cycle[ 8545] = 1'b0;  wr_cycle[ 8545] = 1'b0;  addr_rom[ 8545]='h00000000;  wr_data_rom[ 8545]='h00000000;
    rd_cycle[ 8546] = 1'b0;  wr_cycle[ 8546] = 1'b0;  addr_rom[ 8546]='h00000000;  wr_data_rom[ 8546]='h00000000;
    rd_cycle[ 8547] = 1'b0;  wr_cycle[ 8547] = 1'b0;  addr_rom[ 8547]='h00000000;  wr_data_rom[ 8547]='h00000000;
    rd_cycle[ 8548] = 1'b0;  wr_cycle[ 8548] = 1'b0;  addr_rom[ 8548]='h00000000;  wr_data_rom[ 8548]='h00000000;
    rd_cycle[ 8549] = 1'b0;  wr_cycle[ 8549] = 1'b0;  addr_rom[ 8549]='h00000000;  wr_data_rom[ 8549]='h00000000;
    rd_cycle[ 8550] = 1'b0;  wr_cycle[ 8550] = 1'b0;  addr_rom[ 8550]='h00000000;  wr_data_rom[ 8550]='h00000000;
    rd_cycle[ 8551] = 1'b0;  wr_cycle[ 8551] = 1'b0;  addr_rom[ 8551]='h00000000;  wr_data_rom[ 8551]='h00000000;
    rd_cycle[ 8552] = 1'b0;  wr_cycle[ 8552] = 1'b0;  addr_rom[ 8552]='h00000000;  wr_data_rom[ 8552]='h00000000;
    rd_cycle[ 8553] = 1'b0;  wr_cycle[ 8553] = 1'b0;  addr_rom[ 8553]='h00000000;  wr_data_rom[ 8553]='h00000000;
    rd_cycle[ 8554] = 1'b0;  wr_cycle[ 8554] = 1'b0;  addr_rom[ 8554]='h00000000;  wr_data_rom[ 8554]='h00000000;
    rd_cycle[ 8555] = 1'b0;  wr_cycle[ 8555] = 1'b0;  addr_rom[ 8555]='h00000000;  wr_data_rom[ 8555]='h00000000;
    rd_cycle[ 8556] = 1'b0;  wr_cycle[ 8556] = 1'b0;  addr_rom[ 8556]='h00000000;  wr_data_rom[ 8556]='h00000000;
    rd_cycle[ 8557] = 1'b0;  wr_cycle[ 8557] = 1'b0;  addr_rom[ 8557]='h00000000;  wr_data_rom[ 8557]='h00000000;
    rd_cycle[ 8558] = 1'b0;  wr_cycle[ 8558] = 1'b0;  addr_rom[ 8558]='h00000000;  wr_data_rom[ 8558]='h00000000;
    rd_cycle[ 8559] = 1'b0;  wr_cycle[ 8559] = 1'b0;  addr_rom[ 8559]='h00000000;  wr_data_rom[ 8559]='h00000000;
    rd_cycle[ 8560] = 1'b0;  wr_cycle[ 8560] = 1'b0;  addr_rom[ 8560]='h00000000;  wr_data_rom[ 8560]='h00000000;
    rd_cycle[ 8561] = 1'b0;  wr_cycle[ 8561] = 1'b0;  addr_rom[ 8561]='h00000000;  wr_data_rom[ 8561]='h00000000;
    rd_cycle[ 8562] = 1'b0;  wr_cycle[ 8562] = 1'b0;  addr_rom[ 8562]='h00000000;  wr_data_rom[ 8562]='h00000000;
    rd_cycle[ 8563] = 1'b0;  wr_cycle[ 8563] = 1'b0;  addr_rom[ 8563]='h00000000;  wr_data_rom[ 8563]='h00000000;
    rd_cycle[ 8564] = 1'b0;  wr_cycle[ 8564] = 1'b0;  addr_rom[ 8564]='h00000000;  wr_data_rom[ 8564]='h00000000;
    rd_cycle[ 8565] = 1'b0;  wr_cycle[ 8565] = 1'b0;  addr_rom[ 8565]='h00000000;  wr_data_rom[ 8565]='h00000000;
    rd_cycle[ 8566] = 1'b0;  wr_cycle[ 8566] = 1'b0;  addr_rom[ 8566]='h00000000;  wr_data_rom[ 8566]='h00000000;
    rd_cycle[ 8567] = 1'b0;  wr_cycle[ 8567] = 1'b0;  addr_rom[ 8567]='h00000000;  wr_data_rom[ 8567]='h00000000;
    rd_cycle[ 8568] = 1'b0;  wr_cycle[ 8568] = 1'b0;  addr_rom[ 8568]='h00000000;  wr_data_rom[ 8568]='h00000000;
    rd_cycle[ 8569] = 1'b0;  wr_cycle[ 8569] = 1'b0;  addr_rom[ 8569]='h00000000;  wr_data_rom[ 8569]='h00000000;
    rd_cycle[ 8570] = 1'b0;  wr_cycle[ 8570] = 1'b0;  addr_rom[ 8570]='h00000000;  wr_data_rom[ 8570]='h00000000;
    rd_cycle[ 8571] = 1'b0;  wr_cycle[ 8571] = 1'b0;  addr_rom[ 8571]='h00000000;  wr_data_rom[ 8571]='h00000000;
    rd_cycle[ 8572] = 1'b0;  wr_cycle[ 8572] = 1'b0;  addr_rom[ 8572]='h00000000;  wr_data_rom[ 8572]='h00000000;
    rd_cycle[ 8573] = 1'b0;  wr_cycle[ 8573] = 1'b0;  addr_rom[ 8573]='h00000000;  wr_data_rom[ 8573]='h00000000;
    rd_cycle[ 8574] = 1'b0;  wr_cycle[ 8574] = 1'b0;  addr_rom[ 8574]='h00000000;  wr_data_rom[ 8574]='h00000000;
    rd_cycle[ 8575] = 1'b0;  wr_cycle[ 8575] = 1'b0;  addr_rom[ 8575]='h00000000;  wr_data_rom[ 8575]='h00000000;
    rd_cycle[ 8576] = 1'b0;  wr_cycle[ 8576] = 1'b0;  addr_rom[ 8576]='h00000000;  wr_data_rom[ 8576]='h00000000;
    rd_cycle[ 8577] = 1'b0;  wr_cycle[ 8577] = 1'b0;  addr_rom[ 8577]='h00000000;  wr_data_rom[ 8577]='h00000000;
    rd_cycle[ 8578] = 1'b0;  wr_cycle[ 8578] = 1'b0;  addr_rom[ 8578]='h00000000;  wr_data_rom[ 8578]='h00000000;
    rd_cycle[ 8579] = 1'b0;  wr_cycle[ 8579] = 1'b0;  addr_rom[ 8579]='h00000000;  wr_data_rom[ 8579]='h00000000;
    rd_cycle[ 8580] = 1'b0;  wr_cycle[ 8580] = 1'b0;  addr_rom[ 8580]='h00000000;  wr_data_rom[ 8580]='h00000000;
    rd_cycle[ 8581] = 1'b0;  wr_cycle[ 8581] = 1'b0;  addr_rom[ 8581]='h00000000;  wr_data_rom[ 8581]='h00000000;
    rd_cycle[ 8582] = 1'b0;  wr_cycle[ 8582] = 1'b0;  addr_rom[ 8582]='h00000000;  wr_data_rom[ 8582]='h00000000;
    rd_cycle[ 8583] = 1'b0;  wr_cycle[ 8583] = 1'b0;  addr_rom[ 8583]='h00000000;  wr_data_rom[ 8583]='h00000000;
    rd_cycle[ 8584] = 1'b0;  wr_cycle[ 8584] = 1'b0;  addr_rom[ 8584]='h00000000;  wr_data_rom[ 8584]='h00000000;
    rd_cycle[ 8585] = 1'b0;  wr_cycle[ 8585] = 1'b0;  addr_rom[ 8585]='h00000000;  wr_data_rom[ 8585]='h00000000;
    rd_cycle[ 8586] = 1'b0;  wr_cycle[ 8586] = 1'b0;  addr_rom[ 8586]='h00000000;  wr_data_rom[ 8586]='h00000000;
    rd_cycle[ 8587] = 1'b0;  wr_cycle[ 8587] = 1'b0;  addr_rom[ 8587]='h00000000;  wr_data_rom[ 8587]='h00000000;
    rd_cycle[ 8588] = 1'b0;  wr_cycle[ 8588] = 1'b0;  addr_rom[ 8588]='h00000000;  wr_data_rom[ 8588]='h00000000;
    rd_cycle[ 8589] = 1'b0;  wr_cycle[ 8589] = 1'b0;  addr_rom[ 8589]='h00000000;  wr_data_rom[ 8589]='h00000000;
    rd_cycle[ 8590] = 1'b0;  wr_cycle[ 8590] = 1'b0;  addr_rom[ 8590]='h00000000;  wr_data_rom[ 8590]='h00000000;
    rd_cycle[ 8591] = 1'b0;  wr_cycle[ 8591] = 1'b0;  addr_rom[ 8591]='h00000000;  wr_data_rom[ 8591]='h00000000;
    rd_cycle[ 8592] = 1'b0;  wr_cycle[ 8592] = 1'b0;  addr_rom[ 8592]='h00000000;  wr_data_rom[ 8592]='h00000000;
    rd_cycle[ 8593] = 1'b0;  wr_cycle[ 8593] = 1'b0;  addr_rom[ 8593]='h00000000;  wr_data_rom[ 8593]='h00000000;
    rd_cycle[ 8594] = 1'b0;  wr_cycle[ 8594] = 1'b0;  addr_rom[ 8594]='h00000000;  wr_data_rom[ 8594]='h00000000;
    rd_cycle[ 8595] = 1'b0;  wr_cycle[ 8595] = 1'b0;  addr_rom[ 8595]='h00000000;  wr_data_rom[ 8595]='h00000000;
    rd_cycle[ 8596] = 1'b0;  wr_cycle[ 8596] = 1'b0;  addr_rom[ 8596]='h00000000;  wr_data_rom[ 8596]='h00000000;
    rd_cycle[ 8597] = 1'b0;  wr_cycle[ 8597] = 1'b0;  addr_rom[ 8597]='h00000000;  wr_data_rom[ 8597]='h00000000;
    rd_cycle[ 8598] = 1'b0;  wr_cycle[ 8598] = 1'b0;  addr_rom[ 8598]='h00000000;  wr_data_rom[ 8598]='h00000000;
    rd_cycle[ 8599] = 1'b0;  wr_cycle[ 8599] = 1'b0;  addr_rom[ 8599]='h00000000;  wr_data_rom[ 8599]='h00000000;
    rd_cycle[ 8600] = 1'b0;  wr_cycle[ 8600] = 1'b0;  addr_rom[ 8600]='h00000000;  wr_data_rom[ 8600]='h00000000;
    rd_cycle[ 8601] = 1'b0;  wr_cycle[ 8601] = 1'b0;  addr_rom[ 8601]='h00000000;  wr_data_rom[ 8601]='h00000000;
    rd_cycle[ 8602] = 1'b0;  wr_cycle[ 8602] = 1'b0;  addr_rom[ 8602]='h00000000;  wr_data_rom[ 8602]='h00000000;
    rd_cycle[ 8603] = 1'b0;  wr_cycle[ 8603] = 1'b0;  addr_rom[ 8603]='h00000000;  wr_data_rom[ 8603]='h00000000;
    rd_cycle[ 8604] = 1'b0;  wr_cycle[ 8604] = 1'b0;  addr_rom[ 8604]='h00000000;  wr_data_rom[ 8604]='h00000000;
    rd_cycle[ 8605] = 1'b0;  wr_cycle[ 8605] = 1'b0;  addr_rom[ 8605]='h00000000;  wr_data_rom[ 8605]='h00000000;
    rd_cycle[ 8606] = 1'b0;  wr_cycle[ 8606] = 1'b0;  addr_rom[ 8606]='h00000000;  wr_data_rom[ 8606]='h00000000;
    rd_cycle[ 8607] = 1'b0;  wr_cycle[ 8607] = 1'b0;  addr_rom[ 8607]='h00000000;  wr_data_rom[ 8607]='h00000000;
    rd_cycle[ 8608] = 1'b0;  wr_cycle[ 8608] = 1'b0;  addr_rom[ 8608]='h00000000;  wr_data_rom[ 8608]='h00000000;
    rd_cycle[ 8609] = 1'b0;  wr_cycle[ 8609] = 1'b0;  addr_rom[ 8609]='h00000000;  wr_data_rom[ 8609]='h00000000;
    rd_cycle[ 8610] = 1'b0;  wr_cycle[ 8610] = 1'b0;  addr_rom[ 8610]='h00000000;  wr_data_rom[ 8610]='h00000000;
    rd_cycle[ 8611] = 1'b0;  wr_cycle[ 8611] = 1'b0;  addr_rom[ 8611]='h00000000;  wr_data_rom[ 8611]='h00000000;
    rd_cycle[ 8612] = 1'b0;  wr_cycle[ 8612] = 1'b0;  addr_rom[ 8612]='h00000000;  wr_data_rom[ 8612]='h00000000;
    rd_cycle[ 8613] = 1'b0;  wr_cycle[ 8613] = 1'b0;  addr_rom[ 8613]='h00000000;  wr_data_rom[ 8613]='h00000000;
    rd_cycle[ 8614] = 1'b0;  wr_cycle[ 8614] = 1'b0;  addr_rom[ 8614]='h00000000;  wr_data_rom[ 8614]='h00000000;
    rd_cycle[ 8615] = 1'b0;  wr_cycle[ 8615] = 1'b0;  addr_rom[ 8615]='h00000000;  wr_data_rom[ 8615]='h00000000;
    rd_cycle[ 8616] = 1'b0;  wr_cycle[ 8616] = 1'b0;  addr_rom[ 8616]='h00000000;  wr_data_rom[ 8616]='h00000000;
    rd_cycle[ 8617] = 1'b0;  wr_cycle[ 8617] = 1'b0;  addr_rom[ 8617]='h00000000;  wr_data_rom[ 8617]='h00000000;
    rd_cycle[ 8618] = 1'b0;  wr_cycle[ 8618] = 1'b0;  addr_rom[ 8618]='h00000000;  wr_data_rom[ 8618]='h00000000;
    rd_cycle[ 8619] = 1'b0;  wr_cycle[ 8619] = 1'b0;  addr_rom[ 8619]='h00000000;  wr_data_rom[ 8619]='h00000000;
    rd_cycle[ 8620] = 1'b0;  wr_cycle[ 8620] = 1'b0;  addr_rom[ 8620]='h00000000;  wr_data_rom[ 8620]='h00000000;
    rd_cycle[ 8621] = 1'b0;  wr_cycle[ 8621] = 1'b0;  addr_rom[ 8621]='h00000000;  wr_data_rom[ 8621]='h00000000;
    rd_cycle[ 8622] = 1'b0;  wr_cycle[ 8622] = 1'b0;  addr_rom[ 8622]='h00000000;  wr_data_rom[ 8622]='h00000000;
    rd_cycle[ 8623] = 1'b0;  wr_cycle[ 8623] = 1'b0;  addr_rom[ 8623]='h00000000;  wr_data_rom[ 8623]='h00000000;
    rd_cycle[ 8624] = 1'b0;  wr_cycle[ 8624] = 1'b0;  addr_rom[ 8624]='h00000000;  wr_data_rom[ 8624]='h00000000;
    rd_cycle[ 8625] = 1'b0;  wr_cycle[ 8625] = 1'b0;  addr_rom[ 8625]='h00000000;  wr_data_rom[ 8625]='h00000000;
    rd_cycle[ 8626] = 1'b0;  wr_cycle[ 8626] = 1'b0;  addr_rom[ 8626]='h00000000;  wr_data_rom[ 8626]='h00000000;
    rd_cycle[ 8627] = 1'b0;  wr_cycle[ 8627] = 1'b0;  addr_rom[ 8627]='h00000000;  wr_data_rom[ 8627]='h00000000;
    rd_cycle[ 8628] = 1'b0;  wr_cycle[ 8628] = 1'b0;  addr_rom[ 8628]='h00000000;  wr_data_rom[ 8628]='h00000000;
    rd_cycle[ 8629] = 1'b0;  wr_cycle[ 8629] = 1'b0;  addr_rom[ 8629]='h00000000;  wr_data_rom[ 8629]='h00000000;
    rd_cycle[ 8630] = 1'b0;  wr_cycle[ 8630] = 1'b0;  addr_rom[ 8630]='h00000000;  wr_data_rom[ 8630]='h00000000;
    rd_cycle[ 8631] = 1'b0;  wr_cycle[ 8631] = 1'b0;  addr_rom[ 8631]='h00000000;  wr_data_rom[ 8631]='h00000000;
    rd_cycle[ 8632] = 1'b0;  wr_cycle[ 8632] = 1'b0;  addr_rom[ 8632]='h00000000;  wr_data_rom[ 8632]='h00000000;
    rd_cycle[ 8633] = 1'b0;  wr_cycle[ 8633] = 1'b0;  addr_rom[ 8633]='h00000000;  wr_data_rom[ 8633]='h00000000;
    rd_cycle[ 8634] = 1'b0;  wr_cycle[ 8634] = 1'b0;  addr_rom[ 8634]='h00000000;  wr_data_rom[ 8634]='h00000000;
    rd_cycle[ 8635] = 1'b0;  wr_cycle[ 8635] = 1'b0;  addr_rom[ 8635]='h00000000;  wr_data_rom[ 8635]='h00000000;
    rd_cycle[ 8636] = 1'b0;  wr_cycle[ 8636] = 1'b0;  addr_rom[ 8636]='h00000000;  wr_data_rom[ 8636]='h00000000;
    rd_cycle[ 8637] = 1'b0;  wr_cycle[ 8637] = 1'b0;  addr_rom[ 8637]='h00000000;  wr_data_rom[ 8637]='h00000000;
    rd_cycle[ 8638] = 1'b0;  wr_cycle[ 8638] = 1'b0;  addr_rom[ 8638]='h00000000;  wr_data_rom[ 8638]='h00000000;
    rd_cycle[ 8639] = 1'b0;  wr_cycle[ 8639] = 1'b0;  addr_rom[ 8639]='h00000000;  wr_data_rom[ 8639]='h00000000;
    rd_cycle[ 8640] = 1'b0;  wr_cycle[ 8640] = 1'b0;  addr_rom[ 8640]='h00000000;  wr_data_rom[ 8640]='h00000000;
    rd_cycle[ 8641] = 1'b0;  wr_cycle[ 8641] = 1'b0;  addr_rom[ 8641]='h00000000;  wr_data_rom[ 8641]='h00000000;
    rd_cycle[ 8642] = 1'b0;  wr_cycle[ 8642] = 1'b0;  addr_rom[ 8642]='h00000000;  wr_data_rom[ 8642]='h00000000;
    rd_cycle[ 8643] = 1'b0;  wr_cycle[ 8643] = 1'b0;  addr_rom[ 8643]='h00000000;  wr_data_rom[ 8643]='h00000000;
    rd_cycle[ 8644] = 1'b0;  wr_cycle[ 8644] = 1'b0;  addr_rom[ 8644]='h00000000;  wr_data_rom[ 8644]='h00000000;
    rd_cycle[ 8645] = 1'b0;  wr_cycle[ 8645] = 1'b0;  addr_rom[ 8645]='h00000000;  wr_data_rom[ 8645]='h00000000;
    rd_cycle[ 8646] = 1'b0;  wr_cycle[ 8646] = 1'b0;  addr_rom[ 8646]='h00000000;  wr_data_rom[ 8646]='h00000000;
    rd_cycle[ 8647] = 1'b0;  wr_cycle[ 8647] = 1'b0;  addr_rom[ 8647]='h00000000;  wr_data_rom[ 8647]='h00000000;
    rd_cycle[ 8648] = 1'b0;  wr_cycle[ 8648] = 1'b0;  addr_rom[ 8648]='h00000000;  wr_data_rom[ 8648]='h00000000;
    rd_cycle[ 8649] = 1'b0;  wr_cycle[ 8649] = 1'b0;  addr_rom[ 8649]='h00000000;  wr_data_rom[ 8649]='h00000000;
    rd_cycle[ 8650] = 1'b0;  wr_cycle[ 8650] = 1'b0;  addr_rom[ 8650]='h00000000;  wr_data_rom[ 8650]='h00000000;
    rd_cycle[ 8651] = 1'b0;  wr_cycle[ 8651] = 1'b0;  addr_rom[ 8651]='h00000000;  wr_data_rom[ 8651]='h00000000;
    rd_cycle[ 8652] = 1'b0;  wr_cycle[ 8652] = 1'b0;  addr_rom[ 8652]='h00000000;  wr_data_rom[ 8652]='h00000000;
    rd_cycle[ 8653] = 1'b0;  wr_cycle[ 8653] = 1'b0;  addr_rom[ 8653]='h00000000;  wr_data_rom[ 8653]='h00000000;
    rd_cycle[ 8654] = 1'b0;  wr_cycle[ 8654] = 1'b0;  addr_rom[ 8654]='h00000000;  wr_data_rom[ 8654]='h00000000;
    rd_cycle[ 8655] = 1'b0;  wr_cycle[ 8655] = 1'b0;  addr_rom[ 8655]='h00000000;  wr_data_rom[ 8655]='h00000000;
    rd_cycle[ 8656] = 1'b0;  wr_cycle[ 8656] = 1'b0;  addr_rom[ 8656]='h00000000;  wr_data_rom[ 8656]='h00000000;
    rd_cycle[ 8657] = 1'b0;  wr_cycle[ 8657] = 1'b0;  addr_rom[ 8657]='h00000000;  wr_data_rom[ 8657]='h00000000;
    rd_cycle[ 8658] = 1'b0;  wr_cycle[ 8658] = 1'b0;  addr_rom[ 8658]='h00000000;  wr_data_rom[ 8658]='h00000000;
    rd_cycle[ 8659] = 1'b0;  wr_cycle[ 8659] = 1'b0;  addr_rom[ 8659]='h00000000;  wr_data_rom[ 8659]='h00000000;
    rd_cycle[ 8660] = 1'b0;  wr_cycle[ 8660] = 1'b0;  addr_rom[ 8660]='h00000000;  wr_data_rom[ 8660]='h00000000;
    rd_cycle[ 8661] = 1'b0;  wr_cycle[ 8661] = 1'b0;  addr_rom[ 8661]='h00000000;  wr_data_rom[ 8661]='h00000000;
    rd_cycle[ 8662] = 1'b0;  wr_cycle[ 8662] = 1'b0;  addr_rom[ 8662]='h00000000;  wr_data_rom[ 8662]='h00000000;
    rd_cycle[ 8663] = 1'b0;  wr_cycle[ 8663] = 1'b0;  addr_rom[ 8663]='h00000000;  wr_data_rom[ 8663]='h00000000;
    rd_cycle[ 8664] = 1'b0;  wr_cycle[ 8664] = 1'b0;  addr_rom[ 8664]='h00000000;  wr_data_rom[ 8664]='h00000000;
    rd_cycle[ 8665] = 1'b0;  wr_cycle[ 8665] = 1'b0;  addr_rom[ 8665]='h00000000;  wr_data_rom[ 8665]='h00000000;
    rd_cycle[ 8666] = 1'b0;  wr_cycle[ 8666] = 1'b0;  addr_rom[ 8666]='h00000000;  wr_data_rom[ 8666]='h00000000;
    rd_cycle[ 8667] = 1'b0;  wr_cycle[ 8667] = 1'b0;  addr_rom[ 8667]='h00000000;  wr_data_rom[ 8667]='h00000000;
    rd_cycle[ 8668] = 1'b0;  wr_cycle[ 8668] = 1'b0;  addr_rom[ 8668]='h00000000;  wr_data_rom[ 8668]='h00000000;
    rd_cycle[ 8669] = 1'b0;  wr_cycle[ 8669] = 1'b0;  addr_rom[ 8669]='h00000000;  wr_data_rom[ 8669]='h00000000;
    rd_cycle[ 8670] = 1'b0;  wr_cycle[ 8670] = 1'b0;  addr_rom[ 8670]='h00000000;  wr_data_rom[ 8670]='h00000000;
    rd_cycle[ 8671] = 1'b0;  wr_cycle[ 8671] = 1'b0;  addr_rom[ 8671]='h00000000;  wr_data_rom[ 8671]='h00000000;
    rd_cycle[ 8672] = 1'b0;  wr_cycle[ 8672] = 1'b0;  addr_rom[ 8672]='h00000000;  wr_data_rom[ 8672]='h00000000;
    rd_cycle[ 8673] = 1'b0;  wr_cycle[ 8673] = 1'b0;  addr_rom[ 8673]='h00000000;  wr_data_rom[ 8673]='h00000000;
    rd_cycle[ 8674] = 1'b0;  wr_cycle[ 8674] = 1'b0;  addr_rom[ 8674]='h00000000;  wr_data_rom[ 8674]='h00000000;
    rd_cycle[ 8675] = 1'b0;  wr_cycle[ 8675] = 1'b0;  addr_rom[ 8675]='h00000000;  wr_data_rom[ 8675]='h00000000;
    rd_cycle[ 8676] = 1'b0;  wr_cycle[ 8676] = 1'b0;  addr_rom[ 8676]='h00000000;  wr_data_rom[ 8676]='h00000000;
    rd_cycle[ 8677] = 1'b0;  wr_cycle[ 8677] = 1'b0;  addr_rom[ 8677]='h00000000;  wr_data_rom[ 8677]='h00000000;
    rd_cycle[ 8678] = 1'b0;  wr_cycle[ 8678] = 1'b0;  addr_rom[ 8678]='h00000000;  wr_data_rom[ 8678]='h00000000;
    rd_cycle[ 8679] = 1'b0;  wr_cycle[ 8679] = 1'b0;  addr_rom[ 8679]='h00000000;  wr_data_rom[ 8679]='h00000000;
    rd_cycle[ 8680] = 1'b0;  wr_cycle[ 8680] = 1'b0;  addr_rom[ 8680]='h00000000;  wr_data_rom[ 8680]='h00000000;
    rd_cycle[ 8681] = 1'b0;  wr_cycle[ 8681] = 1'b0;  addr_rom[ 8681]='h00000000;  wr_data_rom[ 8681]='h00000000;
    rd_cycle[ 8682] = 1'b0;  wr_cycle[ 8682] = 1'b0;  addr_rom[ 8682]='h00000000;  wr_data_rom[ 8682]='h00000000;
    rd_cycle[ 8683] = 1'b0;  wr_cycle[ 8683] = 1'b0;  addr_rom[ 8683]='h00000000;  wr_data_rom[ 8683]='h00000000;
    rd_cycle[ 8684] = 1'b0;  wr_cycle[ 8684] = 1'b0;  addr_rom[ 8684]='h00000000;  wr_data_rom[ 8684]='h00000000;
    rd_cycle[ 8685] = 1'b0;  wr_cycle[ 8685] = 1'b0;  addr_rom[ 8685]='h00000000;  wr_data_rom[ 8685]='h00000000;
    rd_cycle[ 8686] = 1'b0;  wr_cycle[ 8686] = 1'b0;  addr_rom[ 8686]='h00000000;  wr_data_rom[ 8686]='h00000000;
    rd_cycle[ 8687] = 1'b0;  wr_cycle[ 8687] = 1'b0;  addr_rom[ 8687]='h00000000;  wr_data_rom[ 8687]='h00000000;
    rd_cycle[ 8688] = 1'b0;  wr_cycle[ 8688] = 1'b0;  addr_rom[ 8688]='h00000000;  wr_data_rom[ 8688]='h00000000;
    rd_cycle[ 8689] = 1'b0;  wr_cycle[ 8689] = 1'b0;  addr_rom[ 8689]='h00000000;  wr_data_rom[ 8689]='h00000000;
    rd_cycle[ 8690] = 1'b0;  wr_cycle[ 8690] = 1'b0;  addr_rom[ 8690]='h00000000;  wr_data_rom[ 8690]='h00000000;
    rd_cycle[ 8691] = 1'b0;  wr_cycle[ 8691] = 1'b0;  addr_rom[ 8691]='h00000000;  wr_data_rom[ 8691]='h00000000;
    rd_cycle[ 8692] = 1'b0;  wr_cycle[ 8692] = 1'b0;  addr_rom[ 8692]='h00000000;  wr_data_rom[ 8692]='h00000000;
    rd_cycle[ 8693] = 1'b0;  wr_cycle[ 8693] = 1'b0;  addr_rom[ 8693]='h00000000;  wr_data_rom[ 8693]='h00000000;
    rd_cycle[ 8694] = 1'b0;  wr_cycle[ 8694] = 1'b0;  addr_rom[ 8694]='h00000000;  wr_data_rom[ 8694]='h00000000;
    rd_cycle[ 8695] = 1'b0;  wr_cycle[ 8695] = 1'b0;  addr_rom[ 8695]='h00000000;  wr_data_rom[ 8695]='h00000000;
    rd_cycle[ 8696] = 1'b0;  wr_cycle[ 8696] = 1'b0;  addr_rom[ 8696]='h00000000;  wr_data_rom[ 8696]='h00000000;
    rd_cycle[ 8697] = 1'b0;  wr_cycle[ 8697] = 1'b0;  addr_rom[ 8697]='h00000000;  wr_data_rom[ 8697]='h00000000;
    rd_cycle[ 8698] = 1'b0;  wr_cycle[ 8698] = 1'b0;  addr_rom[ 8698]='h00000000;  wr_data_rom[ 8698]='h00000000;
    rd_cycle[ 8699] = 1'b0;  wr_cycle[ 8699] = 1'b0;  addr_rom[ 8699]='h00000000;  wr_data_rom[ 8699]='h00000000;
    rd_cycle[ 8700] = 1'b0;  wr_cycle[ 8700] = 1'b0;  addr_rom[ 8700]='h00000000;  wr_data_rom[ 8700]='h00000000;
    rd_cycle[ 8701] = 1'b0;  wr_cycle[ 8701] = 1'b0;  addr_rom[ 8701]='h00000000;  wr_data_rom[ 8701]='h00000000;
    rd_cycle[ 8702] = 1'b0;  wr_cycle[ 8702] = 1'b0;  addr_rom[ 8702]='h00000000;  wr_data_rom[ 8702]='h00000000;
    rd_cycle[ 8703] = 1'b0;  wr_cycle[ 8703] = 1'b0;  addr_rom[ 8703]='h00000000;  wr_data_rom[ 8703]='h00000000;
    rd_cycle[ 8704] = 1'b0;  wr_cycle[ 8704] = 1'b0;  addr_rom[ 8704]='h00000000;  wr_data_rom[ 8704]='h00000000;
    rd_cycle[ 8705] = 1'b0;  wr_cycle[ 8705] = 1'b0;  addr_rom[ 8705]='h00000000;  wr_data_rom[ 8705]='h00000000;
    rd_cycle[ 8706] = 1'b0;  wr_cycle[ 8706] = 1'b0;  addr_rom[ 8706]='h00000000;  wr_data_rom[ 8706]='h00000000;
    rd_cycle[ 8707] = 1'b0;  wr_cycle[ 8707] = 1'b0;  addr_rom[ 8707]='h00000000;  wr_data_rom[ 8707]='h00000000;
    rd_cycle[ 8708] = 1'b0;  wr_cycle[ 8708] = 1'b0;  addr_rom[ 8708]='h00000000;  wr_data_rom[ 8708]='h00000000;
    rd_cycle[ 8709] = 1'b0;  wr_cycle[ 8709] = 1'b0;  addr_rom[ 8709]='h00000000;  wr_data_rom[ 8709]='h00000000;
    rd_cycle[ 8710] = 1'b0;  wr_cycle[ 8710] = 1'b0;  addr_rom[ 8710]='h00000000;  wr_data_rom[ 8710]='h00000000;
    rd_cycle[ 8711] = 1'b0;  wr_cycle[ 8711] = 1'b0;  addr_rom[ 8711]='h00000000;  wr_data_rom[ 8711]='h00000000;
    rd_cycle[ 8712] = 1'b0;  wr_cycle[ 8712] = 1'b0;  addr_rom[ 8712]='h00000000;  wr_data_rom[ 8712]='h00000000;
    rd_cycle[ 8713] = 1'b0;  wr_cycle[ 8713] = 1'b0;  addr_rom[ 8713]='h00000000;  wr_data_rom[ 8713]='h00000000;
    rd_cycle[ 8714] = 1'b0;  wr_cycle[ 8714] = 1'b0;  addr_rom[ 8714]='h00000000;  wr_data_rom[ 8714]='h00000000;
    rd_cycle[ 8715] = 1'b0;  wr_cycle[ 8715] = 1'b0;  addr_rom[ 8715]='h00000000;  wr_data_rom[ 8715]='h00000000;
    rd_cycle[ 8716] = 1'b0;  wr_cycle[ 8716] = 1'b0;  addr_rom[ 8716]='h00000000;  wr_data_rom[ 8716]='h00000000;
    rd_cycle[ 8717] = 1'b0;  wr_cycle[ 8717] = 1'b0;  addr_rom[ 8717]='h00000000;  wr_data_rom[ 8717]='h00000000;
    rd_cycle[ 8718] = 1'b0;  wr_cycle[ 8718] = 1'b0;  addr_rom[ 8718]='h00000000;  wr_data_rom[ 8718]='h00000000;
    rd_cycle[ 8719] = 1'b0;  wr_cycle[ 8719] = 1'b0;  addr_rom[ 8719]='h00000000;  wr_data_rom[ 8719]='h00000000;
    rd_cycle[ 8720] = 1'b0;  wr_cycle[ 8720] = 1'b0;  addr_rom[ 8720]='h00000000;  wr_data_rom[ 8720]='h00000000;
    rd_cycle[ 8721] = 1'b0;  wr_cycle[ 8721] = 1'b0;  addr_rom[ 8721]='h00000000;  wr_data_rom[ 8721]='h00000000;
    rd_cycle[ 8722] = 1'b0;  wr_cycle[ 8722] = 1'b0;  addr_rom[ 8722]='h00000000;  wr_data_rom[ 8722]='h00000000;
    rd_cycle[ 8723] = 1'b0;  wr_cycle[ 8723] = 1'b0;  addr_rom[ 8723]='h00000000;  wr_data_rom[ 8723]='h00000000;
    rd_cycle[ 8724] = 1'b0;  wr_cycle[ 8724] = 1'b0;  addr_rom[ 8724]='h00000000;  wr_data_rom[ 8724]='h00000000;
    rd_cycle[ 8725] = 1'b0;  wr_cycle[ 8725] = 1'b0;  addr_rom[ 8725]='h00000000;  wr_data_rom[ 8725]='h00000000;
    rd_cycle[ 8726] = 1'b0;  wr_cycle[ 8726] = 1'b0;  addr_rom[ 8726]='h00000000;  wr_data_rom[ 8726]='h00000000;
    rd_cycle[ 8727] = 1'b0;  wr_cycle[ 8727] = 1'b0;  addr_rom[ 8727]='h00000000;  wr_data_rom[ 8727]='h00000000;
    rd_cycle[ 8728] = 1'b0;  wr_cycle[ 8728] = 1'b0;  addr_rom[ 8728]='h00000000;  wr_data_rom[ 8728]='h00000000;
    rd_cycle[ 8729] = 1'b0;  wr_cycle[ 8729] = 1'b0;  addr_rom[ 8729]='h00000000;  wr_data_rom[ 8729]='h00000000;
    rd_cycle[ 8730] = 1'b0;  wr_cycle[ 8730] = 1'b0;  addr_rom[ 8730]='h00000000;  wr_data_rom[ 8730]='h00000000;
    rd_cycle[ 8731] = 1'b0;  wr_cycle[ 8731] = 1'b0;  addr_rom[ 8731]='h00000000;  wr_data_rom[ 8731]='h00000000;
    rd_cycle[ 8732] = 1'b0;  wr_cycle[ 8732] = 1'b0;  addr_rom[ 8732]='h00000000;  wr_data_rom[ 8732]='h00000000;
    rd_cycle[ 8733] = 1'b0;  wr_cycle[ 8733] = 1'b0;  addr_rom[ 8733]='h00000000;  wr_data_rom[ 8733]='h00000000;
    rd_cycle[ 8734] = 1'b0;  wr_cycle[ 8734] = 1'b0;  addr_rom[ 8734]='h00000000;  wr_data_rom[ 8734]='h00000000;
    rd_cycle[ 8735] = 1'b0;  wr_cycle[ 8735] = 1'b0;  addr_rom[ 8735]='h00000000;  wr_data_rom[ 8735]='h00000000;
    rd_cycle[ 8736] = 1'b0;  wr_cycle[ 8736] = 1'b0;  addr_rom[ 8736]='h00000000;  wr_data_rom[ 8736]='h00000000;
    rd_cycle[ 8737] = 1'b0;  wr_cycle[ 8737] = 1'b0;  addr_rom[ 8737]='h00000000;  wr_data_rom[ 8737]='h00000000;
    rd_cycle[ 8738] = 1'b0;  wr_cycle[ 8738] = 1'b0;  addr_rom[ 8738]='h00000000;  wr_data_rom[ 8738]='h00000000;
    rd_cycle[ 8739] = 1'b0;  wr_cycle[ 8739] = 1'b0;  addr_rom[ 8739]='h00000000;  wr_data_rom[ 8739]='h00000000;
    rd_cycle[ 8740] = 1'b0;  wr_cycle[ 8740] = 1'b0;  addr_rom[ 8740]='h00000000;  wr_data_rom[ 8740]='h00000000;
    rd_cycle[ 8741] = 1'b0;  wr_cycle[ 8741] = 1'b0;  addr_rom[ 8741]='h00000000;  wr_data_rom[ 8741]='h00000000;
    rd_cycle[ 8742] = 1'b0;  wr_cycle[ 8742] = 1'b0;  addr_rom[ 8742]='h00000000;  wr_data_rom[ 8742]='h00000000;
    rd_cycle[ 8743] = 1'b0;  wr_cycle[ 8743] = 1'b0;  addr_rom[ 8743]='h00000000;  wr_data_rom[ 8743]='h00000000;
    rd_cycle[ 8744] = 1'b0;  wr_cycle[ 8744] = 1'b0;  addr_rom[ 8744]='h00000000;  wr_data_rom[ 8744]='h00000000;
    rd_cycle[ 8745] = 1'b0;  wr_cycle[ 8745] = 1'b0;  addr_rom[ 8745]='h00000000;  wr_data_rom[ 8745]='h00000000;
    rd_cycle[ 8746] = 1'b0;  wr_cycle[ 8746] = 1'b0;  addr_rom[ 8746]='h00000000;  wr_data_rom[ 8746]='h00000000;
    rd_cycle[ 8747] = 1'b0;  wr_cycle[ 8747] = 1'b0;  addr_rom[ 8747]='h00000000;  wr_data_rom[ 8747]='h00000000;
    rd_cycle[ 8748] = 1'b0;  wr_cycle[ 8748] = 1'b0;  addr_rom[ 8748]='h00000000;  wr_data_rom[ 8748]='h00000000;
    rd_cycle[ 8749] = 1'b0;  wr_cycle[ 8749] = 1'b0;  addr_rom[ 8749]='h00000000;  wr_data_rom[ 8749]='h00000000;
    rd_cycle[ 8750] = 1'b0;  wr_cycle[ 8750] = 1'b0;  addr_rom[ 8750]='h00000000;  wr_data_rom[ 8750]='h00000000;
    rd_cycle[ 8751] = 1'b0;  wr_cycle[ 8751] = 1'b0;  addr_rom[ 8751]='h00000000;  wr_data_rom[ 8751]='h00000000;
    rd_cycle[ 8752] = 1'b0;  wr_cycle[ 8752] = 1'b0;  addr_rom[ 8752]='h00000000;  wr_data_rom[ 8752]='h00000000;
    rd_cycle[ 8753] = 1'b0;  wr_cycle[ 8753] = 1'b0;  addr_rom[ 8753]='h00000000;  wr_data_rom[ 8753]='h00000000;
    rd_cycle[ 8754] = 1'b0;  wr_cycle[ 8754] = 1'b0;  addr_rom[ 8754]='h00000000;  wr_data_rom[ 8754]='h00000000;
    rd_cycle[ 8755] = 1'b0;  wr_cycle[ 8755] = 1'b0;  addr_rom[ 8755]='h00000000;  wr_data_rom[ 8755]='h00000000;
    rd_cycle[ 8756] = 1'b0;  wr_cycle[ 8756] = 1'b0;  addr_rom[ 8756]='h00000000;  wr_data_rom[ 8756]='h00000000;
    rd_cycle[ 8757] = 1'b0;  wr_cycle[ 8757] = 1'b0;  addr_rom[ 8757]='h00000000;  wr_data_rom[ 8757]='h00000000;
    rd_cycle[ 8758] = 1'b0;  wr_cycle[ 8758] = 1'b0;  addr_rom[ 8758]='h00000000;  wr_data_rom[ 8758]='h00000000;
    rd_cycle[ 8759] = 1'b0;  wr_cycle[ 8759] = 1'b0;  addr_rom[ 8759]='h00000000;  wr_data_rom[ 8759]='h00000000;
    rd_cycle[ 8760] = 1'b0;  wr_cycle[ 8760] = 1'b0;  addr_rom[ 8760]='h00000000;  wr_data_rom[ 8760]='h00000000;
    rd_cycle[ 8761] = 1'b0;  wr_cycle[ 8761] = 1'b0;  addr_rom[ 8761]='h00000000;  wr_data_rom[ 8761]='h00000000;
    rd_cycle[ 8762] = 1'b0;  wr_cycle[ 8762] = 1'b0;  addr_rom[ 8762]='h00000000;  wr_data_rom[ 8762]='h00000000;
    rd_cycle[ 8763] = 1'b0;  wr_cycle[ 8763] = 1'b0;  addr_rom[ 8763]='h00000000;  wr_data_rom[ 8763]='h00000000;
    rd_cycle[ 8764] = 1'b0;  wr_cycle[ 8764] = 1'b0;  addr_rom[ 8764]='h00000000;  wr_data_rom[ 8764]='h00000000;
    rd_cycle[ 8765] = 1'b0;  wr_cycle[ 8765] = 1'b0;  addr_rom[ 8765]='h00000000;  wr_data_rom[ 8765]='h00000000;
    rd_cycle[ 8766] = 1'b0;  wr_cycle[ 8766] = 1'b0;  addr_rom[ 8766]='h00000000;  wr_data_rom[ 8766]='h00000000;
    rd_cycle[ 8767] = 1'b0;  wr_cycle[ 8767] = 1'b0;  addr_rom[ 8767]='h00000000;  wr_data_rom[ 8767]='h00000000;
    rd_cycle[ 8768] = 1'b0;  wr_cycle[ 8768] = 1'b0;  addr_rom[ 8768]='h00000000;  wr_data_rom[ 8768]='h00000000;
    rd_cycle[ 8769] = 1'b0;  wr_cycle[ 8769] = 1'b0;  addr_rom[ 8769]='h00000000;  wr_data_rom[ 8769]='h00000000;
    rd_cycle[ 8770] = 1'b0;  wr_cycle[ 8770] = 1'b0;  addr_rom[ 8770]='h00000000;  wr_data_rom[ 8770]='h00000000;
    rd_cycle[ 8771] = 1'b0;  wr_cycle[ 8771] = 1'b0;  addr_rom[ 8771]='h00000000;  wr_data_rom[ 8771]='h00000000;
    rd_cycle[ 8772] = 1'b0;  wr_cycle[ 8772] = 1'b0;  addr_rom[ 8772]='h00000000;  wr_data_rom[ 8772]='h00000000;
    rd_cycle[ 8773] = 1'b0;  wr_cycle[ 8773] = 1'b0;  addr_rom[ 8773]='h00000000;  wr_data_rom[ 8773]='h00000000;
    rd_cycle[ 8774] = 1'b0;  wr_cycle[ 8774] = 1'b0;  addr_rom[ 8774]='h00000000;  wr_data_rom[ 8774]='h00000000;
    rd_cycle[ 8775] = 1'b0;  wr_cycle[ 8775] = 1'b0;  addr_rom[ 8775]='h00000000;  wr_data_rom[ 8775]='h00000000;
    rd_cycle[ 8776] = 1'b0;  wr_cycle[ 8776] = 1'b0;  addr_rom[ 8776]='h00000000;  wr_data_rom[ 8776]='h00000000;
    rd_cycle[ 8777] = 1'b0;  wr_cycle[ 8777] = 1'b0;  addr_rom[ 8777]='h00000000;  wr_data_rom[ 8777]='h00000000;
    rd_cycle[ 8778] = 1'b0;  wr_cycle[ 8778] = 1'b0;  addr_rom[ 8778]='h00000000;  wr_data_rom[ 8778]='h00000000;
    rd_cycle[ 8779] = 1'b0;  wr_cycle[ 8779] = 1'b0;  addr_rom[ 8779]='h00000000;  wr_data_rom[ 8779]='h00000000;
    rd_cycle[ 8780] = 1'b0;  wr_cycle[ 8780] = 1'b0;  addr_rom[ 8780]='h00000000;  wr_data_rom[ 8780]='h00000000;
    rd_cycle[ 8781] = 1'b0;  wr_cycle[ 8781] = 1'b0;  addr_rom[ 8781]='h00000000;  wr_data_rom[ 8781]='h00000000;
    rd_cycle[ 8782] = 1'b0;  wr_cycle[ 8782] = 1'b0;  addr_rom[ 8782]='h00000000;  wr_data_rom[ 8782]='h00000000;
    rd_cycle[ 8783] = 1'b0;  wr_cycle[ 8783] = 1'b0;  addr_rom[ 8783]='h00000000;  wr_data_rom[ 8783]='h00000000;
    rd_cycle[ 8784] = 1'b0;  wr_cycle[ 8784] = 1'b0;  addr_rom[ 8784]='h00000000;  wr_data_rom[ 8784]='h00000000;
    rd_cycle[ 8785] = 1'b0;  wr_cycle[ 8785] = 1'b0;  addr_rom[ 8785]='h00000000;  wr_data_rom[ 8785]='h00000000;
    rd_cycle[ 8786] = 1'b0;  wr_cycle[ 8786] = 1'b0;  addr_rom[ 8786]='h00000000;  wr_data_rom[ 8786]='h00000000;
    rd_cycle[ 8787] = 1'b0;  wr_cycle[ 8787] = 1'b0;  addr_rom[ 8787]='h00000000;  wr_data_rom[ 8787]='h00000000;
    rd_cycle[ 8788] = 1'b0;  wr_cycle[ 8788] = 1'b0;  addr_rom[ 8788]='h00000000;  wr_data_rom[ 8788]='h00000000;
    rd_cycle[ 8789] = 1'b0;  wr_cycle[ 8789] = 1'b0;  addr_rom[ 8789]='h00000000;  wr_data_rom[ 8789]='h00000000;
    rd_cycle[ 8790] = 1'b0;  wr_cycle[ 8790] = 1'b0;  addr_rom[ 8790]='h00000000;  wr_data_rom[ 8790]='h00000000;
    rd_cycle[ 8791] = 1'b0;  wr_cycle[ 8791] = 1'b0;  addr_rom[ 8791]='h00000000;  wr_data_rom[ 8791]='h00000000;
    rd_cycle[ 8792] = 1'b0;  wr_cycle[ 8792] = 1'b0;  addr_rom[ 8792]='h00000000;  wr_data_rom[ 8792]='h00000000;
    rd_cycle[ 8793] = 1'b0;  wr_cycle[ 8793] = 1'b0;  addr_rom[ 8793]='h00000000;  wr_data_rom[ 8793]='h00000000;
    rd_cycle[ 8794] = 1'b0;  wr_cycle[ 8794] = 1'b0;  addr_rom[ 8794]='h00000000;  wr_data_rom[ 8794]='h00000000;
    rd_cycle[ 8795] = 1'b0;  wr_cycle[ 8795] = 1'b0;  addr_rom[ 8795]='h00000000;  wr_data_rom[ 8795]='h00000000;
    rd_cycle[ 8796] = 1'b0;  wr_cycle[ 8796] = 1'b0;  addr_rom[ 8796]='h00000000;  wr_data_rom[ 8796]='h00000000;
    rd_cycle[ 8797] = 1'b0;  wr_cycle[ 8797] = 1'b0;  addr_rom[ 8797]='h00000000;  wr_data_rom[ 8797]='h00000000;
    rd_cycle[ 8798] = 1'b0;  wr_cycle[ 8798] = 1'b0;  addr_rom[ 8798]='h00000000;  wr_data_rom[ 8798]='h00000000;
    rd_cycle[ 8799] = 1'b0;  wr_cycle[ 8799] = 1'b0;  addr_rom[ 8799]='h00000000;  wr_data_rom[ 8799]='h00000000;
    rd_cycle[ 8800] = 1'b0;  wr_cycle[ 8800] = 1'b0;  addr_rom[ 8800]='h00000000;  wr_data_rom[ 8800]='h00000000;
    rd_cycle[ 8801] = 1'b0;  wr_cycle[ 8801] = 1'b0;  addr_rom[ 8801]='h00000000;  wr_data_rom[ 8801]='h00000000;
    rd_cycle[ 8802] = 1'b0;  wr_cycle[ 8802] = 1'b0;  addr_rom[ 8802]='h00000000;  wr_data_rom[ 8802]='h00000000;
    rd_cycle[ 8803] = 1'b0;  wr_cycle[ 8803] = 1'b0;  addr_rom[ 8803]='h00000000;  wr_data_rom[ 8803]='h00000000;
    rd_cycle[ 8804] = 1'b0;  wr_cycle[ 8804] = 1'b0;  addr_rom[ 8804]='h00000000;  wr_data_rom[ 8804]='h00000000;
    rd_cycle[ 8805] = 1'b0;  wr_cycle[ 8805] = 1'b0;  addr_rom[ 8805]='h00000000;  wr_data_rom[ 8805]='h00000000;
    rd_cycle[ 8806] = 1'b0;  wr_cycle[ 8806] = 1'b0;  addr_rom[ 8806]='h00000000;  wr_data_rom[ 8806]='h00000000;
    rd_cycle[ 8807] = 1'b0;  wr_cycle[ 8807] = 1'b0;  addr_rom[ 8807]='h00000000;  wr_data_rom[ 8807]='h00000000;
    rd_cycle[ 8808] = 1'b0;  wr_cycle[ 8808] = 1'b0;  addr_rom[ 8808]='h00000000;  wr_data_rom[ 8808]='h00000000;
    rd_cycle[ 8809] = 1'b0;  wr_cycle[ 8809] = 1'b0;  addr_rom[ 8809]='h00000000;  wr_data_rom[ 8809]='h00000000;
    rd_cycle[ 8810] = 1'b0;  wr_cycle[ 8810] = 1'b0;  addr_rom[ 8810]='h00000000;  wr_data_rom[ 8810]='h00000000;
    rd_cycle[ 8811] = 1'b0;  wr_cycle[ 8811] = 1'b0;  addr_rom[ 8811]='h00000000;  wr_data_rom[ 8811]='h00000000;
    rd_cycle[ 8812] = 1'b0;  wr_cycle[ 8812] = 1'b0;  addr_rom[ 8812]='h00000000;  wr_data_rom[ 8812]='h00000000;
    rd_cycle[ 8813] = 1'b0;  wr_cycle[ 8813] = 1'b0;  addr_rom[ 8813]='h00000000;  wr_data_rom[ 8813]='h00000000;
    rd_cycle[ 8814] = 1'b0;  wr_cycle[ 8814] = 1'b0;  addr_rom[ 8814]='h00000000;  wr_data_rom[ 8814]='h00000000;
    rd_cycle[ 8815] = 1'b0;  wr_cycle[ 8815] = 1'b0;  addr_rom[ 8815]='h00000000;  wr_data_rom[ 8815]='h00000000;
    rd_cycle[ 8816] = 1'b0;  wr_cycle[ 8816] = 1'b0;  addr_rom[ 8816]='h00000000;  wr_data_rom[ 8816]='h00000000;
    rd_cycle[ 8817] = 1'b0;  wr_cycle[ 8817] = 1'b0;  addr_rom[ 8817]='h00000000;  wr_data_rom[ 8817]='h00000000;
    rd_cycle[ 8818] = 1'b0;  wr_cycle[ 8818] = 1'b0;  addr_rom[ 8818]='h00000000;  wr_data_rom[ 8818]='h00000000;
    rd_cycle[ 8819] = 1'b0;  wr_cycle[ 8819] = 1'b0;  addr_rom[ 8819]='h00000000;  wr_data_rom[ 8819]='h00000000;
    rd_cycle[ 8820] = 1'b0;  wr_cycle[ 8820] = 1'b0;  addr_rom[ 8820]='h00000000;  wr_data_rom[ 8820]='h00000000;
    rd_cycle[ 8821] = 1'b0;  wr_cycle[ 8821] = 1'b0;  addr_rom[ 8821]='h00000000;  wr_data_rom[ 8821]='h00000000;
    rd_cycle[ 8822] = 1'b0;  wr_cycle[ 8822] = 1'b0;  addr_rom[ 8822]='h00000000;  wr_data_rom[ 8822]='h00000000;
    rd_cycle[ 8823] = 1'b0;  wr_cycle[ 8823] = 1'b0;  addr_rom[ 8823]='h00000000;  wr_data_rom[ 8823]='h00000000;
    rd_cycle[ 8824] = 1'b0;  wr_cycle[ 8824] = 1'b0;  addr_rom[ 8824]='h00000000;  wr_data_rom[ 8824]='h00000000;
    rd_cycle[ 8825] = 1'b0;  wr_cycle[ 8825] = 1'b0;  addr_rom[ 8825]='h00000000;  wr_data_rom[ 8825]='h00000000;
    rd_cycle[ 8826] = 1'b0;  wr_cycle[ 8826] = 1'b0;  addr_rom[ 8826]='h00000000;  wr_data_rom[ 8826]='h00000000;
    rd_cycle[ 8827] = 1'b0;  wr_cycle[ 8827] = 1'b0;  addr_rom[ 8827]='h00000000;  wr_data_rom[ 8827]='h00000000;
    rd_cycle[ 8828] = 1'b0;  wr_cycle[ 8828] = 1'b0;  addr_rom[ 8828]='h00000000;  wr_data_rom[ 8828]='h00000000;
    rd_cycle[ 8829] = 1'b0;  wr_cycle[ 8829] = 1'b0;  addr_rom[ 8829]='h00000000;  wr_data_rom[ 8829]='h00000000;
    rd_cycle[ 8830] = 1'b0;  wr_cycle[ 8830] = 1'b0;  addr_rom[ 8830]='h00000000;  wr_data_rom[ 8830]='h00000000;
    rd_cycle[ 8831] = 1'b0;  wr_cycle[ 8831] = 1'b0;  addr_rom[ 8831]='h00000000;  wr_data_rom[ 8831]='h00000000;
    rd_cycle[ 8832] = 1'b0;  wr_cycle[ 8832] = 1'b0;  addr_rom[ 8832]='h00000000;  wr_data_rom[ 8832]='h00000000;
    rd_cycle[ 8833] = 1'b0;  wr_cycle[ 8833] = 1'b0;  addr_rom[ 8833]='h00000000;  wr_data_rom[ 8833]='h00000000;
    rd_cycle[ 8834] = 1'b0;  wr_cycle[ 8834] = 1'b0;  addr_rom[ 8834]='h00000000;  wr_data_rom[ 8834]='h00000000;
    rd_cycle[ 8835] = 1'b0;  wr_cycle[ 8835] = 1'b0;  addr_rom[ 8835]='h00000000;  wr_data_rom[ 8835]='h00000000;
    rd_cycle[ 8836] = 1'b0;  wr_cycle[ 8836] = 1'b0;  addr_rom[ 8836]='h00000000;  wr_data_rom[ 8836]='h00000000;
    rd_cycle[ 8837] = 1'b0;  wr_cycle[ 8837] = 1'b0;  addr_rom[ 8837]='h00000000;  wr_data_rom[ 8837]='h00000000;
    rd_cycle[ 8838] = 1'b0;  wr_cycle[ 8838] = 1'b0;  addr_rom[ 8838]='h00000000;  wr_data_rom[ 8838]='h00000000;
    rd_cycle[ 8839] = 1'b0;  wr_cycle[ 8839] = 1'b0;  addr_rom[ 8839]='h00000000;  wr_data_rom[ 8839]='h00000000;
    rd_cycle[ 8840] = 1'b0;  wr_cycle[ 8840] = 1'b0;  addr_rom[ 8840]='h00000000;  wr_data_rom[ 8840]='h00000000;
    rd_cycle[ 8841] = 1'b0;  wr_cycle[ 8841] = 1'b0;  addr_rom[ 8841]='h00000000;  wr_data_rom[ 8841]='h00000000;
    rd_cycle[ 8842] = 1'b0;  wr_cycle[ 8842] = 1'b0;  addr_rom[ 8842]='h00000000;  wr_data_rom[ 8842]='h00000000;
    rd_cycle[ 8843] = 1'b0;  wr_cycle[ 8843] = 1'b0;  addr_rom[ 8843]='h00000000;  wr_data_rom[ 8843]='h00000000;
    rd_cycle[ 8844] = 1'b0;  wr_cycle[ 8844] = 1'b0;  addr_rom[ 8844]='h00000000;  wr_data_rom[ 8844]='h00000000;
    rd_cycle[ 8845] = 1'b0;  wr_cycle[ 8845] = 1'b0;  addr_rom[ 8845]='h00000000;  wr_data_rom[ 8845]='h00000000;
    rd_cycle[ 8846] = 1'b0;  wr_cycle[ 8846] = 1'b0;  addr_rom[ 8846]='h00000000;  wr_data_rom[ 8846]='h00000000;
    rd_cycle[ 8847] = 1'b0;  wr_cycle[ 8847] = 1'b0;  addr_rom[ 8847]='h00000000;  wr_data_rom[ 8847]='h00000000;
    rd_cycle[ 8848] = 1'b0;  wr_cycle[ 8848] = 1'b0;  addr_rom[ 8848]='h00000000;  wr_data_rom[ 8848]='h00000000;
    rd_cycle[ 8849] = 1'b0;  wr_cycle[ 8849] = 1'b0;  addr_rom[ 8849]='h00000000;  wr_data_rom[ 8849]='h00000000;
    rd_cycle[ 8850] = 1'b0;  wr_cycle[ 8850] = 1'b0;  addr_rom[ 8850]='h00000000;  wr_data_rom[ 8850]='h00000000;
    rd_cycle[ 8851] = 1'b0;  wr_cycle[ 8851] = 1'b0;  addr_rom[ 8851]='h00000000;  wr_data_rom[ 8851]='h00000000;
    rd_cycle[ 8852] = 1'b0;  wr_cycle[ 8852] = 1'b0;  addr_rom[ 8852]='h00000000;  wr_data_rom[ 8852]='h00000000;
    rd_cycle[ 8853] = 1'b0;  wr_cycle[ 8853] = 1'b0;  addr_rom[ 8853]='h00000000;  wr_data_rom[ 8853]='h00000000;
    rd_cycle[ 8854] = 1'b0;  wr_cycle[ 8854] = 1'b0;  addr_rom[ 8854]='h00000000;  wr_data_rom[ 8854]='h00000000;
    rd_cycle[ 8855] = 1'b0;  wr_cycle[ 8855] = 1'b0;  addr_rom[ 8855]='h00000000;  wr_data_rom[ 8855]='h00000000;
    rd_cycle[ 8856] = 1'b0;  wr_cycle[ 8856] = 1'b0;  addr_rom[ 8856]='h00000000;  wr_data_rom[ 8856]='h00000000;
    rd_cycle[ 8857] = 1'b0;  wr_cycle[ 8857] = 1'b0;  addr_rom[ 8857]='h00000000;  wr_data_rom[ 8857]='h00000000;
    rd_cycle[ 8858] = 1'b0;  wr_cycle[ 8858] = 1'b0;  addr_rom[ 8858]='h00000000;  wr_data_rom[ 8858]='h00000000;
    rd_cycle[ 8859] = 1'b0;  wr_cycle[ 8859] = 1'b0;  addr_rom[ 8859]='h00000000;  wr_data_rom[ 8859]='h00000000;
    rd_cycle[ 8860] = 1'b0;  wr_cycle[ 8860] = 1'b0;  addr_rom[ 8860]='h00000000;  wr_data_rom[ 8860]='h00000000;
    rd_cycle[ 8861] = 1'b0;  wr_cycle[ 8861] = 1'b0;  addr_rom[ 8861]='h00000000;  wr_data_rom[ 8861]='h00000000;
    rd_cycle[ 8862] = 1'b0;  wr_cycle[ 8862] = 1'b0;  addr_rom[ 8862]='h00000000;  wr_data_rom[ 8862]='h00000000;
    rd_cycle[ 8863] = 1'b0;  wr_cycle[ 8863] = 1'b0;  addr_rom[ 8863]='h00000000;  wr_data_rom[ 8863]='h00000000;
    rd_cycle[ 8864] = 1'b0;  wr_cycle[ 8864] = 1'b0;  addr_rom[ 8864]='h00000000;  wr_data_rom[ 8864]='h00000000;
    rd_cycle[ 8865] = 1'b0;  wr_cycle[ 8865] = 1'b0;  addr_rom[ 8865]='h00000000;  wr_data_rom[ 8865]='h00000000;
    rd_cycle[ 8866] = 1'b0;  wr_cycle[ 8866] = 1'b0;  addr_rom[ 8866]='h00000000;  wr_data_rom[ 8866]='h00000000;
    rd_cycle[ 8867] = 1'b0;  wr_cycle[ 8867] = 1'b0;  addr_rom[ 8867]='h00000000;  wr_data_rom[ 8867]='h00000000;
    rd_cycle[ 8868] = 1'b0;  wr_cycle[ 8868] = 1'b0;  addr_rom[ 8868]='h00000000;  wr_data_rom[ 8868]='h00000000;
    rd_cycle[ 8869] = 1'b0;  wr_cycle[ 8869] = 1'b0;  addr_rom[ 8869]='h00000000;  wr_data_rom[ 8869]='h00000000;
    rd_cycle[ 8870] = 1'b0;  wr_cycle[ 8870] = 1'b0;  addr_rom[ 8870]='h00000000;  wr_data_rom[ 8870]='h00000000;
    rd_cycle[ 8871] = 1'b0;  wr_cycle[ 8871] = 1'b0;  addr_rom[ 8871]='h00000000;  wr_data_rom[ 8871]='h00000000;
    rd_cycle[ 8872] = 1'b0;  wr_cycle[ 8872] = 1'b0;  addr_rom[ 8872]='h00000000;  wr_data_rom[ 8872]='h00000000;
    rd_cycle[ 8873] = 1'b0;  wr_cycle[ 8873] = 1'b0;  addr_rom[ 8873]='h00000000;  wr_data_rom[ 8873]='h00000000;
    rd_cycle[ 8874] = 1'b0;  wr_cycle[ 8874] = 1'b0;  addr_rom[ 8874]='h00000000;  wr_data_rom[ 8874]='h00000000;
    rd_cycle[ 8875] = 1'b0;  wr_cycle[ 8875] = 1'b0;  addr_rom[ 8875]='h00000000;  wr_data_rom[ 8875]='h00000000;
    rd_cycle[ 8876] = 1'b0;  wr_cycle[ 8876] = 1'b0;  addr_rom[ 8876]='h00000000;  wr_data_rom[ 8876]='h00000000;
    rd_cycle[ 8877] = 1'b0;  wr_cycle[ 8877] = 1'b0;  addr_rom[ 8877]='h00000000;  wr_data_rom[ 8877]='h00000000;
    rd_cycle[ 8878] = 1'b0;  wr_cycle[ 8878] = 1'b0;  addr_rom[ 8878]='h00000000;  wr_data_rom[ 8878]='h00000000;
    rd_cycle[ 8879] = 1'b0;  wr_cycle[ 8879] = 1'b0;  addr_rom[ 8879]='h00000000;  wr_data_rom[ 8879]='h00000000;
    rd_cycle[ 8880] = 1'b0;  wr_cycle[ 8880] = 1'b0;  addr_rom[ 8880]='h00000000;  wr_data_rom[ 8880]='h00000000;
    rd_cycle[ 8881] = 1'b0;  wr_cycle[ 8881] = 1'b0;  addr_rom[ 8881]='h00000000;  wr_data_rom[ 8881]='h00000000;
    rd_cycle[ 8882] = 1'b0;  wr_cycle[ 8882] = 1'b0;  addr_rom[ 8882]='h00000000;  wr_data_rom[ 8882]='h00000000;
    rd_cycle[ 8883] = 1'b0;  wr_cycle[ 8883] = 1'b0;  addr_rom[ 8883]='h00000000;  wr_data_rom[ 8883]='h00000000;
    rd_cycle[ 8884] = 1'b0;  wr_cycle[ 8884] = 1'b0;  addr_rom[ 8884]='h00000000;  wr_data_rom[ 8884]='h00000000;
    rd_cycle[ 8885] = 1'b0;  wr_cycle[ 8885] = 1'b0;  addr_rom[ 8885]='h00000000;  wr_data_rom[ 8885]='h00000000;
    rd_cycle[ 8886] = 1'b0;  wr_cycle[ 8886] = 1'b0;  addr_rom[ 8886]='h00000000;  wr_data_rom[ 8886]='h00000000;
    rd_cycle[ 8887] = 1'b0;  wr_cycle[ 8887] = 1'b0;  addr_rom[ 8887]='h00000000;  wr_data_rom[ 8887]='h00000000;
    rd_cycle[ 8888] = 1'b0;  wr_cycle[ 8888] = 1'b0;  addr_rom[ 8888]='h00000000;  wr_data_rom[ 8888]='h00000000;
    rd_cycle[ 8889] = 1'b0;  wr_cycle[ 8889] = 1'b0;  addr_rom[ 8889]='h00000000;  wr_data_rom[ 8889]='h00000000;
    rd_cycle[ 8890] = 1'b0;  wr_cycle[ 8890] = 1'b0;  addr_rom[ 8890]='h00000000;  wr_data_rom[ 8890]='h00000000;
    rd_cycle[ 8891] = 1'b0;  wr_cycle[ 8891] = 1'b0;  addr_rom[ 8891]='h00000000;  wr_data_rom[ 8891]='h00000000;
    rd_cycle[ 8892] = 1'b0;  wr_cycle[ 8892] = 1'b0;  addr_rom[ 8892]='h00000000;  wr_data_rom[ 8892]='h00000000;
    rd_cycle[ 8893] = 1'b0;  wr_cycle[ 8893] = 1'b0;  addr_rom[ 8893]='h00000000;  wr_data_rom[ 8893]='h00000000;
    rd_cycle[ 8894] = 1'b0;  wr_cycle[ 8894] = 1'b0;  addr_rom[ 8894]='h00000000;  wr_data_rom[ 8894]='h00000000;
    rd_cycle[ 8895] = 1'b0;  wr_cycle[ 8895] = 1'b0;  addr_rom[ 8895]='h00000000;  wr_data_rom[ 8895]='h00000000;
    rd_cycle[ 8896] = 1'b0;  wr_cycle[ 8896] = 1'b0;  addr_rom[ 8896]='h00000000;  wr_data_rom[ 8896]='h00000000;
    rd_cycle[ 8897] = 1'b0;  wr_cycle[ 8897] = 1'b0;  addr_rom[ 8897]='h00000000;  wr_data_rom[ 8897]='h00000000;
    rd_cycle[ 8898] = 1'b0;  wr_cycle[ 8898] = 1'b0;  addr_rom[ 8898]='h00000000;  wr_data_rom[ 8898]='h00000000;
    rd_cycle[ 8899] = 1'b0;  wr_cycle[ 8899] = 1'b0;  addr_rom[ 8899]='h00000000;  wr_data_rom[ 8899]='h00000000;
    rd_cycle[ 8900] = 1'b0;  wr_cycle[ 8900] = 1'b0;  addr_rom[ 8900]='h00000000;  wr_data_rom[ 8900]='h00000000;
    rd_cycle[ 8901] = 1'b0;  wr_cycle[ 8901] = 1'b0;  addr_rom[ 8901]='h00000000;  wr_data_rom[ 8901]='h00000000;
    rd_cycle[ 8902] = 1'b0;  wr_cycle[ 8902] = 1'b0;  addr_rom[ 8902]='h00000000;  wr_data_rom[ 8902]='h00000000;
    rd_cycle[ 8903] = 1'b0;  wr_cycle[ 8903] = 1'b0;  addr_rom[ 8903]='h00000000;  wr_data_rom[ 8903]='h00000000;
    rd_cycle[ 8904] = 1'b0;  wr_cycle[ 8904] = 1'b0;  addr_rom[ 8904]='h00000000;  wr_data_rom[ 8904]='h00000000;
    rd_cycle[ 8905] = 1'b0;  wr_cycle[ 8905] = 1'b0;  addr_rom[ 8905]='h00000000;  wr_data_rom[ 8905]='h00000000;
    rd_cycle[ 8906] = 1'b0;  wr_cycle[ 8906] = 1'b0;  addr_rom[ 8906]='h00000000;  wr_data_rom[ 8906]='h00000000;
    rd_cycle[ 8907] = 1'b0;  wr_cycle[ 8907] = 1'b0;  addr_rom[ 8907]='h00000000;  wr_data_rom[ 8907]='h00000000;
    rd_cycle[ 8908] = 1'b0;  wr_cycle[ 8908] = 1'b0;  addr_rom[ 8908]='h00000000;  wr_data_rom[ 8908]='h00000000;
    rd_cycle[ 8909] = 1'b0;  wr_cycle[ 8909] = 1'b0;  addr_rom[ 8909]='h00000000;  wr_data_rom[ 8909]='h00000000;
    rd_cycle[ 8910] = 1'b0;  wr_cycle[ 8910] = 1'b0;  addr_rom[ 8910]='h00000000;  wr_data_rom[ 8910]='h00000000;
    rd_cycle[ 8911] = 1'b0;  wr_cycle[ 8911] = 1'b0;  addr_rom[ 8911]='h00000000;  wr_data_rom[ 8911]='h00000000;
    rd_cycle[ 8912] = 1'b0;  wr_cycle[ 8912] = 1'b0;  addr_rom[ 8912]='h00000000;  wr_data_rom[ 8912]='h00000000;
    rd_cycle[ 8913] = 1'b0;  wr_cycle[ 8913] = 1'b0;  addr_rom[ 8913]='h00000000;  wr_data_rom[ 8913]='h00000000;
    rd_cycle[ 8914] = 1'b0;  wr_cycle[ 8914] = 1'b0;  addr_rom[ 8914]='h00000000;  wr_data_rom[ 8914]='h00000000;
    rd_cycle[ 8915] = 1'b0;  wr_cycle[ 8915] = 1'b0;  addr_rom[ 8915]='h00000000;  wr_data_rom[ 8915]='h00000000;
    rd_cycle[ 8916] = 1'b0;  wr_cycle[ 8916] = 1'b0;  addr_rom[ 8916]='h00000000;  wr_data_rom[ 8916]='h00000000;
    rd_cycle[ 8917] = 1'b0;  wr_cycle[ 8917] = 1'b0;  addr_rom[ 8917]='h00000000;  wr_data_rom[ 8917]='h00000000;
    rd_cycle[ 8918] = 1'b0;  wr_cycle[ 8918] = 1'b0;  addr_rom[ 8918]='h00000000;  wr_data_rom[ 8918]='h00000000;
    rd_cycle[ 8919] = 1'b0;  wr_cycle[ 8919] = 1'b0;  addr_rom[ 8919]='h00000000;  wr_data_rom[ 8919]='h00000000;
    rd_cycle[ 8920] = 1'b0;  wr_cycle[ 8920] = 1'b0;  addr_rom[ 8920]='h00000000;  wr_data_rom[ 8920]='h00000000;
    rd_cycle[ 8921] = 1'b0;  wr_cycle[ 8921] = 1'b0;  addr_rom[ 8921]='h00000000;  wr_data_rom[ 8921]='h00000000;
    rd_cycle[ 8922] = 1'b0;  wr_cycle[ 8922] = 1'b0;  addr_rom[ 8922]='h00000000;  wr_data_rom[ 8922]='h00000000;
    rd_cycle[ 8923] = 1'b0;  wr_cycle[ 8923] = 1'b0;  addr_rom[ 8923]='h00000000;  wr_data_rom[ 8923]='h00000000;
    rd_cycle[ 8924] = 1'b0;  wr_cycle[ 8924] = 1'b0;  addr_rom[ 8924]='h00000000;  wr_data_rom[ 8924]='h00000000;
    rd_cycle[ 8925] = 1'b0;  wr_cycle[ 8925] = 1'b0;  addr_rom[ 8925]='h00000000;  wr_data_rom[ 8925]='h00000000;
    rd_cycle[ 8926] = 1'b0;  wr_cycle[ 8926] = 1'b0;  addr_rom[ 8926]='h00000000;  wr_data_rom[ 8926]='h00000000;
    rd_cycle[ 8927] = 1'b0;  wr_cycle[ 8927] = 1'b0;  addr_rom[ 8927]='h00000000;  wr_data_rom[ 8927]='h00000000;
    rd_cycle[ 8928] = 1'b0;  wr_cycle[ 8928] = 1'b0;  addr_rom[ 8928]='h00000000;  wr_data_rom[ 8928]='h00000000;
    rd_cycle[ 8929] = 1'b0;  wr_cycle[ 8929] = 1'b0;  addr_rom[ 8929]='h00000000;  wr_data_rom[ 8929]='h00000000;
    rd_cycle[ 8930] = 1'b0;  wr_cycle[ 8930] = 1'b0;  addr_rom[ 8930]='h00000000;  wr_data_rom[ 8930]='h00000000;
    rd_cycle[ 8931] = 1'b0;  wr_cycle[ 8931] = 1'b0;  addr_rom[ 8931]='h00000000;  wr_data_rom[ 8931]='h00000000;
    rd_cycle[ 8932] = 1'b0;  wr_cycle[ 8932] = 1'b0;  addr_rom[ 8932]='h00000000;  wr_data_rom[ 8932]='h00000000;
    rd_cycle[ 8933] = 1'b0;  wr_cycle[ 8933] = 1'b0;  addr_rom[ 8933]='h00000000;  wr_data_rom[ 8933]='h00000000;
    rd_cycle[ 8934] = 1'b0;  wr_cycle[ 8934] = 1'b0;  addr_rom[ 8934]='h00000000;  wr_data_rom[ 8934]='h00000000;
    rd_cycle[ 8935] = 1'b0;  wr_cycle[ 8935] = 1'b0;  addr_rom[ 8935]='h00000000;  wr_data_rom[ 8935]='h00000000;
    rd_cycle[ 8936] = 1'b0;  wr_cycle[ 8936] = 1'b0;  addr_rom[ 8936]='h00000000;  wr_data_rom[ 8936]='h00000000;
    rd_cycle[ 8937] = 1'b0;  wr_cycle[ 8937] = 1'b0;  addr_rom[ 8937]='h00000000;  wr_data_rom[ 8937]='h00000000;
    rd_cycle[ 8938] = 1'b0;  wr_cycle[ 8938] = 1'b0;  addr_rom[ 8938]='h00000000;  wr_data_rom[ 8938]='h00000000;
    rd_cycle[ 8939] = 1'b0;  wr_cycle[ 8939] = 1'b0;  addr_rom[ 8939]='h00000000;  wr_data_rom[ 8939]='h00000000;
    rd_cycle[ 8940] = 1'b0;  wr_cycle[ 8940] = 1'b0;  addr_rom[ 8940]='h00000000;  wr_data_rom[ 8940]='h00000000;
    rd_cycle[ 8941] = 1'b0;  wr_cycle[ 8941] = 1'b0;  addr_rom[ 8941]='h00000000;  wr_data_rom[ 8941]='h00000000;
    rd_cycle[ 8942] = 1'b0;  wr_cycle[ 8942] = 1'b0;  addr_rom[ 8942]='h00000000;  wr_data_rom[ 8942]='h00000000;
    rd_cycle[ 8943] = 1'b0;  wr_cycle[ 8943] = 1'b0;  addr_rom[ 8943]='h00000000;  wr_data_rom[ 8943]='h00000000;
    rd_cycle[ 8944] = 1'b0;  wr_cycle[ 8944] = 1'b0;  addr_rom[ 8944]='h00000000;  wr_data_rom[ 8944]='h00000000;
    rd_cycle[ 8945] = 1'b0;  wr_cycle[ 8945] = 1'b0;  addr_rom[ 8945]='h00000000;  wr_data_rom[ 8945]='h00000000;
    rd_cycle[ 8946] = 1'b0;  wr_cycle[ 8946] = 1'b0;  addr_rom[ 8946]='h00000000;  wr_data_rom[ 8946]='h00000000;
    rd_cycle[ 8947] = 1'b0;  wr_cycle[ 8947] = 1'b0;  addr_rom[ 8947]='h00000000;  wr_data_rom[ 8947]='h00000000;
    rd_cycle[ 8948] = 1'b0;  wr_cycle[ 8948] = 1'b0;  addr_rom[ 8948]='h00000000;  wr_data_rom[ 8948]='h00000000;
    rd_cycle[ 8949] = 1'b0;  wr_cycle[ 8949] = 1'b0;  addr_rom[ 8949]='h00000000;  wr_data_rom[ 8949]='h00000000;
    rd_cycle[ 8950] = 1'b0;  wr_cycle[ 8950] = 1'b0;  addr_rom[ 8950]='h00000000;  wr_data_rom[ 8950]='h00000000;
    rd_cycle[ 8951] = 1'b0;  wr_cycle[ 8951] = 1'b0;  addr_rom[ 8951]='h00000000;  wr_data_rom[ 8951]='h00000000;
    rd_cycle[ 8952] = 1'b0;  wr_cycle[ 8952] = 1'b0;  addr_rom[ 8952]='h00000000;  wr_data_rom[ 8952]='h00000000;
    rd_cycle[ 8953] = 1'b0;  wr_cycle[ 8953] = 1'b0;  addr_rom[ 8953]='h00000000;  wr_data_rom[ 8953]='h00000000;
    rd_cycle[ 8954] = 1'b0;  wr_cycle[ 8954] = 1'b0;  addr_rom[ 8954]='h00000000;  wr_data_rom[ 8954]='h00000000;
    rd_cycle[ 8955] = 1'b0;  wr_cycle[ 8955] = 1'b0;  addr_rom[ 8955]='h00000000;  wr_data_rom[ 8955]='h00000000;
    rd_cycle[ 8956] = 1'b0;  wr_cycle[ 8956] = 1'b0;  addr_rom[ 8956]='h00000000;  wr_data_rom[ 8956]='h00000000;
    rd_cycle[ 8957] = 1'b0;  wr_cycle[ 8957] = 1'b0;  addr_rom[ 8957]='h00000000;  wr_data_rom[ 8957]='h00000000;
    rd_cycle[ 8958] = 1'b0;  wr_cycle[ 8958] = 1'b0;  addr_rom[ 8958]='h00000000;  wr_data_rom[ 8958]='h00000000;
    rd_cycle[ 8959] = 1'b0;  wr_cycle[ 8959] = 1'b0;  addr_rom[ 8959]='h00000000;  wr_data_rom[ 8959]='h00000000;
    rd_cycle[ 8960] = 1'b0;  wr_cycle[ 8960] = 1'b0;  addr_rom[ 8960]='h00000000;  wr_data_rom[ 8960]='h00000000;
    rd_cycle[ 8961] = 1'b0;  wr_cycle[ 8961] = 1'b0;  addr_rom[ 8961]='h00000000;  wr_data_rom[ 8961]='h00000000;
    rd_cycle[ 8962] = 1'b0;  wr_cycle[ 8962] = 1'b0;  addr_rom[ 8962]='h00000000;  wr_data_rom[ 8962]='h00000000;
    rd_cycle[ 8963] = 1'b0;  wr_cycle[ 8963] = 1'b0;  addr_rom[ 8963]='h00000000;  wr_data_rom[ 8963]='h00000000;
    rd_cycle[ 8964] = 1'b0;  wr_cycle[ 8964] = 1'b0;  addr_rom[ 8964]='h00000000;  wr_data_rom[ 8964]='h00000000;
    rd_cycle[ 8965] = 1'b0;  wr_cycle[ 8965] = 1'b0;  addr_rom[ 8965]='h00000000;  wr_data_rom[ 8965]='h00000000;
    rd_cycle[ 8966] = 1'b0;  wr_cycle[ 8966] = 1'b0;  addr_rom[ 8966]='h00000000;  wr_data_rom[ 8966]='h00000000;
    rd_cycle[ 8967] = 1'b0;  wr_cycle[ 8967] = 1'b0;  addr_rom[ 8967]='h00000000;  wr_data_rom[ 8967]='h00000000;
    rd_cycle[ 8968] = 1'b0;  wr_cycle[ 8968] = 1'b0;  addr_rom[ 8968]='h00000000;  wr_data_rom[ 8968]='h00000000;
    rd_cycle[ 8969] = 1'b0;  wr_cycle[ 8969] = 1'b0;  addr_rom[ 8969]='h00000000;  wr_data_rom[ 8969]='h00000000;
    rd_cycle[ 8970] = 1'b0;  wr_cycle[ 8970] = 1'b0;  addr_rom[ 8970]='h00000000;  wr_data_rom[ 8970]='h00000000;
    rd_cycle[ 8971] = 1'b0;  wr_cycle[ 8971] = 1'b0;  addr_rom[ 8971]='h00000000;  wr_data_rom[ 8971]='h00000000;
    rd_cycle[ 8972] = 1'b0;  wr_cycle[ 8972] = 1'b0;  addr_rom[ 8972]='h00000000;  wr_data_rom[ 8972]='h00000000;
    rd_cycle[ 8973] = 1'b0;  wr_cycle[ 8973] = 1'b0;  addr_rom[ 8973]='h00000000;  wr_data_rom[ 8973]='h00000000;
    rd_cycle[ 8974] = 1'b0;  wr_cycle[ 8974] = 1'b0;  addr_rom[ 8974]='h00000000;  wr_data_rom[ 8974]='h00000000;
    rd_cycle[ 8975] = 1'b0;  wr_cycle[ 8975] = 1'b0;  addr_rom[ 8975]='h00000000;  wr_data_rom[ 8975]='h00000000;
    rd_cycle[ 8976] = 1'b0;  wr_cycle[ 8976] = 1'b0;  addr_rom[ 8976]='h00000000;  wr_data_rom[ 8976]='h00000000;
    rd_cycle[ 8977] = 1'b0;  wr_cycle[ 8977] = 1'b0;  addr_rom[ 8977]='h00000000;  wr_data_rom[ 8977]='h00000000;
    rd_cycle[ 8978] = 1'b0;  wr_cycle[ 8978] = 1'b0;  addr_rom[ 8978]='h00000000;  wr_data_rom[ 8978]='h00000000;
    rd_cycle[ 8979] = 1'b0;  wr_cycle[ 8979] = 1'b0;  addr_rom[ 8979]='h00000000;  wr_data_rom[ 8979]='h00000000;
    rd_cycle[ 8980] = 1'b0;  wr_cycle[ 8980] = 1'b0;  addr_rom[ 8980]='h00000000;  wr_data_rom[ 8980]='h00000000;
    rd_cycle[ 8981] = 1'b0;  wr_cycle[ 8981] = 1'b0;  addr_rom[ 8981]='h00000000;  wr_data_rom[ 8981]='h00000000;
    rd_cycle[ 8982] = 1'b0;  wr_cycle[ 8982] = 1'b0;  addr_rom[ 8982]='h00000000;  wr_data_rom[ 8982]='h00000000;
    rd_cycle[ 8983] = 1'b0;  wr_cycle[ 8983] = 1'b0;  addr_rom[ 8983]='h00000000;  wr_data_rom[ 8983]='h00000000;
    rd_cycle[ 8984] = 1'b0;  wr_cycle[ 8984] = 1'b0;  addr_rom[ 8984]='h00000000;  wr_data_rom[ 8984]='h00000000;
    rd_cycle[ 8985] = 1'b0;  wr_cycle[ 8985] = 1'b0;  addr_rom[ 8985]='h00000000;  wr_data_rom[ 8985]='h00000000;
    rd_cycle[ 8986] = 1'b0;  wr_cycle[ 8986] = 1'b0;  addr_rom[ 8986]='h00000000;  wr_data_rom[ 8986]='h00000000;
    rd_cycle[ 8987] = 1'b0;  wr_cycle[ 8987] = 1'b0;  addr_rom[ 8987]='h00000000;  wr_data_rom[ 8987]='h00000000;
    rd_cycle[ 8988] = 1'b0;  wr_cycle[ 8988] = 1'b0;  addr_rom[ 8988]='h00000000;  wr_data_rom[ 8988]='h00000000;
    rd_cycle[ 8989] = 1'b0;  wr_cycle[ 8989] = 1'b0;  addr_rom[ 8989]='h00000000;  wr_data_rom[ 8989]='h00000000;
    rd_cycle[ 8990] = 1'b0;  wr_cycle[ 8990] = 1'b0;  addr_rom[ 8990]='h00000000;  wr_data_rom[ 8990]='h00000000;
    rd_cycle[ 8991] = 1'b0;  wr_cycle[ 8991] = 1'b0;  addr_rom[ 8991]='h00000000;  wr_data_rom[ 8991]='h00000000;
    rd_cycle[ 8992] = 1'b0;  wr_cycle[ 8992] = 1'b0;  addr_rom[ 8992]='h00000000;  wr_data_rom[ 8992]='h00000000;
    rd_cycle[ 8993] = 1'b0;  wr_cycle[ 8993] = 1'b0;  addr_rom[ 8993]='h00000000;  wr_data_rom[ 8993]='h00000000;
    rd_cycle[ 8994] = 1'b0;  wr_cycle[ 8994] = 1'b0;  addr_rom[ 8994]='h00000000;  wr_data_rom[ 8994]='h00000000;
    rd_cycle[ 8995] = 1'b0;  wr_cycle[ 8995] = 1'b0;  addr_rom[ 8995]='h00000000;  wr_data_rom[ 8995]='h00000000;
    rd_cycle[ 8996] = 1'b0;  wr_cycle[ 8996] = 1'b0;  addr_rom[ 8996]='h00000000;  wr_data_rom[ 8996]='h00000000;
    rd_cycle[ 8997] = 1'b0;  wr_cycle[ 8997] = 1'b0;  addr_rom[ 8997]='h00000000;  wr_data_rom[ 8997]='h00000000;
    rd_cycle[ 8998] = 1'b0;  wr_cycle[ 8998] = 1'b0;  addr_rom[ 8998]='h00000000;  wr_data_rom[ 8998]='h00000000;
    rd_cycle[ 8999] = 1'b0;  wr_cycle[ 8999] = 1'b0;  addr_rom[ 8999]='h00000000;  wr_data_rom[ 8999]='h00000000;
    rd_cycle[ 9000] = 1'b0;  wr_cycle[ 9000] = 1'b0;  addr_rom[ 9000]='h00000000;  wr_data_rom[ 9000]='h00000000;
    rd_cycle[ 9001] = 1'b0;  wr_cycle[ 9001] = 1'b0;  addr_rom[ 9001]='h00000000;  wr_data_rom[ 9001]='h00000000;
    rd_cycle[ 9002] = 1'b0;  wr_cycle[ 9002] = 1'b0;  addr_rom[ 9002]='h00000000;  wr_data_rom[ 9002]='h00000000;
    rd_cycle[ 9003] = 1'b0;  wr_cycle[ 9003] = 1'b0;  addr_rom[ 9003]='h00000000;  wr_data_rom[ 9003]='h00000000;
    rd_cycle[ 9004] = 1'b0;  wr_cycle[ 9004] = 1'b0;  addr_rom[ 9004]='h00000000;  wr_data_rom[ 9004]='h00000000;
    rd_cycle[ 9005] = 1'b0;  wr_cycle[ 9005] = 1'b0;  addr_rom[ 9005]='h00000000;  wr_data_rom[ 9005]='h00000000;
    rd_cycle[ 9006] = 1'b0;  wr_cycle[ 9006] = 1'b0;  addr_rom[ 9006]='h00000000;  wr_data_rom[ 9006]='h00000000;
    rd_cycle[ 9007] = 1'b0;  wr_cycle[ 9007] = 1'b0;  addr_rom[ 9007]='h00000000;  wr_data_rom[ 9007]='h00000000;
    rd_cycle[ 9008] = 1'b0;  wr_cycle[ 9008] = 1'b0;  addr_rom[ 9008]='h00000000;  wr_data_rom[ 9008]='h00000000;
    rd_cycle[ 9009] = 1'b0;  wr_cycle[ 9009] = 1'b0;  addr_rom[ 9009]='h00000000;  wr_data_rom[ 9009]='h00000000;
    rd_cycle[ 9010] = 1'b0;  wr_cycle[ 9010] = 1'b0;  addr_rom[ 9010]='h00000000;  wr_data_rom[ 9010]='h00000000;
    rd_cycle[ 9011] = 1'b0;  wr_cycle[ 9011] = 1'b0;  addr_rom[ 9011]='h00000000;  wr_data_rom[ 9011]='h00000000;
    rd_cycle[ 9012] = 1'b0;  wr_cycle[ 9012] = 1'b0;  addr_rom[ 9012]='h00000000;  wr_data_rom[ 9012]='h00000000;
    rd_cycle[ 9013] = 1'b0;  wr_cycle[ 9013] = 1'b0;  addr_rom[ 9013]='h00000000;  wr_data_rom[ 9013]='h00000000;
    rd_cycle[ 9014] = 1'b0;  wr_cycle[ 9014] = 1'b0;  addr_rom[ 9014]='h00000000;  wr_data_rom[ 9014]='h00000000;
    rd_cycle[ 9015] = 1'b0;  wr_cycle[ 9015] = 1'b0;  addr_rom[ 9015]='h00000000;  wr_data_rom[ 9015]='h00000000;
    rd_cycle[ 9016] = 1'b0;  wr_cycle[ 9016] = 1'b0;  addr_rom[ 9016]='h00000000;  wr_data_rom[ 9016]='h00000000;
    rd_cycle[ 9017] = 1'b0;  wr_cycle[ 9017] = 1'b0;  addr_rom[ 9017]='h00000000;  wr_data_rom[ 9017]='h00000000;
    rd_cycle[ 9018] = 1'b0;  wr_cycle[ 9018] = 1'b0;  addr_rom[ 9018]='h00000000;  wr_data_rom[ 9018]='h00000000;
    rd_cycle[ 9019] = 1'b0;  wr_cycle[ 9019] = 1'b0;  addr_rom[ 9019]='h00000000;  wr_data_rom[ 9019]='h00000000;
    rd_cycle[ 9020] = 1'b0;  wr_cycle[ 9020] = 1'b0;  addr_rom[ 9020]='h00000000;  wr_data_rom[ 9020]='h00000000;
    rd_cycle[ 9021] = 1'b0;  wr_cycle[ 9021] = 1'b0;  addr_rom[ 9021]='h00000000;  wr_data_rom[ 9021]='h00000000;
    rd_cycle[ 9022] = 1'b0;  wr_cycle[ 9022] = 1'b0;  addr_rom[ 9022]='h00000000;  wr_data_rom[ 9022]='h00000000;
    rd_cycle[ 9023] = 1'b0;  wr_cycle[ 9023] = 1'b0;  addr_rom[ 9023]='h00000000;  wr_data_rom[ 9023]='h00000000;
    rd_cycle[ 9024] = 1'b0;  wr_cycle[ 9024] = 1'b0;  addr_rom[ 9024]='h00000000;  wr_data_rom[ 9024]='h00000000;
    rd_cycle[ 9025] = 1'b0;  wr_cycle[ 9025] = 1'b0;  addr_rom[ 9025]='h00000000;  wr_data_rom[ 9025]='h00000000;
    rd_cycle[ 9026] = 1'b0;  wr_cycle[ 9026] = 1'b0;  addr_rom[ 9026]='h00000000;  wr_data_rom[ 9026]='h00000000;
    rd_cycle[ 9027] = 1'b0;  wr_cycle[ 9027] = 1'b0;  addr_rom[ 9027]='h00000000;  wr_data_rom[ 9027]='h00000000;
    rd_cycle[ 9028] = 1'b0;  wr_cycle[ 9028] = 1'b0;  addr_rom[ 9028]='h00000000;  wr_data_rom[ 9028]='h00000000;
    rd_cycle[ 9029] = 1'b0;  wr_cycle[ 9029] = 1'b0;  addr_rom[ 9029]='h00000000;  wr_data_rom[ 9029]='h00000000;
    rd_cycle[ 9030] = 1'b0;  wr_cycle[ 9030] = 1'b0;  addr_rom[ 9030]='h00000000;  wr_data_rom[ 9030]='h00000000;
    rd_cycle[ 9031] = 1'b0;  wr_cycle[ 9031] = 1'b0;  addr_rom[ 9031]='h00000000;  wr_data_rom[ 9031]='h00000000;
    rd_cycle[ 9032] = 1'b0;  wr_cycle[ 9032] = 1'b0;  addr_rom[ 9032]='h00000000;  wr_data_rom[ 9032]='h00000000;
    rd_cycle[ 9033] = 1'b0;  wr_cycle[ 9033] = 1'b0;  addr_rom[ 9033]='h00000000;  wr_data_rom[ 9033]='h00000000;
    rd_cycle[ 9034] = 1'b0;  wr_cycle[ 9034] = 1'b0;  addr_rom[ 9034]='h00000000;  wr_data_rom[ 9034]='h00000000;
    rd_cycle[ 9035] = 1'b0;  wr_cycle[ 9035] = 1'b0;  addr_rom[ 9035]='h00000000;  wr_data_rom[ 9035]='h00000000;
    rd_cycle[ 9036] = 1'b0;  wr_cycle[ 9036] = 1'b0;  addr_rom[ 9036]='h00000000;  wr_data_rom[ 9036]='h00000000;
    rd_cycle[ 9037] = 1'b0;  wr_cycle[ 9037] = 1'b0;  addr_rom[ 9037]='h00000000;  wr_data_rom[ 9037]='h00000000;
    rd_cycle[ 9038] = 1'b0;  wr_cycle[ 9038] = 1'b0;  addr_rom[ 9038]='h00000000;  wr_data_rom[ 9038]='h00000000;
    rd_cycle[ 9039] = 1'b0;  wr_cycle[ 9039] = 1'b0;  addr_rom[ 9039]='h00000000;  wr_data_rom[ 9039]='h00000000;
    rd_cycle[ 9040] = 1'b0;  wr_cycle[ 9040] = 1'b0;  addr_rom[ 9040]='h00000000;  wr_data_rom[ 9040]='h00000000;
    rd_cycle[ 9041] = 1'b0;  wr_cycle[ 9041] = 1'b0;  addr_rom[ 9041]='h00000000;  wr_data_rom[ 9041]='h00000000;
    rd_cycle[ 9042] = 1'b0;  wr_cycle[ 9042] = 1'b0;  addr_rom[ 9042]='h00000000;  wr_data_rom[ 9042]='h00000000;
    rd_cycle[ 9043] = 1'b0;  wr_cycle[ 9043] = 1'b0;  addr_rom[ 9043]='h00000000;  wr_data_rom[ 9043]='h00000000;
    rd_cycle[ 9044] = 1'b0;  wr_cycle[ 9044] = 1'b0;  addr_rom[ 9044]='h00000000;  wr_data_rom[ 9044]='h00000000;
    rd_cycle[ 9045] = 1'b0;  wr_cycle[ 9045] = 1'b0;  addr_rom[ 9045]='h00000000;  wr_data_rom[ 9045]='h00000000;
    rd_cycle[ 9046] = 1'b0;  wr_cycle[ 9046] = 1'b0;  addr_rom[ 9046]='h00000000;  wr_data_rom[ 9046]='h00000000;
    rd_cycle[ 9047] = 1'b0;  wr_cycle[ 9047] = 1'b0;  addr_rom[ 9047]='h00000000;  wr_data_rom[ 9047]='h00000000;
    rd_cycle[ 9048] = 1'b0;  wr_cycle[ 9048] = 1'b0;  addr_rom[ 9048]='h00000000;  wr_data_rom[ 9048]='h00000000;
    rd_cycle[ 9049] = 1'b0;  wr_cycle[ 9049] = 1'b0;  addr_rom[ 9049]='h00000000;  wr_data_rom[ 9049]='h00000000;
    rd_cycle[ 9050] = 1'b0;  wr_cycle[ 9050] = 1'b0;  addr_rom[ 9050]='h00000000;  wr_data_rom[ 9050]='h00000000;
    rd_cycle[ 9051] = 1'b0;  wr_cycle[ 9051] = 1'b0;  addr_rom[ 9051]='h00000000;  wr_data_rom[ 9051]='h00000000;
    rd_cycle[ 9052] = 1'b0;  wr_cycle[ 9052] = 1'b0;  addr_rom[ 9052]='h00000000;  wr_data_rom[ 9052]='h00000000;
    rd_cycle[ 9053] = 1'b0;  wr_cycle[ 9053] = 1'b0;  addr_rom[ 9053]='h00000000;  wr_data_rom[ 9053]='h00000000;
    rd_cycle[ 9054] = 1'b0;  wr_cycle[ 9054] = 1'b0;  addr_rom[ 9054]='h00000000;  wr_data_rom[ 9054]='h00000000;
    rd_cycle[ 9055] = 1'b0;  wr_cycle[ 9055] = 1'b0;  addr_rom[ 9055]='h00000000;  wr_data_rom[ 9055]='h00000000;
    rd_cycle[ 9056] = 1'b0;  wr_cycle[ 9056] = 1'b0;  addr_rom[ 9056]='h00000000;  wr_data_rom[ 9056]='h00000000;
    rd_cycle[ 9057] = 1'b0;  wr_cycle[ 9057] = 1'b0;  addr_rom[ 9057]='h00000000;  wr_data_rom[ 9057]='h00000000;
    rd_cycle[ 9058] = 1'b0;  wr_cycle[ 9058] = 1'b0;  addr_rom[ 9058]='h00000000;  wr_data_rom[ 9058]='h00000000;
    rd_cycle[ 9059] = 1'b0;  wr_cycle[ 9059] = 1'b0;  addr_rom[ 9059]='h00000000;  wr_data_rom[ 9059]='h00000000;
    rd_cycle[ 9060] = 1'b0;  wr_cycle[ 9060] = 1'b0;  addr_rom[ 9060]='h00000000;  wr_data_rom[ 9060]='h00000000;
    rd_cycle[ 9061] = 1'b0;  wr_cycle[ 9061] = 1'b0;  addr_rom[ 9061]='h00000000;  wr_data_rom[ 9061]='h00000000;
    rd_cycle[ 9062] = 1'b0;  wr_cycle[ 9062] = 1'b0;  addr_rom[ 9062]='h00000000;  wr_data_rom[ 9062]='h00000000;
    rd_cycle[ 9063] = 1'b0;  wr_cycle[ 9063] = 1'b0;  addr_rom[ 9063]='h00000000;  wr_data_rom[ 9063]='h00000000;
    rd_cycle[ 9064] = 1'b0;  wr_cycle[ 9064] = 1'b0;  addr_rom[ 9064]='h00000000;  wr_data_rom[ 9064]='h00000000;
    rd_cycle[ 9065] = 1'b0;  wr_cycle[ 9065] = 1'b0;  addr_rom[ 9065]='h00000000;  wr_data_rom[ 9065]='h00000000;
    rd_cycle[ 9066] = 1'b0;  wr_cycle[ 9066] = 1'b0;  addr_rom[ 9066]='h00000000;  wr_data_rom[ 9066]='h00000000;
    rd_cycle[ 9067] = 1'b0;  wr_cycle[ 9067] = 1'b0;  addr_rom[ 9067]='h00000000;  wr_data_rom[ 9067]='h00000000;
    rd_cycle[ 9068] = 1'b0;  wr_cycle[ 9068] = 1'b0;  addr_rom[ 9068]='h00000000;  wr_data_rom[ 9068]='h00000000;
    rd_cycle[ 9069] = 1'b0;  wr_cycle[ 9069] = 1'b0;  addr_rom[ 9069]='h00000000;  wr_data_rom[ 9069]='h00000000;
    rd_cycle[ 9070] = 1'b0;  wr_cycle[ 9070] = 1'b0;  addr_rom[ 9070]='h00000000;  wr_data_rom[ 9070]='h00000000;
    rd_cycle[ 9071] = 1'b0;  wr_cycle[ 9071] = 1'b0;  addr_rom[ 9071]='h00000000;  wr_data_rom[ 9071]='h00000000;
    rd_cycle[ 9072] = 1'b0;  wr_cycle[ 9072] = 1'b0;  addr_rom[ 9072]='h00000000;  wr_data_rom[ 9072]='h00000000;
    rd_cycle[ 9073] = 1'b0;  wr_cycle[ 9073] = 1'b0;  addr_rom[ 9073]='h00000000;  wr_data_rom[ 9073]='h00000000;
    rd_cycle[ 9074] = 1'b0;  wr_cycle[ 9074] = 1'b0;  addr_rom[ 9074]='h00000000;  wr_data_rom[ 9074]='h00000000;
    rd_cycle[ 9075] = 1'b0;  wr_cycle[ 9075] = 1'b0;  addr_rom[ 9075]='h00000000;  wr_data_rom[ 9075]='h00000000;
    rd_cycle[ 9076] = 1'b0;  wr_cycle[ 9076] = 1'b0;  addr_rom[ 9076]='h00000000;  wr_data_rom[ 9076]='h00000000;
    rd_cycle[ 9077] = 1'b0;  wr_cycle[ 9077] = 1'b0;  addr_rom[ 9077]='h00000000;  wr_data_rom[ 9077]='h00000000;
    rd_cycle[ 9078] = 1'b0;  wr_cycle[ 9078] = 1'b0;  addr_rom[ 9078]='h00000000;  wr_data_rom[ 9078]='h00000000;
    rd_cycle[ 9079] = 1'b0;  wr_cycle[ 9079] = 1'b0;  addr_rom[ 9079]='h00000000;  wr_data_rom[ 9079]='h00000000;
    rd_cycle[ 9080] = 1'b0;  wr_cycle[ 9080] = 1'b0;  addr_rom[ 9080]='h00000000;  wr_data_rom[ 9080]='h00000000;
    rd_cycle[ 9081] = 1'b0;  wr_cycle[ 9081] = 1'b0;  addr_rom[ 9081]='h00000000;  wr_data_rom[ 9081]='h00000000;
    rd_cycle[ 9082] = 1'b0;  wr_cycle[ 9082] = 1'b0;  addr_rom[ 9082]='h00000000;  wr_data_rom[ 9082]='h00000000;
    rd_cycle[ 9083] = 1'b0;  wr_cycle[ 9083] = 1'b0;  addr_rom[ 9083]='h00000000;  wr_data_rom[ 9083]='h00000000;
    rd_cycle[ 9084] = 1'b0;  wr_cycle[ 9084] = 1'b0;  addr_rom[ 9084]='h00000000;  wr_data_rom[ 9084]='h00000000;
    rd_cycle[ 9085] = 1'b0;  wr_cycle[ 9085] = 1'b0;  addr_rom[ 9085]='h00000000;  wr_data_rom[ 9085]='h00000000;
    rd_cycle[ 9086] = 1'b0;  wr_cycle[ 9086] = 1'b0;  addr_rom[ 9086]='h00000000;  wr_data_rom[ 9086]='h00000000;
    rd_cycle[ 9087] = 1'b0;  wr_cycle[ 9087] = 1'b0;  addr_rom[ 9087]='h00000000;  wr_data_rom[ 9087]='h00000000;
    rd_cycle[ 9088] = 1'b0;  wr_cycle[ 9088] = 1'b0;  addr_rom[ 9088]='h00000000;  wr_data_rom[ 9088]='h00000000;
    rd_cycle[ 9089] = 1'b0;  wr_cycle[ 9089] = 1'b0;  addr_rom[ 9089]='h00000000;  wr_data_rom[ 9089]='h00000000;
    rd_cycle[ 9090] = 1'b0;  wr_cycle[ 9090] = 1'b0;  addr_rom[ 9090]='h00000000;  wr_data_rom[ 9090]='h00000000;
    rd_cycle[ 9091] = 1'b0;  wr_cycle[ 9091] = 1'b0;  addr_rom[ 9091]='h00000000;  wr_data_rom[ 9091]='h00000000;
    rd_cycle[ 9092] = 1'b0;  wr_cycle[ 9092] = 1'b0;  addr_rom[ 9092]='h00000000;  wr_data_rom[ 9092]='h00000000;
    rd_cycle[ 9093] = 1'b0;  wr_cycle[ 9093] = 1'b0;  addr_rom[ 9093]='h00000000;  wr_data_rom[ 9093]='h00000000;
    rd_cycle[ 9094] = 1'b0;  wr_cycle[ 9094] = 1'b0;  addr_rom[ 9094]='h00000000;  wr_data_rom[ 9094]='h00000000;
    rd_cycle[ 9095] = 1'b0;  wr_cycle[ 9095] = 1'b0;  addr_rom[ 9095]='h00000000;  wr_data_rom[ 9095]='h00000000;
    rd_cycle[ 9096] = 1'b0;  wr_cycle[ 9096] = 1'b0;  addr_rom[ 9096]='h00000000;  wr_data_rom[ 9096]='h00000000;
    rd_cycle[ 9097] = 1'b0;  wr_cycle[ 9097] = 1'b0;  addr_rom[ 9097]='h00000000;  wr_data_rom[ 9097]='h00000000;
    rd_cycle[ 9098] = 1'b0;  wr_cycle[ 9098] = 1'b0;  addr_rom[ 9098]='h00000000;  wr_data_rom[ 9098]='h00000000;
    rd_cycle[ 9099] = 1'b0;  wr_cycle[ 9099] = 1'b0;  addr_rom[ 9099]='h00000000;  wr_data_rom[ 9099]='h00000000;
    rd_cycle[ 9100] = 1'b0;  wr_cycle[ 9100] = 1'b0;  addr_rom[ 9100]='h00000000;  wr_data_rom[ 9100]='h00000000;
    rd_cycle[ 9101] = 1'b0;  wr_cycle[ 9101] = 1'b0;  addr_rom[ 9101]='h00000000;  wr_data_rom[ 9101]='h00000000;
    rd_cycle[ 9102] = 1'b0;  wr_cycle[ 9102] = 1'b0;  addr_rom[ 9102]='h00000000;  wr_data_rom[ 9102]='h00000000;
    rd_cycle[ 9103] = 1'b0;  wr_cycle[ 9103] = 1'b0;  addr_rom[ 9103]='h00000000;  wr_data_rom[ 9103]='h00000000;
    rd_cycle[ 9104] = 1'b0;  wr_cycle[ 9104] = 1'b0;  addr_rom[ 9104]='h00000000;  wr_data_rom[ 9104]='h00000000;
    rd_cycle[ 9105] = 1'b0;  wr_cycle[ 9105] = 1'b0;  addr_rom[ 9105]='h00000000;  wr_data_rom[ 9105]='h00000000;
    rd_cycle[ 9106] = 1'b0;  wr_cycle[ 9106] = 1'b0;  addr_rom[ 9106]='h00000000;  wr_data_rom[ 9106]='h00000000;
    rd_cycle[ 9107] = 1'b0;  wr_cycle[ 9107] = 1'b0;  addr_rom[ 9107]='h00000000;  wr_data_rom[ 9107]='h00000000;
    rd_cycle[ 9108] = 1'b0;  wr_cycle[ 9108] = 1'b0;  addr_rom[ 9108]='h00000000;  wr_data_rom[ 9108]='h00000000;
    rd_cycle[ 9109] = 1'b0;  wr_cycle[ 9109] = 1'b0;  addr_rom[ 9109]='h00000000;  wr_data_rom[ 9109]='h00000000;
    rd_cycle[ 9110] = 1'b0;  wr_cycle[ 9110] = 1'b0;  addr_rom[ 9110]='h00000000;  wr_data_rom[ 9110]='h00000000;
    rd_cycle[ 9111] = 1'b0;  wr_cycle[ 9111] = 1'b0;  addr_rom[ 9111]='h00000000;  wr_data_rom[ 9111]='h00000000;
    rd_cycle[ 9112] = 1'b0;  wr_cycle[ 9112] = 1'b0;  addr_rom[ 9112]='h00000000;  wr_data_rom[ 9112]='h00000000;
    rd_cycle[ 9113] = 1'b0;  wr_cycle[ 9113] = 1'b0;  addr_rom[ 9113]='h00000000;  wr_data_rom[ 9113]='h00000000;
    rd_cycle[ 9114] = 1'b0;  wr_cycle[ 9114] = 1'b0;  addr_rom[ 9114]='h00000000;  wr_data_rom[ 9114]='h00000000;
    rd_cycle[ 9115] = 1'b0;  wr_cycle[ 9115] = 1'b0;  addr_rom[ 9115]='h00000000;  wr_data_rom[ 9115]='h00000000;
    rd_cycle[ 9116] = 1'b0;  wr_cycle[ 9116] = 1'b0;  addr_rom[ 9116]='h00000000;  wr_data_rom[ 9116]='h00000000;
    rd_cycle[ 9117] = 1'b0;  wr_cycle[ 9117] = 1'b0;  addr_rom[ 9117]='h00000000;  wr_data_rom[ 9117]='h00000000;
    rd_cycle[ 9118] = 1'b0;  wr_cycle[ 9118] = 1'b0;  addr_rom[ 9118]='h00000000;  wr_data_rom[ 9118]='h00000000;
    rd_cycle[ 9119] = 1'b0;  wr_cycle[ 9119] = 1'b0;  addr_rom[ 9119]='h00000000;  wr_data_rom[ 9119]='h00000000;
    rd_cycle[ 9120] = 1'b0;  wr_cycle[ 9120] = 1'b0;  addr_rom[ 9120]='h00000000;  wr_data_rom[ 9120]='h00000000;
    rd_cycle[ 9121] = 1'b0;  wr_cycle[ 9121] = 1'b0;  addr_rom[ 9121]='h00000000;  wr_data_rom[ 9121]='h00000000;
    rd_cycle[ 9122] = 1'b0;  wr_cycle[ 9122] = 1'b0;  addr_rom[ 9122]='h00000000;  wr_data_rom[ 9122]='h00000000;
    rd_cycle[ 9123] = 1'b0;  wr_cycle[ 9123] = 1'b0;  addr_rom[ 9123]='h00000000;  wr_data_rom[ 9123]='h00000000;
    rd_cycle[ 9124] = 1'b0;  wr_cycle[ 9124] = 1'b0;  addr_rom[ 9124]='h00000000;  wr_data_rom[ 9124]='h00000000;
    rd_cycle[ 9125] = 1'b0;  wr_cycle[ 9125] = 1'b0;  addr_rom[ 9125]='h00000000;  wr_data_rom[ 9125]='h00000000;
    rd_cycle[ 9126] = 1'b0;  wr_cycle[ 9126] = 1'b0;  addr_rom[ 9126]='h00000000;  wr_data_rom[ 9126]='h00000000;
    rd_cycle[ 9127] = 1'b0;  wr_cycle[ 9127] = 1'b0;  addr_rom[ 9127]='h00000000;  wr_data_rom[ 9127]='h00000000;
    rd_cycle[ 9128] = 1'b0;  wr_cycle[ 9128] = 1'b0;  addr_rom[ 9128]='h00000000;  wr_data_rom[ 9128]='h00000000;
    rd_cycle[ 9129] = 1'b0;  wr_cycle[ 9129] = 1'b0;  addr_rom[ 9129]='h00000000;  wr_data_rom[ 9129]='h00000000;
    rd_cycle[ 9130] = 1'b0;  wr_cycle[ 9130] = 1'b0;  addr_rom[ 9130]='h00000000;  wr_data_rom[ 9130]='h00000000;
    rd_cycle[ 9131] = 1'b0;  wr_cycle[ 9131] = 1'b0;  addr_rom[ 9131]='h00000000;  wr_data_rom[ 9131]='h00000000;
    rd_cycle[ 9132] = 1'b0;  wr_cycle[ 9132] = 1'b0;  addr_rom[ 9132]='h00000000;  wr_data_rom[ 9132]='h00000000;
    rd_cycle[ 9133] = 1'b0;  wr_cycle[ 9133] = 1'b0;  addr_rom[ 9133]='h00000000;  wr_data_rom[ 9133]='h00000000;
    rd_cycle[ 9134] = 1'b0;  wr_cycle[ 9134] = 1'b0;  addr_rom[ 9134]='h00000000;  wr_data_rom[ 9134]='h00000000;
    rd_cycle[ 9135] = 1'b0;  wr_cycle[ 9135] = 1'b0;  addr_rom[ 9135]='h00000000;  wr_data_rom[ 9135]='h00000000;
    rd_cycle[ 9136] = 1'b0;  wr_cycle[ 9136] = 1'b0;  addr_rom[ 9136]='h00000000;  wr_data_rom[ 9136]='h00000000;
    rd_cycle[ 9137] = 1'b0;  wr_cycle[ 9137] = 1'b0;  addr_rom[ 9137]='h00000000;  wr_data_rom[ 9137]='h00000000;
    rd_cycle[ 9138] = 1'b0;  wr_cycle[ 9138] = 1'b0;  addr_rom[ 9138]='h00000000;  wr_data_rom[ 9138]='h00000000;
    rd_cycle[ 9139] = 1'b0;  wr_cycle[ 9139] = 1'b0;  addr_rom[ 9139]='h00000000;  wr_data_rom[ 9139]='h00000000;
    rd_cycle[ 9140] = 1'b0;  wr_cycle[ 9140] = 1'b0;  addr_rom[ 9140]='h00000000;  wr_data_rom[ 9140]='h00000000;
    rd_cycle[ 9141] = 1'b0;  wr_cycle[ 9141] = 1'b0;  addr_rom[ 9141]='h00000000;  wr_data_rom[ 9141]='h00000000;
    rd_cycle[ 9142] = 1'b0;  wr_cycle[ 9142] = 1'b0;  addr_rom[ 9142]='h00000000;  wr_data_rom[ 9142]='h00000000;
    rd_cycle[ 9143] = 1'b0;  wr_cycle[ 9143] = 1'b0;  addr_rom[ 9143]='h00000000;  wr_data_rom[ 9143]='h00000000;
    rd_cycle[ 9144] = 1'b0;  wr_cycle[ 9144] = 1'b0;  addr_rom[ 9144]='h00000000;  wr_data_rom[ 9144]='h00000000;
    rd_cycle[ 9145] = 1'b0;  wr_cycle[ 9145] = 1'b0;  addr_rom[ 9145]='h00000000;  wr_data_rom[ 9145]='h00000000;
    rd_cycle[ 9146] = 1'b0;  wr_cycle[ 9146] = 1'b0;  addr_rom[ 9146]='h00000000;  wr_data_rom[ 9146]='h00000000;
    rd_cycle[ 9147] = 1'b0;  wr_cycle[ 9147] = 1'b0;  addr_rom[ 9147]='h00000000;  wr_data_rom[ 9147]='h00000000;
    rd_cycle[ 9148] = 1'b0;  wr_cycle[ 9148] = 1'b0;  addr_rom[ 9148]='h00000000;  wr_data_rom[ 9148]='h00000000;
    rd_cycle[ 9149] = 1'b0;  wr_cycle[ 9149] = 1'b0;  addr_rom[ 9149]='h00000000;  wr_data_rom[ 9149]='h00000000;
    rd_cycle[ 9150] = 1'b0;  wr_cycle[ 9150] = 1'b0;  addr_rom[ 9150]='h00000000;  wr_data_rom[ 9150]='h00000000;
    rd_cycle[ 9151] = 1'b0;  wr_cycle[ 9151] = 1'b0;  addr_rom[ 9151]='h00000000;  wr_data_rom[ 9151]='h00000000;
    rd_cycle[ 9152] = 1'b0;  wr_cycle[ 9152] = 1'b0;  addr_rom[ 9152]='h00000000;  wr_data_rom[ 9152]='h00000000;
    rd_cycle[ 9153] = 1'b0;  wr_cycle[ 9153] = 1'b0;  addr_rom[ 9153]='h00000000;  wr_data_rom[ 9153]='h00000000;
    rd_cycle[ 9154] = 1'b0;  wr_cycle[ 9154] = 1'b0;  addr_rom[ 9154]='h00000000;  wr_data_rom[ 9154]='h00000000;
    rd_cycle[ 9155] = 1'b0;  wr_cycle[ 9155] = 1'b0;  addr_rom[ 9155]='h00000000;  wr_data_rom[ 9155]='h00000000;
    rd_cycle[ 9156] = 1'b0;  wr_cycle[ 9156] = 1'b0;  addr_rom[ 9156]='h00000000;  wr_data_rom[ 9156]='h00000000;
    rd_cycle[ 9157] = 1'b0;  wr_cycle[ 9157] = 1'b0;  addr_rom[ 9157]='h00000000;  wr_data_rom[ 9157]='h00000000;
    rd_cycle[ 9158] = 1'b0;  wr_cycle[ 9158] = 1'b0;  addr_rom[ 9158]='h00000000;  wr_data_rom[ 9158]='h00000000;
    rd_cycle[ 9159] = 1'b0;  wr_cycle[ 9159] = 1'b0;  addr_rom[ 9159]='h00000000;  wr_data_rom[ 9159]='h00000000;
    rd_cycle[ 9160] = 1'b0;  wr_cycle[ 9160] = 1'b0;  addr_rom[ 9160]='h00000000;  wr_data_rom[ 9160]='h00000000;
    rd_cycle[ 9161] = 1'b0;  wr_cycle[ 9161] = 1'b0;  addr_rom[ 9161]='h00000000;  wr_data_rom[ 9161]='h00000000;
    rd_cycle[ 9162] = 1'b0;  wr_cycle[ 9162] = 1'b0;  addr_rom[ 9162]='h00000000;  wr_data_rom[ 9162]='h00000000;
    rd_cycle[ 9163] = 1'b0;  wr_cycle[ 9163] = 1'b0;  addr_rom[ 9163]='h00000000;  wr_data_rom[ 9163]='h00000000;
    rd_cycle[ 9164] = 1'b0;  wr_cycle[ 9164] = 1'b0;  addr_rom[ 9164]='h00000000;  wr_data_rom[ 9164]='h00000000;
    rd_cycle[ 9165] = 1'b0;  wr_cycle[ 9165] = 1'b0;  addr_rom[ 9165]='h00000000;  wr_data_rom[ 9165]='h00000000;
    rd_cycle[ 9166] = 1'b0;  wr_cycle[ 9166] = 1'b0;  addr_rom[ 9166]='h00000000;  wr_data_rom[ 9166]='h00000000;
    rd_cycle[ 9167] = 1'b0;  wr_cycle[ 9167] = 1'b0;  addr_rom[ 9167]='h00000000;  wr_data_rom[ 9167]='h00000000;
    rd_cycle[ 9168] = 1'b0;  wr_cycle[ 9168] = 1'b0;  addr_rom[ 9168]='h00000000;  wr_data_rom[ 9168]='h00000000;
    rd_cycle[ 9169] = 1'b0;  wr_cycle[ 9169] = 1'b0;  addr_rom[ 9169]='h00000000;  wr_data_rom[ 9169]='h00000000;
    rd_cycle[ 9170] = 1'b0;  wr_cycle[ 9170] = 1'b0;  addr_rom[ 9170]='h00000000;  wr_data_rom[ 9170]='h00000000;
    rd_cycle[ 9171] = 1'b0;  wr_cycle[ 9171] = 1'b0;  addr_rom[ 9171]='h00000000;  wr_data_rom[ 9171]='h00000000;
    rd_cycle[ 9172] = 1'b0;  wr_cycle[ 9172] = 1'b0;  addr_rom[ 9172]='h00000000;  wr_data_rom[ 9172]='h00000000;
    rd_cycle[ 9173] = 1'b0;  wr_cycle[ 9173] = 1'b0;  addr_rom[ 9173]='h00000000;  wr_data_rom[ 9173]='h00000000;
    rd_cycle[ 9174] = 1'b0;  wr_cycle[ 9174] = 1'b0;  addr_rom[ 9174]='h00000000;  wr_data_rom[ 9174]='h00000000;
    rd_cycle[ 9175] = 1'b0;  wr_cycle[ 9175] = 1'b0;  addr_rom[ 9175]='h00000000;  wr_data_rom[ 9175]='h00000000;
    rd_cycle[ 9176] = 1'b0;  wr_cycle[ 9176] = 1'b0;  addr_rom[ 9176]='h00000000;  wr_data_rom[ 9176]='h00000000;
    rd_cycle[ 9177] = 1'b0;  wr_cycle[ 9177] = 1'b0;  addr_rom[ 9177]='h00000000;  wr_data_rom[ 9177]='h00000000;
    rd_cycle[ 9178] = 1'b0;  wr_cycle[ 9178] = 1'b0;  addr_rom[ 9178]='h00000000;  wr_data_rom[ 9178]='h00000000;
    rd_cycle[ 9179] = 1'b0;  wr_cycle[ 9179] = 1'b0;  addr_rom[ 9179]='h00000000;  wr_data_rom[ 9179]='h00000000;
    rd_cycle[ 9180] = 1'b0;  wr_cycle[ 9180] = 1'b0;  addr_rom[ 9180]='h00000000;  wr_data_rom[ 9180]='h00000000;
    rd_cycle[ 9181] = 1'b0;  wr_cycle[ 9181] = 1'b0;  addr_rom[ 9181]='h00000000;  wr_data_rom[ 9181]='h00000000;
    rd_cycle[ 9182] = 1'b0;  wr_cycle[ 9182] = 1'b0;  addr_rom[ 9182]='h00000000;  wr_data_rom[ 9182]='h00000000;
    rd_cycle[ 9183] = 1'b0;  wr_cycle[ 9183] = 1'b0;  addr_rom[ 9183]='h00000000;  wr_data_rom[ 9183]='h00000000;
    rd_cycle[ 9184] = 1'b0;  wr_cycle[ 9184] = 1'b0;  addr_rom[ 9184]='h00000000;  wr_data_rom[ 9184]='h00000000;
    rd_cycle[ 9185] = 1'b0;  wr_cycle[ 9185] = 1'b0;  addr_rom[ 9185]='h00000000;  wr_data_rom[ 9185]='h00000000;
    rd_cycle[ 9186] = 1'b0;  wr_cycle[ 9186] = 1'b0;  addr_rom[ 9186]='h00000000;  wr_data_rom[ 9186]='h00000000;
    rd_cycle[ 9187] = 1'b0;  wr_cycle[ 9187] = 1'b0;  addr_rom[ 9187]='h00000000;  wr_data_rom[ 9187]='h00000000;
    rd_cycle[ 9188] = 1'b0;  wr_cycle[ 9188] = 1'b0;  addr_rom[ 9188]='h00000000;  wr_data_rom[ 9188]='h00000000;
    rd_cycle[ 9189] = 1'b0;  wr_cycle[ 9189] = 1'b0;  addr_rom[ 9189]='h00000000;  wr_data_rom[ 9189]='h00000000;
    rd_cycle[ 9190] = 1'b0;  wr_cycle[ 9190] = 1'b0;  addr_rom[ 9190]='h00000000;  wr_data_rom[ 9190]='h00000000;
    rd_cycle[ 9191] = 1'b0;  wr_cycle[ 9191] = 1'b0;  addr_rom[ 9191]='h00000000;  wr_data_rom[ 9191]='h00000000;
    rd_cycle[ 9192] = 1'b0;  wr_cycle[ 9192] = 1'b0;  addr_rom[ 9192]='h00000000;  wr_data_rom[ 9192]='h00000000;
    rd_cycle[ 9193] = 1'b0;  wr_cycle[ 9193] = 1'b0;  addr_rom[ 9193]='h00000000;  wr_data_rom[ 9193]='h00000000;
    rd_cycle[ 9194] = 1'b0;  wr_cycle[ 9194] = 1'b0;  addr_rom[ 9194]='h00000000;  wr_data_rom[ 9194]='h00000000;
    rd_cycle[ 9195] = 1'b0;  wr_cycle[ 9195] = 1'b0;  addr_rom[ 9195]='h00000000;  wr_data_rom[ 9195]='h00000000;
    rd_cycle[ 9196] = 1'b0;  wr_cycle[ 9196] = 1'b0;  addr_rom[ 9196]='h00000000;  wr_data_rom[ 9196]='h00000000;
    rd_cycle[ 9197] = 1'b0;  wr_cycle[ 9197] = 1'b0;  addr_rom[ 9197]='h00000000;  wr_data_rom[ 9197]='h00000000;
    rd_cycle[ 9198] = 1'b0;  wr_cycle[ 9198] = 1'b0;  addr_rom[ 9198]='h00000000;  wr_data_rom[ 9198]='h00000000;
    rd_cycle[ 9199] = 1'b0;  wr_cycle[ 9199] = 1'b0;  addr_rom[ 9199]='h00000000;  wr_data_rom[ 9199]='h00000000;
    rd_cycle[ 9200] = 1'b0;  wr_cycle[ 9200] = 1'b0;  addr_rom[ 9200]='h00000000;  wr_data_rom[ 9200]='h00000000;
    rd_cycle[ 9201] = 1'b0;  wr_cycle[ 9201] = 1'b0;  addr_rom[ 9201]='h00000000;  wr_data_rom[ 9201]='h00000000;
    rd_cycle[ 9202] = 1'b0;  wr_cycle[ 9202] = 1'b0;  addr_rom[ 9202]='h00000000;  wr_data_rom[ 9202]='h00000000;
    rd_cycle[ 9203] = 1'b0;  wr_cycle[ 9203] = 1'b0;  addr_rom[ 9203]='h00000000;  wr_data_rom[ 9203]='h00000000;
    rd_cycle[ 9204] = 1'b0;  wr_cycle[ 9204] = 1'b0;  addr_rom[ 9204]='h00000000;  wr_data_rom[ 9204]='h00000000;
    rd_cycle[ 9205] = 1'b0;  wr_cycle[ 9205] = 1'b0;  addr_rom[ 9205]='h00000000;  wr_data_rom[ 9205]='h00000000;
    rd_cycle[ 9206] = 1'b0;  wr_cycle[ 9206] = 1'b0;  addr_rom[ 9206]='h00000000;  wr_data_rom[ 9206]='h00000000;
    rd_cycle[ 9207] = 1'b0;  wr_cycle[ 9207] = 1'b0;  addr_rom[ 9207]='h00000000;  wr_data_rom[ 9207]='h00000000;
    rd_cycle[ 9208] = 1'b0;  wr_cycle[ 9208] = 1'b0;  addr_rom[ 9208]='h00000000;  wr_data_rom[ 9208]='h00000000;
    rd_cycle[ 9209] = 1'b0;  wr_cycle[ 9209] = 1'b0;  addr_rom[ 9209]='h00000000;  wr_data_rom[ 9209]='h00000000;
    rd_cycle[ 9210] = 1'b0;  wr_cycle[ 9210] = 1'b0;  addr_rom[ 9210]='h00000000;  wr_data_rom[ 9210]='h00000000;
    rd_cycle[ 9211] = 1'b0;  wr_cycle[ 9211] = 1'b0;  addr_rom[ 9211]='h00000000;  wr_data_rom[ 9211]='h00000000;
    rd_cycle[ 9212] = 1'b0;  wr_cycle[ 9212] = 1'b0;  addr_rom[ 9212]='h00000000;  wr_data_rom[ 9212]='h00000000;
    rd_cycle[ 9213] = 1'b0;  wr_cycle[ 9213] = 1'b0;  addr_rom[ 9213]='h00000000;  wr_data_rom[ 9213]='h00000000;
    rd_cycle[ 9214] = 1'b0;  wr_cycle[ 9214] = 1'b0;  addr_rom[ 9214]='h00000000;  wr_data_rom[ 9214]='h00000000;
    rd_cycle[ 9215] = 1'b0;  wr_cycle[ 9215] = 1'b0;  addr_rom[ 9215]='h00000000;  wr_data_rom[ 9215]='h00000000;
    rd_cycle[ 9216] = 1'b0;  wr_cycle[ 9216] = 1'b0;  addr_rom[ 9216]='h00000000;  wr_data_rom[ 9216]='h00000000;
    rd_cycle[ 9217] = 1'b0;  wr_cycle[ 9217] = 1'b0;  addr_rom[ 9217]='h00000000;  wr_data_rom[ 9217]='h00000000;
    rd_cycle[ 9218] = 1'b0;  wr_cycle[ 9218] = 1'b0;  addr_rom[ 9218]='h00000000;  wr_data_rom[ 9218]='h00000000;
    rd_cycle[ 9219] = 1'b0;  wr_cycle[ 9219] = 1'b0;  addr_rom[ 9219]='h00000000;  wr_data_rom[ 9219]='h00000000;
    rd_cycle[ 9220] = 1'b0;  wr_cycle[ 9220] = 1'b0;  addr_rom[ 9220]='h00000000;  wr_data_rom[ 9220]='h00000000;
    rd_cycle[ 9221] = 1'b0;  wr_cycle[ 9221] = 1'b0;  addr_rom[ 9221]='h00000000;  wr_data_rom[ 9221]='h00000000;
    rd_cycle[ 9222] = 1'b0;  wr_cycle[ 9222] = 1'b0;  addr_rom[ 9222]='h00000000;  wr_data_rom[ 9222]='h00000000;
    rd_cycle[ 9223] = 1'b0;  wr_cycle[ 9223] = 1'b0;  addr_rom[ 9223]='h00000000;  wr_data_rom[ 9223]='h00000000;
    rd_cycle[ 9224] = 1'b0;  wr_cycle[ 9224] = 1'b0;  addr_rom[ 9224]='h00000000;  wr_data_rom[ 9224]='h00000000;
    rd_cycle[ 9225] = 1'b0;  wr_cycle[ 9225] = 1'b0;  addr_rom[ 9225]='h00000000;  wr_data_rom[ 9225]='h00000000;
    rd_cycle[ 9226] = 1'b0;  wr_cycle[ 9226] = 1'b0;  addr_rom[ 9226]='h00000000;  wr_data_rom[ 9226]='h00000000;
    rd_cycle[ 9227] = 1'b0;  wr_cycle[ 9227] = 1'b0;  addr_rom[ 9227]='h00000000;  wr_data_rom[ 9227]='h00000000;
    rd_cycle[ 9228] = 1'b0;  wr_cycle[ 9228] = 1'b0;  addr_rom[ 9228]='h00000000;  wr_data_rom[ 9228]='h00000000;
    rd_cycle[ 9229] = 1'b0;  wr_cycle[ 9229] = 1'b0;  addr_rom[ 9229]='h00000000;  wr_data_rom[ 9229]='h00000000;
    rd_cycle[ 9230] = 1'b0;  wr_cycle[ 9230] = 1'b0;  addr_rom[ 9230]='h00000000;  wr_data_rom[ 9230]='h00000000;
    rd_cycle[ 9231] = 1'b0;  wr_cycle[ 9231] = 1'b0;  addr_rom[ 9231]='h00000000;  wr_data_rom[ 9231]='h00000000;
    rd_cycle[ 9232] = 1'b0;  wr_cycle[ 9232] = 1'b0;  addr_rom[ 9232]='h00000000;  wr_data_rom[ 9232]='h00000000;
    rd_cycle[ 9233] = 1'b0;  wr_cycle[ 9233] = 1'b0;  addr_rom[ 9233]='h00000000;  wr_data_rom[ 9233]='h00000000;
    rd_cycle[ 9234] = 1'b0;  wr_cycle[ 9234] = 1'b0;  addr_rom[ 9234]='h00000000;  wr_data_rom[ 9234]='h00000000;
    rd_cycle[ 9235] = 1'b0;  wr_cycle[ 9235] = 1'b0;  addr_rom[ 9235]='h00000000;  wr_data_rom[ 9235]='h00000000;
    rd_cycle[ 9236] = 1'b0;  wr_cycle[ 9236] = 1'b0;  addr_rom[ 9236]='h00000000;  wr_data_rom[ 9236]='h00000000;
    rd_cycle[ 9237] = 1'b0;  wr_cycle[ 9237] = 1'b0;  addr_rom[ 9237]='h00000000;  wr_data_rom[ 9237]='h00000000;
    rd_cycle[ 9238] = 1'b0;  wr_cycle[ 9238] = 1'b0;  addr_rom[ 9238]='h00000000;  wr_data_rom[ 9238]='h00000000;
    rd_cycle[ 9239] = 1'b0;  wr_cycle[ 9239] = 1'b0;  addr_rom[ 9239]='h00000000;  wr_data_rom[ 9239]='h00000000;
    rd_cycle[ 9240] = 1'b0;  wr_cycle[ 9240] = 1'b0;  addr_rom[ 9240]='h00000000;  wr_data_rom[ 9240]='h00000000;
    rd_cycle[ 9241] = 1'b0;  wr_cycle[ 9241] = 1'b0;  addr_rom[ 9241]='h00000000;  wr_data_rom[ 9241]='h00000000;
    rd_cycle[ 9242] = 1'b0;  wr_cycle[ 9242] = 1'b0;  addr_rom[ 9242]='h00000000;  wr_data_rom[ 9242]='h00000000;
    rd_cycle[ 9243] = 1'b0;  wr_cycle[ 9243] = 1'b0;  addr_rom[ 9243]='h00000000;  wr_data_rom[ 9243]='h00000000;
    rd_cycle[ 9244] = 1'b0;  wr_cycle[ 9244] = 1'b0;  addr_rom[ 9244]='h00000000;  wr_data_rom[ 9244]='h00000000;
    rd_cycle[ 9245] = 1'b0;  wr_cycle[ 9245] = 1'b0;  addr_rom[ 9245]='h00000000;  wr_data_rom[ 9245]='h00000000;
    rd_cycle[ 9246] = 1'b0;  wr_cycle[ 9246] = 1'b0;  addr_rom[ 9246]='h00000000;  wr_data_rom[ 9246]='h00000000;
    rd_cycle[ 9247] = 1'b0;  wr_cycle[ 9247] = 1'b0;  addr_rom[ 9247]='h00000000;  wr_data_rom[ 9247]='h00000000;
    rd_cycle[ 9248] = 1'b0;  wr_cycle[ 9248] = 1'b0;  addr_rom[ 9248]='h00000000;  wr_data_rom[ 9248]='h00000000;
    rd_cycle[ 9249] = 1'b0;  wr_cycle[ 9249] = 1'b0;  addr_rom[ 9249]='h00000000;  wr_data_rom[ 9249]='h00000000;
    rd_cycle[ 9250] = 1'b0;  wr_cycle[ 9250] = 1'b0;  addr_rom[ 9250]='h00000000;  wr_data_rom[ 9250]='h00000000;
    rd_cycle[ 9251] = 1'b0;  wr_cycle[ 9251] = 1'b0;  addr_rom[ 9251]='h00000000;  wr_data_rom[ 9251]='h00000000;
    rd_cycle[ 9252] = 1'b0;  wr_cycle[ 9252] = 1'b0;  addr_rom[ 9252]='h00000000;  wr_data_rom[ 9252]='h00000000;
    rd_cycle[ 9253] = 1'b0;  wr_cycle[ 9253] = 1'b0;  addr_rom[ 9253]='h00000000;  wr_data_rom[ 9253]='h00000000;
    rd_cycle[ 9254] = 1'b0;  wr_cycle[ 9254] = 1'b0;  addr_rom[ 9254]='h00000000;  wr_data_rom[ 9254]='h00000000;
    rd_cycle[ 9255] = 1'b0;  wr_cycle[ 9255] = 1'b0;  addr_rom[ 9255]='h00000000;  wr_data_rom[ 9255]='h00000000;
    rd_cycle[ 9256] = 1'b0;  wr_cycle[ 9256] = 1'b0;  addr_rom[ 9256]='h00000000;  wr_data_rom[ 9256]='h00000000;
    rd_cycle[ 9257] = 1'b0;  wr_cycle[ 9257] = 1'b0;  addr_rom[ 9257]='h00000000;  wr_data_rom[ 9257]='h00000000;
    rd_cycle[ 9258] = 1'b0;  wr_cycle[ 9258] = 1'b0;  addr_rom[ 9258]='h00000000;  wr_data_rom[ 9258]='h00000000;
    rd_cycle[ 9259] = 1'b0;  wr_cycle[ 9259] = 1'b0;  addr_rom[ 9259]='h00000000;  wr_data_rom[ 9259]='h00000000;
    rd_cycle[ 9260] = 1'b0;  wr_cycle[ 9260] = 1'b0;  addr_rom[ 9260]='h00000000;  wr_data_rom[ 9260]='h00000000;
    rd_cycle[ 9261] = 1'b0;  wr_cycle[ 9261] = 1'b0;  addr_rom[ 9261]='h00000000;  wr_data_rom[ 9261]='h00000000;
    rd_cycle[ 9262] = 1'b0;  wr_cycle[ 9262] = 1'b0;  addr_rom[ 9262]='h00000000;  wr_data_rom[ 9262]='h00000000;
    rd_cycle[ 9263] = 1'b0;  wr_cycle[ 9263] = 1'b0;  addr_rom[ 9263]='h00000000;  wr_data_rom[ 9263]='h00000000;
    rd_cycle[ 9264] = 1'b0;  wr_cycle[ 9264] = 1'b0;  addr_rom[ 9264]='h00000000;  wr_data_rom[ 9264]='h00000000;
    rd_cycle[ 9265] = 1'b0;  wr_cycle[ 9265] = 1'b0;  addr_rom[ 9265]='h00000000;  wr_data_rom[ 9265]='h00000000;
    rd_cycle[ 9266] = 1'b0;  wr_cycle[ 9266] = 1'b0;  addr_rom[ 9266]='h00000000;  wr_data_rom[ 9266]='h00000000;
    rd_cycle[ 9267] = 1'b0;  wr_cycle[ 9267] = 1'b0;  addr_rom[ 9267]='h00000000;  wr_data_rom[ 9267]='h00000000;
    rd_cycle[ 9268] = 1'b0;  wr_cycle[ 9268] = 1'b0;  addr_rom[ 9268]='h00000000;  wr_data_rom[ 9268]='h00000000;
    rd_cycle[ 9269] = 1'b0;  wr_cycle[ 9269] = 1'b0;  addr_rom[ 9269]='h00000000;  wr_data_rom[ 9269]='h00000000;
    rd_cycle[ 9270] = 1'b0;  wr_cycle[ 9270] = 1'b0;  addr_rom[ 9270]='h00000000;  wr_data_rom[ 9270]='h00000000;
    rd_cycle[ 9271] = 1'b0;  wr_cycle[ 9271] = 1'b0;  addr_rom[ 9271]='h00000000;  wr_data_rom[ 9271]='h00000000;
    rd_cycle[ 9272] = 1'b0;  wr_cycle[ 9272] = 1'b0;  addr_rom[ 9272]='h00000000;  wr_data_rom[ 9272]='h00000000;
    rd_cycle[ 9273] = 1'b0;  wr_cycle[ 9273] = 1'b0;  addr_rom[ 9273]='h00000000;  wr_data_rom[ 9273]='h00000000;
    rd_cycle[ 9274] = 1'b0;  wr_cycle[ 9274] = 1'b0;  addr_rom[ 9274]='h00000000;  wr_data_rom[ 9274]='h00000000;
    rd_cycle[ 9275] = 1'b0;  wr_cycle[ 9275] = 1'b0;  addr_rom[ 9275]='h00000000;  wr_data_rom[ 9275]='h00000000;
    rd_cycle[ 9276] = 1'b0;  wr_cycle[ 9276] = 1'b0;  addr_rom[ 9276]='h00000000;  wr_data_rom[ 9276]='h00000000;
    rd_cycle[ 9277] = 1'b0;  wr_cycle[ 9277] = 1'b0;  addr_rom[ 9277]='h00000000;  wr_data_rom[ 9277]='h00000000;
    rd_cycle[ 9278] = 1'b0;  wr_cycle[ 9278] = 1'b0;  addr_rom[ 9278]='h00000000;  wr_data_rom[ 9278]='h00000000;
    rd_cycle[ 9279] = 1'b0;  wr_cycle[ 9279] = 1'b0;  addr_rom[ 9279]='h00000000;  wr_data_rom[ 9279]='h00000000;
    rd_cycle[ 9280] = 1'b0;  wr_cycle[ 9280] = 1'b0;  addr_rom[ 9280]='h00000000;  wr_data_rom[ 9280]='h00000000;
    rd_cycle[ 9281] = 1'b0;  wr_cycle[ 9281] = 1'b0;  addr_rom[ 9281]='h00000000;  wr_data_rom[ 9281]='h00000000;
    rd_cycle[ 9282] = 1'b0;  wr_cycle[ 9282] = 1'b0;  addr_rom[ 9282]='h00000000;  wr_data_rom[ 9282]='h00000000;
    rd_cycle[ 9283] = 1'b0;  wr_cycle[ 9283] = 1'b0;  addr_rom[ 9283]='h00000000;  wr_data_rom[ 9283]='h00000000;
    rd_cycle[ 9284] = 1'b0;  wr_cycle[ 9284] = 1'b0;  addr_rom[ 9284]='h00000000;  wr_data_rom[ 9284]='h00000000;
    rd_cycle[ 9285] = 1'b0;  wr_cycle[ 9285] = 1'b0;  addr_rom[ 9285]='h00000000;  wr_data_rom[ 9285]='h00000000;
    rd_cycle[ 9286] = 1'b0;  wr_cycle[ 9286] = 1'b0;  addr_rom[ 9286]='h00000000;  wr_data_rom[ 9286]='h00000000;
    rd_cycle[ 9287] = 1'b0;  wr_cycle[ 9287] = 1'b0;  addr_rom[ 9287]='h00000000;  wr_data_rom[ 9287]='h00000000;
    rd_cycle[ 9288] = 1'b0;  wr_cycle[ 9288] = 1'b0;  addr_rom[ 9288]='h00000000;  wr_data_rom[ 9288]='h00000000;
    rd_cycle[ 9289] = 1'b0;  wr_cycle[ 9289] = 1'b0;  addr_rom[ 9289]='h00000000;  wr_data_rom[ 9289]='h00000000;
    rd_cycle[ 9290] = 1'b0;  wr_cycle[ 9290] = 1'b0;  addr_rom[ 9290]='h00000000;  wr_data_rom[ 9290]='h00000000;
    rd_cycle[ 9291] = 1'b0;  wr_cycle[ 9291] = 1'b0;  addr_rom[ 9291]='h00000000;  wr_data_rom[ 9291]='h00000000;
    rd_cycle[ 9292] = 1'b0;  wr_cycle[ 9292] = 1'b0;  addr_rom[ 9292]='h00000000;  wr_data_rom[ 9292]='h00000000;
    rd_cycle[ 9293] = 1'b0;  wr_cycle[ 9293] = 1'b0;  addr_rom[ 9293]='h00000000;  wr_data_rom[ 9293]='h00000000;
    rd_cycle[ 9294] = 1'b0;  wr_cycle[ 9294] = 1'b0;  addr_rom[ 9294]='h00000000;  wr_data_rom[ 9294]='h00000000;
    rd_cycle[ 9295] = 1'b0;  wr_cycle[ 9295] = 1'b0;  addr_rom[ 9295]='h00000000;  wr_data_rom[ 9295]='h00000000;
    rd_cycle[ 9296] = 1'b0;  wr_cycle[ 9296] = 1'b0;  addr_rom[ 9296]='h00000000;  wr_data_rom[ 9296]='h00000000;
    rd_cycle[ 9297] = 1'b0;  wr_cycle[ 9297] = 1'b0;  addr_rom[ 9297]='h00000000;  wr_data_rom[ 9297]='h00000000;
    rd_cycle[ 9298] = 1'b0;  wr_cycle[ 9298] = 1'b0;  addr_rom[ 9298]='h00000000;  wr_data_rom[ 9298]='h00000000;
    rd_cycle[ 9299] = 1'b0;  wr_cycle[ 9299] = 1'b0;  addr_rom[ 9299]='h00000000;  wr_data_rom[ 9299]='h00000000;
    rd_cycle[ 9300] = 1'b0;  wr_cycle[ 9300] = 1'b0;  addr_rom[ 9300]='h00000000;  wr_data_rom[ 9300]='h00000000;
    rd_cycle[ 9301] = 1'b0;  wr_cycle[ 9301] = 1'b0;  addr_rom[ 9301]='h00000000;  wr_data_rom[ 9301]='h00000000;
    rd_cycle[ 9302] = 1'b0;  wr_cycle[ 9302] = 1'b0;  addr_rom[ 9302]='h00000000;  wr_data_rom[ 9302]='h00000000;
    rd_cycle[ 9303] = 1'b0;  wr_cycle[ 9303] = 1'b0;  addr_rom[ 9303]='h00000000;  wr_data_rom[ 9303]='h00000000;
    rd_cycle[ 9304] = 1'b0;  wr_cycle[ 9304] = 1'b0;  addr_rom[ 9304]='h00000000;  wr_data_rom[ 9304]='h00000000;
    rd_cycle[ 9305] = 1'b0;  wr_cycle[ 9305] = 1'b0;  addr_rom[ 9305]='h00000000;  wr_data_rom[ 9305]='h00000000;
    rd_cycle[ 9306] = 1'b0;  wr_cycle[ 9306] = 1'b0;  addr_rom[ 9306]='h00000000;  wr_data_rom[ 9306]='h00000000;
    rd_cycle[ 9307] = 1'b0;  wr_cycle[ 9307] = 1'b0;  addr_rom[ 9307]='h00000000;  wr_data_rom[ 9307]='h00000000;
    rd_cycle[ 9308] = 1'b0;  wr_cycle[ 9308] = 1'b0;  addr_rom[ 9308]='h00000000;  wr_data_rom[ 9308]='h00000000;
    rd_cycle[ 9309] = 1'b0;  wr_cycle[ 9309] = 1'b0;  addr_rom[ 9309]='h00000000;  wr_data_rom[ 9309]='h00000000;
    rd_cycle[ 9310] = 1'b0;  wr_cycle[ 9310] = 1'b0;  addr_rom[ 9310]='h00000000;  wr_data_rom[ 9310]='h00000000;
    rd_cycle[ 9311] = 1'b0;  wr_cycle[ 9311] = 1'b0;  addr_rom[ 9311]='h00000000;  wr_data_rom[ 9311]='h00000000;
    rd_cycle[ 9312] = 1'b0;  wr_cycle[ 9312] = 1'b0;  addr_rom[ 9312]='h00000000;  wr_data_rom[ 9312]='h00000000;
    rd_cycle[ 9313] = 1'b0;  wr_cycle[ 9313] = 1'b0;  addr_rom[ 9313]='h00000000;  wr_data_rom[ 9313]='h00000000;
    rd_cycle[ 9314] = 1'b0;  wr_cycle[ 9314] = 1'b0;  addr_rom[ 9314]='h00000000;  wr_data_rom[ 9314]='h00000000;
    rd_cycle[ 9315] = 1'b0;  wr_cycle[ 9315] = 1'b0;  addr_rom[ 9315]='h00000000;  wr_data_rom[ 9315]='h00000000;
    rd_cycle[ 9316] = 1'b0;  wr_cycle[ 9316] = 1'b0;  addr_rom[ 9316]='h00000000;  wr_data_rom[ 9316]='h00000000;
    rd_cycle[ 9317] = 1'b0;  wr_cycle[ 9317] = 1'b0;  addr_rom[ 9317]='h00000000;  wr_data_rom[ 9317]='h00000000;
    rd_cycle[ 9318] = 1'b0;  wr_cycle[ 9318] = 1'b0;  addr_rom[ 9318]='h00000000;  wr_data_rom[ 9318]='h00000000;
    rd_cycle[ 9319] = 1'b0;  wr_cycle[ 9319] = 1'b0;  addr_rom[ 9319]='h00000000;  wr_data_rom[ 9319]='h00000000;
    rd_cycle[ 9320] = 1'b0;  wr_cycle[ 9320] = 1'b0;  addr_rom[ 9320]='h00000000;  wr_data_rom[ 9320]='h00000000;
    rd_cycle[ 9321] = 1'b0;  wr_cycle[ 9321] = 1'b0;  addr_rom[ 9321]='h00000000;  wr_data_rom[ 9321]='h00000000;
    rd_cycle[ 9322] = 1'b0;  wr_cycle[ 9322] = 1'b0;  addr_rom[ 9322]='h00000000;  wr_data_rom[ 9322]='h00000000;
    rd_cycle[ 9323] = 1'b0;  wr_cycle[ 9323] = 1'b0;  addr_rom[ 9323]='h00000000;  wr_data_rom[ 9323]='h00000000;
    rd_cycle[ 9324] = 1'b0;  wr_cycle[ 9324] = 1'b0;  addr_rom[ 9324]='h00000000;  wr_data_rom[ 9324]='h00000000;
    rd_cycle[ 9325] = 1'b0;  wr_cycle[ 9325] = 1'b0;  addr_rom[ 9325]='h00000000;  wr_data_rom[ 9325]='h00000000;
    rd_cycle[ 9326] = 1'b0;  wr_cycle[ 9326] = 1'b0;  addr_rom[ 9326]='h00000000;  wr_data_rom[ 9326]='h00000000;
    rd_cycle[ 9327] = 1'b0;  wr_cycle[ 9327] = 1'b0;  addr_rom[ 9327]='h00000000;  wr_data_rom[ 9327]='h00000000;
    rd_cycle[ 9328] = 1'b0;  wr_cycle[ 9328] = 1'b0;  addr_rom[ 9328]='h00000000;  wr_data_rom[ 9328]='h00000000;
    rd_cycle[ 9329] = 1'b0;  wr_cycle[ 9329] = 1'b0;  addr_rom[ 9329]='h00000000;  wr_data_rom[ 9329]='h00000000;
    rd_cycle[ 9330] = 1'b0;  wr_cycle[ 9330] = 1'b0;  addr_rom[ 9330]='h00000000;  wr_data_rom[ 9330]='h00000000;
    rd_cycle[ 9331] = 1'b0;  wr_cycle[ 9331] = 1'b0;  addr_rom[ 9331]='h00000000;  wr_data_rom[ 9331]='h00000000;
    rd_cycle[ 9332] = 1'b0;  wr_cycle[ 9332] = 1'b0;  addr_rom[ 9332]='h00000000;  wr_data_rom[ 9332]='h00000000;
    rd_cycle[ 9333] = 1'b0;  wr_cycle[ 9333] = 1'b0;  addr_rom[ 9333]='h00000000;  wr_data_rom[ 9333]='h00000000;
    rd_cycle[ 9334] = 1'b0;  wr_cycle[ 9334] = 1'b0;  addr_rom[ 9334]='h00000000;  wr_data_rom[ 9334]='h00000000;
    rd_cycle[ 9335] = 1'b0;  wr_cycle[ 9335] = 1'b0;  addr_rom[ 9335]='h00000000;  wr_data_rom[ 9335]='h00000000;
    rd_cycle[ 9336] = 1'b0;  wr_cycle[ 9336] = 1'b0;  addr_rom[ 9336]='h00000000;  wr_data_rom[ 9336]='h00000000;
    rd_cycle[ 9337] = 1'b0;  wr_cycle[ 9337] = 1'b0;  addr_rom[ 9337]='h00000000;  wr_data_rom[ 9337]='h00000000;
    rd_cycle[ 9338] = 1'b0;  wr_cycle[ 9338] = 1'b0;  addr_rom[ 9338]='h00000000;  wr_data_rom[ 9338]='h00000000;
    rd_cycle[ 9339] = 1'b0;  wr_cycle[ 9339] = 1'b0;  addr_rom[ 9339]='h00000000;  wr_data_rom[ 9339]='h00000000;
    rd_cycle[ 9340] = 1'b0;  wr_cycle[ 9340] = 1'b0;  addr_rom[ 9340]='h00000000;  wr_data_rom[ 9340]='h00000000;
    rd_cycle[ 9341] = 1'b0;  wr_cycle[ 9341] = 1'b0;  addr_rom[ 9341]='h00000000;  wr_data_rom[ 9341]='h00000000;
    rd_cycle[ 9342] = 1'b0;  wr_cycle[ 9342] = 1'b0;  addr_rom[ 9342]='h00000000;  wr_data_rom[ 9342]='h00000000;
    rd_cycle[ 9343] = 1'b0;  wr_cycle[ 9343] = 1'b0;  addr_rom[ 9343]='h00000000;  wr_data_rom[ 9343]='h00000000;
    rd_cycle[ 9344] = 1'b0;  wr_cycle[ 9344] = 1'b0;  addr_rom[ 9344]='h00000000;  wr_data_rom[ 9344]='h00000000;
    rd_cycle[ 9345] = 1'b0;  wr_cycle[ 9345] = 1'b0;  addr_rom[ 9345]='h00000000;  wr_data_rom[ 9345]='h00000000;
    rd_cycle[ 9346] = 1'b0;  wr_cycle[ 9346] = 1'b0;  addr_rom[ 9346]='h00000000;  wr_data_rom[ 9346]='h00000000;
    rd_cycle[ 9347] = 1'b0;  wr_cycle[ 9347] = 1'b0;  addr_rom[ 9347]='h00000000;  wr_data_rom[ 9347]='h00000000;
    rd_cycle[ 9348] = 1'b0;  wr_cycle[ 9348] = 1'b0;  addr_rom[ 9348]='h00000000;  wr_data_rom[ 9348]='h00000000;
    rd_cycle[ 9349] = 1'b0;  wr_cycle[ 9349] = 1'b0;  addr_rom[ 9349]='h00000000;  wr_data_rom[ 9349]='h00000000;
    rd_cycle[ 9350] = 1'b0;  wr_cycle[ 9350] = 1'b0;  addr_rom[ 9350]='h00000000;  wr_data_rom[ 9350]='h00000000;
    rd_cycle[ 9351] = 1'b0;  wr_cycle[ 9351] = 1'b0;  addr_rom[ 9351]='h00000000;  wr_data_rom[ 9351]='h00000000;
    rd_cycle[ 9352] = 1'b0;  wr_cycle[ 9352] = 1'b0;  addr_rom[ 9352]='h00000000;  wr_data_rom[ 9352]='h00000000;
    rd_cycle[ 9353] = 1'b0;  wr_cycle[ 9353] = 1'b0;  addr_rom[ 9353]='h00000000;  wr_data_rom[ 9353]='h00000000;
    rd_cycle[ 9354] = 1'b0;  wr_cycle[ 9354] = 1'b0;  addr_rom[ 9354]='h00000000;  wr_data_rom[ 9354]='h00000000;
    rd_cycle[ 9355] = 1'b0;  wr_cycle[ 9355] = 1'b0;  addr_rom[ 9355]='h00000000;  wr_data_rom[ 9355]='h00000000;
    rd_cycle[ 9356] = 1'b0;  wr_cycle[ 9356] = 1'b0;  addr_rom[ 9356]='h00000000;  wr_data_rom[ 9356]='h00000000;
    rd_cycle[ 9357] = 1'b0;  wr_cycle[ 9357] = 1'b0;  addr_rom[ 9357]='h00000000;  wr_data_rom[ 9357]='h00000000;
    rd_cycle[ 9358] = 1'b0;  wr_cycle[ 9358] = 1'b0;  addr_rom[ 9358]='h00000000;  wr_data_rom[ 9358]='h00000000;
    rd_cycle[ 9359] = 1'b0;  wr_cycle[ 9359] = 1'b0;  addr_rom[ 9359]='h00000000;  wr_data_rom[ 9359]='h00000000;
    rd_cycle[ 9360] = 1'b0;  wr_cycle[ 9360] = 1'b0;  addr_rom[ 9360]='h00000000;  wr_data_rom[ 9360]='h00000000;
    rd_cycle[ 9361] = 1'b0;  wr_cycle[ 9361] = 1'b0;  addr_rom[ 9361]='h00000000;  wr_data_rom[ 9361]='h00000000;
    rd_cycle[ 9362] = 1'b0;  wr_cycle[ 9362] = 1'b0;  addr_rom[ 9362]='h00000000;  wr_data_rom[ 9362]='h00000000;
    rd_cycle[ 9363] = 1'b0;  wr_cycle[ 9363] = 1'b0;  addr_rom[ 9363]='h00000000;  wr_data_rom[ 9363]='h00000000;
    rd_cycle[ 9364] = 1'b0;  wr_cycle[ 9364] = 1'b0;  addr_rom[ 9364]='h00000000;  wr_data_rom[ 9364]='h00000000;
    rd_cycle[ 9365] = 1'b0;  wr_cycle[ 9365] = 1'b0;  addr_rom[ 9365]='h00000000;  wr_data_rom[ 9365]='h00000000;
    rd_cycle[ 9366] = 1'b0;  wr_cycle[ 9366] = 1'b0;  addr_rom[ 9366]='h00000000;  wr_data_rom[ 9366]='h00000000;
    rd_cycle[ 9367] = 1'b0;  wr_cycle[ 9367] = 1'b0;  addr_rom[ 9367]='h00000000;  wr_data_rom[ 9367]='h00000000;
    rd_cycle[ 9368] = 1'b0;  wr_cycle[ 9368] = 1'b0;  addr_rom[ 9368]='h00000000;  wr_data_rom[ 9368]='h00000000;
    rd_cycle[ 9369] = 1'b0;  wr_cycle[ 9369] = 1'b0;  addr_rom[ 9369]='h00000000;  wr_data_rom[ 9369]='h00000000;
    rd_cycle[ 9370] = 1'b0;  wr_cycle[ 9370] = 1'b0;  addr_rom[ 9370]='h00000000;  wr_data_rom[ 9370]='h00000000;
    rd_cycle[ 9371] = 1'b0;  wr_cycle[ 9371] = 1'b0;  addr_rom[ 9371]='h00000000;  wr_data_rom[ 9371]='h00000000;
    rd_cycle[ 9372] = 1'b0;  wr_cycle[ 9372] = 1'b0;  addr_rom[ 9372]='h00000000;  wr_data_rom[ 9372]='h00000000;
    rd_cycle[ 9373] = 1'b0;  wr_cycle[ 9373] = 1'b0;  addr_rom[ 9373]='h00000000;  wr_data_rom[ 9373]='h00000000;
    rd_cycle[ 9374] = 1'b0;  wr_cycle[ 9374] = 1'b0;  addr_rom[ 9374]='h00000000;  wr_data_rom[ 9374]='h00000000;
    rd_cycle[ 9375] = 1'b0;  wr_cycle[ 9375] = 1'b0;  addr_rom[ 9375]='h00000000;  wr_data_rom[ 9375]='h00000000;
    rd_cycle[ 9376] = 1'b0;  wr_cycle[ 9376] = 1'b0;  addr_rom[ 9376]='h00000000;  wr_data_rom[ 9376]='h00000000;
    rd_cycle[ 9377] = 1'b0;  wr_cycle[ 9377] = 1'b0;  addr_rom[ 9377]='h00000000;  wr_data_rom[ 9377]='h00000000;
    rd_cycle[ 9378] = 1'b0;  wr_cycle[ 9378] = 1'b0;  addr_rom[ 9378]='h00000000;  wr_data_rom[ 9378]='h00000000;
    rd_cycle[ 9379] = 1'b0;  wr_cycle[ 9379] = 1'b0;  addr_rom[ 9379]='h00000000;  wr_data_rom[ 9379]='h00000000;
    rd_cycle[ 9380] = 1'b0;  wr_cycle[ 9380] = 1'b0;  addr_rom[ 9380]='h00000000;  wr_data_rom[ 9380]='h00000000;
    rd_cycle[ 9381] = 1'b0;  wr_cycle[ 9381] = 1'b0;  addr_rom[ 9381]='h00000000;  wr_data_rom[ 9381]='h00000000;
    rd_cycle[ 9382] = 1'b0;  wr_cycle[ 9382] = 1'b0;  addr_rom[ 9382]='h00000000;  wr_data_rom[ 9382]='h00000000;
    rd_cycle[ 9383] = 1'b0;  wr_cycle[ 9383] = 1'b0;  addr_rom[ 9383]='h00000000;  wr_data_rom[ 9383]='h00000000;
    rd_cycle[ 9384] = 1'b0;  wr_cycle[ 9384] = 1'b0;  addr_rom[ 9384]='h00000000;  wr_data_rom[ 9384]='h00000000;
    rd_cycle[ 9385] = 1'b0;  wr_cycle[ 9385] = 1'b0;  addr_rom[ 9385]='h00000000;  wr_data_rom[ 9385]='h00000000;
    rd_cycle[ 9386] = 1'b0;  wr_cycle[ 9386] = 1'b0;  addr_rom[ 9386]='h00000000;  wr_data_rom[ 9386]='h00000000;
    rd_cycle[ 9387] = 1'b0;  wr_cycle[ 9387] = 1'b0;  addr_rom[ 9387]='h00000000;  wr_data_rom[ 9387]='h00000000;
    rd_cycle[ 9388] = 1'b0;  wr_cycle[ 9388] = 1'b0;  addr_rom[ 9388]='h00000000;  wr_data_rom[ 9388]='h00000000;
    rd_cycle[ 9389] = 1'b0;  wr_cycle[ 9389] = 1'b0;  addr_rom[ 9389]='h00000000;  wr_data_rom[ 9389]='h00000000;
    rd_cycle[ 9390] = 1'b0;  wr_cycle[ 9390] = 1'b0;  addr_rom[ 9390]='h00000000;  wr_data_rom[ 9390]='h00000000;
    rd_cycle[ 9391] = 1'b0;  wr_cycle[ 9391] = 1'b0;  addr_rom[ 9391]='h00000000;  wr_data_rom[ 9391]='h00000000;
    rd_cycle[ 9392] = 1'b0;  wr_cycle[ 9392] = 1'b0;  addr_rom[ 9392]='h00000000;  wr_data_rom[ 9392]='h00000000;
    rd_cycle[ 9393] = 1'b0;  wr_cycle[ 9393] = 1'b0;  addr_rom[ 9393]='h00000000;  wr_data_rom[ 9393]='h00000000;
    rd_cycle[ 9394] = 1'b0;  wr_cycle[ 9394] = 1'b0;  addr_rom[ 9394]='h00000000;  wr_data_rom[ 9394]='h00000000;
    rd_cycle[ 9395] = 1'b0;  wr_cycle[ 9395] = 1'b0;  addr_rom[ 9395]='h00000000;  wr_data_rom[ 9395]='h00000000;
    rd_cycle[ 9396] = 1'b0;  wr_cycle[ 9396] = 1'b0;  addr_rom[ 9396]='h00000000;  wr_data_rom[ 9396]='h00000000;
    rd_cycle[ 9397] = 1'b0;  wr_cycle[ 9397] = 1'b0;  addr_rom[ 9397]='h00000000;  wr_data_rom[ 9397]='h00000000;
    rd_cycle[ 9398] = 1'b0;  wr_cycle[ 9398] = 1'b0;  addr_rom[ 9398]='h00000000;  wr_data_rom[ 9398]='h00000000;
    rd_cycle[ 9399] = 1'b0;  wr_cycle[ 9399] = 1'b0;  addr_rom[ 9399]='h00000000;  wr_data_rom[ 9399]='h00000000;
    rd_cycle[ 9400] = 1'b0;  wr_cycle[ 9400] = 1'b0;  addr_rom[ 9400]='h00000000;  wr_data_rom[ 9400]='h00000000;
    rd_cycle[ 9401] = 1'b0;  wr_cycle[ 9401] = 1'b0;  addr_rom[ 9401]='h00000000;  wr_data_rom[ 9401]='h00000000;
    rd_cycle[ 9402] = 1'b0;  wr_cycle[ 9402] = 1'b0;  addr_rom[ 9402]='h00000000;  wr_data_rom[ 9402]='h00000000;
    rd_cycle[ 9403] = 1'b0;  wr_cycle[ 9403] = 1'b0;  addr_rom[ 9403]='h00000000;  wr_data_rom[ 9403]='h00000000;
    rd_cycle[ 9404] = 1'b0;  wr_cycle[ 9404] = 1'b0;  addr_rom[ 9404]='h00000000;  wr_data_rom[ 9404]='h00000000;
    rd_cycle[ 9405] = 1'b0;  wr_cycle[ 9405] = 1'b0;  addr_rom[ 9405]='h00000000;  wr_data_rom[ 9405]='h00000000;
    rd_cycle[ 9406] = 1'b0;  wr_cycle[ 9406] = 1'b0;  addr_rom[ 9406]='h00000000;  wr_data_rom[ 9406]='h00000000;
    rd_cycle[ 9407] = 1'b0;  wr_cycle[ 9407] = 1'b0;  addr_rom[ 9407]='h00000000;  wr_data_rom[ 9407]='h00000000;
    rd_cycle[ 9408] = 1'b0;  wr_cycle[ 9408] = 1'b0;  addr_rom[ 9408]='h00000000;  wr_data_rom[ 9408]='h00000000;
    rd_cycle[ 9409] = 1'b0;  wr_cycle[ 9409] = 1'b0;  addr_rom[ 9409]='h00000000;  wr_data_rom[ 9409]='h00000000;
    rd_cycle[ 9410] = 1'b0;  wr_cycle[ 9410] = 1'b0;  addr_rom[ 9410]='h00000000;  wr_data_rom[ 9410]='h00000000;
    rd_cycle[ 9411] = 1'b0;  wr_cycle[ 9411] = 1'b0;  addr_rom[ 9411]='h00000000;  wr_data_rom[ 9411]='h00000000;
    rd_cycle[ 9412] = 1'b0;  wr_cycle[ 9412] = 1'b0;  addr_rom[ 9412]='h00000000;  wr_data_rom[ 9412]='h00000000;
    rd_cycle[ 9413] = 1'b0;  wr_cycle[ 9413] = 1'b0;  addr_rom[ 9413]='h00000000;  wr_data_rom[ 9413]='h00000000;
    rd_cycle[ 9414] = 1'b0;  wr_cycle[ 9414] = 1'b0;  addr_rom[ 9414]='h00000000;  wr_data_rom[ 9414]='h00000000;
    rd_cycle[ 9415] = 1'b0;  wr_cycle[ 9415] = 1'b0;  addr_rom[ 9415]='h00000000;  wr_data_rom[ 9415]='h00000000;
    rd_cycle[ 9416] = 1'b0;  wr_cycle[ 9416] = 1'b0;  addr_rom[ 9416]='h00000000;  wr_data_rom[ 9416]='h00000000;
    rd_cycle[ 9417] = 1'b0;  wr_cycle[ 9417] = 1'b0;  addr_rom[ 9417]='h00000000;  wr_data_rom[ 9417]='h00000000;
    rd_cycle[ 9418] = 1'b0;  wr_cycle[ 9418] = 1'b0;  addr_rom[ 9418]='h00000000;  wr_data_rom[ 9418]='h00000000;
    rd_cycle[ 9419] = 1'b0;  wr_cycle[ 9419] = 1'b0;  addr_rom[ 9419]='h00000000;  wr_data_rom[ 9419]='h00000000;
    rd_cycle[ 9420] = 1'b0;  wr_cycle[ 9420] = 1'b0;  addr_rom[ 9420]='h00000000;  wr_data_rom[ 9420]='h00000000;
    rd_cycle[ 9421] = 1'b0;  wr_cycle[ 9421] = 1'b0;  addr_rom[ 9421]='h00000000;  wr_data_rom[ 9421]='h00000000;
    rd_cycle[ 9422] = 1'b0;  wr_cycle[ 9422] = 1'b0;  addr_rom[ 9422]='h00000000;  wr_data_rom[ 9422]='h00000000;
    rd_cycle[ 9423] = 1'b0;  wr_cycle[ 9423] = 1'b0;  addr_rom[ 9423]='h00000000;  wr_data_rom[ 9423]='h00000000;
    rd_cycle[ 9424] = 1'b0;  wr_cycle[ 9424] = 1'b0;  addr_rom[ 9424]='h00000000;  wr_data_rom[ 9424]='h00000000;
    rd_cycle[ 9425] = 1'b0;  wr_cycle[ 9425] = 1'b0;  addr_rom[ 9425]='h00000000;  wr_data_rom[ 9425]='h00000000;
    rd_cycle[ 9426] = 1'b0;  wr_cycle[ 9426] = 1'b0;  addr_rom[ 9426]='h00000000;  wr_data_rom[ 9426]='h00000000;
    rd_cycle[ 9427] = 1'b0;  wr_cycle[ 9427] = 1'b0;  addr_rom[ 9427]='h00000000;  wr_data_rom[ 9427]='h00000000;
    rd_cycle[ 9428] = 1'b0;  wr_cycle[ 9428] = 1'b0;  addr_rom[ 9428]='h00000000;  wr_data_rom[ 9428]='h00000000;
    rd_cycle[ 9429] = 1'b0;  wr_cycle[ 9429] = 1'b0;  addr_rom[ 9429]='h00000000;  wr_data_rom[ 9429]='h00000000;
    rd_cycle[ 9430] = 1'b0;  wr_cycle[ 9430] = 1'b0;  addr_rom[ 9430]='h00000000;  wr_data_rom[ 9430]='h00000000;
    rd_cycle[ 9431] = 1'b0;  wr_cycle[ 9431] = 1'b0;  addr_rom[ 9431]='h00000000;  wr_data_rom[ 9431]='h00000000;
    rd_cycle[ 9432] = 1'b0;  wr_cycle[ 9432] = 1'b0;  addr_rom[ 9432]='h00000000;  wr_data_rom[ 9432]='h00000000;
    rd_cycle[ 9433] = 1'b0;  wr_cycle[ 9433] = 1'b0;  addr_rom[ 9433]='h00000000;  wr_data_rom[ 9433]='h00000000;
    rd_cycle[ 9434] = 1'b0;  wr_cycle[ 9434] = 1'b0;  addr_rom[ 9434]='h00000000;  wr_data_rom[ 9434]='h00000000;
    rd_cycle[ 9435] = 1'b0;  wr_cycle[ 9435] = 1'b0;  addr_rom[ 9435]='h00000000;  wr_data_rom[ 9435]='h00000000;
    rd_cycle[ 9436] = 1'b0;  wr_cycle[ 9436] = 1'b0;  addr_rom[ 9436]='h00000000;  wr_data_rom[ 9436]='h00000000;
    rd_cycle[ 9437] = 1'b0;  wr_cycle[ 9437] = 1'b0;  addr_rom[ 9437]='h00000000;  wr_data_rom[ 9437]='h00000000;
    rd_cycle[ 9438] = 1'b0;  wr_cycle[ 9438] = 1'b0;  addr_rom[ 9438]='h00000000;  wr_data_rom[ 9438]='h00000000;
    rd_cycle[ 9439] = 1'b0;  wr_cycle[ 9439] = 1'b0;  addr_rom[ 9439]='h00000000;  wr_data_rom[ 9439]='h00000000;
    rd_cycle[ 9440] = 1'b0;  wr_cycle[ 9440] = 1'b0;  addr_rom[ 9440]='h00000000;  wr_data_rom[ 9440]='h00000000;
    rd_cycle[ 9441] = 1'b0;  wr_cycle[ 9441] = 1'b0;  addr_rom[ 9441]='h00000000;  wr_data_rom[ 9441]='h00000000;
    rd_cycle[ 9442] = 1'b0;  wr_cycle[ 9442] = 1'b0;  addr_rom[ 9442]='h00000000;  wr_data_rom[ 9442]='h00000000;
    rd_cycle[ 9443] = 1'b0;  wr_cycle[ 9443] = 1'b0;  addr_rom[ 9443]='h00000000;  wr_data_rom[ 9443]='h00000000;
    rd_cycle[ 9444] = 1'b0;  wr_cycle[ 9444] = 1'b0;  addr_rom[ 9444]='h00000000;  wr_data_rom[ 9444]='h00000000;
    rd_cycle[ 9445] = 1'b0;  wr_cycle[ 9445] = 1'b0;  addr_rom[ 9445]='h00000000;  wr_data_rom[ 9445]='h00000000;
    rd_cycle[ 9446] = 1'b0;  wr_cycle[ 9446] = 1'b0;  addr_rom[ 9446]='h00000000;  wr_data_rom[ 9446]='h00000000;
    rd_cycle[ 9447] = 1'b0;  wr_cycle[ 9447] = 1'b0;  addr_rom[ 9447]='h00000000;  wr_data_rom[ 9447]='h00000000;
    rd_cycle[ 9448] = 1'b0;  wr_cycle[ 9448] = 1'b0;  addr_rom[ 9448]='h00000000;  wr_data_rom[ 9448]='h00000000;
    rd_cycle[ 9449] = 1'b0;  wr_cycle[ 9449] = 1'b0;  addr_rom[ 9449]='h00000000;  wr_data_rom[ 9449]='h00000000;
    rd_cycle[ 9450] = 1'b0;  wr_cycle[ 9450] = 1'b0;  addr_rom[ 9450]='h00000000;  wr_data_rom[ 9450]='h00000000;
    rd_cycle[ 9451] = 1'b0;  wr_cycle[ 9451] = 1'b0;  addr_rom[ 9451]='h00000000;  wr_data_rom[ 9451]='h00000000;
    rd_cycle[ 9452] = 1'b0;  wr_cycle[ 9452] = 1'b0;  addr_rom[ 9452]='h00000000;  wr_data_rom[ 9452]='h00000000;
    rd_cycle[ 9453] = 1'b0;  wr_cycle[ 9453] = 1'b0;  addr_rom[ 9453]='h00000000;  wr_data_rom[ 9453]='h00000000;
    rd_cycle[ 9454] = 1'b0;  wr_cycle[ 9454] = 1'b0;  addr_rom[ 9454]='h00000000;  wr_data_rom[ 9454]='h00000000;
    rd_cycle[ 9455] = 1'b0;  wr_cycle[ 9455] = 1'b0;  addr_rom[ 9455]='h00000000;  wr_data_rom[ 9455]='h00000000;
    rd_cycle[ 9456] = 1'b0;  wr_cycle[ 9456] = 1'b0;  addr_rom[ 9456]='h00000000;  wr_data_rom[ 9456]='h00000000;
    rd_cycle[ 9457] = 1'b0;  wr_cycle[ 9457] = 1'b0;  addr_rom[ 9457]='h00000000;  wr_data_rom[ 9457]='h00000000;
    rd_cycle[ 9458] = 1'b0;  wr_cycle[ 9458] = 1'b0;  addr_rom[ 9458]='h00000000;  wr_data_rom[ 9458]='h00000000;
    rd_cycle[ 9459] = 1'b0;  wr_cycle[ 9459] = 1'b0;  addr_rom[ 9459]='h00000000;  wr_data_rom[ 9459]='h00000000;
    rd_cycle[ 9460] = 1'b0;  wr_cycle[ 9460] = 1'b0;  addr_rom[ 9460]='h00000000;  wr_data_rom[ 9460]='h00000000;
    rd_cycle[ 9461] = 1'b0;  wr_cycle[ 9461] = 1'b0;  addr_rom[ 9461]='h00000000;  wr_data_rom[ 9461]='h00000000;
    rd_cycle[ 9462] = 1'b0;  wr_cycle[ 9462] = 1'b0;  addr_rom[ 9462]='h00000000;  wr_data_rom[ 9462]='h00000000;
    rd_cycle[ 9463] = 1'b0;  wr_cycle[ 9463] = 1'b0;  addr_rom[ 9463]='h00000000;  wr_data_rom[ 9463]='h00000000;
    rd_cycle[ 9464] = 1'b0;  wr_cycle[ 9464] = 1'b0;  addr_rom[ 9464]='h00000000;  wr_data_rom[ 9464]='h00000000;
    rd_cycle[ 9465] = 1'b0;  wr_cycle[ 9465] = 1'b0;  addr_rom[ 9465]='h00000000;  wr_data_rom[ 9465]='h00000000;
    rd_cycle[ 9466] = 1'b0;  wr_cycle[ 9466] = 1'b0;  addr_rom[ 9466]='h00000000;  wr_data_rom[ 9466]='h00000000;
    rd_cycle[ 9467] = 1'b0;  wr_cycle[ 9467] = 1'b0;  addr_rom[ 9467]='h00000000;  wr_data_rom[ 9467]='h00000000;
    rd_cycle[ 9468] = 1'b0;  wr_cycle[ 9468] = 1'b0;  addr_rom[ 9468]='h00000000;  wr_data_rom[ 9468]='h00000000;
    rd_cycle[ 9469] = 1'b0;  wr_cycle[ 9469] = 1'b0;  addr_rom[ 9469]='h00000000;  wr_data_rom[ 9469]='h00000000;
    rd_cycle[ 9470] = 1'b0;  wr_cycle[ 9470] = 1'b0;  addr_rom[ 9470]='h00000000;  wr_data_rom[ 9470]='h00000000;
    rd_cycle[ 9471] = 1'b0;  wr_cycle[ 9471] = 1'b0;  addr_rom[ 9471]='h00000000;  wr_data_rom[ 9471]='h00000000;
    rd_cycle[ 9472] = 1'b0;  wr_cycle[ 9472] = 1'b0;  addr_rom[ 9472]='h00000000;  wr_data_rom[ 9472]='h00000000;
    rd_cycle[ 9473] = 1'b0;  wr_cycle[ 9473] = 1'b0;  addr_rom[ 9473]='h00000000;  wr_data_rom[ 9473]='h00000000;
    rd_cycle[ 9474] = 1'b0;  wr_cycle[ 9474] = 1'b0;  addr_rom[ 9474]='h00000000;  wr_data_rom[ 9474]='h00000000;
    rd_cycle[ 9475] = 1'b0;  wr_cycle[ 9475] = 1'b0;  addr_rom[ 9475]='h00000000;  wr_data_rom[ 9475]='h00000000;
    rd_cycle[ 9476] = 1'b0;  wr_cycle[ 9476] = 1'b0;  addr_rom[ 9476]='h00000000;  wr_data_rom[ 9476]='h00000000;
    rd_cycle[ 9477] = 1'b0;  wr_cycle[ 9477] = 1'b0;  addr_rom[ 9477]='h00000000;  wr_data_rom[ 9477]='h00000000;
    rd_cycle[ 9478] = 1'b0;  wr_cycle[ 9478] = 1'b0;  addr_rom[ 9478]='h00000000;  wr_data_rom[ 9478]='h00000000;
    rd_cycle[ 9479] = 1'b0;  wr_cycle[ 9479] = 1'b0;  addr_rom[ 9479]='h00000000;  wr_data_rom[ 9479]='h00000000;
    rd_cycle[ 9480] = 1'b0;  wr_cycle[ 9480] = 1'b0;  addr_rom[ 9480]='h00000000;  wr_data_rom[ 9480]='h00000000;
    rd_cycle[ 9481] = 1'b0;  wr_cycle[ 9481] = 1'b0;  addr_rom[ 9481]='h00000000;  wr_data_rom[ 9481]='h00000000;
    rd_cycle[ 9482] = 1'b0;  wr_cycle[ 9482] = 1'b0;  addr_rom[ 9482]='h00000000;  wr_data_rom[ 9482]='h00000000;
    rd_cycle[ 9483] = 1'b0;  wr_cycle[ 9483] = 1'b0;  addr_rom[ 9483]='h00000000;  wr_data_rom[ 9483]='h00000000;
    rd_cycle[ 9484] = 1'b0;  wr_cycle[ 9484] = 1'b0;  addr_rom[ 9484]='h00000000;  wr_data_rom[ 9484]='h00000000;
    rd_cycle[ 9485] = 1'b0;  wr_cycle[ 9485] = 1'b0;  addr_rom[ 9485]='h00000000;  wr_data_rom[ 9485]='h00000000;
    rd_cycle[ 9486] = 1'b0;  wr_cycle[ 9486] = 1'b0;  addr_rom[ 9486]='h00000000;  wr_data_rom[ 9486]='h00000000;
    rd_cycle[ 9487] = 1'b0;  wr_cycle[ 9487] = 1'b0;  addr_rom[ 9487]='h00000000;  wr_data_rom[ 9487]='h00000000;
    rd_cycle[ 9488] = 1'b0;  wr_cycle[ 9488] = 1'b0;  addr_rom[ 9488]='h00000000;  wr_data_rom[ 9488]='h00000000;
    rd_cycle[ 9489] = 1'b0;  wr_cycle[ 9489] = 1'b0;  addr_rom[ 9489]='h00000000;  wr_data_rom[ 9489]='h00000000;
    rd_cycle[ 9490] = 1'b0;  wr_cycle[ 9490] = 1'b0;  addr_rom[ 9490]='h00000000;  wr_data_rom[ 9490]='h00000000;
    rd_cycle[ 9491] = 1'b0;  wr_cycle[ 9491] = 1'b0;  addr_rom[ 9491]='h00000000;  wr_data_rom[ 9491]='h00000000;
    rd_cycle[ 9492] = 1'b0;  wr_cycle[ 9492] = 1'b0;  addr_rom[ 9492]='h00000000;  wr_data_rom[ 9492]='h00000000;
    rd_cycle[ 9493] = 1'b0;  wr_cycle[ 9493] = 1'b0;  addr_rom[ 9493]='h00000000;  wr_data_rom[ 9493]='h00000000;
    rd_cycle[ 9494] = 1'b0;  wr_cycle[ 9494] = 1'b0;  addr_rom[ 9494]='h00000000;  wr_data_rom[ 9494]='h00000000;
    rd_cycle[ 9495] = 1'b0;  wr_cycle[ 9495] = 1'b0;  addr_rom[ 9495]='h00000000;  wr_data_rom[ 9495]='h00000000;
    rd_cycle[ 9496] = 1'b0;  wr_cycle[ 9496] = 1'b0;  addr_rom[ 9496]='h00000000;  wr_data_rom[ 9496]='h00000000;
    rd_cycle[ 9497] = 1'b0;  wr_cycle[ 9497] = 1'b0;  addr_rom[ 9497]='h00000000;  wr_data_rom[ 9497]='h00000000;
    rd_cycle[ 9498] = 1'b0;  wr_cycle[ 9498] = 1'b0;  addr_rom[ 9498]='h00000000;  wr_data_rom[ 9498]='h00000000;
    rd_cycle[ 9499] = 1'b0;  wr_cycle[ 9499] = 1'b0;  addr_rom[ 9499]='h00000000;  wr_data_rom[ 9499]='h00000000;
    rd_cycle[ 9500] = 1'b0;  wr_cycle[ 9500] = 1'b0;  addr_rom[ 9500]='h00000000;  wr_data_rom[ 9500]='h00000000;
    rd_cycle[ 9501] = 1'b0;  wr_cycle[ 9501] = 1'b0;  addr_rom[ 9501]='h00000000;  wr_data_rom[ 9501]='h00000000;
    rd_cycle[ 9502] = 1'b0;  wr_cycle[ 9502] = 1'b0;  addr_rom[ 9502]='h00000000;  wr_data_rom[ 9502]='h00000000;
    rd_cycle[ 9503] = 1'b0;  wr_cycle[ 9503] = 1'b0;  addr_rom[ 9503]='h00000000;  wr_data_rom[ 9503]='h00000000;
    rd_cycle[ 9504] = 1'b0;  wr_cycle[ 9504] = 1'b0;  addr_rom[ 9504]='h00000000;  wr_data_rom[ 9504]='h00000000;
    rd_cycle[ 9505] = 1'b0;  wr_cycle[ 9505] = 1'b0;  addr_rom[ 9505]='h00000000;  wr_data_rom[ 9505]='h00000000;
    rd_cycle[ 9506] = 1'b0;  wr_cycle[ 9506] = 1'b0;  addr_rom[ 9506]='h00000000;  wr_data_rom[ 9506]='h00000000;
    rd_cycle[ 9507] = 1'b0;  wr_cycle[ 9507] = 1'b0;  addr_rom[ 9507]='h00000000;  wr_data_rom[ 9507]='h00000000;
    rd_cycle[ 9508] = 1'b0;  wr_cycle[ 9508] = 1'b0;  addr_rom[ 9508]='h00000000;  wr_data_rom[ 9508]='h00000000;
    rd_cycle[ 9509] = 1'b0;  wr_cycle[ 9509] = 1'b0;  addr_rom[ 9509]='h00000000;  wr_data_rom[ 9509]='h00000000;
    rd_cycle[ 9510] = 1'b0;  wr_cycle[ 9510] = 1'b0;  addr_rom[ 9510]='h00000000;  wr_data_rom[ 9510]='h00000000;
    rd_cycle[ 9511] = 1'b0;  wr_cycle[ 9511] = 1'b0;  addr_rom[ 9511]='h00000000;  wr_data_rom[ 9511]='h00000000;
    rd_cycle[ 9512] = 1'b0;  wr_cycle[ 9512] = 1'b0;  addr_rom[ 9512]='h00000000;  wr_data_rom[ 9512]='h00000000;
    rd_cycle[ 9513] = 1'b0;  wr_cycle[ 9513] = 1'b0;  addr_rom[ 9513]='h00000000;  wr_data_rom[ 9513]='h00000000;
    rd_cycle[ 9514] = 1'b0;  wr_cycle[ 9514] = 1'b0;  addr_rom[ 9514]='h00000000;  wr_data_rom[ 9514]='h00000000;
    rd_cycle[ 9515] = 1'b0;  wr_cycle[ 9515] = 1'b0;  addr_rom[ 9515]='h00000000;  wr_data_rom[ 9515]='h00000000;
    rd_cycle[ 9516] = 1'b0;  wr_cycle[ 9516] = 1'b0;  addr_rom[ 9516]='h00000000;  wr_data_rom[ 9516]='h00000000;
    rd_cycle[ 9517] = 1'b0;  wr_cycle[ 9517] = 1'b0;  addr_rom[ 9517]='h00000000;  wr_data_rom[ 9517]='h00000000;
    rd_cycle[ 9518] = 1'b0;  wr_cycle[ 9518] = 1'b0;  addr_rom[ 9518]='h00000000;  wr_data_rom[ 9518]='h00000000;
    rd_cycle[ 9519] = 1'b0;  wr_cycle[ 9519] = 1'b0;  addr_rom[ 9519]='h00000000;  wr_data_rom[ 9519]='h00000000;
    rd_cycle[ 9520] = 1'b0;  wr_cycle[ 9520] = 1'b0;  addr_rom[ 9520]='h00000000;  wr_data_rom[ 9520]='h00000000;
    rd_cycle[ 9521] = 1'b0;  wr_cycle[ 9521] = 1'b0;  addr_rom[ 9521]='h00000000;  wr_data_rom[ 9521]='h00000000;
    rd_cycle[ 9522] = 1'b0;  wr_cycle[ 9522] = 1'b0;  addr_rom[ 9522]='h00000000;  wr_data_rom[ 9522]='h00000000;
    rd_cycle[ 9523] = 1'b0;  wr_cycle[ 9523] = 1'b0;  addr_rom[ 9523]='h00000000;  wr_data_rom[ 9523]='h00000000;
    rd_cycle[ 9524] = 1'b0;  wr_cycle[ 9524] = 1'b0;  addr_rom[ 9524]='h00000000;  wr_data_rom[ 9524]='h00000000;
    rd_cycle[ 9525] = 1'b0;  wr_cycle[ 9525] = 1'b0;  addr_rom[ 9525]='h00000000;  wr_data_rom[ 9525]='h00000000;
    rd_cycle[ 9526] = 1'b0;  wr_cycle[ 9526] = 1'b0;  addr_rom[ 9526]='h00000000;  wr_data_rom[ 9526]='h00000000;
    rd_cycle[ 9527] = 1'b0;  wr_cycle[ 9527] = 1'b0;  addr_rom[ 9527]='h00000000;  wr_data_rom[ 9527]='h00000000;
    rd_cycle[ 9528] = 1'b0;  wr_cycle[ 9528] = 1'b0;  addr_rom[ 9528]='h00000000;  wr_data_rom[ 9528]='h00000000;
    rd_cycle[ 9529] = 1'b0;  wr_cycle[ 9529] = 1'b0;  addr_rom[ 9529]='h00000000;  wr_data_rom[ 9529]='h00000000;
    rd_cycle[ 9530] = 1'b0;  wr_cycle[ 9530] = 1'b0;  addr_rom[ 9530]='h00000000;  wr_data_rom[ 9530]='h00000000;
    rd_cycle[ 9531] = 1'b0;  wr_cycle[ 9531] = 1'b0;  addr_rom[ 9531]='h00000000;  wr_data_rom[ 9531]='h00000000;
    rd_cycle[ 9532] = 1'b0;  wr_cycle[ 9532] = 1'b0;  addr_rom[ 9532]='h00000000;  wr_data_rom[ 9532]='h00000000;
    rd_cycle[ 9533] = 1'b0;  wr_cycle[ 9533] = 1'b0;  addr_rom[ 9533]='h00000000;  wr_data_rom[ 9533]='h00000000;
    rd_cycle[ 9534] = 1'b0;  wr_cycle[ 9534] = 1'b0;  addr_rom[ 9534]='h00000000;  wr_data_rom[ 9534]='h00000000;
    rd_cycle[ 9535] = 1'b0;  wr_cycle[ 9535] = 1'b0;  addr_rom[ 9535]='h00000000;  wr_data_rom[ 9535]='h00000000;
    rd_cycle[ 9536] = 1'b0;  wr_cycle[ 9536] = 1'b0;  addr_rom[ 9536]='h00000000;  wr_data_rom[ 9536]='h00000000;
    rd_cycle[ 9537] = 1'b0;  wr_cycle[ 9537] = 1'b0;  addr_rom[ 9537]='h00000000;  wr_data_rom[ 9537]='h00000000;
    rd_cycle[ 9538] = 1'b0;  wr_cycle[ 9538] = 1'b0;  addr_rom[ 9538]='h00000000;  wr_data_rom[ 9538]='h00000000;
    rd_cycle[ 9539] = 1'b0;  wr_cycle[ 9539] = 1'b0;  addr_rom[ 9539]='h00000000;  wr_data_rom[ 9539]='h00000000;
    rd_cycle[ 9540] = 1'b0;  wr_cycle[ 9540] = 1'b0;  addr_rom[ 9540]='h00000000;  wr_data_rom[ 9540]='h00000000;
    rd_cycle[ 9541] = 1'b0;  wr_cycle[ 9541] = 1'b0;  addr_rom[ 9541]='h00000000;  wr_data_rom[ 9541]='h00000000;
    rd_cycle[ 9542] = 1'b0;  wr_cycle[ 9542] = 1'b0;  addr_rom[ 9542]='h00000000;  wr_data_rom[ 9542]='h00000000;
    rd_cycle[ 9543] = 1'b0;  wr_cycle[ 9543] = 1'b0;  addr_rom[ 9543]='h00000000;  wr_data_rom[ 9543]='h00000000;
    rd_cycle[ 9544] = 1'b0;  wr_cycle[ 9544] = 1'b0;  addr_rom[ 9544]='h00000000;  wr_data_rom[ 9544]='h00000000;
    rd_cycle[ 9545] = 1'b0;  wr_cycle[ 9545] = 1'b0;  addr_rom[ 9545]='h00000000;  wr_data_rom[ 9545]='h00000000;
    rd_cycle[ 9546] = 1'b0;  wr_cycle[ 9546] = 1'b0;  addr_rom[ 9546]='h00000000;  wr_data_rom[ 9546]='h00000000;
    rd_cycle[ 9547] = 1'b0;  wr_cycle[ 9547] = 1'b0;  addr_rom[ 9547]='h00000000;  wr_data_rom[ 9547]='h00000000;
    rd_cycle[ 9548] = 1'b0;  wr_cycle[ 9548] = 1'b0;  addr_rom[ 9548]='h00000000;  wr_data_rom[ 9548]='h00000000;
    rd_cycle[ 9549] = 1'b0;  wr_cycle[ 9549] = 1'b0;  addr_rom[ 9549]='h00000000;  wr_data_rom[ 9549]='h00000000;
    rd_cycle[ 9550] = 1'b0;  wr_cycle[ 9550] = 1'b0;  addr_rom[ 9550]='h00000000;  wr_data_rom[ 9550]='h00000000;
    rd_cycle[ 9551] = 1'b0;  wr_cycle[ 9551] = 1'b0;  addr_rom[ 9551]='h00000000;  wr_data_rom[ 9551]='h00000000;
    rd_cycle[ 9552] = 1'b0;  wr_cycle[ 9552] = 1'b0;  addr_rom[ 9552]='h00000000;  wr_data_rom[ 9552]='h00000000;
    rd_cycle[ 9553] = 1'b0;  wr_cycle[ 9553] = 1'b0;  addr_rom[ 9553]='h00000000;  wr_data_rom[ 9553]='h00000000;
    rd_cycle[ 9554] = 1'b0;  wr_cycle[ 9554] = 1'b0;  addr_rom[ 9554]='h00000000;  wr_data_rom[ 9554]='h00000000;
    rd_cycle[ 9555] = 1'b0;  wr_cycle[ 9555] = 1'b0;  addr_rom[ 9555]='h00000000;  wr_data_rom[ 9555]='h00000000;
    rd_cycle[ 9556] = 1'b0;  wr_cycle[ 9556] = 1'b0;  addr_rom[ 9556]='h00000000;  wr_data_rom[ 9556]='h00000000;
    rd_cycle[ 9557] = 1'b0;  wr_cycle[ 9557] = 1'b0;  addr_rom[ 9557]='h00000000;  wr_data_rom[ 9557]='h00000000;
    rd_cycle[ 9558] = 1'b0;  wr_cycle[ 9558] = 1'b0;  addr_rom[ 9558]='h00000000;  wr_data_rom[ 9558]='h00000000;
    rd_cycle[ 9559] = 1'b0;  wr_cycle[ 9559] = 1'b0;  addr_rom[ 9559]='h00000000;  wr_data_rom[ 9559]='h00000000;
    rd_cycle[ 9560] = 1'b0;  wr_cycle[ 9560] = 1'b0;  addr_rom[ 9560]='h00000000;  wr_data_rom[ 9560]='h00000000;
    rd_cycle[ 9561] = 1'b0;  wr_cycle[ 9561] = 1'b0;  addr_rom[ 9561]='h00000000;  wr_data_rom[ 9561]='h00000000;
    rd_cycle[ 9562] = 1'b0;  wr_cycle[ 9562] = 1'b0;  addr_rom[ 9562]='h00000000;  wr_data_rom[ 9562]='h00000000;
    rd_cycle[ 9563] = 1'b0;  wr_cycle[ 9563] = 1'b0;  addr_rom[ 9563]='h00000000;  wr_data_rom[ 9563]='h00000000;
    rd_cycle[ 9564] = 1'b0;  wr_cycle[ 9564] = 1'b0;  addr_rom[ 9564]='h00000000;  wr_data_rom[ 9564]='h00000000;
    rd_cycle[ 9565] = 1'b0;  wr_cycle[ 9565] = 1'b0;  addr_rom[ 9565]='h00000000;  wr_data_rom[ 9565]='h00000000;
    rd_cycle[ 9566] = 1'b0;  wr_cycle[ 9566] = 1'b0;  addr_rom[ 9566]='h00000000;  wr_data_rom[ 9566]='h00000000;
    rd_cycle[ 9567] = 1'b0;  wr_cycle[ 9567] = 1'b0;  addr_rom[ 9567]='h00000000;  wr_data_rom[ 9567]='h00000000;
    rd_cycle[ 9568] = 1'b0;  wr_cycle[ 9568] = 1'b0;  addr_rom[ 9568]='h00000000;  wr_data_rom[ 9568]='h00000000;
    rd_cycle[ 9569] = 1'b0;  wr_cycle[ 9569] = 1'b0;  addr_rom[ 9569]='h00000000;  wr_data_rom[ 9569]='h00000000;
    rd_cycle[ 9570] = 1'b0;  wr_cycle[ 9570] = 1'b0;  addr_rom[ 9570]='h00000000;  wr_data_rom[ 9570]='h00000000;
    rd_cycle[ 9571] = 1'b0;  wr_cycle[ 9571] = 1'b0;  addr_rom[ 9571]='h00000000;  wr_data_rom[ 9571]='h00000000;
    rd_cycle[ 9572] = 1'b0;  wr_cycle[ 9572] = 1'b0;  addr_rom[ 9572]='h00000000;  wr_data_rom[ 9572]='h00000000;
    rd_cycle[ 9573] = 1'b0;  wr_cycle[ 9573] = 1'b0;  addr_rom[ 9573]='h00000000;  wr_data_rom[ 9573]='h00000000;
    rd_cycle[ 9574] = 1'b0;  wr_cycle[ 9574] = 1'b0;  addr_rom[ 9574]='h00000000;  wr_data_rom[ 9574]='h00000000;
    rd_cycle[ 9575] = 1'b0;  wr_cycle[ 9575] = 1'b0;  addr_rom[ 9575]='h00000000;  wr_data_rom[ 9575]='h00000000;
    rd_cycle[ 9576] = 1'b0;  wr_cycle[ 9576] = 1'b0;  addr_rom[ 9576]='h00000000;  wr_data_rom[ 9576]='h00000000;
    rd_cycle[ 9577] = 1'b0;  wr_cycle[ 9577] = 1'b0;  addr_rom[ 9577]='h00000000;  wr_data_rom[ 9577]='h00000000;
    rd_cycle[ 9578] = 1'b0;  wr_cycle[ 9578] = 1'b0;  addr_rom[ 9578]='h00000000;  wr_data_rom[ 9578]='h00000000;
    rd_cycle[ 9579] = 1'b0;  wr_cycle[ 9579] = 1'b0;  addr_rom[ 9579]='h00000000;  wr_data_rom[ 9579]='h00000000;
    rd_cycle[ 9580] = 1'b0;  wr_cycle[ 9580] = 1'b0;  addr_rom[ 9580]='h00000000;  wr_data_rom[ 9580]='h00000000;
    rd_cycle[ 9581] = 1'b0;  wr_cycle[ 9581] = 1'b0;  addr_rom[ 9581]='h00000000;  wr_data_rom[ 9581]='h00000000;
    rd_cycle[ 9582] = 1'b0;  wr_cycle[ 9582] = 1'b0;  addr_rom[ 9582]='h00000000;  wr_data_rom[ 9582]='h00000000;
    rd_cycle[ 9583] = 1'b0;  wr_cycle[ 9583] = 1'b0;  addr_rom[ 9583]='h00000000;  wr_data_rom[ 9583]='h00000000;
    rd_cycle[ 9584] = 1'b0;  wr_cycle[ 9584] = 1'b0;  addr_rom[ 9584]='h00000000;  wr_data_rom[ 9584]='h00000000;
    rd_cycle[ 9585] = 1'b0;  wr_cycle[ 9585] = 1'b0;  addr_rom[ 9585]='h00000000;  wr_data_rom[ 9585]='h00000000;
    rd_cycle[ 9586] = 1'b0;  wr_cycle[ 9586] = 1'b0;  addr_rom[ 9586]='h00000000;  wr_data_rom[ 9586]='h00000000;
    rd_cycle[ 9587] = 1'b0;  wr_cycle[ 9587] = 1'b0;  addr_rom[ 9587]='h00000000;  wr_data_rom[ 9587]='h00000000;
    rd_cycle[ 9588] = 1'b0;  wr_cycle[ 9588] = 1'b0;  addr_rom[ 9588]='h00000000;  wr_data_rom[ 9588]='h00000000;
    rd_cycle[ 9589] = 1'b0;  wr_cycle[ 9589] = 1'b0;  addr_rom[ 9589]='h00000000;  wr_data_rom[ 9589]='h00000000;
    rd_cycle[ 9590] = 1'b0;  wr_cycle[ 9590] = 1'b0;  addr_rom[ 9590]='h00000000;  wr_data_rom[ 9590]='h00000000;
    rd_cycle[ 9591] = 1'b0;  wr_cycle[ 9591] = 1'b0;  addr_rom[ 9591]='h00000000;  wr_data_rom[ 9591]='h00000000;
    rd_cycle[ 9592] = 1'b0;  wr_cycle[ 9592] = 1'b0;  addr_rom[ 9592]='h00000000;  wr_data_rom[ 9592]='h00000000;
    rd_cycle[ 9593] = 1'b0;  wr_cycle[ 9593] = 1'b0;  addr_rom[ 9593]='h00000000;  wr_data_rom[ 9593]='h00000000;
    rd_cycle[ 9594] = 1'b0;  wr_cycle[ 9594] = 1'b0;  addr_rom[ 9594]='h00000000;  wr_data_rom[ 9594]='h00000000;
    rd_cycle[ 9595] = 1'b0;  wr_cycle[ 9595] = 1'b0;  addr_rom[ 9595]='h00000000;  wr_data_rom[ 9595]='h00000000;
    rd_cycle[ 9596] = 1'b0;  wr_cycle[ 9596] = 1'b0;  addr_rom[ 9596]='h00000000;  wr_data_rom[ 9596]='h00000000;
    rd_cycle[ 9597] = 1'b0;  wr_cycle[ 9597] = 1'b0;  addr_rom[ 9597]='h00000000;  wr_data_rom[ 9597]='h00000000;
    rd_cycle[ 9598] = 1'b0;  wr_cycle[ 9598] = 1'b0;  addr_rom[ 9598]='h00000000;  wr_data_rom[ 9598]='h00000000;
    rd_cycle[ 9599] = 1'b0;  wr_cycle[ 9599] = 1'b0;  addr_rom[ 9599]='h00000000;  wr_data_rom[ 9599]='h00000000;
    rd_cycle[ 9600] = 1'b0;  wr_cycle[ 9600] = 1'b0;  addr_rom[ 9600]='h00000000;  wr_data_rom[ 9600]='h00000000;
    rd_cycle[ 9601] = 1'b0;  wr_cycle[ 9601] = 1'b0;  addr_rom[ 9601]='h00000000;  wr_data_rom[ 9601]='h00000000;
    rd_cycle[ 9602] = 1'b0;  wr_cycle[ 9602] = 1'b0;  addr_rom[ 9602]='h00000000;  wr_data_rom[ 9602]='h00000000;
    rd_cycle[ 9603] = 1'b0;  wr_cycle[ 9603] = 1'b0;  addr_rom[ 9603]='h00000000;  wr_data_rom[ 9603]='h00000000;
    rd_cycle[ 9604] = 1'b0;  wr_cycle[ 9604] = 1'b0;  addr_rom[ 9604]='h00000000;  wr_data_rom[ 9604]='h00000000;
    rd_cycle[ 9605] = 1'b0;  wr_cycle[ 9605] = 1'b0;  addr_rom[ 9605]='h00000000;  wr_data_rom[ 9605]='h00000000;
    rd_cycle[ 9606] = 1'b0;  wr_cycle[ 9606] = 1'b0;  addr_rom[ 9606]='h00000000;  wr_data_rom[ 9606]='h00000000;
    rd_cycle[ 9607] = 1'b0;  wr_cycle[ 9607] = 1'b0;  addr_rom[ 9607]='h00000000;  wr_data_rom[ 9607]='h00000000;
    rd_cycle[ 9608] = 1'b0;  wr_cycle[ 9608] = 1'b0;  addr_rom[ 9608]='h00000000;  wr_data_rom[ 9608]='h00000000;
    rd_cycle[ 9609] = 1'b0;  wr_cycle[ 9609] = 1'b0;  addr_rom[ 9609]='h00000000;  wr_data_rom[ 9609]='h00000000;
    rd_cycle[ 9610] = 1'b0;  wr_cycle[ 9610] = 1'b0;  addr_rom[ 9610]='h00000000;  wr_data_rom[ 9610]='h00000000;
    rd_cycle[ 9611] = 1'b0;  wr_cycle[ 9611] = 1'b0;  addr_rom[ 9611]='h00000000;  wr_data_rom[ 9611]='h00000000;
    rd_cycle[ 9612] = 1'b0;  wr_cycle[ 9612] = 1'b0;  addr_rom[ 9612]='h00000000;  wr_data_rom[ 9612]='h00000000;
    rd_cycle[ 9613] = 1'b0;  wr_cycle[ 9613] = 1'b0;  addr_rom[ 9613]='h00000000;  wr_data_rom[ 9613]='h00000000;
    rd_cycle[ 9614] = 1'b0;  wr_cycle[ 9614] = 1'b0;  addr_rom[ 9614]='h00000000;  wr_data_rom[ 9614]='h00000000;
    rd_cycle[ 9615] = 1'b0;  wr_cycle[ 9615] = 1'b0;  addr_rom[ 9615]='h00000000;  wr_data_rom[ 9615]='h00000000;
    rd_cycle[ 9616] = 1'b0;  wr_cycle[ 9616] = 1'b0;  addr_rom[ 9616]='h00000000;  wr_data_rom[ 9616]='h00000000;
    rd_cycle[ 9617] = 1'b0;  wr_cycle[ 9617] = 1'b0;  addr_rom[ 9617]='h00000000;  wr_data_rom[ 9617]='h00000000;
    rd_cycle[ 9618] = 1'b0;  wr_cycle[ 9618] = 1'b0;  addr_rom[ 9618]='h00000000;  wr_data_rom[ 9618]='h00000000;
    rd_cycle[ 9619] = 1'b0;  wr_cycle[ 9619] = 1'b0;  addr_rom[ 9619]='h00000000;  wr_data_rom[ 9619]='h00000000;
    rd_cycle[ 9620] = 1'b0;  wr_cycle[ 9620] = 1'b0;  addr_rom[ 9620]='h00000000;  wr_data_rom[ 9620]='h00000000;
    rd_cycle[ 9621] = 1'b0;  wr_cycle[ 9621] = 1'b0;  addr_rom[ 9621]='h00000000;  wr_data_rom[ 9621]='h00000000;
    rd_cycle[ 9622] = 1'b0;  wr_cycle[ 9622] = 1'b0;  addr_rom[ 9622]='h00000000;  wr_data_rom[ 9622]='h00000000;
    rd_cycle[ 9623] = 1'b0;  wr_cycle[ 9623] = 1'b0;  addr_rom[ 9623]='h00000000;  wr_data_rom[ 9623]='h00000000;
    rd_cycle[ 9624] = 1'b0;  wr_cycle[ 9624] = 1'b0;  addr_rom[ 9624]='h00000000;  wr_data_rom[ 9624]='h00000000;
    rd_cycle[ 9625] = 1'b0;  wr_cycle[ 9625] = 1'b0;  addr_rom[ 9625]='h00000000;  wr_data_rom[ 9625]='h00000000;
    rd_cycle[ 9626] = 1'b0;  wr_cycle[ 9626] = 1'b0;  addr_rom[ 9626]='h00000000;  wr_data_rom[ 9626]='h00000000;
    rd_cycle[ 9627] = 1'b0;  wr_cycle[ 9627] = 1'b0;  addr_rom[ 9627]='h00000000;  wr_data_rom[ 9627]='h00000000;
    rd_cycle[ 9628] = 1'b0;  wr_cycle[ 9628] = 1'b0;  addr_rom[ 9628]='h00000000;  wr_data_rom[ 9628]='h00000000;
    rd_cycle[ 9629] = 1'b0;  wr_cycle[ 9629] = 1'b0;  addr_rom[ 9629]='h00000000;  wr_data_rom[ 9629]='h00000000;
    rd_cycle[ 9630] = 1'b0;  wr_cycle[ 9630] = 1'b0;  addr_rom[ 9630]='h00000000;  wr_data_rom[ 9630]='h00000000;
    rd_cycle[ 9631] = 1'b0;  wr_cycle[ 9631] = 1'b0;  addr_rom[ 9631]='h00000000;  wr_data_rom[ 9631]='h00000000;
    rd_cycle[ 9632] = 1'b0;  wr_cycle[ 9632] = 1'b0;  addr_rom[ 9632]='h00000000;  wr_data_rom[ 9632]='h00000000;
    rd_cycle[ 9633] = 1'b0;  wr_cycle[ 9633] = 1'b0;  addr_rom[ 9633]='h00000000;  wr_data_rom[ 9633]='h00000000;
    rd_cycle[ 9634] = 1'b0;  wr_cycle[ 9634] = 1'b0;  addr_rom[ 9634]='h00000000;  wr_data_rom[ 9634]='h00000000;
    rd_cycle[ 9635] = 1'b0;  wr_cycle[ 9635] = 1'b0;  addr_rom[ 9635]='h00000000;  wr_data_rom[ 9635]='h00000000;
    rd_cycle[ 9636] = 1'b0;  wr_cycle[ 9636] = 1'b0;  addr_rom[ 9636]='h00000000;  wr_data_rom[ 9636]='h00000000;
    rd_cycle[ 9637] = 1'b0;  wr_cycle[ 9637] = 1'b0;  addr_rom[ 9637]='h00000000;  wr_data_rom[ 9637]='h00000000;
    rd_cycle[ 9638] = 1'b0;  wr_cycle[ 9638] = 1'b0;  addr_rom[ 9638]='h00000000;  wr_data_rom[ 9638]='h00000000;
    rd_cycle[ 9639] = 1'b0;  wr_cycle[ 9639] = 1'b0;  addr_rom[ 9639]='h00000000;  wr_data_rom[ 9639]='h00000000;
    rd_cycle[ 9640] = 1'b0;  wr_cycle[ 9640] = 1'b0;  addr_rom[ 9640]='h00000000;  wr_data_rom[ 9640]='h00000000;
    rd_cycle[ 9641] = 1'b0;  wr_cycle[ 9641] = 1'b0;  addr_rom[ 9641]='h00000000;  wr_data_rom[ 9641]='h00000000;
    rd_cycle[ 9642] = 1'b0;  wr_cycle[ 9642] = 1'b0;  addr_rom[ 9642]='h00000000;  wr_data_rom[ 9642]='h00000000;
    rd_cycle[ 9643] = 1'b0;  wr_cycle[ 9643] = 1'b0;  addr_rom[ 9643]='h00000000;  wr_data_rom[ 9643]='h00000000;
    rd_cycle[ 9644] = 1'b0;  wr_cycle[ 9644] = 1'b0;  addr_rom[ 9644]='h00000000;  wr_data_rom[ 9644]='h00000000;
    rd_cycle[ 9645] = 1'b0;  wr_cycle[ 9645] = 1'b0;  addr_rom[ 9645]='h00000000;  wr_data_rom[ 9645]='h00000000;
    rd_cycle[ 9646] = 1'b0;  wr_cycle[ 9646] = 1'b0;  addr_rom[ 9646]='h00000000;  wr_data_rom[ 9646]='h00000000;
    rd_cycle[ 9647] = 1'b0;  wr_cycle[ 9647] = 1'b0;  addr_rom[ 9647]='h00000000;  wr_data_rom[ 9647]='h00000000;
    rd_cycle[ 9648] = 1'b0;  wr_cycle[ 9648] = 1'b0;  addr_rom[ 9648]='h00000000;  wr_data_rom[ 9648]='h00000000;
    rd_cycle[ 9649] = 1'b0;  wr_cycle[ 9649] = 1'b0;  addr_rom[ 9649]='h00000000;  wr_data_rom[ 9649]='h00000000;
    rd_cycle[ 9650] = 1'b0;  wr_cycle[ 9650] = 1'b0;  addr_rom[ 9650]='h00000000;  wr_data_rom[ 9650]='h00000000;
    rd_cycle[ 9651] = 1'b0;  wr_cycle[ 9651] = 1'b0;  addr_rom[ 9651]='h00000000;  wr_data_rom[ 9651]='h00000000;
    rd_cycle[ 9652] = 1'b0;  wr_cycle[ 9652] = 1'b0;  addr_rom[ 9652]='h00000000;  wr_data_rom[ 9652]='h00000000;
    rd_cycle[ 9653] = 1'b0;  wr_cycle[ 9653] = 1'b0;  addr_rom[ 9653]='h00000000;  wr_data_rom[ 9653]='h00000000;
    rd_cycle[ 9654] = 1'b0;  wr_cycle[ 9654] = 1'b0;  addr_rom[ 9654]='h00000000;  wr_data_rom[ 9654]='h00000000;
    rd_cycle[ 9655] = 1'b0;  wr_cycle[ 9655] = 1'b0;  addr_rom[ 9655]='h00000000;  wr_data_rom[ 9655]='h00000000;
    rd_cycle[ 9656] = 1'b0;  wr_cycle[ 9656] = 1'b0;  addr_rom[ 9656]='h00000000;  wr_data_rom[ 9656]='h00000000;
    rd_cycle[ 9657] = 1'b0;  wr_cycle[ 9657] = 1'b0;  addr_rom[ 9657]='h00000000;  wr_data_rom[ 9657]='h00000000;
    rd_cycle[ 9658] = 1'b0;  wr_cycle[ 9658] = 1'b0;  addr_rom[ 9658]='h00000000;  wr_data_rom[ 9658]='h00000000;
    rd_cycle[ 9659] = 1'b0;  wr_cycle[ 9659] = 1'b0;  addr_rom[ 9659]='h00000000;  wr_data_rom[ 9659]='h00000000;
    rd_cycle[ 9660] = 1'b0;  wr_cycle[ 9660] = 1'b0;  addr_rom[ 9660]='h00000000;  wr_data_rom[ 9660]='h00000000;
    rd_cycle[ 9661] = 1'b0;  wr_cycle[ 9661] = 1'b0;  addr_rom[ 9661]='h00000000;  wr_data_rom[ 9661]='h00000000;
    rd_cycle[ 9662] = 1'b0;  wr_cycle[ 9662] = 1'b0;  addr_rom[ 9662]='h00000000;  wr_data_rom[ 9662]='h00000000;
    rd_cycle[ 9663] = 1'b0;  wr_cycle[ 9663] = 1'b0;  addr_rom[ 9663]='h00000000;  wr_data_rom[ 9663]='h00000000;
    rd_cycle[ 9664] = 1'b0;  wr_cycle[ 9664] = 1'b0;  addr_rom[ 9664]='h00000000;  wr_data_rom[ 9664]='h00000000;
    rd_cycle[ 9665] = 1'b0;  wr_cycle[ 9665] = 1'b0;  addr_rom[ 9665]='h00000000;  wr_data_rom[ 9665]='h00000000;
    rd_cycle[ 9666] = 1'b0;  wr_cycle[ 9666] = 1'b0;  addr_rom[ 9666]='h00000000;  wr_data_rom[ 9666]='h00000000;
    rd_cycle[ 9667] = 1'b0;  wr_cycle[ 9667] = 1'b0;  addr_rom[ 9667]='h00000000;  wr_data_rom[ 9667]='h00000000;
    rd_cycle[ 9668] = 1'b0;  wr_cycle[ 9668] = 1'b0;  addr_rom[ 9668]='h00000000;  wr_data_rom[ 9668]='h00000000;
    rd_cycle[ 9669] = 1'b0;  wr_cycle[ 9669] = 1'b0;  addr_rom[ 9669]='h00000000;  wr_data_rom[ 9669]='h00000000;
    rd_cycle[ 9670] = 1'b0;  wr_cycle[ 9670] = 1'b0;  addr_rom[ 9670]='h00000000;  wr_data_rom[ 9670]='h00000000;
    rd_cycle[ 9671] = 1'b0;  wr_cycle[ 9671] = 1'b0;  addr_rom[ 9671]='h00000000;  wr_data_rom[ 9671]='h00000000;
    rd_cycle[ 9672] = 1'b0;  wr_cycle[ 9672] = 1'b0;  addr_rom[ 9672]='h00000000;  wr_data_rom[ 9672]='h00000000;
    rd_cycle[ 9673] = 1'b0;  wr_cycle[ 9673] = 1'b0;  addr_rom[ 9673]='h00000000;  wr_data_rom[ 9673]='h00000000;
    rd_cycle[ 9674] = 1'b0;  wr_cycle[ 9674] = 1'b0;  addr_rom[ 9674]='h00000000;  wr_data_rom[ 9674]='h00000000;
    rd_cycle[ 9675] = 1'b0;  wr_cycle[ 9675] = 1'b0;  addr_rom[ 9675]='h00000000;  wr_data_rom[ 9675]='h00000000;
    rd_cycle[ 9676] = 1'b0;  wr_cycle[ 9676] = 1'b0;  addr_rom[ 9676]='h00000000;  wr_data_rom[ 9676]='h00000000;
    rd_cycle[ 9677] = 1'b0;  wr_cycle[ 9677] = 1'b0;  addr_rom[ 9677]='h00000000;  wr_data_rom[ 9677]='h00000000;
    rd_cycle[ 9678] = 1'b0;  wr_cycle[ 9678] = 1'b0;  addr_rom[ 9678]='h00000000;  wr_data_rom[ 9678]='h00000000;
    rd_cycle[ 9679] = 1'b0;  wr_cycle[ 9679] = 1'b0;  addr_rom[ 9679]='h00000000;  wr_data_rom[ 9679]='h00000000;
    rd_cycle[ 9680] = 1'b0;  wr_cycle[ 9680] = 1'b0;  addr_rom[ 9680]='h00000000;  wr_data_rom[ 9680]='h00000000;
    rd_cycle[ 9681] = 1'b0;  wr_cycle[ 9681] = 1'b0;  addr_rom[ 9681]='h00000000;  wr_data_rom[ 9681]='h00000000;
    rd_cycle[ 9682] = 1'b0;  wr_cycle[ 9682] = 1'b0;  addr_rom[ 9682]='h00000000;  wr_data_rom[ 9682]='h00000000;
    rd_cycle[ 9683] = 1'b0;  wr_cycle[ 9683] = 1'b0;  addr_rom[ 9683]='h00000000;  wr_data_rom[ 9683]='h00000000;
    rd_cycle[ 9684] = 1'b0;  wr_cycle[ 9684] = 1'b0;  addr_rom[ 9684]='h00000000;  wr_data_rom[ 9684]='h00000000;
    rd_cycle[ 9685] = 1'b0;  wr_cycle[ 9685] = 1'b0;  addr_rom[ 9685]='h00000000;  wr_data_rom[ 9685]='h00000000;
    rd_cycle[ 9686] = 1'b0;  wr_cycle[ 9686] = 1'b0;  addr_rom[ 9686]='h00000000;  wr_data_rom[ 9686]='h00000000;
    rd_cycle[ 9687] = 1'b0;  wr_cycle[ 9687] = 1'b0;  addr_rom[ 9687]='h00000000;  wr_data_rom[ 9687]='h00000000;
    rd_cycle[ 9688] = 1'b0;  wr_cycle[ 9688] = 1'b0;  addr_rom[ 9688]='h00000000;  wr_data_rom[ 9688]='h00000000;
    rd_cycle[ 9689] = 1'b0;  wr_cycle[ 9689] = 1'b0;  addr_rom[ 9689]='h00000000;  wr_data_rom[ 9689]='h00000000;
    rd_cycle[ 9690] = 1'b0;  wr_cycle[ 9690] = 1'b0;  addr_rom[ 9690]='h00000000;  wr_data_rom[ 9690]='h00000000;
    rd_cycle[ 9691] = 1'b0;  wr_cycle[ 9691] = 1'b0;  addr_rom[ 9691]='h00000000;  wr_data_rom[ 9691]='h00000000;
    rd_cycle[ 9692] = 1'b0;  wr_cycle[ 9692] = 1'b0;  addr_rom[ 9692]='h00000000;  wr_data_rom[ 9692]='h00000000;
    rd_cycle[ 9693] = 1'b0;  wr_cycle[ 9693] = 1'b0;  addr_rom[ 9693]='h00000000;  wr_data_rom[ 9693]='h00000000;
    rd_cycle[ 9694] = 1'b0;  wr_cycle[ 9694] = 1'b0;  addr_rom[ 9694]='h00000000;  wr_data_rom[ 9694]='h00000000;
    rd_cycle[ 9695] = 1'b0;  wr_cycle[ 9695] = 1'b0;  addr_rom[ 9695]='h00000000;  wr_data_rom[ 9695]='h00000000;
    rd_cycle[ 9696] = 1'b0;  wr_cycle[ 9696] = 1'b0;  addr_rom[ 9696]='h00000000;  wr_data_rom[ 9696]='h00000000;
    rd_cycle[ 9697] = 1'b0;  wr_cycle[ 9697] = 1'b0;  addr_rom[ 9697]='h00000000;  wr_data_rom[ 9697]='h00000000;
    rd_cycle[ 9698] = 1'b0;  wr_cycle[ 9698] = 1'b0;  addr_rom[ 9698]='h00000000;  wr_data_rom[ 9698]='h00000000;
    rd_cycle[ 9699] = 1'b0;  wr_cycle[ 9699] = 1'b0;  addr_rom[ 9699]='h00000000;  wr_data_rom[ 9699]='h00000000;
    rd_cycle[ 9700] = 1'b0;  wr_cycle[ 9700] = 1'b0;  addr_rom[ 9700]='h00000000;  wr_data_rom[ 9700]='h00000000;
    rd_cycle[ 9701] = 1'b0;  wr_cycle[ 9701] = 1'b0;  addr_rom[ 9701]='h00000000;  wr_data_rom[ 9701]='h00000000;
    rd_cycle[ 9702] = 1'b0;  wr_cycle[ 9702] = 1'b0;  addr_rom[ 9702]='h00000000;  wr_data_rom[ 9702]='h00000000;
    rd_cycle[ 9703] = 1'b0;  wr_cycle[ 9703] = 1'b0;  addr_rom[ 9703]='h00000000;  wr_data_rom[ 9703]='h00000000;
    rd_cycle[ 9704] = 1'b0;  wr_cycle[ 9704] = 1'b0;  addr_rom[ 9704]='h00000000;  wr_data_rom[ 9704]='h00000000;
    rd_cycle[ 9705] = 1'b0;  wr_cycle[ 9705] = 1'b0;  addr_rom[ 9705]='h00000000;  wr_data_rom[ 9705]='h00000000;
    rd_cycle[ 9706] = 1'b0;  wr_cycle[ 9706] = 1'b0;  addr_rom[ 9706]='h00000000;  wr_data_rom[ 9706]='h00000000;
    rd_cycle[ 9707] = 1'b0;  wr_cycle[ 9707] = 1'b0;  addr_rom[ 9707]='h00000000;  wr_data_rom[ 9707]='h00000000;
    rd_cycle[ 9708] = 1'b0;  wr_cycle[ 9708] = 1'b0;  addr_rom[ 9708]='h00000000;  wr_data_rom[ 9708]='h00000000;
    rd_cycle[ 9709] = 1'b0;  wr_cycle[ 9709] = 1'b0;  addr_rom[ 9709]='h00000000;  wr_data_rom[ 9709]='h00000000;
    rd_cycle[ 9710] = 1'b0;  wr_cycle[ 9710] = 1'b0;  addr_rom[ 9710]='h00000000;  wr_data_rom[ 9710]='h00000000;
    rd_cycle[ 9711] = 1'b0;  wr_cycle[ 9711] = 1'b0;  addr_rom[ 9711]='h00000000;  wr_data_rom[ 9711]='h00000000;
    rd_cycle[ 9712] = 1'b0;  wr_cycle[ 9712] = 1'b0;  addr_rom[ 9712]='h00000000;  wr_data_rom[ 9712]='h00000000;
    rd_cycle[ 9713] = 1'b0;  wr_cycle[ 9713] = 1'b0;  addr_rom[ 9713]='h00000000;  wr_data_rom[ 9713]='h00000000;
    rd_cycle[ 9714] = 1'b0;  wr_cycle[ 9714] = 1'b0;  addr_rom[ 9714]='h00000000;  wr_data_rom[ 9714]='h00000000;
    rd_cycle[ 9715] = 1'b0;  wr_cycle[ 9715] = 1'b0;  addr_rom[ 9715]='h00000000;  wr_data_rom[ 9715]='h00000000;
    rd_cycle[ 9716] = 1'b0;  wr_cycle[ 9716] = 1'b0;  addr_rom[ 9716]='h00000000;  wr_data_rom[ 9716]='h00000000;
    rd_cycle[ 9717] = 1'b0;  wr_cycle[ 9717] = 1'b0;  addr_rom[ 9717]='h00000000;  wr_data_rom[ 9717]='h00000000;
    rd_cycle[ 9718] = 1'b0;  wr_cycle[ 9718] = 1'b0;  addr_rom[ 9718]='h00000000;  wr_data_rom[ 9718]='h00000000;
    rd_cycle[ 9719] = 1'b0;  wr_cycle[ 9719] = 1'b0;  addr_rom[ 9719]='h00000000;  wr_data_rom[ 9719]='h00000000;
    rd_cycle[ 9720] = 1'b0;  wr_cycle[ 9720] = 1'b0;  addr_rom[ 9720]='h00000000;  wr_data_rom[ 9720]='h00000000;
    rd_cycle[ 9721] = 1'b0;  wr_cycle[ 9721] = 1'b0;  addr_rom[ 9721]='h00000000;  wr_data_rom[ 9721]='h00000000;
    rd_cycle[ 9722] = 1'b0;  wr_cycle[ 9722] = 1'b0;  addr_rom[ 9722]='h00000000;  wr_data_rom[ 9722]='h00000000;
    rd_cycle[ 9723] = 1'b0;  wr_cycle[ 9723] = 1'b0;  addr_rom[ 9723]='h00000000;  wr_data_rom[ 9723]='h00000000;
    rd_cycle[ 9724] = 1'b0;  wr_cycle[ 9724] = 1'b0;  addr_rom[ 9724]='h00000000;  wr_data_rom[ 9724]='h00000000;
    rd_cycle[ 9725] = 1'b0;  wr_cycle[ 9725] = 1'b0;  addr_rom[ 9725]='h00000000;  wr_data_rom[ 9725]='h00000000;
    rd_cycle[ 9726] = 1'b0;  wr_cycle[ 9726] = 1'b0;  addr_rom[ 9726]='h00000000;  wr_data_rom[ 9726]='h00000000;
    rd_cycle[ 9727] = 1'b0;  wr_cycle[ 9727] = 1'b0;  addr_rom[ 9727]='h00000000;  wr_data_rom[ 9727]='h00000000;
    rd_cycle[ 9728] = 1'b0;  wr_cycle[ 9728] = 1'b0;  addr_rom[ 9728]='h00000000;  wr_data_rom[ 9728]='h00000000;
    rd_cycle[ 9729] = 1'b0;  wr_cycle[ 9729] = 1'b0;  addr_rom[ 9729]='h00000000;  wr_data_rom[ 9729]='h00000000;
    rd_cycle[ 9730] = 1'b0;  wr_cycle[ 9730] = 1'b0;  addr_rom[ 9730]='h00000000;  wr_data_rom[ 9730]='h00000000;
    rd_cycle[ 9731] = 1'b0;  wr_cycle[ 9731] = 1'b0;  addr_rom[ 9731]='h00000000;  wr_data_rom[ 9731]='h00000000;
    rd_cycle[ 9732] = 1'b0;  wr_cycle[ 9732] = 1'b0;  addr_rom[ 9732]='h00000000;  wr_data_rom[ 9732]='h00000000;
    rd_cycle[ 9733] = 1'b0;  wr_cycle[ 9733] = 1'b0;  addr_rom[ 9733]='h00000000;  wr_data_rom[ 9733]='h00000000;
    rd_cycle[ 9734] = 1'b0;  wr_cycle[ 9734] = 1'b0;  addr_rom[ 9734]='h00000000;  wr_data_rom[ 9734]='h00000000;
    rd_cycle[ 9735] = 1'b0;  wr_cycle[ 9735] = 1'b0;  addr_rom[ 9735]='h00000000;  wr_data_rom[ 9735]='h00000000;
    rd_cycle[ 9736] = 1'b0;  wr_cycle[ 9736] = 1'b0;  addr_rom[ 9736]='h00000000;  wr_data_rom[ 9736]='h00000000;
    rd_cycle[ 9737] = 1'b0;  wr_cycle[ 9737] = 1'b0;  addr_rom[ 9737]='h00000000;  wr_data_rom[ 9737]='h00000000;
    rd_cycle[ 9738] = 1'b0;  wr_cycle[ 9738] = 1'b0;  addr_rom[ 9738]='h00000000;  wr_data_rom[ 9738]='h00000000;
    rd_cycle[ 9739] = 1'b0;  wr_cycle[ 9739] = 1'b0;  addr_rom[ 9739]='h00000000;  wr_data_rom[ 9739]='h00000000;
    rd_cycle[ 9740] = 1'b0;  wr_cycle[ 9740] = 1'b0;  addr_rom[ 9740]='h00000000;  wr_data_rom[ 9740]='h00000000;
    rd_cycle[ 9741] = 1'b0;  wr_cycle[ 9741] = 1'b0;  addr_rom[ 9741]='h00000000;  wr_data_rom[ 9741]='h00000000;
    rd_cycle[ 9742] = 1'b0;  wr_cycle[ 9742] = 1'b0;  addr_rom[ 9742]='h00000000;  wr_data_rom[ 9742]='h00000000;
    rd_cycle[ 9743] = 1'b0;  wr_cycle[ 9743] = 1'b0;  addr_rom[ 9743]='h00000000;  wr_data_rom[ 9743]='h00000000;
    rd_cycle[ 9744] = 1'b0;  wr_cycle[ 9744] = 1'b0;  addr_rom[ 9744]='h00000000;  wr_data_rom[ 9744]='h00000000;
    rd_cycle[ 9745] = 1'b0;  wr_cycle[ 9745] = 1'b0;  addr_rom[ 9745]='h00000000;  wr_data_rom[ 9745]='h00000000;
    rd_cycle[ 9746] = 1'b0;  wr_cycle[ 9746] = 1'b0;  addr_rom[ 9746]='h00000000;  wr_data_rom[ 9746]='h00000000;
    rd_cycle[ 9747] = 1'b0;  wr_cycle[ 9747] = 1'b0;  addr_rom[ 9747]='h00000000;  wr_data_rom[ 9747]='h00000000;
    rd_cycle[ 9748] = 1'b0;  wr_cycle[ 9748] = 1'b0;  addr_rom[ 9748]='h00000000;  wr_data_rom[ 9748]='h00000000;
    rd_cycle[ 9749] = 1'b0;  wr_cycle[ 9749] = 1'b0;  addr_rom[ 9749]='h00000000;  wr_data_rom[ 9749]='h00000000;
    rd_cycle[ 9750] = 1'b0;  wr_cycle[ 9750] = 1'b0;  addr_rom[ 9750]='h00000000;  wr_data_rom[ 9750]='h00000000;
    rd_cycle[ 9751] = 1'b0;  wr_cycle[ 9751] = 1'b0;  addr_rom[ 9751]='h00000000;  wr_data_rom[ 9751]='h00000000;
    rd_cycle[ 9752] = 1'b0;  wr_cycle[ 9752] = 1'b0;  addr_rom[ 9752]='h00000000;  wr_data_rom[ 9752]='h00000000;
    rd_cycle[ 9753] = 1'b0;  wr_cycle[ 9753] = 1'b0;  addr_rom[ 9753]='h00000000;  wr_data_rom[ 9753]='h00000000;
    rd_cycle[ 9754] = 1'b0;  wr_cycle[ 9754] = 1'b0;  addr_rom[ 9754]='h00000000;  wr_data_rom[ 9754]='h00000000;
    rd_cycle[ 9755] = 1'b0;  wr_cycle[ 9755] = 1'b0;  addr_rom[ 9755]='h00000000;  wr_data_rom[ 9755]='h00000000;
    rd_cycle[ 9756] = 1'b0;  wr_cycle[ 9756] = 1'b0;  addr_rom[ 9756]='h00000000;  wr_data_rom[ 9756]='h00000000;
    rd_cycle[ 9757] = 1'b0;  wr_cycle[ 9757] = 1'b0;  addr_rom[ 9757]='h00000000;  wr_data_rom[ 9757]='h00000000;
    rd_cycle[ 9758] = 1'b0;  wr_cycle[ 9758] = 1'b0;  addr_rom[ 9758]='h00000000;  wr_data_rom[ 9758]='h00000000;
    rd_cycle[ 9759] = 1'b0;  wr_cycle[ 9759] = 1'b0;  addr_rom[ 9759]='h00000000;  wr_data_rom[ 9759]='h00000000;
    rd_cycle[ 9760] = 1'b0;  wr_cycle[ 9760] = 1'b0;  addr_rom[ 9760]='h00000000;  wr_data_rom[ 9760]='h00000000;
    rd_cycle[ 9761] = 1'b0;  wr_cycle[ 9761] = 1'b0;  addr_rom[ 9761]='h00000000;  wr_data_rom[ 9761]='h00000000;
    rd_cycle[ 9762] = 1'b0;  wr_cycle[ 9762] = 1'b0;  addr_rom[ 9762]='h00000000;  wr_data_rom[ 9762]='h00000000;
    rd_cycle[ 9763] = 1'b0;  wr_cycle[ 9763] = 1'b0;  addr_rom[ 9763]='h00000000;  wr_data_rom[ 9763]='h00000000;
    rd_cycle[ 9764] = 1'b0;  wr_cycle[ 9764] = 1'b0;  addr_rom[ 9764]='h00000000;  wr_data_rom[ 9764]='h00000000;
    rd_cycle[ 9765] = 1'b0;  wr_cycle[ 9765] = 1'b0;  addr_rom[ 9765]='h00000000;  wr_data_rom[ 9765]='h00000000;
    rd_cycle[ 9766] = 1'b0;  wr_cycle[ 9766] = 1'b0;  addr_rom[ 9766]='h00000000;  wr_data_rom[ 9766]='h00000000;
    rd_cycle[ 9767] = 1'b0;  wr_cycle[ 9767] = 1'b0;  addr_rom[ 9767]='h00000000;  wr_data_rom[ 9767]='h00000000;
    rd_cycle[ 9768] = 1'b0;  wr_cycle[ 9768] = 1'b0;  addr_rom[ 9768]='h00000000;  wr_data_rom[ 9768]='h00000000;
    rd_cycle[ 9769] = 1'b0;  wr_cycle[ 9769] = 1'b0;  addr_rom[ 9769]='h00000000;  wr_data_rom[ 9769]='h00000000;
    rd_cycle[ 9770] = 1'b0;  wr_cycle[ 9770] = 1'b0;  addr_rom[ 9770]='h00000000;  wr_data_rom[ 9770]='h00000000;
    rd_cycle[ 9771] = 1'b0;  wr_cycle[ 9771] = 1'b0;  addr_rom[ 9771]='h00000000;  wr_data_rom[ 9771]='h00000000;
    rd_cycle[ 9772] = 1'b0;  wr_cycle[ 9772] = 1'b0;  addr_rom[ 9772]='h00000000;  wr_data_rom[ 9772]='h00000000;
    rd_cycle[ 9773] = 1'b0;  wr_cycle[ 9773] = 1'b0;  addr_rom[ 9773]='h00000000;  wr_data_rom[ 9773]='h00000000;
    rd_cycle[ 9774] = 1'b0;  wr_cycle[ 9774] = 1'b0;  addr_rom[ 9774]='h00000000;  wr_data_rom[ 9774]='h00000000;
    rd_cycle[ 9775] = 1'b0;  wr_cycle[ 9775] = 1'b0;  addr_rom[ 9775]='h00000000;  wr_data_rom[ 9775]='h00000000;
    rd_cycle[ 9776] = 1'b0;  wr_cycle[ 9776] = 1'b0;  addr_rom[ 9776]='h00000000;  wr_data_rom[ 9776]='h00000000;
    rd_cycle[ 9777] = 1'b0;  wr_cycle[ 9777] = 1'b0;  addr_rom[ 9777]='h00000000;  wr_data_rom[ 9777]='h00000000;
    rd_cycle[ 9778] = 1'b0;  wr_cycle[ 9778] = 1'b0;  addr_rom[ 9778]='h00000000;  wr_data_rom[ 9778]='h00000000;
    rd_cycle[ 9779] = 1'b0;  wr_cycle[ 9779] = 1'b0;  addr_rom[ 9779]='h00000000;  wr_data_rom[ 9779]='h00000000;
    rd_cycle[ 9780] = 1'b0;  wr_cycle[ 9780] = 1'b0;  addr_rom[ 9780]='h00000000;  wr_data_rom[ 9780]='h00000000;
    rd_cycle[ 9781] = 1'b0;  wr_cycle[ 9781] = 1'b0;  addr_rom[ 9781]='h00000000;  wr_data_rom[ 9781]='h00000000;
    rd_cycle[ 9782] = 1'b0;  wr_cycle[ 9782] = 1'b0;  addr_rom[ 9782]='h00000000;  wr_data_rom[ 9782]='h00000000;
    rd_cycle[ 9783] = 1'b0;  wr_cycle[ 9783] = 1'b0;  addr_rom[ 9783]='h00000000;  wr_data_rom[ 9783]='h00000000;
    rd_cycle[ 9784] = 1'b0;  wr_cycle[ 9784] = 1'b0;  addr_rom[ 9784]='h00000000;  wr_data_rom[ 9784]='h00000000;
    rd_cycle[ 9785] = 1'b0;  wr_cycle[ 9785] = 1'b0;  addr_rom[ 9785]='h00000000;  wr_data_rom[ 9785]='h00000000;
    rd_cycle[ 9786] = 1'b0;  wr_cycle[ 9786] = 1'b0;  addr_rom[ 9786]='h00000000;  wr_data_rom[ 9786]='h00000000;
    rd_cycle[ 9787] = 1'b0;  wr_cycle[ 9787] = 1'b0;  addr_rom[ 9787]='h00000000;  wr_data_rom[ 9787]='h00000000;
    rd_cycle[ 9788] = 1'b0;  wr_cycle[ 9788] = 1'b0;  addr_rom[ 9788]='h00000000;  wr_data_rom[ 9788]='h00000000;
    rd_cycle[ 9789] = 1'b0;  wr_cycle[ 9789] = 1'b0;  addr_rom[ 9789]='h00000000;  wr_data_rom[ 9789]='h00000000;
    rd_cycle[ 9790] = 1'b0;  wr_cycle[ 9790] = 1'b0;  addr_rom[ 9790]='h00000000;  wr_data_rom[ 9790]='h00000000;
    rd_cycle[ 9791] = 1'b0;  wr_cycle[ 9791] = 1'b0;  addr_rom[ 9791]='h00000000;  wr_data_rom[ 9791]='h00000000;
    rd_cycle[ 9792] = 1'b0;  wr_cycle[ 9792] = 1'b0;  addr_rom[ 9792]='h00000000;  wr_data_rom[ 9792]='h00000000;
    rd_cycle[ 9793] = 1'b0;  wr_cycle[ 9793] = 1'b0;  addr_rom[ 9793]='h00000000;  wr_data_rom[ 9793]='h00000000;
    rd_cycle[ 9794] = 1'b0;  wr_cycle[ 9794] = 1'b0;  addr_rom[ 9794]='h00000000;  wr_data_rom[ 9794]='h00000000;
    rd_cycle[ 9795] = 1'b0;  wr_cycle[ 9795] = 1'b0;  addr_rom[ 9795]='h00000000;  wr_data_rom[ 9795]='h00000000;
    rd_cycle[ 9796] = 1'b0;  wr_cycle[ 9796] = 1'b0;  addr_rom[ 9796]='h00000000;  wr_data_rom[ 9796]='h00000000;
    rd_cycle[ 9797] = 1'b0;  wr_cycle[ 9797] = 1'b0;  addr_rom[ 9797]='h00000000;  wr_data_rom[ 9797]='h00000000;
    rd_cycle[ 9798] = 1'b0;  wr_cycle[ 9798] = 1'b0;  addr_rom[ 9798]='h00000000;  wr_data_rom[ 9798]='h00000000;
    rd_cycle[ 9799] = 1'b0;  wr_cycle[ 9799] = 1'b0;  addr_rom[ 9799]='h00000000;  wr_data_rom[ 9799]='h00000000;
    rd_cycle[ 9800] = 1'b0;  wr_cycle[ 9800] = 1'b0;  addr_rom[ 9800]='h00000000;  wr_data_rom[ 9800]='h00000000;
    rd_cycle[ 9801] = 1'b0;  wr_cycle[ 9801] = 1'b0;  addr_rom[ 9801]='h00000000;  wr_data_rom[ 9801]='h00000000;
    rd_cycle[ 9802] = 1'b0;  wr_cycle[ 9802] = 1'b0;  addr_rom[ 9802]='h00000000;  wr_data_rom[ 9802]='h00000000;
    rd_cycle[ 9803] = 1'b0;  wr_cycle[ 9803] = 1'b0;  addr_rom[ 9803]='h00000000;  wr_data_rom[ 9803]='h00000000;
    rd_cycle[ 9804] = 1'b0;  wr_cycle[ 9804] = 1'b0;  addr_rom[ 9804]='h00000000;  wr_data_rom[ 9804]='h00000000;
    rd_cycle[ 9805] = 1'b0;  wr_cycle[ 9805] = 1'b0;  addr_rom[ 9805]='h00000000;  wr_data_rom[ 9805]='h00000000;
    rd_cycle[ 9806] = 1'b0;  wr_cycle[ 9806] = 1'b0;  addr_rom[ 9806]='h00000000;  wr_data_rom[ 9806]='h00000000;
    rd_cycle[ 9807] = 1'b0;  wr_cycle[ 9807] = 1'b0;  addr_rom[ 9807]='h00000000;  wr_data_rom[ 9807]='h00000000;
    rd_cycle[ 9808] = 1'b0;  wr_cycle[ 9808] = 1'b0;  addr_rom[ 9808]='h00000000;  wr_data_rom[ 9808]='h00000000;
    rd_cycle[ 9809] = 1'b0;  wr_cycle[ 9809] = 1'b0;  addr_rom[ 9809]='h00000000;  wr_data_rom[ 9809]='h00000000;
    rd_cycle[ 9810] = 1'b0;  wr_cycle[ 9810] = 1'b0;  addr_rom[ 9810]='h00000000;  wr_data_rom[ 9810]='h00000000;
    rd_cycle[ 9811] = 1'b0;  wr_cycle[ 9811] = 1'b0;  addr_rom[ 9811]='h00000000;  wr_data_rom[ 9811]='h00000000;
    rd_cycle[ 9812] = 1'b0;  wr_cycle[ 9812] = 1'b0;  addr_rom[ 9812]='h00000000;  wr_data_rom[ 9812]='h00000000;
    rd_cycle[ 9813] = 1'b0;  wr_cycle[ 9813] = 1'b0;  addr_rom[ 9813]='h00000000;  wr_data_rom[ 9813]='h00000000;
    rd_cycle[ 9814] = 1'b0;  wr_cycle[ 9814] = 1'b0;  addr_rom[ 9814]='h00000000;  wr_data_rom[ 9814]='h00000000;
    rd_cycle[ 9815] = 1'b0;  wr_cycle[ 9815] = 1'b0;  addr_rom[ 9815]='h00000000;  wr_data_rom[ 9815]='h00000000;
    rd_cycle[ 9816] = 1'b0;  wr_cycle[ 9816] = 1'b0;  addr_rom[ 9816]='h00000000;  wr_data_rom[ 9816]='h00000000;
    rd_cycle[ 9817] = 1'b0;  wr_cycle[ 9817] = 1'b0;  addr_rom[ 9817]='h00000000;  wr_data_rom[ 9817]='h00000000;
    rd_cycle[ 9818] = 1'b0;  wr_cycle[ 9818] = 1'b0;  addr_rom[ 9818]='h00000000;  wr_data_rom[ 9818]='h00000000;
    rd_cycle[ 9819] = 1'b0;  wr_cycle[ 9819] = 1'b0;  addr_rom[ 9819]='h00000000;  wr_data_rom[ 9819]='h00000000;
    rd_cycle[ 9820] = 1'b0;  wr_cycle[ 9820] = 1'b0;  addr_rom[ 9820]='h00000000;  wr_data_rom[ 9820]='h00000000;
    rd_cycle[ 9821] = 1'b0;  wr_cycle[ 9821] = 1'b0;  addr_rom[ 9821]='h00000000;  wr_data_rom[ 9821]='h00000000;
    rd_cycle[ 9822] = 1'b0;  wr_cycle[ 9822] = 1'b0;  addr_rom[ 9822]='h00000000;  wr_data_rom[ 9822]='h00000000;
    rd_cycle[ 9823] = 1'b0;  wr_cycle[ 9823] = 1'b0;  addr_rom[ 9823]='h00000000;  wr_data_rom[ 9823]='h00000000;
    rd_cycle[ 9824] = 1'b0;  wr_cycle[ 9824] = 1'b0;  addr_rom[ 9824]='h00000000;  wr_data_rom[ 9824]='h00000000;
    rd_cycle[ 9825] = 1'b0;  wr_cycle[ 9825] = 1'b0;  addr_rom[ 9825]='h00000000;  wr_data_rom[ 9825]='h00000000;
    rd_cycle[ 9826] = 1'b0;  wr_cycle[ 9826] = 1'b0;  addr_rom[ 9826]='h00000000;  wr_data_rom[ 9826]='h00000000;
    rd_cycle[ 9827] = 1'b0;  wr_cycle[ 9827] = 1'b0;  addr_rom[ 9827]='h00000000;  wr_data_rom[ 9827]='h00000000;
    rd_cycle[ 9828] = 1'b0;  wr_cycle[ 9828] = 1'b0;  addr_rom[ 9828]='h00000000;  wr_data_rom[ 9828]='h00000000;
    rd_cycle[ 9829] = 1'b0;  wr_cycle[ 9829] = 1'b0;  addr_rom[ 9829]='h00000000;  wr_data_rom[ 9829]='h00000000;
    rd_cycle[ 9830] = 1'b0;  wr_cycle[ 9830] = 1'b0;  addr_rom[ 9830]='h00000000;  wr_data_rom[ 9830]='h00000000;
    rd_cycle[ 9831] = 1'b0;  wr_cycle[ 9831] = 1'b0;  addr_rom[ 9831]='h00000000;  wr_data_rom[ 9831]='h00000000;
    rd_cycle[ 9832] = 1'b0;  wr_cycle[ 9832] = 1'b0;  addr_rom[ 9832]='h00000000;  wr_data_rom[ 9832]='h00000000;
    rd_cycle[ 9833] = 1'b0;  wr_cycle[ 9833] = 1'b0;  addr_rom[ 9833]='h00000000;  wr_data_rom[ 9833]='h00000000;
    rd_cycle[ 9834] = 1'b0;  wr_cycle[ 9834] = 1'b0;  addr_rom[ 9834]='h00000000;  wr_data_rom[ 9834]='h00000000;
    rd_cycle[ 9835] = 1'b0;  wr_cycle[ 9835] = 1'b0;  addr_rom[ 9835]='h00000000;  wr_data_rom[ 9835]='h00000000;
    rd_cycle[ 9836] = 1'b0;  wr_cycle[ 9836] = 1'b0;  addr_rom[ 9836]='h00000000;  wr_data_rom[ 9836]='h00000000;
    rd_cycle[ 9837] = 1'b0;  wr_cycle[ 9837] = 1'b0;  addr_rom[ 9837]='h00000000;  wr_data_rom[ 9837]='h00000000;
    rd_cycle[ 9838] = 1'b0;  wr_cycle[ 9838] = 1'b0;  addr_rom[ 9838]='h00000000;  wr_data_rom[ 9838]='h00000000;
    rd_cycle[ 9839] = 1'b0;  wr_cycle[ 9839] = 1'b0;  addr_rom[ 9839]='h00000000;  wr_data_rom[ 9839]='h00000000;
    rd_cycle[ 9840] = 1'b0;  wr_cycle[ 9840] = 1'b0;  addr_rom[ 9840]='h00000000;  wr_data_rom[ 9840]='h00000000;
    rd_cycle[ 9841] = 1'b0;  wr_cycle[ 9841] = 1'b0;  addr_rom[ 9841]='h00000000;  wr_data_rom[ 9841]='h00000000;
    rd_cycle[ 9842] = 1'b0;  wr_cycle[ 9842] = 1'b0;  addr_rom[ 9842]='h00000000;  wr_data_rom[ 9842]='h00000000;
    rd_cycle[ 9843] = 1'b0;  wr_cycle[ 9843] = 1'b0;  addr_rom[ 9843]='h00000000;  wr_data_rom[ 9843]='h00000000;
    rd_cycle[ 9844] = 1'b0;  wr_cycle[ 9844] = 1'b0;  addr_rom[ 9844]='h00000000;  wr_data_rom[ 9844]='h00000000;
    rd_cycle[ 9845] = 1'b0;  wr_cycle[ 9845] = 1'b0;  addr_rom[ 9845]='h00000000;  wr_data_rom[ 9845]='h00000000;
    rd_cycle[ 9846] = 1'b0;  wr_cycle[ 9846] = 1'b0;  addr_rom[ 9846]='h00000000;  wr_data_rom[ 9846]='h00000000;
    rd_cycle[ 9847] = 1'b0;  wr_cycle[ 9847] = 1'b0;  addr_rom[ 9847]='h00000000;  wr_data_rom[ 9847]='h00000000;
    rd_cycle[ 9848] = 1'b0;  wr_cycle[ 9848] = 1'b0;  addr_rom[ 9848]='h00000000;  wr_data_rom[ 9848]='h00000000;
    rd_cycle[ 9849] = 1'b0;  wr_cycle[ 9849] = 1'b0;  addr_rom[ 9849]='h00000000;  wr_data_rom[ 9849]='h00000000;
    rd_cycle[ 9850] = 1'b0;  wr_cycle[ 9850] = 1'b0;  addr_rom[ 9850]='h00000000;  wr_data_rom[ 9850]='h00000000;
    rd_cycle[ 9851] = 1'b0;  wr_cycle[ 9851] = 1'b0;  addr_rom[ 9851]='h00000000;  wr_data_rom[ 9851]='h00000000;
    rd_cycle[ 9852] = 1'b0;  wr_cycle[ 9852] = 1'b0;  addr_rom[ 9852]='h00000000;  wr_data_rom[ 9852]='h00000000;
    rd_cycle[ 9853] = 1'b0;  wr_cycle[ 9853] = 1'b0;  addr_rom[ 9853]='h00000000;  wr_data_rom[ 9853]='h00000000;
    rd_cycle[ 9854] = 1'b0;  wr_cycle[ 9854] = 1'b0;  addr_rom[ 9854]='h00000000;  wr_data_rom[ 9854]='h00000000;
    rd_cycle[ 9855] = 1'b0;  wr_cycle[ 9855] = 1'b0;  addr_rom[ 9855]='h00000000;  wr_data_rom[ 9855]='h00000000;
    rd_cycle[ 9856] = 1'b0;  wr_cycle[ 9856] = 1'b0;  addr_rom[ 9856]='h00000000;  wr_data_rom[ 9856]='h00000000;
    rd_cycle[ 9857] = 1'b0;  wr_cycle[ 9857] = 1'b0;  addr_rom[ 9857]='h00000000;  wr_data_rom[ 9857]='h00000000;
    rd_cycle[ 9858] = 1'b0;  wr_cycle[ 9858] = 1'b0;  addr_rom[ 9858]='h00000000;  wr_data_rom[ 9858]='h00000000;
    rd_cycle[ 9859] = 1'b0;  wr_cycle[ 9859] = 1'b0;  addr_rom[ 9859]='h00000000;  wr_data_rom[ 9859]='h00000000;
    rd_cycle[ 9860] = 1'b0;  wr_cycle[ 9860] = 1'b0;  addr_rom[ 9860]='h00000000;  wr_data_rom[ 9860]='h00000000;
    rd_cycle[ 9861] = 1'b0;  wr_cycle[ 9861] = 1'b0;  addr_rom[ 9861]='h00000000;  wr_data_rom[ 9861]='h00000000;
    rd_cycle[ 9862] = 1'b0;  wr_cycle[ 9862] = 1'b0;  addr_rom[ 9862]='h00000000;  wr_data_rom[ 9862]='h00000000;
    rd_cycle[ 9863] = 1'b0;  wr_cycle[ 9863] = 1'b0;  addr_rom[ 9863]='h00000000;  wr_data_rom[ 9863]='h00000000;
    rd_cycle[ 9864] = 1'b0;  wr_cycle[ 9864] = 1'b0;  addr_rom[ 9864]='h00000000;  wr_data_rom[ 9864]='h00000000;
    rd_cycle[ 9865] = 1'b0;  wr_cycle[ 9865] = 1'b0;  addr_rom[ 9865]='h00000000;  wr_data_rom[ 9865]='h00000000;
    rd_cycle[ 9866] = 1'b0;  wr_cycle[ 9866] = 1'b0;  addr_rom[ 9866]='h00000000;  wr_data_rom[ 9866]='h00000000;
    rd_cycle[ 9867] = 1'b0;  wr_cycle[ 9867] = 1'b0;  addr_rom[ 9867]='h00000000;  wr_data_rom[ 9867]='h00000000;
    rd_cycle[ 9868] = 1'b0;  wr_cycle[ 9868] = 1'b0;  addr_rom[ 9868]='h00000000;  wr_data_rom[ 9868]='h00000000;
    rd_cycle[ 9869] = 1'b0;  wr_cycle[ 9869] = 1'b0;  addr_rom[ 9869]='h00000000;  wr_data_rom[ 9869]='h00000000;
    rd_cycle[ 9870] = 1'b0;  wr_cycle[ 9870] = 1'b0;  addr_rom[ 9870]='h00000000;  wr_data_rom[ 9870]='h00000000;
    rd_cycle[ 9871] = 1'b0;  wr_cycle[ 9871] = 1'b0;  addr_rom[ 9871]='h00000000;  wr_data_rom[ 9871]='h00000000;
    rd_cycle[ 9872] = 1'b0;  wr_cycle[ 9872] = 1'b0;  addr_rom[ 9872]='h00000000;  wr_data_rom[ 9872]='h00000000;
    rd_cycle[ 9873] = 1'b0;  wr_cycle[ 9873] = 1'b0;  addr_rom[ 9873]='h00000000;  wr_data_rom[ 9873]='h00000000;
    rd_cycle[ 9874] = 1'b0;  wr_cycle[ 9874] = 1'b0;  addr_rom[ 9874]='h00000000;  wr_data_rom[ 9874]='h00000000;
    rd_cycle[ 9875] = 1'b0;  wr_cycle[ 9875] = 1'b0;  addr_rom[ 9875]='h00000000;  wr_data_rom[ 9875]='h00000000;
    rd_cycle[ 9876] = 1'b0;  wr_cycle[ 9876] = 1'b0;  addr_rom[ 9876]='h00000000;  wr_data_rom[ 9876]='h00000000;
    rd_cycle[ 9877] = 1'b0;  wr_cycle[ 9877] = 1'b0;  addr_rom[ 9877]='h00000000;  wr_data_rom[ 9877]='h00000000;
    rd_cycle[ 9878] = 1'b0;  wr_cycle[ 9878] = 1'b0;  addr_rom[ 9878]='h00000000;  wr_data_rom[ 9878]='h00000000;
    rd_cycle[ 9879] = 1'b0;  wr_cycle[ 9879] = 1'b0;  addr_rom[ 9879]='h00000000;  wr_data_rom[ 9879]='h00000000;
    rd_cycle[ 9880] = 1'b0;  wr_cycle[ 9880] = 1'b0;  addr_rom[ 9880]='h00000000;  wr_data_rom[ 9880]='h00000000;
    rd_cycle[ 9881] = 1'b0;  wr_cycle[ 9881] = 1'b0;  addr_rom[ 9881]='h00000000;  wr_data_rom[ 9881]='h00000000;
    rd_cycle[ 9882] = 1'b0;  wr_cycle[ 9882] = 1'b0;  addr_rom[ 9882]='h00000000;  wr_data_rom[ 9882]='h00000000;
    rd_cycle[ 9883] = 1'b0;  wr_cycle[ 9883] = 1'b0;  addr_rom[ 9883]='h00000000;  wr_data_rom[ 9883]='h00000000;
    rd_cycle[ 9884] = 1'b0;  wr_cycle[ 9884] = 1'b0;  addr_rom[ 9884]='h00000000;  wr_data_rom[ 9884]='h00000000;
    rd_cycle[ 9885] = 1'b0;  wr_cycle[ 9885] = 1'b0;  addr_rom[ 9885]='h00000000;  wr_data_rom[ 9885]='h00000000;
    rd_cycle[ 9886] = 1'b0;  wr_cycle[ 9886] = 1'b0;  addr_rom[ 9886]='h00000000;  wr_data_rom[ 9886]='h00000000;
    rd_cycle[ 9887] = 1'b0;  wr_cycle[ 9887] = 1'b0;  addr_rom[ 9887]='h00000000;  wr_data_rom[ 9887]='h00000000;
    rd_cycle[ 9888] = 1'b0;  wr_cycle[ 9888] = 1'b0;  addr_rom[ 9888]='h00000000;  wr_data_rom[ 9888]='h00000000;
    rd_cycle[ 9889] = 1'b0;  wr_cycle[ 9889] = 1'b0;  addr_rom[ 9889]='h00000000;  wr_data_rom[ 9889]='h00000000;
    rd_cycle[ 9890] = 1'b0;  wr_cycle[ 9890] = 1'b0;  addr_rom[ 9890]='h00000000;  wr_data_rom[ 9890]='h00000000;
    rd_cycle[ 9891] = 1'b0;  wr_cycle[ 9891] = 1'b0;  addr_rom[ 9891]='h00000000;  wr_data_rom[ 9891]='h00000000;
    rd_cycle[ 9892] = 1'b0;  wr_cycle[ 9892] = 1'b0;  addr_rom[ 9892]='h00000000;  wr_data_rom[ 9892]='h00000000;
    rd_cycle[ 9893] = 1'b0;  wr_cycle[ 9893] = 1'b0;  addr_rom[ 9893]='h00000000;  wr_data_rom[ 9893]='h00000000;
    rd_cycle[ 9894] = 1'b0;  wr_cycle[ 9894] = 1'b0;  addr_rom[ 9894]='h00000000;  wr_data_rom[ 9894]='h00000000;
    rd_cycle[ 9895] = 1'b0;  wr_cycle[ 9895] = 1'b0;  addr_rom[ 9895]='h00000000;  wr_data_rom[ 9895]='h00000000;
    rd_cycle[ 9896] = 1'b0;  wr_cycle[ 9896] = 1'b0;  addr_rom[ 9896]='h00000000;  wr_data_rom[ 9896]='h00000000;
    rd_cycle[ 9897] = 1'b0;  wr_cycle[ 9897] = 1'b0;  addr_rom[ 9897]='h00000000;  wr_data_rom[ 9897]='h00000000;
    rd_cycle[ 9898] = 1'b0;  wr_cycle[ 9898] = 1'b0;  addr_rom[ 9898]='h00000000;  wr_data_rom[ 9898]='h00000000;
    rd_cycle[ 9899] = 1'b0;  wr_cycle[ 9899] = 1'b0;  addr_rom[ 9899]='h00000000;  wr_data_rom[ 9899]='h00000000;
    rd_cycle[ 9900] = 1'b0;  wr_cycle[ 9900] = 1'b0;  addr_rom[ 9900]='h00000000;  wr_data_rom[ 9900]='h00000000;
    rd_cycle[ 9901] = 1'b0;  wr_cycle[ 9901] = 1'b0;  addr_rom[ 9901]='h00000000;  wr_data_rom[ 9901]='h00000000;
    rd_cycle[ 9902] = 1'b0;  wr_cycle[ 9902] = 1'b0;  addr_rom[ 9902]='h00000000;  wr_data_rom[ 9902]='h00000000;
    rd_cycle[ 9903] = 1'b0;  wr_cycle[ 9903] = 1'b0;  addr_rom[ 9903]='h00000000;  wr_data_rom[ 9903]='h00000000;
    rd_cycle[ 9904] = 1'b0;  wr_cycle[ 9904] = 1'b0;  addr_rom[ 9904]='h00000000;  wr_data_rom[ 9904]='h00000000;
    rd_cycle[ 9905] = 1'b0;  wr_cycle[ 9905] = 1'b0;  addr_rom[ 9905]='h00000000;  wr_data_rom[ 9905]='h00000000;
    rd_cycle[ 9906] = 1'b0;  wr_cycle[ 9906] = 1'b0;  addr_rom[ 9906]='h00000000;  wr_data_rom[ 9906]='h00000000;
    rd_cycle[ 9907] = 1'b0;  wr_cycle[ 9907] = 1'b0;  addr_rom[ 9907]='h00000000;  wr_data_rom[ 9907]='h00000000;
    rd_cycle[ 9908] = 1'b0;  wr_cycle[ 9908] = 1'b0;  addr_rom[ 9908]='h00000000;  wr_data_rom[ 9908]='h00000000;
    rd_cycle[ 9909] = 1'b0;  wr_cycle[ 9909] = 1'b0;  addr_rom[ 9909]='h00000000;  wr_data_rom[ 9909]='h00000000;
    rd_cycle[ 9910] = 1'b0;  wr_cycle[ 9910] = 1'b0;  addr_rom[ 9910]='h00000000;  wr_data_rom[ 9910]='h00000000;
    rd_cycle[ 9911] = 1'b0;  wr_cycle[ 9911] = 1'b0;  addr_rom[ 9911]='h00000000;  wr_data_rom[ 9911]='h00000000;
    rd_cycle[ 9912] = 1'b0;  wr_cycle[ 9912] = 1'b0;  addr_rom[ 9912]='h00000000;  wr_data_rom[ 9912]='h00000000;
    rd_cycle[ 9913] = 1'b0;  wr_cycle[ 9913] = 1'b0;  addr_rom[ 9913]='h00000000;  wr_data_rom[ 9913]='h00000000;
    rd_cycle[ 9914] = 1'b0;  wr_cycle[ 9914] = 1'b0;  addr_rom[ 9914]='h00000000;  wr_data_rom[ 9914]='h00000000;
    rd_cycle[ 9915] = 1'b0;  wr_cycle[ 9915] = 1'b0;  addr_rom[ 9915]='h00000000;  wr_data_rom[ 9915]='h00000000;
    rd_cycle[ 9916] = 1'b0;  wr_cycle[ 9916] = 1'b0;  addr_rom[ 9916]='h00000000;  wr_data_rom[ 9916]='h00000000;
    rd_cycle[ 9917] = 1'b0;  wr_cycle[ 9917] = 1'b0;  addr_rom[ 9917]='h00000000;  wr_data_rom[ 9917]='h00000000;
    rd_cycle[ 9918] = 1'b0;  wr_cycle[ 9918] = 1'b0;  addr_rom[ 9918]='h00000000;  wr_data_rom[ 9918]='h00000000;
    rd_cycle[ 9919] = 1'b0;  wr_cycle[ 9919] = 1'b0;  addr_rom[ 9919]='h00000000;  wr_data_rom[ 9919]='h00000000;
    rd_cycle[ 9920] = 1'b0;  wr_cycle[ 9920] = 1'b0;  addr_rom[ 9920]='h00000000;  wr_data_rom[ 9920]='h00000000;
    rd_cycle[ 9921] = 1'b0;  wr_cycle[ 9921] = 1'b0;  addr_rom[ 9921]='h00000000;  wr_data_rom[ 9921]='h00000000;
    rd_cycle[ 9922] = 1'b0;  wr_cycle[ 9922] = 1'b0;  addr_rom[ 9922]='h00000000;  wr_data_rom[ 9922]='h00000000;
    rd_cycle[ 9923] = 1'b0;  wr_cycle[ 9923] = 1'b0;  addr_rom[ 9923]='h00000000;  wr_data_rom[ 9923]='h00000000;
    rd_cycle[ 9924] = 1'b0;  wr_cycle[ 9924] = 1'b0;  addr_rom[ 9924]='h00000000;  wr_data_rom[ 9924]='h00000000;
    rd_cycle[ 9925] = 1'b0;  wr_cycle[ 9925] = 1'b0;  addr_rom[ 9925]='h00000000;  wr_data_rom[ 9925]='h00000000;
    rd_cycle[ 9926] = 1'b0;  wr_cycle[ 9926] = 1'b0;  addr_rom[ 9926]='h00000000;  wr_data_rom[ 9926]='h00000000;
    rd_cycle[ 9927] = 1'b0;  wr_cycle[ 9927] = 1'b0;  addr_rom[ 9927]='h00000000;  wr_data_rom[ 9927]='h00000000;
    rd_cycle[ 9928] = 1'b0;  wr_cycle[ 9928] = 1'b0;  addr_rom[ 9928]='h00000000;  wr_data_rom[ 9928]='h00000000;
    rd_cycle[ 9929] = 1'b0;  wr_cycle[ 9929] = 1'b0;  addr_rom[ 9929]='h00000000;  wr_data_rom[ 9929]='h00000000;
    rd_cycle[ 9930] = 1'b0;  wr_cycle[ 9930] = 1'b0;  addr_rom[ 9930]='h00000000;  wr_data_rom[ 9930]='h00000000;
    rd_cycle[ 9931] = 1'b0;  wr_cycle[ 9931] = 1'b0;  addr_rom[ 9931]='h00000000;  wr_data_rom[ 9931]='h00000000;
    rd_cycle[ 9932] = 1'b0;  wr_cycle[ 9932] = 1'b0;  addr_rom[ 9932]='h00000000;  wr_data_rom[ 9932]='h00000000;
    rd_cycle[ 9933] = 1'b0;  wr_cycle[ 9933] = 1'b0;  addr_rom[ 9933]='h00000000;  wr_data_rom[ 9933]='h00000000;
    rd_cycle[ 9934] = 1'b0;  wr_cycle[ 9934] = 1'b0;  addr_rom[ 9934]='h00000000;  wr_data_rom[ 9934]='h00000000;
    rd_cycle[ 9935] = 1'b0;  wr_cycle[ 9935] = 1'b0;  addr_rom[ 9935]='h00000000;  wr_data_rom[ 9935]='h00000000;
    rd_cycle[ 9936] = 1'b0;  wr_cycle[ 9936] = 1'b0;  addr_rom[ 9936]='h00000000;  wr_data_rom[ 9936]='h00000000;
    rd_cycle[ 9937] = 1'b0;  wr_cycle[ 9937] = 1'b0;  addr_rom[ 9937]='h00000000;  wr_data_rom[ 9937]='h00000000;
    rd_cycle[ 9938] = 1'b0;  wr_cycle[ 9938] = 1'b0;  addr_rom[ 9938]='h00000000;  wr_data_rom[ 9938]='h00000000;
    rd_cycle[ 9939] = 1'b0;  wr_cycle[ 9939] = 1'b0;  addr_rom[ 9939]='h00000000;  wr_data_rom[ 9939]='h00000000;
    rd_cycle[ 9940] = 1'b0;  wr_cycle[ 9940] = 1'b0;  addr_rom[ 9940]='h00000000;  wr_data_rom[ 9940]='h00000000;
    rd_cycle[ 9941] = 1'b0;  wr_cycle[ 9941] = 1'b0;  addr_rom[ 9941]='h00000000;  wr_data_rom[ 9941]='h00000000;
    rd_cycle[ 9942] = 1'b0;  wr_cycle[ 9942] = 1'b0;  addr_rom[ 9942]='h00000000;  wr_data_rom[ 9942]='h00000000;
    rd_cycle[ 9943] = 1'b0;  wr_cycle[ 9943] = 1'b0;  addr_rom[ 9943]='h00000000;  wr_data_rom[ 9943]='h00000000;
    rd_cycle[ 9944] = 1'b0;  wr_cycle[ 9944] = 1'b0;  addr_rom[ 9944]='h00000000;  wr_data_rom[ 9944]='h00000000;
    rd_cycle[ 9945] = 1'b0;  wr_cycle[ 9945] = 1'b0;  addr_rom[ 9945]='h00000000;  wr_data_rom[ 9945]='h00000000;
    rd_cycle[ 9946] = 1'b0;  wr_cycle[ 9946] = 1'b0;  addr_rom[ 9946]='h00000000;  wr_data_rom[ 9946]='h00000000;
    rd_cycle[ 9947] = 1'b0;  wr_cycle[ 9947] = 1'b0;  addr_rom[ 9947]='h00000000;  wr_data_rom[ 9947]='h00000000;
    rd_cycle[ 9948] = 1'b0;  wr_cycle[ 9948] = 1'b0;  addr_rom[ 9948]='h00000000;  wr_data_rom[ 9948]='h00000000;
    rd_cycle[ 9949] = 1'b0;  wr_cycle[ 9949] = 1'b0;  addr_rom[ 9949]='h00000000;  wr_data_rom[ 9949]='h00000000;
    rd_cycle[ 9950] = 1'b0;  wr_cycle[ 9950] = 1'b0;  addr_rom[ 9950]='h00000000;  wr_data_rom[ 9950]='h00000000;
    rd_cycle[ 9951] = 1'b0;  wr_cycle[ 9951] = 1'b0;  addr_rom[ 9951]='h00000000;  wr_data_rom[ 9951]='h00000000;
    rd_cycle[ 9952] = 1'b0;  wr_cycle[ 9952] = 1'b0;  addr_rom[ 9952]='h00000000;  wr_data_rom[ 9952]='h00000000;
    rd_cycle[ 9953] = 1'b0;  wr_cycle[ 9953] = 1'b0;  addr_rom[ 9953]='h00000000;  wr_data_rom[ 9953]='h00000000;
    rd_cycle[ 9954] = 1'b0;  wr_cycle[ 9954] = 1'b0;  addr_rom[ 9954]='h00000000;  wr_data_rom[ 9954]='h00000000;
    rd_cycle[ 9955] = 1'b0;  wr_cycle[ 9955] = 1'b0;  addr_rom[ 9955]='h00000000;  wr_data_rom[ 9955]='h00000000;
    rd_cycle[ 9956] = 1'b0;  wr_cycle[ 9956] = 1'b0;  addr_rom[ 9956]='h00000000;  wr_data_rom[ 9956]='h00000000;
    rd_cycle[ 9957] = 1'b0;  wr_cycle[ 9957] = 1'b0;  addr_rom[ 9957]='h00000000;  wr_data_rom[ 9957]='h00000000;
    rd_cycle[ 9958] = 1'b0;  wr_cycle[ 9958] = 1'b0;  addr_rom[ 9958]='h00000000;  wr_data_rom[ 9958]='h00000000;
    rd_cycle[ 9959] = 1'b0;  wr_cycle[ 9959] = 1'b0;  addr_rom[ 9959]='h00000000;  wr_data_rom[ 9959]='h00000000;
    rd_cycle[ 9960] = 1'b0;  wr_cycle[ 9960] = 1'b0;  addr_rom[ 9960]='h00000000;  wr_data_rom[ 9960]='h00000000;
    rd_cycle[ 9961] = 1'b0;  wr_cycle[ 9961] = 1'b0;  addr_rom[ 9961]='h00000000;  wr_data_rom[ 9961]='h00000000;
    rd_cycle[ 9962] = 1'b0;  wr_cycle[ 9962] = 1'b0;  addr_rom[ 9962]='h00000000;  wr_data_rom[ 9962]='h00000000;
    rd_cycle[ 9963] = 1'b0;  wr_cycle[ 9963] = 1'b0;  addr_rom[ 9963]='h00000000;  wr_data_rom[ 9963]='h00000000;
    rd_cycle[ 9964] = 1'b0;  wr_cycle[ 9964] = 1'b0;  addr_rom[ 9964]='h00000000;  wr_data_rom[ 9964]='h00000000;
    rd_cycle[ 9965] = 1'b0;  wr_cycle[ 9965] = 1'b0;  addr_rom[ 9965]='h00000000;  wr_data_rom[ 9965]='h00000000;
    rd_cycle[ 9966] = 1'b0;  wr_cycle[ 9966] = 1'b0;  addr_rom[ 9966]='h00000000;  wr_data_rom[ 9966]='h00000000;
    rd_cycle[ 9967] = 1'b0;  wr_cycle[ 9967] = 1'b0;  addr_rom[ 9967]='h00000000;  wr_data_rom[ 9967]='h00000000;
    rd_cycle[ 9968] = 1'b0;  wr_cycle[ 9968] = 1'b0;  addr_rom[ 9968]='h00000000;  wr_data_rom[ 9968]='h00000000;
    rd_cycle[ 9969] = 1'b0;  wr_cycle[ 9969] = 1'b0;  addr_rom[ 9969]='h00000000;  wr_data_rom[ 9969]='h00000000;
    rd_cycle[ 9970] = 1'b0;  wr_cycle[ 9970] = 1'b0;  addr_rom[ 9970]='h00000000;  wr_data_rom[ 9970]='h00000000;
    rd_cycle[ 9971] = 1'b0;  wr_cycle[ 9971] = 1'b0;  addr_rom[ 9971]='h00000000;  wr_data_rom[ 9971]='h00000000;
    rd_cycle[ 9972] = 1'b0;  wr_cycle[ 9972] = 1'b0;  addr_rom[ 9972]='h00000000;  wr_data_rom[ 9972]='h00000000;
    rd_cycle[ 9973] = 1'b0;  wr_cycle[ 9973] = 1'b0;  addr_rom[ 9973]='h00000000;  wr_data_rom[ 9973]='h00000000;
    rd_cycle[ 9974] = 1'b0;  wr_cycle[ 9974] = 1'b0;  addr_rom[ 9974]='h00000000;  wr_data_rom[ 9974]='h00000000;
    rd_cycle[ 9975] = 1'b0;  wr_cycle[ 9975] = 1'b0;  addr_rom[ 9975]='h00000000;  wr_data_rom[ 9975]='h00000000;
    rd_cycle[ 9976] = 1'b0;  wr_cycle[ 9976] = 1'b0;  addr_rom[ 9976]='h00000000;  wr_data_rom[ 9976]='h00000000;
    rd_cycle[ 9977] = 1'b0;  wr_cycle[ 9977] = 1'b0;  addr_rom[ 9977]='h00000000;  wr_data_rom[ 9977]='h00000000;
    rd_cycle[ 9978] = 1'b0;  wr_cycle[ 9978] = 1'b0;  addr_rom[ 9978]='h00000000;  wr_data_rom[ 9978]='h00000000;
    rd_cycle[ 9979] = 1'b0;  wr_cycle[ 9979] = 1'b0;  addr_rom[ 9979]='h00000000;  wr_data_rom[ 9979]='h00000000;
    rd_cycle[ 9980] = 1'b0;  wr_cycle[ 9980] = 1'b0;  addr_rom[ 9980]='h00000000;  wr_data_rom[ 9980]='h00000000;
    rd_cycle[ 9981] = 1'b0;  wr_cycle[ 9981] = 1'b0;  addr_rom[ 9981]='h00000000;  wr_data_rom[ 9981]='h00000000;
    rd_cycle[ 9982] = 1'b0;  wr_cycle[ 9982] = 1'b0;  addr_rom[ 9982]='h00000000;  wr_data_rom[ 9982]='h00000000;
    rd_cycle[ 9983] = 1'b0;  wr_cycle[ 9983] = 1'b0;  addr_rom[ 9983]='h00000000;  wr_data_rom[ 9983]='h00000000;
    rd_cycle[ 9984] = 1'b0;  wr_cycle[ 9984] = 1'b0;  addr_rom[ 9984]='h00000000;  wr_data_rom[ 9984]='h00000000;
    rd_cycle[ 9985] = 1'b0;  wr_cycle[ 9985] = 1'b0;  addr_rom[ 9985]='h00000000;  wr_data_rom[ 9985]='h00000000;
    rd_cycle[ 9986] = 1'b0;  wr_cycle[ 9986] = 1'b0;  addr_rom[ 9986]='h00000000;  wr_data_rom[ 9986]='h00000000;
    rd_cycle[ 9987] = 1'b0;  wr_cycle[ 9987] = 1'b0;  addr_rom[ 9987]='h00000000;  wr_data_rom[ 9987]='h00000000;
    rd_cycle[ 9988] = 1'b0;  wr_cycle[ 9988] = 1'b0;  addr_rom[ 9988]='h00000000;  wr_data_rom[ 9988]='h00000000;
    rd_cycle[ 9989] = 1'b0;  wr_cycle[ 9989] = 1'b0;  addr_rom[ 9989]='h00000000;  wr_data_rom[ 9989]='h00000000;
    rd_cycle[ 9990] = 1'b0;  wr_cycle[ 9990] = 1'b0;  addr_rom[ 9990]='h00000000;  wr_data_rom[ 9990]='h00000000;
    rd_cycle[ 9991] = 1'b0;  wr_cycle[ 9991] = 1'b0;  addr_rom[ 9991]='h00000000;  wr_data_rom[ 9991]='h00000000;
    rd_cycle[ 9992] = 1'b0;  wr_cycle[ 9992] = 1'b0;  addr_rom[ 9992]='h00000000;  wr_data_rom[ 9992]='h00000000;
    rd_cycle[ 9993] = 1'b0;  wr_cycle[ 9993] = 1'b0;  addr_rom[ 9993]='h00000000;  wr_data_rom[ 9993]='h00000000;
    rd_cycle[ 9994] = 1'b0;  wr_cycle[ 9994] = 1'b0;  addr_rom[ 9994]='h00000000;  wr_data_rom[ 9994]='h00000000;
    rd_cycle[ 9995] = 1'b0;  wr_cycle[ 9995] = 1'b0;  addr_rom[ 9995]='h00000000;  wr_data_rom[ 9995]='h00000000;
    rd_cycle[ 9996] = 1'b0;  wr_cycle[ 9996] = 1'b0;  addr_rom[ 9996]='h00000000;  wr_data_rom[ 9996]='h00000000;
    rd_cycle[ 9997] = 1'b0;  wr_cycle[ 9997] = 1'b0;  addr_rom[ 9997]='h00000000;  wr_data_rom[ 9997]='h00000000;
    rd_cycle[ 9998] = 1'b0;  wr_cycle[ 9998] = 1'b0;  addr_rom[ 9998]='h00000000;  wr_data_rom[ 9998]='h00000000;
    rd_cycle[ 9999] = 1'b0;  wr_cycle[ 9999] = 1'b0;  addr_rom[ 9999]='h00000000;  wr_data_rom[ 9999]='h00000000;
    // 2000 sequence read cycles
    rd_cycle[10000] = 1'b1;  wr_cycle[10000] = 1'b0;  addr_rom[10000]='h00000000;  wr_data_rom[10000]='h00000000;
    rd_cycle[10001] = 1'b1;  wr_cycle[10001] = 1'b0;  addr_rom[10001]='h00000004;  wr_data_rom[10001]='h00000000;
    rd_cycle[10002] = 1'b1;  wr_cycle[10002] = 1'b0;  addr_rom[10002]='h00000008;  wr_data_rom[10002]='h00000000;
    rd_cycle[10003] = 1'b1;  wr_cycle[10003] = 1'b0;  addr_rom[10003]='h0000000c;  wr_data_rom[10003]='h00000000;
    rd_cycle[10004] = 1'b1;  wr_cycle[10004] = 1'b0;  addr_rom[10004]='h00000010;  wr_data_rom[10004]='h00000000;
    rd_cycle[10005] = 1'b1;  wr_cycle[10005] = 1'b0;  addr_rom[10005]='h00000014;  wr_data_rom[10005]='h00000000;
    rd_cycle[10006] = 1'b1;  wr_cycle[10006] = 1'b0;  addr_rom[10006]='h00000018;  wr_data_rom[10006]='h00000000;
    rd_cycle[10007] = 1'b1;  wr_cycle[10007] = 1'b0;  addr_rom[10007]='h0000001c;  wr_data_rom[10007]='h00000000;
    rd_cycle[10008] = 1'b1;  wr_cycle[10008] = 1'b0;  addr_rom[10008]='h00000020;  wr_data_rom[10008]='h00000000;
    rd_cycle[10009] = 1'b1;  wr_cycle[10009] = 1'b0;  addr_rom[10009]='h00000024;  wr_data_rom[10009]='h00000000;
    rd_cycle[10010] = 1'b1;  wr_cycle[10010] = 1'b0;  addr_rom[10010]='h00000028;  wr_data_rom[10010]='h00000000;
    rd_cycle[10011] = 1'b1;  wr_cycle[10011] = 1'b0;  addr_rom[10011]='h0000002c;  wr_data_rom[10011]='h00000000;
    rd_cycle[10012] = 1'b1;  wr_cycle[10012] = 1'b0;  addr_rom[10012]='h00000030;  wr_data_rom[10012]='h00000000;
    rd_cycle[10013] = 1'b1;  wr_cycle[10013] = 1'b0;  addr_rom[10013]='h00000034;  wr_data_rom[10013]='h00000000;
    rd_cycle[10014] = 1'b1;  wr_cycle[10014] = 1'b0;  addr_rom[10014]='h00000038;  wr_data_rom[10014]='h00000000;
    rd_cycle[10015] = 1'b1;  wr_cycle[10015] = 1'b0;  addr_rom[10015]='h0000003c;  wr_data_rom[10015]='h00000000;
    rd_cycle[10016] = 1'b1;  wr_cycle[10016] = 1'b0;  addr_rom[10016]='h00000040;  wr_data_rom[10016]='h00000000;
    rd_cycle[10017] = 1'b1;  wr_cycle[10017] = 1'b0;  addr_rom[10017]='h00000044;  wr_data_rom[10017]='h00000000;
    rd_cycle[10018] = 1'b1;  wr_cycle[10018] = 1'b0;  addr_rom[10018]='h00000048;  wr_data_rom[10018]='h00000000;
    rd_cycle[10019] = 1'b1;  wr_cycle[10019] = 1'b0;  addr_rom[10019]='h0000004c;  wr_data_rom[10019]='h00000000;
    rd_cycle[10020] = 1'b1;  wr_cycle[10020] = 1'b0;  addr_rom[10020]='h00000050;  wr_data_rom[10020]='h00000000;
    rd_cycle[10021] = 1'b1;  wr_cycle[10021] = 1'b0;  addr_rom[10021]='h00000054;  wr_data_rom[10021]='h00000000;
    rd_cycle[10022] = 1'b1;  wr_cycle[10022] = 1'b0;  addr_rom[10022]='h00000058;  wr_data_rom[10022]='h00000000;
    rd_cycle[10023] = 1'b1;  wr_cycle[10023] = 1'b0;  addr_rom[10023]='h0000005c;  wr_data_rom[10023]='h00000000;
    rd_cycle[10024] = 1'b1;  wr_cycle[10024] = 1'b0;  addr_rom[10024]='h00000060;  wr_data_rom[10024]='h00000000;
    rd_cycle[10025] = 1'b1;  wr_cycle[10025] = 1'b0;  addr_rom[10025]='h00000064;  wr_data_rom[10025]='h00000000;
    rd_cycle[10026] = 1'b1;  wr_cycle[10026] = 1'b0;  addr_rom[10026]='h00000068;  wr_data_rom[10026]='h00000000;
    rd_cycle[10027] = 1'b1;  wr_cycle[10027] = 1'b0;  addr_rom[10027]='h0000006c;  wr_data_rom[10027]='h00000000;
    rd_cycle[10028] = 1'b1;  wr_cycle[10028] = 1'b0;  addr_rom[10028]='h00000070;  wr_data_rom[10028]='h00000000;
    rd_cycle[10029] = 1'b1;  wr_cycle[10029] = 1'b0;  addr_rom[10029]='h00000074;  wr_data_rom[10029]='h00000000;
    rd_cycle[10030] = 1'b1;  wr_cycle[10030] = 1'b0;  addr_rom[10030]='h00000078;  wr_data_rom[10030]='h00000000;
    rd_cycle[10031] = 1'b1;  wr_cycle[10031] = 1'b0;  addr_rom[10031]='h0000007c;  wr_data_rom[10031]='h00000000;
    rd_cycle[10032] = 1'b1;  wr_cycle[10032] = 1'b0;  addr_rom[10032]='h00000080;  wr_data_rom[10032]='h00000000;
    rd_cycle[10033] = 1'b1;  wr_cycle[10033] = 1'b0;  addr_rom[10033]='h00000084;  wr_data_rom[10033]='h00000000;
    rd_cycle[10034] = 1'b1;  wr_cycle[10034] = 1'b0;  addr_rom[10034]='h00000088;  wr_data_rom[10034]='h00000000;
    rd_cycle[10035] = 1'b1;  wr_cycle[10035] = 1'b0;  addr_rom[10035]='h0000008c;  wr_data_rom[10035]='h00000000;
    rd_cycle[10036] = 1'b1;  wr_cycle[10036] = 1'b0;  addr_rom[10036]='h00000090;  wr_data_rom[10036]='h00000000;
    rd_cycle[10037] = 1'b1;  wr_cycle[10037] = 1'b0;  addr_rom[10037]='h00000094;  wr_data_rom[10037]='h00000000;
    rd_cycle[10038] = 1'b1;  wr_cycle[10038] = 1'b0;  addr_rom[10038]='h00000098;  wr_data_rom[10038]='h00000000;
    rd_cycle[10039] = 1'b1;  wr_cycle[10039] = 1'b0;  addr_rom[10039]='h0000009c;  wr_data_rom[10039]='h00000000;
    rd_cycle[10040] = 1'b1;  wr_cycle[10040] = 1'b0;  addr_rom[10040]='h000000a0;  wr_data_rom[10040]='h00000000;
    rd_cycle[10041] = 1'b1;  wr_cycle[10041] = 1'b0;  addr_rom[10041]='h000000a4;  wr_data_rom[10041]='h00000000;
    rd_cycle[10042] = 1'b1;  wr_cycle[10042] = 1'b0;  addr_rom[10042]='h000000a8;  wr_data_rom[10042]='h00000000;
    rd_cycle[10043] = 1'b1;  wr_cycle[10043] = 1'b0;  addr_rom[10043]='h000000ac;  wr_data_rom[10043]='h00000000;
    rd_cycle[10044] = 1'b1;  wr_cycle[10044] = 1'b0;  addr_rom[10044]='h000000b0;  wr_data_rom[10044]='h00000000;
    rd_cycle[10045] = 1'b1;  wr_cycle[10045] = 1'b0;  addr_rom[10045]='h000000b4;  wr_data_rom[10045]='h00000000;
    rd_cycle[10046] = 1'b1;  wr_cycle[10046] = 1'b0;  addr_rom[10046]='h000000b8;  wr_data_rom[10046]='h00000000;
    rd_cycle[10047] = 1'b1;  wr_cycle[10047] = 1'b0;  addr_rom[10047]='h000000bc;  wr_data_rom[10047]='h00000000;
    rd_cycle[10048] = 1'b1;  wr_cycle[10048] = 1'b0;  addr_rom[10048]='h000000c0;  wr_data_rom[10048]='h00000000;
    rd_cycle[10049] = 1'b1;  wr_cycle[10049] = 1'b0;  addr_rom[10049]='h000000c4;  wr_data_rom[10049]='h00000000;
    rd_cycle[10050] = 1'b1;  wr_cycle[10050] = 1'b0;  addr_rom[10050]='h000000c8;  wr_data_rom[10050]='h00000000;
    rd_cycle[10051] = 1'b1;  wr_cycle[10051] = 1'b0;  addr_rom[10051]='h000000cc;  wr_data_rom[10051]='h00000000;
    rd_cycle[10052] = 1'b1;  wr_cycle[10052] = 1'b0;  addr_rom[10052]='h000000d0;  wr_data_rom[10052]='h00000000;
    rd_cycle[10053] = 1'b1;  wr_cycle[10053] = 1'b0;  addr_rom[10053]='h000000d4;  wr_data_rom[10053]='h00000000;
    rd_cycle[10054] = 1'b1;  wr_cycle[10054] = 1'b0;  addr_rom[10054]='h000000d8;  wr_data_rom[10054]='h00000000;
    rd_cycle[10055] = 1'b1;  wr_cycle[10055] = 1'b0;  addr_rom[10055]='h000000dc;  wr_data_rom[10055]='h00000000;
    rd_cycle[10056] = 1'b1;  wr_cycle[10056] = 1'b0;  addr_rom[10056]='h000000e0;  wr_data_rom[10056]='h00000000;
    rd_cycle[10057] = 1'b1;  wr_cycle[10057] = 1'b0;  addr_rom[10057]='h000000e4;  wr_data_rom[10057]='h00000000;
    rd_cycle[10058] = 1'b1;  wr_cycle[10058] = 1'b0;  addr_rom[10058]='h000000e8;  wr_data_rom[10058]='h00000000;
    rd_cycle[10059] = 1'b1;  wr_cycle[10059] = 1'b0;  addr_rom[10059]='h000000ec;  wr_data_rom[10059]='h00000000;
    rd_cycle[10060] = 1'b1;  wr_cycle[10060] = 1'b0;  addr_rom[10060]='h000000f0;  wr_data_rom[10060]='h00000000;
    rd_cycle[10061] = 1'b1;  wr_cycle[10061] = 1'b0;  addr_rom[10061]='h000000f4;  wr_data_rom[10061]='h00000000;
    rd_cycle[10062] = 1'b1;  wr_cycle[10062] = 1'b0;  addr_rom[10062]='h000000f8;  wr_data_rom[10062]='h00000000;
    rd_cycle[10063] = 1'b1;  wr_cycle[10063] = 1'b0;  addr_rom[10063]='h000000fc;  wr_data_rom[10063]='h00000000;
    rd_cycle[10064] = 1'b1;  wr_cycle[10064] = 1'b0;  addr_rom[10064]='h00000100;  wr_data_rom[10064]='h00000000;
    rd_cycle[10065] = 1'b1;  wr_cycle[10065] = 1'b0;  addr_rom[10065]='h00000104;  wr_data_rom[10065]='h00000000;
    rd_cycle[10066] = 1'b1;  wr_cycle[10066] = 1'b0;  addr_rom[10066]='h00000108;  wr_data_rom[10066]='h00000000;
    rd_cycle[10067] = 1'b1;  wr_cycle[10067] = 1'b0;  addr_rom[10067]='h0000010c;  wr_data_rom[10067]='h00000000;
    rd_cycle[10068] = 1'b1;  wr_cycle[10068] = 1'b0;  addr_rom[10068]='h00000110;  wr_data_rom[10068]='h00000000;
    rd_cycle[10069] = 1'b1;  wr_cycle[10069] = 1'b0;  addr_rom[10069]='h00000114;  wr_data_rom[10069]='h00000000;
    rd_cycle[10070] = 1'b1;  wr_cycle[10070] = 1'b0;  addr_rom[10070]='h00000118;  wr_data_rom[10070]='h00000000;
    rd_cycle[10071] = 1'b1;  wr_cycle[10071] = 1'b0;  addr_rom[10071]='h0000011c;  wr_data_rom[10071]='h00000000;
    rd_cycle[10072] = 1'b1;  wr_cycle[10072] = 1'b0;  addr_rom[10072]='h00000120;  wr_data_rom[10072]='h00000000;
    rd_cycle[10073] = 1'b1;  wr_cycle[10073] = 1'b0;  addr_rom[10073]='h00000124;  wr_data_rom[10073]='h00000000;
    rd_cycle[10074] = 1'b1;  wr_cycle[10074] = 1'b0;  addr_rom[10074]='h00000128;  wr_data_rom[10074]='h00000000;
    rd_cycle[10075] = 1'b1;  wr_cycle[10075] = 1'b0;  addr_rom[10075]='h0000012c;  wr_data_rom[10075]='h00000000;
    rd_cycle[10076] = 1'b1;  wr_cycle[10076] = 1'b0;  addr_rom[10076]='h00000130;  wr_data_rom[10076]='h00000000;
    rd_cycle[10077] = 1'b1;  wr_cycle[10077] = 1'b0;  addr_rom[10077]='h00000134;  wr_data_rom[10077]='h00000000;
    rd_cycle[10078] = 1'b1;  wr_cycle[10078] = 1'b0;  addr_rom[10078]='h00000138;  wr_data_rom[10078]='h00000000;
    rd_cycle[10079] = 1'b1;  wr_cycle[10079] = 1'b0;  addr_rom[10079]='h0000013c;  wr_data_rom[10079]='h00000000;
    rd_cycle[10080] = 1'b1;  wr_cycle[10080] = 1'b0;  addr_rom[10080]='h00000140;  wr_data_rom[10080]='h00000000;
    rd_cycle[10081] = 1'b1;  wr_cycle[10081] = 1'b0;  addr_rom[10081]='h00000144;  wr_data_rom[10081]='h00000000;
    rd_cycle[10082] = 1'b1;  wr_cycle[10082] = 1'b0;  addr_rom[10082]='h00000148;  wr_data_rom[10082]='h00000000;
    rd_cycle[10083] = 1'b1;  wr_cycle[10083] = 1'b0;  addr_rom[10083]='h0000014c;  wr_data_rom[10083]='h00000000;
    rd_cycle[10084] = 1'b1;  wr_cycle[10084] = 1'b0;  addr_rom[10084]='h00000150;  wr_data_rom[10084]='h00000000;
    rd_cycle[10085] = 1'b1;  wr_cycle[10085] = 1'b0;  addr_rom[10085]='h00000154;  wr_data_rom[10085]='h00000000;
    rd_cycle[10086] = 1'b1;  wr_cycle[10086] = 1'b0;  addr_rom[10086]='h00000158;  wr_data_rom[10086]='h00000000;
    rd_cycle[10087] = 1'b1;  wr_cycle[10087] = 1'b0;  addr_rom[10087]='h0000015c;  wr_data_rom[10087]='h00000000;
    rd_cycle[10088] = 1'b1;  wr_cycle[10088] = 1'b0;  addr_rom[10088]='h00000160;  wr_data_rom[10088]='h00000000;
    rd_cycle[10089] = 1'b1;  wr_cycle[10089] = 1'b0;  addr_rom[10089]='h00000164;  wr_data_rom[10089]='h00000000;
    rd_cycle[10090] = 1'b1;  wr_cycle[10090] = 1'b0;  addr_rom[10090]='h00000168;  wr_data_rom[10090]='h00000000;
    rd_cycle[10091] = 1'b1;  wr_cycle[10091] = 1'b0;  addr_rom[10091]='h0000016c;  wr_data_rom[10091]='h00000000;
    rd_cycle[10092] = 1'b1;  wr_cycle[10092] = 1'b0;  addr_rom[10092]='h00000170;  wr_data_rom[10092]='h00000000;
    rd_cycle[10093] = 1'b1;  wr_cycle[10093] = 1'b0;  addr_rom[10093]='h00000174;  wr_data_rom[10093]='h00000000;
    rd_cycle[10094] = 1'b1;  wr_cycle[10094] = 1'b0;  addr_rom[10094]='h00000178;  wr_data_rom[10094]='h00000000;
    rd_cycle[10095] = 1'b1;  wr_cycle[10095] = 1'b0;  addr_rom[10095]='h0000017c;  wr_data_rom[10095]='h00000000;
    rd_cycle[10096] = 1'b1;  wr_cycle[10096] = 1'b0;  addr_rom[10096]='h00000180;  wr_data_rom[10096]='h00000000;
    rd_cycle[10097] = 1'b1;  wr_cycle[10097] = 1'b0;  addr_rom[10097]='h00000184;  wr_data_rom[10097]='h00000000;
    rd_cycle[10098] = 1'b1;  wr_cycle[10098] = 1'b0;  addr_rom[10098]='h00000188;  wr_data_rom[10098]='h00000000;
    rd_cycle[10099] = 1'b1;  wr_cycle[10099] = 1'b0;  addr_rom[10099]='h0000018c;  wr_data_rom[10099]='h00000000;
    rd_cycle[10100] = 1'b1;  wr_cycle[10100] = 1'b0;  addr_rom[10100]='h00000190;  wr_data_rom[10100]='h00000000;
    rd_cycle[10101] = 1'b1;  wr_cycle[10101] = 1'b0;  addr_rom[10101]='h00000194;  wr_data_rom[10101]='h00000000;
    rd_cycle[10102] = 1'b1;  wr_cycle[10102] = 1'b0;  addr_rom[10102]='h00000198;  wr_data_rom[10102]='h00000000;
    rd_cycle[10103] = 1'b1;  wr_cycle[10103] = 1'b0;  addr_rom[10103]='h0000019c;  wr_data_rom[10103]='h00000000;
    rd_cycle[10104] = 1'b1;  wr_cycle[10104] = 1'b0;  addr_rom[10104]='h000001a0;  wr_data_rom[10104]='h00000000;
    rd_cycle[10105] = 1'b1;  wr_cycle[10105] = 1'b0;  addr_rom[10105]='h000001a4;  wr_data_rom[10105]='h00000000;
    rd_cycle[10106] = 1'b1;  wr_cycle[10106] = 1'b0;  addr_rom[10106]='h000001a8;  wr_data_rom[10106]='h00000000;
    rd_cycle[10107] = 1'b1;  wr_cycle[10107] = 1'b0;  addr_rom[10107]='h000001ac;  wr_data_rom[10107]='h00000000;
    rd_cycle[10108] = 1'b1;  wr_cycle[10108] = 1'b0;  addr_rom[10108]='h000001b0;  wr_data_rom[10108]='h00000000;
    rd_cycle[10109] = 1'b1;  wr_cycle[10109] = 1'b0;  addr_rom[10109]='h000001b4;  wr_data_rom[10109]='h00000000;
    rd_cycle[10110] = 1'b1;  wr_cycle[10110] = 1'b0;  addr_rom[10110]='h000001b8;  wr_data_rom[10110]='h00000000;
    rd_cycle[10111] = 1'b1;  wr_cycle[10111] = 1'b0;  addr_rom[10111]='h000001bc;  wr_data_rom[10111]='h00000000;
    rd_cycle[10112] = 1'b1;  wr_cycle[10112] = 1'b0;  addr_rom[10112]='h000001c0;  wr_data_rom[10112]='h00000000;
    rd_cycle[10113] = 1'b1;  wr_cycle[10113] = 1'b0;  addr_rom[10113]='h000001c4;  wr_data_rom[10113]='h00000000;
    rd_cycle[10114] = 1'b1;  wr_cycle[10114] = 1'b0;  addr_rom[10114]='h000001c8;  wr_data_rom[10114]='h00000000;
    rd_cycle[10115] = 1'b1;  wr_cycle[10115] = 1'b0;  addr_rom[10115]='h000001cc;  wr_data_rom[10115]='h00000000;
    rd_cycle[10116] = 1'b1;  wr_cycle[10116] = 1'b0;  addr_rom[10116]='h000001d0;  wr_data_rom[10116]='h00000000;
    rd_cycle[10117] = 1'b1;  wr_cycle[10117] = 1'b0;  addr_rom[10117]='h000001d4;  wr_data_rom[10117]='h00000000;
    rd_cycle[10118] = 1'b1;  wr_cycle[10118] = 1'b0;  addr_rom[10118]='h000001d8;  wr_data_rom[10118]='h00000000;
    rd_cycle[10119] = 1'b1;  wr_cycle[10119] = 1'b0;  addr_rom[10119]='h000001dc;  wr_data_rom[10119]='h00000000;
    rd_cycle[10120] = 1'b1;  wr_cycle[10120] = 1'b0;  addr_rom[10120]='h000001e0;  wr_data_rom[10120]='h00000000;
    rd_cycle[10121] = 1'b1;  wr_cycle[10121] = 1'b0;  addr_rom[10121]='h000001e4;  wr_data_rom[10121]='h00000000;
    rd_cycle[10122] = 1'b1;  wr_cycle[10122] = 1'b0;  addr_rom[10122]='h000001e8;  wr_data_rom[10122]='h00000000;
    rd_cycle[10123] = 1'b1;  wr_cycle[10123] = 1'b0;  addr_rom[10123]='h000001ec;  wr_data_rom[10123]='h00000000;
    rd_cycle[10124] = 1'b1;  wr_cycle[10124] = 1'b0;  addr_rom[10124]='h000001f0;  wr_data_rom[10124]='h00000000;
    rd_cycle[10125] = 1'b1;  wr_cycle[10125] = 1'b0;  addr_rom[10125]='h000001f4;  wr_data_rom[10125]='h00000000;
    rd_cycle[10126] = 1'b1;  wr_cycle[10126] = 1'b0;  addr_rom[10126]='h000001f8;  wr_data_rom[10126]='h00000000;
    rd_cycle[10127] = 1'b1;  wr_cycle[10127] = 1'b0;  addr_rom[10127]='h000001fc;  wr_data_rom[10127]='h00000000;
    rd_cycle[10128] = 1'b1;  wr_cycle[10128] = 1'b0;  addr_rom[10128]='h00000200;  wr_data_rom[10128]='h00000000;
    rd_cycle[10129] = 1'b1;  wr_cycle[10129] = 1'b0;  addr_rom[10129]='h00000204;  wr_data_rom[10129]='h00000000;
    rd_cycle[10130] = 1'b1;  wr_cycle[10130] = 1'b0;  addr_rom[10130]='h00000208;  wr_data_rom[10130]='h00000000;
    rd_cycle[10131] = 1'b1;  wr_cycle[10131] = 1'b0;  addr_rom[10131]='h0000020c;  wr_data_rom[10131]='h00000000;
    rd_cycle[10132] = 1'b1;  wr_cycle[10132] = 1'b0;  addr_rom[10132]='h00000210;  wr_data_rom[10132]='h00000000;
    rd_cycle[10133] = 1'b1;  wr_cycle[10133] = 1'b0;  addr_rom[10133]='h00000214;  wr_data_rom[10133]='h00000000;
    rd_cycle[10134] = 1'b1;  wr_cycle[10134] = 1'b0;  addr_rom[10134]='h00000218;  wr_data_rom[10134]='h00000000;
    rd_cycle[10135] = 1'b1;  wr_cycle[10135] = 1'b0;  addr_rom[10135]='h0000021c;  wr_data_rom[10135]='h00000000;
    rd_cycle[10136] = 1'b1;  wr_cycle[10136] = 1'b0;  addr_rom[10136]='h00000220;  wr_data_rom[10136]='h00000000;
    rd_cycle[10137] = 1'b1;  wr_cycle[10137] = 1'b0;  addr_rom[10137]='h00000224;  wr_data_rom[10137]='h00000000;
    rd_cycle[10138] = 1'b1;  wr_cycle[10138] = 1'b0;  addr_rom[10138]='h00000228;  wr_data_rom[10138]='h00000000;
    rd_cycle[10139] = 1'b1;  wr_cycle[10139] = 1'b0;  addr_rom[10139]='h0000022c;  wr_data_rom[10139]='h00000000;
    rd_cycle[10140] = 1'b1;  wr_cycle[10140] = 1'b0;  addr_rom[10140]='h00000230;  wr_data_rom[10140]='h00000000;
    rd_cycle[10141] = 1'b1;  wr_cycle[10141] = 1'b0;  addr_rom[10141]='h00000234;  wr_data_rom[10141]='h00000000;
    rd_cycle[10142] = 1'b1;  wr_cycle[10142] = 1'b0;  addr_rom[10142]='h00000238;  wr_data_rom[10142]='h00000000;
    rd_cycle[10143] = 1'b1;  wr_cycle[10143] = 1'b0;  addr_rom[10143]='h0000023c;  wr_data_rom[10143]='h00000000;
    rd_cycle[10144] = 1'b1;  wr_cycle[10144] = 1'b0;  addr_rom[10144]='h00000240;  wr_data_rom[10144]='h00000000;
    rd_cycle[10145] = 1'b1;  wr_cycle[10145] = 1'b0;  addr_rom[10145]='h00000244;  wr_data_rom[10145]='h00000000;
    rd_cycle[10146] = 1'b1;  wr_cycle[10146] = 1'b0;  addr_rom[10146]='h00000248;  wr_data_rom[10146]='h00000000;
    rd_cycle[10147] = 1'b1;  wr_cycle[10147] = 1'b0;  addr_rom[10147]='h0000024c;  wr_data_rom[10147]='h00000000;
    rd_cycle[10148] = 1'b1;  wr_cycle[10148] = 1'b0;  addr_rom[10148]='h00000250;  wr_data_rom[10148]='h00000000;
    rd_cycle[10149] = 1'b1;  wr_cycle[10149] = 1'b0;  addr_rom[10149]='h00000254;  wr_data_rom[10149]='h00000000;
    rd_cycle[10150] = 1'b1;  wr_cycle[10150] = 1'b0;  addr_rom[10150]='h00000258;  wr_data_rom[10150]='h00000000;
    rd_cycle[10151] = 1'b1;  wr_cycle[10151] = 1'b0;  addr_rom[10151]='h0000025c;  wr_data_rom[10151]='h00000000;
    rd_cycle[10152] = 1'b1;  wr_cycle[10152] = 1'b0;  addr_rom[10152]='h00000260;  wr_data_rom[10152]='h00000000;
    rd_cycle[10153] = 1'b1;  wr_cycle[10153] = 1'b0;  addr_rom[10153]='h00000264;  wr_data_rom[10153]='h00000000;
    rd_cycle[10154] = 1'b1;  wr_cycle[10154] = 1'b0;  addr_rom[10154]='h00000268;  wr_data_rom[10154]='h00000000;
    rd_cycle[10155] = 1'b1;  wr_cycle[10155] = 1'b0;  addr_rom[10155]='h0000026c;  wr_data_rom[10155]='h00000000;
    rd_cycle[10156] = 1'b1;  wr_cycle[10156] = 1'b0;  addr_rom[10156]='h00000270;  wr_data_rom[10156]='h00000000;
    rd_cycle[10157] = 1'b1;  wr_cycle[10157] = 1'b0;  addr_rom[10157]='h00000274;  wr_data_rom[10157]='h00000000;
    rd_cycle[10158] = 1'b1;  wr_cycle[10158] = 1'b0;  addr_rom[10158]='h00000278;  wr_data_rom[10158]='h00000000;
    rd_cycle[10159] = 1'b1;  wr_cycle[10159] = 1'b0;  addr_rom[10159]='h0000027c;  wr_data_rom[10159]='h00000000;
    rd_cycle[10160] = 1'b1;  wr_cycle[10160] = 1'b0;  addr_rom[10160]='h00000280;  wr_data_rom[10160]='h00000000;
    rd_cycle[10161] = 1'b1;  wr_cycle[10161] = 1'b0;  addr_rom[10161]='h00000284;  wr_data_rom[10161]='h00000000;
    rd_cycle[10162] = 1'b1;  wr_cycle[10162] = 1'b0;  addr_rom[10162]='h00000288;  wr_data_rom[10162]='h00000000;
    rd_cycle[10163] = 1'b1;  wr_cycle[10163] = 1'b0;  addr_rom[10163]='h0000028c;  wr_data_rom[10163]='h00000000;
    rd_cycle[10164] = 1'b1;  wr_cycle[10164] = 1'b0;  addr_rom[10164]='h00000290;  wr_data_rom[10164]='h00000000;
    rd_cycle[10165] = 1'b1;  wr_cycle[10165] = 1'b0;  addr_rom[10165]='h00000294;  wr_data_rom[10165]='h00000000;
    rd_cycle[10166] = 1'b1;  wr_cycle[10166] = 1'b0;  addr_rom[10166]='h00000298;  wr_data_rom[10166]='h00000000;
    rd_cycle[10167] = 1'b1;  wr_cycle[10167] = 1'b0;  addr_rom[10167]='h0000029c;  wr_data_rom[10167]='h00000000;
    rd_cycle[10168] = 1'b1;  wr_cycle[10168] = 1'b0;  addr_rom[10168]='h000002a0;  wr_data_rom[10168]='h00000000;
    rd_cycle[10169] = 1'b1;  wr_cycle[10169] = 1'b0;  addr_rom[10169]='h000002a4;  wr_data_rom[10169]='h00000000;
    rd_cycle[10170] = 1'b1;  wr_cycle[10170] = 1'b0;  addr_rom[10170]='h000002a8;  wr_data_rom[10170]='h00000000;
    rd_cycle[10171] = 1'b1;  wr_cycle[10171] = 1'b0;  addr_rom[10171]='h000002ac;  wr_data_rom[10171]='h00000000;
    rd_cycle[10172] = 1'b1;  wr_cycle[10172] = 1'b0;  addr_rom[10172]='h000002b0;  wr_data_rom[10172]='h00000000;
    rd_cycle[10173] = 1'b1;  wr_cycle[10173] = 1'b0;  addr_rom[10173]='h000002b4;  wr_data_rom[10173]='h00000000;
    rd_cycle[10174] = 1'b1;  wr_cycle[10174] = 1'b0;  addr_rom[10174]='h000002b8;  wr_data_rom[10174]='h00000000;
    rd_cycle[10175] = 1'b1;  wr_cycle[10175] = 1'b0;  addr_rom[10175]='h000002bc;  wr_data_rom[10175]='h00000000;
    rd_cycle[10176] = 1'b1;  wr_cycle[10176] = 1'b0;  addr_rom[10176]='h000002c0;  wr_data_rom[10176]='h00000000;
    rd_cycle[10177] = 1'b1;  wr_cycle[10177] = 1'b0;  addr_rom[10177]='h000002c4;  wr_data_rom[10177]='h00000000;
    rd_cycle[10178] = 1'b1;  wr_cycle[10178] = 1'b0;  addr_rom[10178]='h000002c8;  wr_data_rom[10178]='h00000000;
    rd_cycle[10179] = 1'b1;  wr_cycle[10179] = 1'b0;  addr_rom[10179]='h000002cc;  wr_data_rom[10179]='h00000000;
    rd_cycle[10180] = 1'b1;  wr_cycle[10180] = 1'b0;  addr_rom[10180]='h000002d0;  wr_data_rom[10180]='h00000000;
    rd_cycle[10181] = 1'b1;  wr_cycle[10181] = 1'b0;  addr_rom[10181]='h000002d4;  wr_data_rom[10181]='h00000000;
    rd_cycle[10182] = 1'b1;  wr_cycle[10182] = 1'b0;  addr_rom[10182]='h000002d8;  wr_data_rom[10182]='h00000000;
    rd_cycle[10183] = 1'b1;  wr_cycle[10183] = 1'b0;  addr_rom[10183]='h000002dc;  wr_data_rom[10183]='h00000000;
    rd_cycle[10184] = 1'b1;  wr_cycle[10184] = 1'b0;  addr_rom[10184]='h000002e0;  wr_data_rom[10184]='h00000000;
    rd_cycle[10185] = 1'b1;  wr_cycle[10185] = 1'b0;  addr_rom[10185]='h000002e4;  wr_data_rom[10185]='h00000000;
    rd_cycle[10186] = 1'b1;  wr_cycle[10186] = 1'b0;  addr_rom[10186]='h000002e8;  wr_data_rom[10186]='h00000000;
    rd_cycle[10187] = 1'b1;  wr_cycle[10187] = 1'b0;  addr_rom[10187]='h000002ec;  wr_data_rom[10187]='h00000000;
    rd_cycle[10188] = 1'b1;  wr_cycle[10188] = 1'b0;  addr_rom[10188]='h000002f0;  wr_data_rom[10188]='h00000000;
    rd_cycle[10189] = 1'b1;  wr_cycle[10189] = 1'b0;  addr_rom[10189]='h000002f4;  wr_data_rom[10189]='h00000000;
    rd_cycle[10190] = 1'b1;  wr_cycle[10190] = 1'b0;  addr_rom[10190]='h000002f8;  wr_data_rom[10190]='h00000000;
    rd_cycle[10191] = 1'b1;  wr_cycle[10191] = 1'b0;  addr_rom[10191]='h000002fc;  wr_data_rom[10191]='h00000000;
    rd_cycle[10192] = 1'b1;  wr_cycle[10192] = 1'b0;  addr_rom[10192]='h00000300;  wr_data_rom[10192]='h00000000;
    rd_cycle[10193] = 1'b1;  wr_cycle[10193] = 1'b0;  addr_rom[10193]='h00000304;  wr_data_rom[10193]='h00000000;
    rd_cycle[10194] = 1'b1;  wr_cycle[10194] = 1'b0;  addr_rom[10194]='h00000308;  wr_data_rom[10194]='h00000000;
    rd_cycle[10195] = 1'b1;  wr_cycle[10195] = 1'b0;  addr_rom[10195]='h0000030c;  wr_data_rom[10195]='h00000000;
    rd_cycle[10196] = 1'b1;  wr_cycle[10196] = 1'b0;  addr_rom[10196]='h00000310;  wr_data_rom[10196]='h00000000;
    rd_cycle[10197] = 1'b1;  wr_cycle[10197] = 1'b0;  addr_rom[10197]='h00000314;  wr_data_rom[10197]='h00000000;
    rd_cycle[10198] = 1'b1;  wr_cycle[10198] = 1'b0;  addr_rom[10198]='h00000318;  wr_data_rom[10198]='h00000000;
    rd_cycle[10199] = 1'b1;  wr_cycle[10199] = 1'b0;  addr_rom[10199]='h0000031c;  wr_data_rom[10199]='h00000000;
    rd_cycle[10200] = 1'b1;  wr_cycle[10200] = 1'b0;  addr_rom[10200]='h00000320;  wr_data_rom[10200]='h00000000;
    rd_cycle[10201] = 1'b1;  wr_cycle[10201] = 1'b0;  addr_rom[10201]='h00000324;  wr_data_rom[10201]='h00000000;
    rd_cycle[10202] = 1'b1;  wr_cycle[10202] = 1'b0;  addr_rom[10202]='h00000328;  wr_data_rom[10202]='h00000000;
    rd_cycle[10203] = 1'b1;  wr_cycle[10203] = 1'b0;  addr_rom[10203]='h0000032c;  wr_data_rom[10203]='h00000000;
    rd_cycle[10204] = 1'b1;  wr_cycle[10204] = 1'b0;  addr_rom[10204]='h00000330;  wr_data_rom[10204]='h00000000;
    rd_cycle[10205] = 1'b1;  wr_cycle[10205] = 1'b0;  addr_rom[10205]='h00000334;  wr_data_rom[10205]='h00000000;
    rd_cycle[10206] = 1'b1;  wr_cycle[10206] = 1'b0;  addr_rom[10206]='h00000338;  wr_data_rom[10206]='h00000000;
    rd_cycle[10207] = 1'b1;  wr_cycle[10207] = 1'b0;  addr_rom[10207]='h0000033c;  wr_data_rom[10207]='h00000000;
    rd_cycle[10208] = 1'b1;  wr_cycle[10208] = 1'b0;  addr_rom[10208]='h00000340;  wr_data_rom[10208]='h00000000;
    rd_cycle[10209] = 1'b1;  wr_cycle[10209] = 1'b0;  addr_rom[10209]='h00000344;  wr_data_rom[10209]='h00000000;
    rd_cycle[10210] = 1'b1;  wr_cycle[10210] = 1'b0;  addr_rom[10210]='h00000348;  wr_data_rom[10210]='h00000000;
    rd_cycle[10211] = 1'b1;  wr_cycle[10211] = 1'b0;  addr_rom[10211]='h0000034c;  wr_data_rom[10211]='h00000000;
    rd_cycle[10212] = 1'b1;  wr_cycle[10212] = 1'b0;  addr_rom[10212]='h00000350;  wr_data_rom[10212]='h00000000;
    rd_cycle[10213] = 1'b1;  wr_cycle[10213] = 1'b0;  addr_rom[10213]='h00000354;  wr_data_rom[10213]='h00000000;
    rd_cycle[10214] = 1'b1;  wr_cycle[10214] = 1'b0;  addr_rom[10214]='h00000358;  wr_data_rom[10214]='h00000000;
    rd_cycle[10215] = 1'b1;  wr_cycle[10215] = 1'b0;  addr_rom[10215]='h0000035c;  wr_data_rom[10215]='h00000000;
    rd_cycle[10216] = 1'b1;  wr_cycle[10216] = 1'b0;  addr_rom[10216]='h00000360;  wr_data_rom[10216]='h00000000;
    rd_cycle[10217] = 1'b1;  wr_cycle[10217] = 1'b0;  addr_rom[10217]='h00000364;  wr_data_rom[10217]='h00000000;
    rd_cycle[10218] = 1'b1;  wr_cycle[10218] = 1'b0;  addr_rom[10218]='h00000368;  wr_data_rom[10218]='h00000000;
    rd_cycle[10219] = 1'b1;  wr_cycle[10219] = 1'b0;  addr_rom[10219]='h0000036c;  wr_data_rom[10219]='h00000000;
    rd_cycle[10220] = 1'b1;  wr_cycle[10220] = 1'b0;  addr_rom[10220]='h00000370;  wr_data_rom[10220]='h00000000;
    rd_cycle[10221] = 1'b1;  wr_cycle[10221] = 1'b0;  addr_rom[10221]='h00000374;  wr_data_rom[10221]='h00000000;
    rd_cycle[10222] = 1'b1;  wr_cycle[10222] = 1'b0;  addr_rom[10222]='h00000378;  wr_data_rom[10222]='h00000000;
    rd_cycle[10223] = 1'b1;  wr_cycle[10223] = 1'b0;  addr_rom[10223]='h0000037c;  wr_data_rom[10223]='h00000000;
    rd_cycle[10224] = 1'b1;  wr_cycle[10224] = 1'b0;  addr_rom[10224]='h00000380;  wr_data_rom[10224]='h00000000;
    rd_cycle[10225] = 1'b1;  wr_cycle[10225] = 1'b0;  addr_rom[10225]='h00000384;  wr_data_rom[10225]='h00000000;
    rd_cycle[10226] = 1'b1;  wr_cycle[10226] = 1'b0;  addr_rom[10226]='h00000388;  wr_data_rom[10226]='h00000000;
    rd_cycle[10227] = 1'b1;  wr_cycle[10227] = 1'b0;  addr_rom[10227]='h0000038c;  wr_data_rom[10227]='h00000000;
    rd_cycle[10228] = 1'b1;  wr_cycle[10228] = 1'b0;  addr_rom[10228]='h00000390;  wr_data_rom[10228]='h00000000;
    rd_cycle[10229] = 1'b1;  wr_cycle[10229] = 1'b0;  addr_rom[10229]='h00000394;  wr_data_rom[10229]='h00000000;
    rd_cycle[10230] = 1'b1;  wr_cycle[10230] = 1'b0;  addr_rom[10230]='h00000398;  wr_data_rom[10230]='h00000000;
    rd_cycle[10231] = 1'b1;  wr_cycle[10231] = 1'b0;  addr_rom[10231]='h0000039c;  wr_data_rom[10231]='h00000000;
    rd_cycle[10232] = 1'b1;  wr_cycle[10232] = 1'b0;  addr_rom[10232]='h000003a0;  wr_data_rom[10232]='h00000000;
    rd_cycle[10233] = 1'b1;  wr_cycle[10233] = 1'b0;  addr_rom[10233]='h000003a4;  wr_data_rom[10233]='h00000000;
    rd_cycle[10234] = 1'b1;  wr_cycle[10234] = 1'b0;  addr_rom[10234]='h000003a8;  wr_data_rom[10234]='h00000000;
    rd_cycle[10235] = 1'b1;  wr_cycle[10235] = 1'b0;  addr_rom[10235]='h000003ac;  wr_data_rom[10235]='h00000000;
    rd_cycle[10236] = 1'b1;  wr_cycle[10236] = 1'b0;  addr_rom[10236]='h000003b0;  wr_data_rom[10236]='h00000000;
    rd_cycle[10237] = 1'b1;  wr_cycle[10237] = 1'b0;  addr_rom[10237]='h000003b4;  wr_data_rom[10237]='h00000000;
    rd_cycle[10238] = 1'b1;  wr_cycle[10238] = 1'b0;  addr_rom[10238]='h000003b8;  wr_data_rom[10238]='h00000000;
    rd_cycle[10239] = 1'b1;  wr_cycle[10239] = 1'b0;  addr_rom[10239]='h000003bc;  wr_data_rom[10239]='h00000000;
    rd_cycle[10240] = 1'b1;  wr_cycle[10240] = 1'b0;  addr_rom[10240]='h000003c0;  wr_data_rom[10240]='h00000000;
    rd_cycle[10241] = 1'b1;  wr_cycle[10241] = 1'b0;  addr_rom[10241]='h000003c4;  wr_data_rom[10241]='h00000000;
    rd_cycle[10242] = 1'b1;  wr_cycle[10242] = 1'b0;  addr_rom[10242]='h000003c8;  wr_data_rom[10242]='h00000000;
    rd_cycle[10243] = 1'b1;  wr_cycle[10243] = 1'b0;  addr_rom[10243]='h000003cc;  wr_data_rom[10243]='h00000000;
    rd_cycle[10244] = 1'b1;  wr_cycle[10244] = 1'b0;  addr_rom[10244]='h000003d0;  wr_data_rom[10244]='h00000000;
    rd_cycle[10245] = 1'b1;  wr_cycle[10245] = 1'b0;  addr_rom[10245]='h000003d4;  wr_data_rom[10245]='h00000000;
    rd_cycle[10246] = 1'b1;  wr_cycle[10246] = 1'b0;  addr_rom[10246]='h000003d8;  wr_data_rom[10246]='h00000000;
    rd_cycle[10247] = 1'b1;  wr_cycle[10247] = 1'b0;  addr_rom[10247]='h000003dc;  wr_data_rom[10247]='h00000000;
    rd_cycle[10248] = 1'b1;  wr_cycle[10248] = 1'b0;  addr_rom[10248]='h000003e0;  wr_data_rom[10248]='h00000000;
    rd_cycle[10249] = 1'b1;  wr_cycle[10249] = 1'b0;  addr_rom[10249]='h000003e4;  wr_data_rom[10249]='h00000000;
    rd_cycle[10250] = 1'b1;  wr_cycle[10250] = 1'b0;  addr_rom[10250]='h000003e8;  wr_data_rom[10250]='h00000000;
    rd_cycle[10251] = 1'b1;  wr_cycle[10251] = 1'b0;  addr_rom[10251]='h000003ec;  wr_data_rom[10251]='h00000000;
    rd_cycle[10252] = 1'b1;  wr_cycle[10252] = 1'b0;  addr_rom[10252]='h000003f0;  wr_data_rom[10252]='h00000000;
    rd_cycle[10253] = 1'b1;  wr_cycle[10253] = 1'b0;  addr_rom[10253]='h000003f4;  wr_data_rom[10253]='h00000000;
    rd_cycle[10254] = 1'b1;  wr_cycle[10254] = 1'b0;  addr_rom[10254]='h000003f8;  wr_data_rom[10254]='h00000000;
    rd_cycle[10255] = 1'b1;  wr_cycle[10255] = 1'b0;  addr_rom[10255]='h000003fc;  wr_data_rom[10255]='h00000000;
    rd_cycle[10256] = 1'b1;  wr_cycle[10256] = 1'b0;  addr_rom[10256]='h00000400;  wr_data_rom[10256]='h00000000;
    rd_cycle[10257] = 1'b1;  wr_cycle[10257] = 1'b0;  addr_rom[10257]='h00000404;  wr_data_rom[10257]='h00000000;
    rd_cycle[10258] = 1'b1;  wr_cycle[10258] = 1'b0;  addr_rom[10258]='h00000408;  wr_data_rom[10258]='h00000000;
    rd_cycle[10259] = 1'b1;  wr_cycle[10259] = 1'b0;  addr_rom[10259]='h0000040c;  wr_data_rom[10259]='h00000000;
    rd_cycle[10260] = 1'b1;  wr_cycle[10260] = 1'b0;  addr_rom[10260]='h00000410;  wr_data_rom[10260]='h00000000;
    rd_cycle[10261] = 1'b1;  wr_cycle[10261] = 1'b0;  addr_rom[10261]='h00000414;  wr_data_rom[10261]='h00000000;
    rd_cycle[10262] = 1'b1;  wr_cycle[10262] = 1'b0;  addr_rom[10262]='h00000418;  wr_data_rom[10262]='h00000000;
    rd_cycle[10263] = 1'b1;  wr_cycle[10263] = 1'b0;  addr_rom[10263]='h0000041c;  wr_data_rom[10263]='h00000000;
    rd_cycle[10264] = 1'b1;  wr_cycle[10264] = 1'b0;  addr_rom[10264]='h00000420;  wr_data_rom[10264]='h00000000;
    rd_cycle[10265] = 1'b1;  wr_cycle[10265] = 1'b0;  addr_rom[10265]='h00000424;  wr_data_rom[10265]='h00000000;
    rd_cycle[10266] = 1'b1;  wr_cycle[10266] = 1'b0;  addr_rom[10266]='h00000428;  wr_data_rom[10266]='h00000000;
    rd_cycle[10267] = 1'b1;  wr_cycle[10267] = 1'b0;  addr_rom[10267]='h0000042c;  wr_data_rom[10267]='h00000000;
    rd_cycle[10268] = 1'b1;  wr_cycle[10268] = 1'b0;  addr_rom[10268]='h00000430;  wr_data_rom[10268]='h00000000;
    rd_cycle[10269] = 1'b1;  wr_cycle[10269] = 1'b0;  addr_rom[10269]='h00000434;  wr_data_rom[10269]='h00000000;
    rd_cycle[10270] = 1'b1;  wr_cycle[10270] = 1'b0;  addr_rom[10270]='h00000438;  wr_data_rom[10270]='h00000000;
    rd_cycle[10271] = 1'b1;  wr_cycle[10271] = 1'b0;  addr_rom[10271]='h0000043c;  wr_data_rom[10271]='h00000000;
    rd_cycle[10272] = 1'b1;  wr_cycle[10272] = 1'b0;  addr_rom[10272]='h00000440;  wr_data_rom[10272]='h00000000;
    rd_cycle[10273] = 1'b1;  wr_cycle[10273] = 1'b0;  addr_rom[10273]='h00000444;  wr_data_rom[10273]='h00000000;
    rd_cycle[10274] = 1'b1;  wr_cycle[10274] = 1'b0;  addr_rom[10274]='h00000448;  wr_data_rom[10274]='h00000000;
    rd_cycle[10275] = 1'b1;  wr_cycle[10275] = 1'b0;  addr_rom[10275]='h0000044c;  wr_data_rom[10275]='h00000000;
    rd_cycle[10276] = 1'b1;  wr_cycle[10276] = 1'b0;  addr_rom[10276]='h00000450;  wr_data_rom[10276]='h00000000;
    rd_cycle[10277] = 1'b1;  wr_cycle[10277] = 1'b0;  addr_rom[10277]='h00000454;  wr_data_rom[10277]='h00000000;
    rd_cycle[10278] = 1'b1;  wr_cycle[10278] = 1'b0;  addr_rom[10278]='h00000458;  wr_data_rom[10278]='h00000000;
    rd_cycle[10279] = 1'b1;  wr_cycle[10279] = 1'b0;  addr_rom[10279]='h0000045c;  wr_data_rom[10279]='h00000000;
    rd_cycle[10280] = 1'b1;  wr_cycle[10280] = 1'b0;  addr_rom[10280]='h00000460;  wr_data_rom[10280]='h00000000;
    rd_cycle[10281] = 1'b1;  wr_cycle[10281] = 1'b0;  addr_rom[10281]='h00000464;  wr_data_rom[10281]='h00000000;
    rd_cycle[10282] = 1'b1;  wr_cycle[10282] = 1'b0;  addr_rom[10282]='h00000468;  wr_data_rom[10282]='h00000000;
    rd_cycle[10283] = 1'b1;  wr_cycle[10283] = 1'b0;  addr_rom[10283]='h0000046c;  wr_data_rom[10283]='h00000000;
    rd_cycle[10284] = 1'b1;  wr_cycle[10284] = 1'b0;  addr_rom[10284]='h00000470;  wr_data_rom[10284]='h00000000;
    rd_cycle[10285] = 1'b1;  wr_cycle[10285] = 1'b0;  addr_rom[10285]='h00000474;  wr_data_rom[10285]='h00000000;
    rd_cycle[10286] = 1'b1;  wr_cycle[10286] = 1'b0;  addr_rom[10286]='h00000478;  wr_data_rom[10286]='h00000000;
    rd_cycle[10287] = 1'b1;  wr_cycle[10287] = 1'b0;  addr_rom[10287]='h0000047c;  wr_data_rom[10287]='h00000000;
    rd_cycle[10288] = 1'b1;  wr_cycle[10288] = 1'b0;  addr_rom[10288]='h00000480;  wr_data_rom[10288]='h00000000;
    rd_cycle[10289] = 1'b1;  wr_cycle[10289] = 1'b0;  addr_rom[10289]='h00000484;  wr_data_rom[10289]='h00000000;
    rd_cycle[10290] = 1'b1;  wr_cycle[10290] = 1'b0;  addr_rom[10290]='h00000488;  wr_data_rom[10290]='h00000000;
    rd_cycle[10291] = 1'b1;  wr_cycle[10291] = 1'b0;  addr_rom[10291]='h0000048c;  wr_data_rom[10291]='h00000000;
    rd_cycle[10292] = 1'b1;  wr_cycle[10292] = 1'b0;  addr_rom[10292]='h00000490;  wr_data_rom[10292]='h00000000;
    rd_cycle[10293] = 1'b1;  wr_cycle[10293] = 1'b0;  addr_rom[10293]='h00000494;  wr_data_rom[10293]='h00000000;
    rd_cycle[10294] = 1'b1;  wr_cycle[10294] = 1'b0;  addr_rom[10294]='h00000498;  wr_data_rom[10294]='h00000000;
    rd_cycle[10295] = 1'b1;  wr_cycle[10295] = 1'b0;  addr_rom[10295]='h0000049c;  wr_data_rom[10295]='h00000000;
    rd_cycle[10296] = 1'b1;  wr_cycle[10296] = 1'b0;  addr_rom[10296]='h000004a0;  wr_data_rom[10296]='h00000000;
    rd_cycle[10297] = 1'b1;  wr_cycle[10297] = 1'b0;  addr_rom[10297]='h000004a4;  wr_data_rom[10297]='h00000000;
    rd_cycle[10298] = 1'b1;  wr_cycle[10298] = 1'b0;  addr_rom[10298]='h000004a8;  wr_data_rom[10298]='h00000000;
    rd_cycle[10299] = 1'b1;  wr_cycle[10299] = 1'b0;  addr_rom[10299]='h000004ac;  wr_data_rom[10299]='h00000000;
    rd_cycle[10300] = 1'b1;  wr_cycle[10300] = 1'b0;  addr_rom[10300]='h000004b0;  wr_data_rom[10300]='h00000000;
    rd_cycle[10301] = 1'b1;  wr_cycle[10301] = 1'b0;  addr_rom[10301]='h000004b4;  wr_data_rom[10301]='h00000000;
    rd_cycle[10302] = 1'b1;  wr_cycle[10302] = 1'b0;  addr_rom[10302]='h000004b8;  wr_data_rom[10302]='h00000000;
    rd_cycle[10303] = 1'b1;  wr_cycle[10303] = 1'b0;  addr_rom[10303]='h000004bc;  wr_data_rom[10303]='h00000000;
    rd_cycle[10304] = 1'b1;  wr_cycle[10304] = 1'b0;  addr_rom[10304]='h000004c0;  wr_data_rom[10304]='h00000000;
    rd_cycle[10305] = 1'b1;  wr_cycle[10305] = 1'b0;  addr_rom[10305]='h000004c4;  wr_data_rom[10305]='h00000000;
    rd_cycle[10306] = 1'b1;  wr_cycle[10306] = 1'b0;  addr_rom[10306]='h000004c8;  wr_data_rom[10306]='h00000000;
    rd_cycle[10307] = 1'b1;  wr_cycle[10307] = 1'b0;  addr_rom[10307]='h000004cc;  wr_data_rom[10307]='h00000000;
    rd_cycle[10308] = 1'b1;  wr_cycle[10308] = 1'b0;  addr_rom[10308]='h000004d0;  wr_data_rom[10308]='h00000000;
    rd_cycle[10309] = 1'b1;  wr_cycle[10309] = 1'b0;  addr_rom[10309]='h000004d4;  wr_data_rom[10309]='h00000000;
    rd_cycle[10310] = 1'b1;  wr_cycle[10310] = 1'b0;  addr_rom[10310]='h000004d8;  wr_data_rom[10310]='h00000000;
    rd_cycle[10311] = 1'b1;  wr_cycle[10311] = 1'b0;  addr_rom[10311]='h000004dc;  wr_data_rom[10311]='h00000000;
    rd_cycle[10312] = 1'b1;  wr_cycle[10312] = 1'b0;  addr_rom[10312]='h000004e0;  wr_data_rom[10312]='h00000000;
    rd_cycle[10313] = 1'b1;  wr_cycle[10313] = 1'b0;  addr_rom[10313]='h000004e4;  wr_data_rom[10313]='h00000000;
    rd_cycle[10314] = 1'b1;  wr_cycle[10314] = 1'b0;  addr_rom[10314]='h000004e8;  wr_data_rom[10314]='h00000000;
    rd_cycle[10315] = 1'b1;  wr_cycle[10315] = 1'b0;  addr_rom[10315]='h000004ec;  wr_data_rom[10315]='h00000000;
    rd_cycle[10316] = 1'b1;  wr_cycle[10316] = 1'b0;  addr_rom[10316]='h000004f0;  wr_data_rom[10316]='h00000000;
    rd_cycle[10317] = 1'b1;  wr_cycle[10317] = 1'b0;  addr_rom[10317]='h000004f4;  wr_data_rom[10317]='h00000000;
    rd_cycle[10318] = 1'b1;  wr_cycle[10318] = 1'b0;  addr_rom[10318]='h000004f8;  wr_data_rom[10318]='h00000000;
    rd_cycle[10319] = 1'b1;  wr_cycle[10319] = 1'b0;  addr_rom[10319]='h000004fc;  wr_data_rom[10319]='h00000000;
    rd_cycle[10320] = 1'b1;  wr_cycle[10320] = 1'b0;  addr_rom[10320]='h00000500;  wr_data_rom[10320]='h00000000;
    rd_cycle[10321] = 1'b1;  wr_cycle[10321] = 1'b0;  addr_rom[10321]='h00000504;  wr_data_rom[10321]='h00000000;
    rd_cycle[10322] = 1'b1;  wr_cycle[10322] = 1'b0;  addr_rom[10322]='h00000508;  wr_data_rom[10322]='h00000000;
    rd_cycle[10323] = 1'b1;  wr_cycle[10323] = 1'b0;  addr_rom[10323]='h0000050c;  wr_data_rom[10323]='h00000000;
    rd_cycle[10324] = 1'b1;  wr_cycle[10324] = 1'b0;  addr_rom[10324]='h00000510;  wr_data_rom[10324]='h00000000;
    rd_cycle[10325] = 1'b1;  wr_cycle[10325] = 1'b0;  addr_rom[10325]='h00000514;  wr_data_rom[10325]='h00000000;
    rd_cycle[10326] = 1'b1;  wr_cycle[10326] = 1'b0;  addr_rom[10326]='h00000518;  wr_data_rom[10326]='h00000000;
    rd_cycle[10327] = 1'b1;  wr_cycle[10327] = 1'b0;  addr_rom[10327]='h0000051c;  wr_data_rom[10327]='h00000000;
    rd_cycle[10328] = 1'b1;  wr_cycle[10328] = 1'b0;  addr_rom[10328]='h00000520;  wr_data_rom[10328]='h00000000;
    rd_cycle[10329] = 1'b1;  wr_cycle[10329] = 1'b0;  addr_rom[10329]='h00000524;  wr_data_rom[10329]='h00000000;
    rd_cycle[10330] = 1'b1;  wr_cycle[10330] = 1'b0;  addr_rom[10330]='h00000528;  wr_data_rom[10330]='h00000000;
    rd_cycle[10331] = 1'b1;  wr_cycle[10331] = 1'b0;  addr_rom[10331]='h0000052c;  wr_data_rom[10331]='h00000000;
    rd_cycle[10332] = 1'b1;  wr_cycle[10332] = 1'b0;  addr_rom[10332]='h00000530;  wr_data_rom[10332]='h00000000;
    rd_cycle[10333] = 1'b1;  wr_cycle[10333] = 1'b0;  addr_rom[10333]='h00000534;  wr_data_rom[10333]='h00000000;
    rd_cycle[10334] = 1'b1;  wr_cycle[10334] = 1'b0;  addr_rom[10334]='h00000538;  wr_data_rom[10334]='h00000000;
    rd_cycle[10335] = 1'b1;  wr_cycle[10335] = 1'b0;  addr_rom[10335]='h0000053c;  wr_data_rom[10335]='h00000000;
    rd_cycle[10336] = 1'b1;  wr_cycle[10336] = 1'b0;  addr_rom[10336]='h00000540;  wr_data_rom[10336]='h00000000;
    rd_cycle[10337] = 1'b1;  wr_cycle[10337] = 1'b0;  addr_rom[10337]='h00000544;  wr_data_rom[10337]='h00000000;
    rd_cycle[10338] = 1'b1;  wr_cycle[10338] = 1'b0;  addr_rom[10338]='h00000548;  wr_data_rom[10338]='h00000000;
    rd_cycle[10339] = 1'b1;  wr_cycle[10339] = 1'b0;  addr_rom[10339]='h0000054c;  wr_data_rom[10339]='h00000000;
    rd_cycle[10340] = 1'b1;  wr_cycle[10340] = 1'b0;  addr_rom[10340]='h00000550;  wr_data_rom[10340]='h00000000;
    rd_cycle[10341] = 1'b1;  wr_cycle[10341] = 1'b0;  addr_rom[10341]='h00000554;  wr_data_rom[10341]='h00000000;
    rd_cycle[10342] = 1'b1;  wr_cycle[10342] = 1'b0;  addr_rom[10342]='h00000558;  wr_data_rom[10342]='h00000000;
    rd_cycle[10343] = 1'b1;  wr_cycle[10343] = 1'b0;  addr_rom[10343]='h0000055c;  wr_data_rom[10343]='h00000000;
    rd_cycle[10344] = 1'b1;  wr_cycle[10344] = 1'b0;  addr_rom[10344]='h00000560;  wr_data_rom[10344]='h00000000;
    rd_cycle[10345] = 1'b1;  wr_cycle[10345] = 1'b0;  addr_rom[10345]='h00000564;  wr_data_rom[10345]='h00000000;
    rd_cycle[10346] = 1'b1;  wr_cycle[10346] = 1'b0;  addr_rom[10346]='h00000568;  wr_data_rom[10346]='h00000000;
    rd_cycle[10347] = 1'b1;  wr_cycle[10347] = 1'b0;  addr_rom[10347]='h0000056c;  wr_data_rom[10347]='h00000000;
    rd_cycle[10348] = 1'b1;  wr_cycle[10348] = 1'b0;  addr_rom[10348]='h00000570;  wr_data_rom[10348]='h00000000;
    rd_cycle[10349] = 1'b1;  wr_cycle[10349] = 1'b0;  addr_rom[10349]='h00000574;  wr_data_rom[10349]='h00000000;
    rd_cycle[10350] = 1'b1;  wr_cycle[10350] = 1'b0;  addr_rom[10350]='h00000578;  wr_data_rom[10350]='h00000000;
    rd_cycle[10351] = 1'b1;  wr_cycle[10351] = 1'b0;  addr_rom[10351]='h0000057c;  wr_data_rom[10351]='h00000000;
    rd_cycle[10352] = 1'b1;  wr_cycle[10352] = 1'b0;  addr_rom[10352]='h00000580;  wr_data_rom[10352]='h00000000;
    rd_cycle[10353] = 1'b1;  wr_cycle[10353] = 1'b0;  addr_rom[10353]='h00000584;  wr_data_rom[10353]='h00000000;
    rd_cycle[10354] = 1'b1;  wr_cycle[10354] = 1'b0;  addr_rom[10354]='h00000588;  wr_data_rom[10354]='h00000000;
    rd_cycle[10355] = 1'b1;  wr_cycle[10355] = 1'b0;  addr_rom[10355]='h0000058c;  wr_data_rom[10355]='h00000000;
    rd_cycle[10356] = 1'b1;  wr_cycle[10356] = 1'b0;  addr_rom[10356]='h00000590;  wr_data_rom[10356]='h00000000;
    rd_cycle[10357] = 1'b1;  wr_cycle[10357] = 1'b0;  addr_rom[10357]='h00000594;  wr_data_rom[10357]='h00000000;
    rd_cycle[10358] = 1'b1;  wr_cycle[10358] = 1'b0;  addr_rom[10358]='h00000598;  wr_data_rom[10358]='h00000000;
    rd_cycle[10359] = 1'b1;  wr_cycle[10359] = 1'b0;  addr_rom[10359]='h0000059c;  wr_data_rom[10359]='h00000000;
    rd_cycle[10360] = 1'b1;  wr_cycle[10360] = 1'b0;  addr_rom[10360]='h000005a0;  wr_data_rom[10360]='h00000000;
    rd_cycle[10361] = 1'b1;  wr_cycle[10361] = 1'b0;  addr_rom[10361]='h000005a4;  wr_data_rom[10361]='h00000000;
    rd_cycle[10362] = 1'b1;  wr_cycle[10362] = 1'b0;  addr_rom[10362]='h000005a8;  wr_data_rom[10362]='h00000000;
    rd_cycle[10363] = 1'b1;  wr_cycle[10363] = 1'b0;  addr_rom[10363]='h000005ac;  wr_data_rom[10363]='h00000000;
    rd_cycle[10364] = 1'b1;  wr_cycle[10364] = 1'b0;  addr_rom[10364]='h000005b0;  wr_data_rom[10364]='h00000000;
    rd_cycle[10365] = 1'b1;  wr_cycle[10365] = 1'b0;  addr_rom[10365]='h000005b4;  wr_data_rom[10365]='h00000000;
    rd_cycle[10366] = 1'b1;  wr_cycle[10366] = 1'b0;  addr_rom[10366]='h000005b8;  wr_data_rom[10366]='h00000000;
    rd_cycle[10367] = 1'b1;  wr_cycle[10367] = 1'b0;  addr_rom[10367]='h000005bc;  wr_data_rom[10367]='h00000000;
    rd_cycle[10368] = 1'b1;  wr_cycle[10368] = 1'b0;  addr_rom[10368]='h000005c0;  wr_data_rom[10368]='h00000000;
    rd_cycle[10369] = 1'b1;  wr_cycle[10369] = 1'b0;  addr_rom[10369]='h000005c4;  wr_data_rom[10369]='h00000000;
    rd_cycle[10370] = 1'b1;  wr_cycle[10370] = 1'b0;  addr_rom[10370]='h000005c8;  wr_data_rom[10370]='h00000000;
    rd_cycle[10371] = 1'b1;  wr_cycle[10371] = 1'b0;  addr_rom[10371]='h000005cc;  wr_data_rom[10371]='h00000000;
    rd_cycle[10372] = 1'b1;  wr_cycle[10372] = 1'b0;  addr_rom[10372]='h000005d0;  wr_data_rom[10372]='h00000000;
    rd_cycle[10373] = 1'b1;  wr_cycle[10373] = 1'b0;  addr_rom[10373]='h000005d4;  wr_data_rom[10373]='h00000000;
    rd_cycle[10374] = 1'b1;  wr_cycle[10374] = 1'b0;  addr_rom[10374]='h000005d8;  wr_data_rom[10374]='h00000000;
    rd_cycle[10375] = 1'b1;  wr_cycle[10375] = 1'b0;  addr_rom[10375]='h000005dc;  wr_data_rom[10375]='h00000000;
    rd_cycle[10376] = 1'b1;  wr_cycle[10376] = 1'b0;  addr_rom[10376]='h000005e0;  wr_data_rom[10376]='h00000000;
    rd_cycle[10377] = 1'b1;  wr_cycle[10377] = 1'b0;  addr_rom[10377]='h000005e4;  wr_data_rom[10377]='h00000000;
    rd_cycle[10378] = 1'b1;  wr_cycle[10378] = 1'b0;  addr_rom[10378]='h000005e8;  wr_data_rom[10378]='h00000000;
    rd_cycle[10379] = 1'b1;  wr_cycle[10379] = 1'b0;  addr_rom[10379]='h000005ec;  wr_data_rom[10379]='h00000000;
    rd_cycle[10380] = 1'b1;  wr_cycle[10380] = 1'b0;  addr_rom[10380]='h000005f0;  wr_data_rom[10380]='h00000000;
    rd_cycle[10381] = 1'b1;  wr_cycle[10381] = 1'b0;  addr_rom[10381]='h000005f4;  wr_data_rom[10381]='h00000000;
    rd_cycle[10382] = 1'b1;  wr_cycle[10382] = 1'b0;  addr_rom[10382]='h000005f8;  wr_data_rom[10382]='h00000000;
    rd_cycle[10383] = 1'b1;  wr_cycle[10383] = 1'b0;  addr_rom[10383]='h000005fc;  wr_data_rom[10383]='h00000000;
    rd_cycle[10384] = 1'b1;  wr_cycle[10384] = 1'b0;  addr_rom[10384]='h00000600;  wr_data_rom[10384]='h00000000;
    rd_cycle[10385] = 1'b1;  wr_cycle[10385] = 1'b0;  addr_rom[10385]='h00000604;  wr_data_rom[10385]='h00000000;
    rd_cycle[10386] = 1'b1;  wr_cycle[10386] = 1'b0;  addr_rom[10386]='h00000608;  wr_data_rom[10386]='h00000000;
    rd_cycle[10387] = 1'b1;  wr_cycle[10387] = 1'b0;  addr_rom[10387]='h0000060c;  wr_data_rom[10387]='h00000000;
    rd_cycle[10388] = 1'b1;  wr_cycle[10388] = 1'b0;  addr_rom[10388]='h00000610;  wr_data_rom[10388]='h00000000;
    rd_cycle[10389] = 1'b1;  wr_cycle[10389] = 1'b0;  addr_rom[10389]='h00000614;  wr_data_rom[10389]='h00000000;
    rd_cycle[10390] = 1'b1;  wr_cycle[10390] = 1'b0;  addr_rom[10390]='h00000618;  wr_data_rom[10390]='h00000000;
    rd_cycle[10391] = 1'b1;  wr_cycle[10391] = 1'b0;  addr_rom[10391]='h0000061c;  wr_data_rom[10391]='h00000000;
    rd_cycle[10392] = 1'b1;  wr_cycle[10392] = 1'b0;  addr_rom[10392]='h00000620;  wr_data_rom[10392]='h00000000;
    rd_cycle[10393] = 1'b1;  wr_cycle[10393] = 1'b0;  addr_rom[10393]='h00000624;  wr_data_rom[10393]='h00000000;
    rd_cycle[10394] = 1'b1;  wr_cycle[10394] = 1'b0;  addr_rom[10394]='h00000628;  wr_data_rom[10394]='h00000000;
    rd_cycle[10395] = 1'b1;  wr_cycle[10395] = 1'b0;  addr_rom[10395]='h0000062c;  wr_data_rom[10395]='h00000000;
    rd_cycle[10396] = 1'b1;  wr_cycle[10396] = 1'b0;  addr_rom[10396]='h00000630;  wr_data_rom[10396]='h00000000;
    rd_cycle[10397] = 1'b1;  wr_cycle[10397] = 1'b0;  addr_rom[10397]='h00000634;  wr_data_rom[10397]='h00000000;
    rd_cycle[10398] = 1'b1;  wr_cycle[10398] = 1'b0;  addr_rom[10398]='h00000638;  wr_data_rom[10398]='h00000000;
    rd_cycle[10399] = 1'b1;  wr_cycle[10399] = 1'b0;  addr_rom[10399]='h0000063c;  wr_data_rom[10399]='h00000000;
    rd_cycle[10400] = 1'b1;  wr_cycle[10400] = 1'b0;  addr_rom[10400]='h00000640;  wr_data_rom[10400]='h00000000;
    rd_cycle[10401] = 1'b1;  wr_cycle[10401] = 1'b0;  addr_rom[10401]='h00000644;  wr_data_rom[10401]='h00000000;
    rd_cycle[10402] = 1'b1;  wr_cycle[10402] = 1'b0;  addr_rom[10402]='h00000648;  wr_data_rom[10402]='h00000000;
    rd_cycle[10403] = 1'b1;  wr_cycle[10403] = 1'b0;  addr_rom[10403]='h0000064c;  wr_data_rom[10403]='h00000000;
    rd_cycle[10404] = 1'b1;  wr_cycle[10404] = 1'b0;  addr_rom[10404]='h00000650;  wr_data_rom[10404]='h00000000;
    rd_cycle[10405] = 1'b1;  wr_cycle[10405] = 1'b0;  addr_rom[10405]='h00000654;  wr_data_rom[10405]='h00000000;
    rd_cycle[10406] = 1'b1;  wr_cycle[10406] = 1'b0;  addr_rom[10406]='h00000658;  wr_data_rom[10406]='h00000000;
    rd_cycle[10407] = 1'b1;  wr_cycle[10407] = 1'b0;  addr_rom[10407]='h0000065c;  wr_data_rom[10407]='h00000000;
    rd_cycle[10408] = 1'b1;  wr_cycle[10408] = 1'b0;  addr_rom[10408]='h00000660;  wr_data_rom[10408]='h00000000;
    rd_cycle[10409] = 1'b1;  wr_cycle[10409] = 1'b0;  addr_rom[10409]='h00000664;  wr_data_rom[10409]='h00000000;
    rd_cycle[10410] = 1'b1;  wr_cycle[10410] = 1'b0;  addr_rom[10410]='h00000668;  wr_data_rom[10410]='h00000000;
    rd_cycle[10411] = 1'b1;  wr_cycle[10411] = 1'b0;  addr_rom[10411]='h0000066c;  wr_data_rom[10411]='h00000000;
    rd_cycle[10412] = 1'b1;  wr_cycle[10412] = 1'b0;  addr_rom[10412]='h00000670;  wr_data_rom[10412]='h00000000;
    rd_cycle[10413] = 1'b1;  wr_cycle[10413] = 1'b0;  addr_rom[10413]='h00000674;  wr_data_rom[10413]='h00000000;
    rd_cycle[10414] = 1'b1;  wr_cycle[10414] = 1'b0;  addr_rom[10414]='h00000678;  wr_data_rom[10414]='h00000000;
    rd_cycle[10415] = 1'b1;  wr_cycle[10415] = 1'b0;  addr_rom[10415]='h0000067c;  wr_data_rom[10415]='h00000000;
    rd_cycle[10416] = 1'b1;  wr_cycle[10416] = 1'b0;  addr_rom[10416]='h00000680;  wr_data_rom[10416]='h00000000;
    rd_cycle[10417] = 1'b1;  wr_cycle[10417] = 1'b0;  addr_rom[10417]='h00000684;  wr_data_rom[10417]='h00000000;
    rd_cycle[10418] = 1'b1;  wr_cycle[10418] = 1'b0;  addr_rom[10418]='h00000688;  wr_data_rom[10418]='h00000000;
    rd_cycle[10419] = 1'b1;  wr_cycle[10419] = 1'b0;  addr_rom[10419]='h0000068c;  wr_data_rom[10419]='h00000000;
    rd_cycle[10420] = 1'b1;  wr_cycle[10420] = 1'b0;  addr_rom[10420]='h00000690;  wr_data_rom[10420]='h00000000;
    rd_cycle[10421] = 1'b1;  wr_cycle[10421] = 1'b0;  addr_rom[10421]='h00000694;  wr_data_rom[10421]='h00000000;
    rd_cycle[10422] = 1'b1;  wr_cycle[10422] = 1'b0;  addr_rom[10422]='h00000698;  wr_data_rom[10422]='h00000000;
    rd_cycle[10423] = 1'b1;  wr_cycle[10423] = 1'b0;  addr_rom[10423]='h0000069c;  wr_data_rom[10423]='h00000000;
    rd_cycle[10424] = 1'b1;  wr_cycle[10424] = 1'b0;  addr_rom[10424]='h000006a0;  wr_data_rom[10424]='h00000000;
    rd_cycle[10425] = 1'b1;  wr_cycle[10425] = 1'b0;  addr_rom[10425]='h000006a4;  wr_data_rom[10425]='h00000000;
    rd_cycle[10426] = 1'b1;  wr_cycle[10426] = 1'b0;  addr_rom[10426]='h000006a8;  wr_data_rom[10426]='h00000000;
    rd_cycle[10427] = 1'b1;  wr_cycle[10427] = 1'b0;  addr_rom[10427]='h000006ac;  wr_data_rom[10427]='h00000000;
    rd_cycle[10428] = 1'b1;  wr_cycle[10428] = 1'b0;  addr_rom[10428]='h000006b0;  wr_data_rom[10428]='h00000000;
    rd_cycle[10429] = 1'b1;  wr_cycle[10429] = 1'b0;  addr_rom[10429]='h000006b4;  wr_data_rom[10429]='h00000000;
    rd_cycle[10430] = 1'b1;  wr_cycle[10430] = 1'b0;  addr_rom[10430]='h000006b8;  wr_data_rom[10430]='h00000000;
    rd_cycle[10431] = 1'b1;  wr_cycle[10431] = 1'b0;  addr_rom[10431]='h000006bc;  wr_data_rom[10431]='h00000000;
    rd_cycle[10432] = 1'b1;  wr_cycle[10432] = 1'b0;  addr_rom[10432]='h000006c0;  wr_data_rom[10432]='h00000000;
    rd_cycle[10433] = 1'b1;  wr_cycle[10433] = 1'b0;  addr_rom[10433]='h000006c4;  wr_data_rom[10433]='h00000000;
    rd_cycle[10434] = 1'b1;  wr_cycle[10434] = 1'b0;  addr_rom[10434]='h000006c8;  wr_data_rom[10434]='h00000000;
    rd_cycle[10435] = 1'b1;  wr_cycle[10435] = 1'b0;  addr_rom[10435]='h000006cc;  wr_data_rom[10435]='h00000000;
    rd_cycle[10436] = 1'b1;  wr_cycle[10436] = 1'b0;  addr_rom[10436]='h000006d0;  wr_data_rom[10436]='h00000000;
    rd_cycle[10437] = 1'b1;  wr_cycle[10437] = 1'b0;  addr_rom[10437]='h000006d4;  wr_data_rom[10437]='h00000000;
    rd_cycle[10438] = 1'b1;  wr_cycle[10438] = 1'b0;  addr_rom[10438]='h000006d8;  wr_data_rom[10438]='h00000000;
    rd_cycle[10439] = 1'b1;  wr_cycle[10439] = 1'b0;  addr_rom[10439]='h000006dc;  wr_data_rom[10439]='h00000000;
    rd_cycle[10440] = 1'b1;  wr_cycle[10440] = 1'b0;  addr_rom[10440]='h000006e0;  wr_data_rom[10440]='h00000000;
    rd_cycle[10441] = 1'b1;  wr_cycle[10441] = 1'b0;  addr_rom[10441]='h000006e4;  wr_data_rom[10441]='h00000000;
    rd_cycle[10442] = 1'b1;  wr_cycle[10442] = 1'b0;  addr_rom[10442]='h000006e8;  wr_data_rom[10442]='h00000000;
    rd_cycle[10443] = 1'b1;  wr_cycle[10443] = 1'b0;  addr_rom[10443]='h000006ec;  wr_data_rom[10443]='h00000000;
    rd_cycle[10444] = 1'b1;  wr_cycle[10444] = 1'b0;  addr_rom[10444]='h000006f0;  wr_data_rom[10444]='h00000000;
    rd_cycle[10445] = 1'b1;  wr_cycle[10445] = 1'b0;  addr_rom[10445]='h000006f4;  wr_data_rom[10445]='h00000000;
    rd_cycle[10446] = 1'b1;  wr_cycle[10446] = 1'b0;  addr_rom[10446]='h000006f8;  wr_data_rom[10446]='h00000000;
    rd_cycle[10447] = 1'b1;  wr_cycle[10447] = 1'b0;  addr_rom[10447]='h000006fc;  wr_data_rom[10447]='h00000000;
    rd_cycle[10448] = 1'b1;  wr_cycle[10448] = 1'b0;  addr_rom[10448]='h00000700;  wr_data_rom[10448]='h00000000;
    rd_cycle[10449] = 1'b1;  wr_cycle[10449] = 1'b0;  addr_rom[10449]='h00000704;  wr_data_rom[10449]='h00000000;
    rd_cycle[10450] = 1'b1;  wr_cycle[10450] = 1'b0;  addr_rom[10450]='h00000708;  wr_data_rom[10450]='h00000000;
    rd_cycle[10451] = 1'b1;  wr_cycle[10451] = 1'b0;  addr_rom[10451]='h0000070c;  wr_data_rom[10451]='h00000000;
    rd_cycle[10452] = 1'b1;  wr_cycle[10452] = 1'b0;  addr_rom[10452]='h00000710;  wr_data_rom[10452]='h00000000;
    rd_cycle[10453] = 1'b1;  wr_cycle[10453] = 1'b0;  addr_rom[10453]='h00000714;  wr_data_rom[10453]='h00000000;
    rd_cycle[10454] = 1'b1;  wr_cycle[10454] = 1'b0;  addr_rom[10454]='h00000718;  wr_data_rom[10454]='h00000000;
    rd_cycle[10455] = 1'b1;  wr_cycle[10455] = 1'b0;  addr_rom[10455]='h0000071c;  wr_data_rom[10455]='h00000000;
    rd_cycle[10456] = 1'b1;  wr_cycle[10456] = 1'b0;  addr_rom[10456]='h00000720;  wr_data_rom[10456]='h00000000;
    rd_cycle[10457] = 1'b1;  wr_cycle[10457] = 1'b0;  addr_rom[10457]='h00000724;  wr_data_rom[10457]='h00000000;
    rd_cycle[10458] = 1'b1;  wr_cycle[10458] = 1'b0;  addr_rom[10458]='h00000728;  wr_data_rom[10458]='h00000000;
    rd_cycle[10459] = 1'b1;  wr_cycle[10459] = 1'b0;  addr_rom[10459]='h0000072c;  wr_data_rom[10459]='h00000000;
    rd_cycle[10460] = 1'b1;  wr_cycle[10460] = 1'b0;  addr_rom[10460]='h00000730;  wr_data_rom[10460]='h00000000;
    rd_cycle[10461] = 1'b1;  wr_cycle[10461] = 1'b0;  addr_rom[10461]='h00000734;  wr_data_rom[10461]='h00000000;
    rd_cycle[10462] = 1'b1;  wr_cycle[10462] = 1'b0;  addr_rom[10462]='h00000738;  wr_data_rom[10462]='h00000000;
    rd_cycle[10463] = 1'b1;  wr_cycle[10463] = 1'b0;  addr_rom[10463]='h0000073c;  wr_data_rom[10463]='h00000000;
    rd_cycle[10464] = 1'b1;  wr_cycle[10464] = 1'b0;  addr_rom[10464]='h00000740;  wr_data_rom[10464]='h00000000;
    rd_cycle[10465] = 1'b1;  wr_cycle[10465] = 1'b0;  addr_rom[10465]='h00000744;  wr_data_rom[10465]='h00000000;
    rd_cycle[10466] = 1'b1;  wr_cycle[10466] = 1'b0;  addr_rom[10466]='h00000748;  wr_data_rom[10466]='h00000000;
    rd_cycle[10467] = 1'b1;  wr_cycle[10467] = 1'b0;  addr_rom[10467]='h0000074c;  wr_data_rom[10467]='h00000000;
    rd_cycle[10468] = 1'b1;  wr_cycle[10468] = 1'b0;  addr_rom[10468]='h00000750;  wr_data_rom[10468]='h00000000;
    rd_cycle[10469] = 1'b1;  wr_cycle[10469] = 1'b0;  addr_rom[10469]='h00000754;  wr_data_rom[10469]='h00000000;
    rd_cycle[10470] = 1'b1;  wr_cycle[10470] = 1'b0;  addr_rom[10470]='h00000758;  wr_data_rom[10470]='h00000000;
    rd_cycle[10471] = 1'b1;  wr_cycle[10471] = 1'b0;  addr_rom[10471]='h0000075c;  wr_data_rom[10471]='h00000000;
    rd_cycle[10472] = 1'b1;  wr_cycle[10472] = 1'b0;  addr_rom[10472]='h00000760;  wr_data_rom[10472]='h00000000;
    rd_cycle[10473] = 1'b1;  wr_cycle[10473] = 1'b0;  addr_rom[10473]='h00000764;  wr_data_rom[10473]='h00000000;
    rd_cycle[10474] = 1'b1;  wr_cycle[10474] = 1'b0;  addr_rom[10474]='h00000768;  wr_data_rom[10474]='h00000000;
    rd_cycle[10475] = 1'b1;  wr_cycle[10475] = 1'b0;  addr_rom[10475]='h0000076c;  wr_data_rom[10475]='h00000000;
    rd_cycle[10476] = 1'b1;  wr_cycle[10476] = 1'b0;  addr_rom[10476]='h00000770;  wr_data_rom[10476]='h00000000;
    rd_cycle[10477] = 1'b1;  wr_cycle[10477] = 1'b0;  addr_rom[10477]='h00000774;  wr_data_rom[10477]='h00000000;
    rd_cycle[10478] = 1'b1;  wr_cycle[10478] = 1'b0;  addr_rom[10478]='h00000778;  wr_data_rom[10478]='h00000000;
    rd_cycle[10479] = 1'b1;  wr_cycle[10479] = 1'b0;  addr_rom[10479]='h0000077c;  wr_data_rom[10479]='h00000000;
    rd_cycle[10480] = 1'b1;  wr_cycle[10480] = 1'b0;  addr_rom[10480]='h00000780;  wr_data_rom[10480]='h00000000;
    rd_cycle[10481] = 1'b1;  wr_cycle[10481] = 1'b0;  addr_rom[10481]='h00000784;  wr_data_rom[10481]='h00000000;
    rd_cycle[10482] = 1'b1;  wr_cycle[10482] = 1'b0;  addr_rom[10482]='h00000788;  wr_data_rom[10482]='h00000000;
    rd_cycle[10483] = 1'b1;  wr_cycle[10483] = 1'b0;  addr_rom[10483]='h0000078c;  wr_data_rom[10483]='h00000000;
    rd_cycle[10484] = 1'b1;  wr_cycle[10484] = 1'b0;  addr_rom[10484]='h00000790;  wr_data_rom[10484]='h00000000;
    rd_cycle[10485] = 1'b1;  wr_cycle[10485] = 1'b0;  addr_rom[10485]='h00000794;  wr_data_rom[10485]='h00000000;
    rd_cycle[10486] = 1'b1;  wr_cycle[10486] = 1'b0;  addr_rom[10486]='h00000798;  wr_data_rom[10486]='h00000000;
    rd_cycle[10487] = 1'b1;  wr_cycle[10487] = 1'b0;  addr_rom[10487]='h0000079c;  wr_data_rom[10487]='h00000000;
    rd_cycle[10488] = 1'b1;  wr_cycle[10488] = 1'b0;  addr_rom[10488]='h000007a0;  wr_data_rom[10488]='h00000000;
    rd_cycle[10489] = 1'b1;  wr_cycle[10489] = 1'b0;  addr_rom[10489]='h000007a4;  wr_data_rom[10489]='h00000000;
    rd_cycle[10490] = 1'b1;  wr_cycle[10490] = 1'b0;  addr_rom[10490]='h000007a8;  wr_data_rom[10490]='h00000000;
    rd_cycle[10491] = 1'b1;  wr_cycle[10491] = 1'b0;  addr_rom[10491]='h000007ac;  wr_data_rom[10491]='h00000000;
    rd_cycle[10492] = 1'b1;  wr_cycle[10492] = 1'b0;  addr_rom[10492]='h000007b0;  wr_data_rom[10492]='h00000000;
    rd_cycle[10493] = 1'b1;  wr_cycle[10493] = 1'b0;  addr_rom[10493]='h000007b4;  wr_data_rom[10493]='h00000000;
    rd_cycle[10494] = 1'b1;  wr_cycle[10494] = 1'b0;  addr_rom[10494]='h000007b8;  wr_data_rom[10494]='h00000000;
    rd_cycle[10495] = 1'b1;  wr_cycle[10495] = 1'b0;  addr_rom[10495]='h000007bc;  wr_data_rom[10495]='h00000000;
    rd_cycle[10496] = 1'b1;  wr_cycle[10496] = 1'b0;  addr_rom[10496]='h000007c0;  wr_data_rom[10496]='h00000000;
    rd_cycle[10497] = 1'b1;  wr_cycle[10497] = 1'b0;  addr_rom[10497]='h000007c4;  wr_data_rom[10497]='h00000000;
    rd_cycle[10498] = 1'b1;  wr_cycle[10498] = 1'b0;  addr_rom[10498]='h000007c8;  wr_data_rom[10498]='h00000000;
    rd_cycle[10499] = 1'b1;  wr_cycle[10499] = 1'b0;  addr_rom[10499]='h000007cc;  wr_data_rom[10499]='h00000000;
    rd_cycle[10500] = 1'b1;  wr_cycle[10500] = 1'b0;  addr_rom[10500]='h000007d0;  wr_data_rom[10500]='h00000000;
    rd_cycle[10501] = 1'b1;  wr_cycle[10501] = 1'b0;  addr_rom[10501]='h000007d4;  wr_data_rom[10501]='h00000000;
    rd_cycle[10502] = 1'b1;  wr_cycle[10502] = 1'b0;  addr_rom[10502]='h000007d8;  wr_data_rom[10502]='h00000000;
    rd_cycle[10503] = 1'b1;  wr_cycle[10503] = 1'b0;  addr_rom[10503]='h000007dc;  wr_data_rom[10503]='h00000000;
    rd_cycle[10504] = 1'b1;  wr_cycle[10504] = 1'b0;  addr_rom[10504]='h000007e0;  wr_data_rom[10504]='h00000000;
    rd_cycle[10505] = 1'b1;  wr_cycle[10505] = 1'b0;  addr_rom[10505]='h000007e4;  wr_data_rom[10505]='h00000000;
    rd_cycle[10506] = 1'b1;  wr_cycle[10506] = 1'b0;  addr_rom[10506]='h000007e8;  wr_data_rom[10506]='h00000000;
    rd_cycle[10507] = 1'b1;  wr_cycle[10507] = 1'b0;  addr_rom[10507]='h000007ec;  wr_data_rom[10507]='h00000000;
    rd_cycle[10508] = 1'b1;  wr_cycle[10508] = 1'b0;  addr_rom[10508]='h000007f0;  wr_data_rom[10508]='h00000000;
    rd_cycle[10509] = 1'b1;  wr_cycle[10509] = 1'b0;  addr_rom[10509]='h000007f4;  wr_data_rom[10509]='h00000000;
    rd_cycle[10510] = 1'b1;  wr_cycle[10510] = 1'b0;  addr_rom[10510]='h000007f8;  wr_data_rom[10510]='h00000000;
    rd_cycle[10511] = 1'b1;  wr_cycle[10511] = 1'b0;  addr_rom[10511]='h000007fc;  wr_data_rom[10511]='h00000000;
    rd_cycle[10512] = 1'b1;  wr_cycle[10512] = 1'b0;  addr_rom[10512]='h00000800;  wr_data_rom[10512]='h00000000;
    rd_cycle[10513] = 1'b1;  wr_cycle[10513] = 1'b0;  addr_rom[10513]='h00000804;  wr_data_rom[10513]='h00000000;
    rd_cycle[10514] = 1'b1;  wr_cycle[10514] = 1'b0;  addr_rom[10514]='h00000808;  wr_data_rom[10514]='h00000000;
    rd_cycle[10515] = 1'b1;  wr_cycle[10515] = 1'b0;  addr_rom[10515]='h0000080c;  wr_data_rom[10515]='h00000000;
    rd_cycle[10516] = 1'b1;  wr_cycle[10516] = 1'b0;  addr_rom[10516]='h00000810;  wr_data_rom[10516]='h00000000;
    rd_cycle[10517] = 1'b1;  wr_cycle[10517] = 1'b0;  addr_rom[10517]='h00000814;  wr_data_rom[10517]='h00000000;
    rd_cycle[10518] = 1'b1;  wr_cycle[10518] = 1'b0;  addr_rom[10518]='h00000818;  wr_data_rom[10518]='h00000000;
    rd_cycle[10519] = 1'b1;  wr_cycle[10519] = 1'b0;  addr_rom[10519]='h0000081c;  wr_data_rom[10519]='h00000000;
    rd_cycle[10520] = 1'b1;  wr_cycle[10520] = 1'b0;  addr_rom[10520]='h00000820;  wr_data_rom[10520]='h00000000;
    rd_cycle[10521] = 1'b1;  wr_cycle[10521] = 1'b0;  addr_rom[10521]='h00000824;  wr_data_rom[10521]='h00000000;
    rd_cycle[10522] = 1'b1;  wr_cycle[10522] = 1'b0;  addr_rom[10522]='h00000828;  wr_data_rom[10522]='h00000000;
    rd_cycle[10523] = 1'b1;  wr_cycle[10523] = 1'b0;  addr_rom[10523]='h0000082c;  wr_data_rom[10523]='h00000000;
    rd_cycle[10524] = 1'b1;  wr_cycle[10524] = 1'b0;  addr_rom[10524]='h00000830;  wr_data_rom[10524]='h00000000;
    rd_cycle[10525] = 1'b1;  wr_cycle[10525] = 1'b0;  addr_rom[10525]='h00000834;  wr_data_rom[10525]='h00000000;
    rd_cycle[10526] = 1'b1;  wr_cycle[10526] = 1'b0;  addr_rom[10526]='h00000838;  wr_data_rom[10526]='h00000000;
    rd_cycle[10527] = 1'b1;  wr_cycle[10527] = 1'b0;  addr_rom[10527]='h0000083c;  wr_data_rom[10527]='h00000000;
    rd_cycle[10528] = 1'b1;  wr_cycle[10528] = 1'b0;  addr_rom[10528]='h00000840;  wr_data_rom[10528]='h00000000;
    rd_cycle[10529] = 1'b1;  wr_cycle[10529] = 1'b0;  addr_rom[10529]='h00000844;  wr_data_rom[10529]='h00000000;
    rd_cycle[10530] = 1'b1;  wr_cycle[10530] = 1'b0;  addr_rom[10530]='h00000848;  wr_data_rom[10530]='h00000000;
    rd_cycle[10531] = 1'b1;  wr_cycle[10531] = 1'b0;  addr_rom[10531]='h0000084c;  wr_data_rom[10531]='h00000000;
    rd_cycle[10532] = 1'b1;  wr_cycle[10532] = 1'b0;  addr_rom[10532]='h00000850;  wr_data_rom[10532]='h00000000;
    rd_cycle[10533] = 1'b1;  wr_cycle[10533] = 1'b0;  addr_rom[10533]='h00000854;  wr_data_rom[10533]='h00000000;
    rd_cycle[10534] = 1'b1;  wr_cycle[10534] = 1'b0;  addr_rom[10534]='h00000858;  wr_data_rom[10534]='h00000000;
    rd_cycle[10535] = 1'b1;  wr_cycle[10535] = 1'b0;  addr_rom[10535]='h0000085c;  wr_data_rom[10535]='h00000000;
    rd_cycle[10536] = 1'b1;  wr_cycle[10536] = 1'b0;  addr_rom[10536]='h00000860;  wr_data_rom[10536]='h00000000;
    rd_cycle[10537] = 1'b1;  wr_cycle[10537] = 1'b0;  addr_rom[10537]='h00000864;  wr_data_rom[10537]='h00000000;
    rd_cycle[10538] = 1'b1;  wr_cycle[10538] = 1'b0;  addr_rom[10538]='h00000868;  wr_data_rom[10538]='h00000000;
    rd_cycle[10539] = 1'b1;  wr_cycle[10539] = 1'b0;  addr_rom[10539]='h0000086c;  wr_data_rom[10539]='h00000000;
    rd_cycle[10540] = 1'b1;  wr_cycle[10540] = 1'b0;  addr_rom[10540]='h00000870;  wr_data_rom[10540]='h00000000;
    rd_cycle[10541] = 1'b1;  wr_cycle[10541] = 1'b0;  addr_rom[10541]='h00000874;  wr_data_rom[10541]='h00000000;
    rd_cycle[10542] = 1'b1;  wr_cycle[10542] = 1'b0;  addr_rom[10542]='h00000878;  wr_data_rom[10542]='h00000000;
    rd_cycle[10543] = 1'b1;  wr_cycle[10543] = 1'b0;  addr_rom[10543]='h0000087c;  wr_data_rom[10543]='h00000000;
    rd_cycle[10544] = 1'b1;  wr_cycle[10544] = 1'b0;  addr_rom[10544]='h00000880;  wr_data_rom[10544]='h00000000;
    rd_cycle[10545] = 1'b1;  wr_cycle[10545] = 1'b0;  addr_rom[10545]='h00000884;  wr_data_rom[10545]='h00000000;
    rd_cycle[10546] = 1'b1;  wr_cycle[10546] = 1'b0;  addr_rom[10546]='h00000888;  wr_data_rom[10546]='h00000000;
    rd_cycle[10547] = 1'b1;  wr_cycle[10547] = 1'b0;  addr_rom[10547]='h0000088c;  wr_data_rom[10547]='h00000000;
    rd_cycle[10548] = 1'b1;  wr_cycle[10548] = 1'b0;  addr_rom[10548]='h00000890;  wr_data_rom[10548]='h00000000;
    rd_cycle[10549] = 1'b1;  wr_cycle[10549] = 1'b0;  addr_rom[10549]='h00000894;  wr_data_rom[10549]='h00000000;
    rd_cycle[10550] = 1'b1;  wr_cycle[10550] = 1'b0;  addr_rom[10550]='h00000898;  wr_data_rom[10550]='h00000000;
    rd_cycle[10551] = 1'b1;  wr_cycle[10551] = 1'b0;  addr_rom[10551]='h0000089c;  wr_data_rom[10551]='h00000000;
    rd_cycle[10552] = 1'b1;  wr_cycle[10552] = 1'b0;  addr_rom[10552]='h000008a0;  wr_data_rom[10552]='h00000000;
    rd_cycle[10553] = 1'b1;  wr_cycle[10553] = 1'b0;  addr_rom[10553]='h000008a4;  wr_data_rom[10553]='h00000000;
    rd_cycle[10554] = 1'b1;  wr_cycle[10554] = 1'b0;  addr_rom[10554]='h000008a8;  wr_data_rom[10554]='h00000000;
    rd_cycle[10555] = 1'b1;  wr_cycle[10555] = 1'b0;  addr_rom[10555]='h000008ac;  wr_data_rom[10555]='h00000000;
    rd_cycle[10556] = 1'b1;  wr_cycle[10556] = 1'b0;  addr_rom[10556]='h000008b0;  wr_data_rom[10556]='h00000000;
    rd_cycle[10557] = 1'b1;  wr_cycle[10557] = 1'b0;  addr_rom[10557]='h000008b4;  wr_data_rom[10557]='h00000000;
    rd_cycle[10558] = 1'b1;  wr_cycle[10558] = 1'b0;  addr_rom[10558]='h000008b8;  wr_data_rom[10558]='h00000000;
    rd_cycle[10559] = 1'b1;  wr_cycle[10559] = 1'b0;  addr_rom[10559]='h000008bc;  wr_data_rom[10559]='h00000000;
    rd_cycle[10560] = 1'b1;  wr_cycle[10560] = 1'b0;  addr_rom[10560]='h000008c0;  wr_data_rom[10560]='h00000000;
    rd_cycle[10561] = 1'b1;  wr_cycle[10561] = 1'b0;  addr_rom[10561]='h000008c4;  wr_data_rom[10561]='h00000000;
    rd_cycle[10562] = 1'b1;  wr_cycle[10562] = 1'b0;  addr_rom[10562]='h000008c8;  wr_data_rom[10562]='h00000000;
    rd_cycle[10563] = 1'b1;  wr_cycle[10563] = 1'b0;  addr_rom[10563]='h000008cc;  wr_data_rom[10563]='h00000000;
    rd_cycle[10564] = 1'b1;  wr_cycle[10564] = 1'b0;  addr_rom[10564]='h000008d0;  wr_data_rom[10564]='h00000000;
    rd_cycle[10565] = 1'b1;  wr_cycle[10565] = 1'b0;  addr_rom[10565]='h000008d4;  wr_data_rom[10565]='h00000000;
    rd_cycle[10566] = 1'b1;  wr_cycle[10566] = 1'b0;  addr_rom[10566]='h000008d8;  wr_data_rom[10566]='h00000000;
    rd_cycle[10567] = 1'b1;  wr_cycle[10567] = 1'b0;  addr_rom[10567]='h000008dc;  wr_data_rom[10567]='h00000000;
    rd_cycle[10568] = 1'b1;  wr_cycle[10568] = 1'b0;  addr_rom[10568]='h000008e0;  wr_data_rom[10568]='h00000000;
    rd_cycle[10569] = 1'b1;  wr_cycle[10569] = 1'b0;  addr_rom[10569]='h000008e4;  wr_data_rom[10569]='h00000000;
    rd_cycle[10570] = 1'b1;  wr_cycle[10570] = 1'b0;  addr_rom[10570]='h000008e8;  wr_data_rom[10570]='h00000000;
    rd_cycle[10571] = 1'b1;  wr_cycle[10571] = 1'b0;  addr_rom[10571]='h000008ec;  wr_data_rom[10571]='h00000000;
    rd_cycle[10572] = 1'b1;  wr_cycle[10572] = 1'b0;  addr_rom[10572]='h000008f0;  wr_data_rom[10572]='h00000000;
    rd_cycle[10573] = 1'b1;  wr_cycle[10573] = 1'b0;  addr_rom[10573]='h000008f4;  wr_data_rom[10573]='h00000000;
    rd_cycle[10574] = 1'b1;  wr_cycle[10574] = 1'b0;  addr_rom[10574]='h000008f8;  wr_data_rom[10574]='h00000000;
    rd_cycle[10575] = 1'b1;  wr_cycle[10575] = 1'b0;  addr_rom[10575]='h000008fc;  wr_data_rom[10575]='h00000000;
    rd_cycle[10576] = 1'b1;  wr_cycle[10576] = 1'b0;  addr_rom[10576]='h00000900;  wr_data_rom[10576]='h00000000;
    rd_cycle[10577] = 1'b1;  wr_cycle[10577] = 1'b0;  addr_rom[10577]='h00000904;  wr_data_rom[10577]='h00000000;
    rd_cycle[10578] = 1'b1;  wr_cycle[10578] = 1'b0;  addr_rom[10578]='h00000908;  wr_data_rom[10578]='h00000000;
    rd_cycle[10579] = 1'b1;  wr_cycle[10579] = 1'b0;  addr_rom[10579]='h0000090c;  wr_data_rom[10579]='h00000000;
    rd_cycle[10580] = 1'b1;  wr_cycle[10580] = 1'b0;  addr_rom[10580]='h00000910;  wr_data_rom[10580]='h00000000;
    rd_cycle[10581] = 1'b1;  wr_cycle[10581] = 1'b0;  addr_rom[10581]='h00000914;  wr_data_rom[10581]='h00000000;
    rd_cycle[10582] = 1'b1;  wr_cycle[10582] = 1'b0;  addr_rom[10582]='h00000918;  wr_data_rom[10582]='h00000000;
    rd_cycle[10583] = 1'b1;  wr_cycle[10583] = 1'b0;  addr_rom[10583]='h0000091c;  wr_data_rom[10583]='h00000000;
    rd_cycle[10584] = 1'b1;  wr_cycle[10584] = 1'b0;  addr_rom[10584]='h00000920;  wr_data_rom[10584]='h00000000;
    rd_cycle[10585] = 1'b1;  wr_cycle[10585] = 1'b0;  addr_rom[10585]='h00000924;  wr_data_rom[10585]='h00000000;
    rd_cycle[10586] = 1'b1;  wr_cycle[10586] = 1'b0;  addr_rom[10586]='h00000928;  wr_data_rom[10586]='h00000000;
    rd_cycle[10587] = 1'b1;  wr_cycle[10587] = 1'b0;  addr_rom[10587]='h0000092c;  wr_data_rom[10587]='h00000000;
    rd_cycle[10588] = 1'b1;  wr_cycle[10588] = 1'b0;  addr_rom[10588]='h00000930;  wr_data_rom[10588]='h00000000;
    rd_cycle[10589] = 1'b1;  wr_cycle[10589] = 1'b0;  addr_rom[10589]='h00000934;  wr_data_rom[10589]='h00000000;
    rd_cycle[10590] = 1'b1;  wr_cycle[10590] = 1'b0;  addr_rom[10590]='h00000938;  wr_data_rom[10590]='h00000000;
    rd_cycle[10591] = 1'b1;  wr_cycle[10591] = 1'b0;  addr_rom[10591]='h0000093c;  wr_data_rom[10591]='h00000000;
    rd_cycle[10592] = 1'b1;  wr_cycle[10592] = 1'b0;  addr_rom[10592]='h00000940;  wr_data_rom[10592]='h00000000;
    rd_cycle[10593] = 1'b1;  wr_cycle[10593] = 1'b0;  addr_rom[10593]='h00000944;  wr_data_rom[10593]='h00000000;
    rd_cycle[10594] = 1'b1;  wr_cycle[10594] = 1'b0;  addr_rom[10594]='h00000948;  wr_data_rom[10594]='h00000000;
    rd_cycle[10595] = 1'b1;  wr_cycle[10595] = 1'b0;  addr_rom[10595]='h0000094c;  wr_data_rom[10595]='h00000000;
    rd_cycle[10596] = 1'b1;  wr_cycle[10596] = 1'b0;  addr_rom[10596]='h00000950;  wr_data_rom[10596]='h00000000;
    rd_cycle[10597] = 1'b1;  wr_cycle[10597] = 1'b0;  addr_rom[10597]='h00000954;  wr_data_rom[10597]='h00000000;
    rd_cycle[10598] = 1'b1;  wr_cycle[10598] = 1'b0;  addr_rom[10598]='h00000958;  wr_data_rom[10598]='h00000000;
    rd_cycle[10599] = 1'b1;  wr_cycle[10599] = 1'b0;  addr_rom[10599]='h0000095c;  wr_data_rom[10599]='h00000000;
    rd_cycle[10600] = 1'b1;  wr_cycle[10600] = 1'b0;  addr_rom[10600]='h00000960;  wr_data_rom[10600]='h00000000;
    rd_cycle[10601] = 1'b1;  wr_cycle[10601] = 1'b0;  addr_rom[10601]='h00000964;  wr_data_rom[10601]='h00000000;
    rd_cycle[10602] = 1'b1;  wr_cycle[10602] = 1'b0;  addr_rom[10602]='h00000968;  wr_data_rom[10602]='h00000000;
    rd_cycle[10603] = 1'b1;  wr_cycle[10603] = 1'b0;  addr_rom[10603]='h0000096c;  wr_data_rom[10603]='h00000000;
    rd_cycle[10604] = 1'b1;  wr_cycle[10604] = 1'b0;  addr_rom[10604]='h00000970;  wr_data_rom[10604]='h00000000;
    rd_cycle[10605] = 1'b1;  wr_cycle[10605] = 1'b0;  addr_rom[10605]='h00000974;  wr_data_rom[10605]='h00000000;
    rd_cycle[10606] = 1'b1;  wr_cycle[10606] = 1'b0;  addr_rom[10606]='h00000978;  wr_data_rom[10606]='h00000000;
    rd_cycle[10607] = 1'b1;  wr_cycle[10607] = 1'b0;  addr_rom[10607]='h0000097c;  wr_data_rom[10607]='h00000000;
    rd_cycle[10608] = 1'b1;  wr_cycle[10608] = 1'b0;  addr_rom[10608]='h00000980;  wr_data_rom[10608]='h00000000;
    rd_cycle[10609] = 1'b1;  wr_cycle[10609] = 1'b0;  addr_rom[10609]='h00000984;  wr_data_rom[10609]='h00000000;
    rd_cycle[10610] = 1'b1;  wr_cycle[10610] = 1'b0;  addr_rom[10610]='h00000988;  wr_data_rom[10610]='h00000000;
    rd_cycle[10611] = 1'b1;  wr_cycle[10611] = 1'b0;  addr_rom[10611]='h0000098c;  wr_data_rom[10611]='h00000000;
    rd_cycle[10612] = 1'b1;  wr_cycle[10612] = 1'b0;  addr_rom[10612]='h00000990;  wr_data_rom[10612]='h00000000;
    rd_cycle[10613] = 1'b1;  wr_cycle[10613] = 1'b0;  addr_rom[10613]='h00000994;  wr_data_rom[10613]='h00000000;
    rd_cycle[10614] = 1'b1;  wr_cycle[10614] = 1'b0;  addr_rom[10614]='h00000998;  wr_data_rom[10614]='h00000000;
    rd_cycle[10615] = 1'b1;  wr_cycle[10615] = 1'b0;  addr_rom[10615]='h0000099c;  wr_data_rom[10615]='h00000000;
    rd_cycle[10616] = 1'b1;  wr_cycle[10616] = 1'b0;  addr_rom[10616]='h000009a0;  wr_data_rom[10616]='h00000000;
    rd_cycle[10617] = 1'b1;  wr_cycle[10617] = 1'b0;  addr_rom[10617]='h000009a4;  wr_data_rom[10617]='h00000000;
    rd_cycle[10618] = 1'b1;  wr_cycle[10618] = 1'b0;  addr_rom[10618]='h000009a8;  wr_data_rom[10618]='h00000000;
    rd_cycle[10619] = 1'b1;  wr_cycle[10619] = 1'b0;  addr_rom[10619]='h000009ac;  wr_data_rom[10619]='h00000000;
    rd_cycle[10620] = 1'b1;  wr_cycle[10620] = 1'b0;  addr_rom[10620]='h000009b0;  wr_data_rom[10620]='h00000000;
    rd_cycle[10621] = 1'b1;  wr_cycle[10621] = 1'b0;  addr_rom[10621]='h000009b4;  wr_data_rom[10621]='h00000000;
    rd_cycle[10622] = 1'b1;  wr_cycle[10622] = 1'b0;  addr_rom[10622]='h000009b8;  wr_data_rom[10622]='h00000000;
    rd_cycle[10623] = 1'b1;  wr_cycle[10623] = 1'b0;  addr_rom[10623]='h000009bc;  wr_data_rom[10623]='h00000000;
    rd_cycle[10624] = 1'b1;  wr_cycle[10624] = 1'b0;  addr_rom[10624]='h000009c0;  wr_data_rom[10624]='h00000000;
    rd_cycle[10625] = 1'b1;  wr_cycle[10625] = 1'b0;  addr_rom[10625]='h000009c4;  wr_data_rom[10625]='h00000000;
    rd_cycle[10626] = 1'b1;  wr_cycle[10626] = 1'b0;  addr_rom[10626]='h000009c8;  wr_data_rom[10626]='h00000000;
    rd_cycle[10627] = 1'b1;  wr_cycle[10627] = 1'b0;  addr_rom[10627]='h000009cc;  wr_data_rom[10627]='h00000000;
    rd_cycle[10628] = 1'b1;  wr_cycle[10628] = 1'b0;  addr_rom[10628]='h000009d0;  wr_data_rom[10628]='h00000000;
    rd_cycle[10629] = 1'b1;  wr_cycle[10629] = 1'b0;  addr_rom[10629]='h000009d4;  wr_data_rom[10629]='h00000000;
    rd_cycle[10630] = 1'b1;  wr_cycle[10630] = 1'b0;  addr_rom[10630]='h000009d8;  wr_data_rom[10630]='h00000000;
    rd_cycle[10631] = 1'b1;  wr_cycle[10631] = 1'b0;  addr_rom[10631]='h000009dc;  wr_data_rom[10631]='h00000000;
    rd_cycle[10632] = 1'b1;  wr_cycle[10632] = 1'b0;  addr_rom[10632]='h000009e0;  wr_data_rom[10632]='h00000000;
    rd_cycle[10633] = 1'b1;  wr_cycle[10633] = 1'b0;  addr_rom[10633]='h000009e4;  wr_data_rom[10633]='h00000000;
    rd_cycle[10634] = 1'b1;  wr_cycle[10634] = 1'b0;  addr_rom[10634]='h000009e8;  wr_data_rom[10634]='h00000000;
    rd_cycle[10635] = 1'b1;  wr_cycle[10635] = 1'b0;  addr_rom[10635]='h000009ec;  wr_data_rom[10635]='h00000000;
    rd_cycle[10636] = 1'b1;  wr_cycle[10636] = 1'b0;  addr_rom[10636]='h000009f0;  wr_data_rom[10636]='h00000000;
    rd_cycle[10637] = 1'b1;  wr_cycle[10637] = 1'b0;  addr_rom[10637]='h000009f4;  wr_data_rom[10637]='h00000000;
    rd_cycle[10638] = 1'b1;  wr_cycle[10638] = 1'b0;  addr_rom[10638]='h000009f8;  wr_data_rom[10638]='h00000000;
    rd_cycle[10639] = 1'b1;  wr_cycle[10639] = 1'b0;  addr_rom[10639]='h000009fc;  wr_data_rom[10639]='h00000000;
    rd_cycle[10640] = 1'b1;  wr_cycle[10640] = 1'b0;  addr_rom[10640]='h00000a00;  wr_data_rom[10640]='h00000000;
    rd_cycle[10641] = 1'b1;  wr_cycle[10641] = 1'b0;  addr_rom[10641]='h00000a04;  wr_data_rom[10641]='h00000000;
    rd_cycle[10642] = 1'b1;  wr_cycle[10642] = 1'b0;  addr_rom[10642]='h00000a08;  wr_data_rom[10642]='h00000000;
    rd_cycle[10643] = 1'b1;  wr_cycle[10643] = 1'b0;  addr_rom[10643]='h00000a0c;  wr_data_rom[10643]='h00000000;
    rd_cycle[10644] = 1'b1;  wr_cycle[10644] = 1'b0;  addr_rom[10644]='h00000a10;  wr_data_rom[10644]='h00000000;
    rd_cycle[10645] = 1'b1;  wr_cycle[10645] = 1'b0;  addr_rom[10645]='h00000a14;  wr_data_rom[10645]='h00000000;
    rd_cycle[10646] = 1'b1;  wr_cycle[10646] = 1'b0;  addr_rom[10646]='h00000a18;  wr_data_rom[10646]='h00000000;
    rd_cycle[10647] = 1'b1;  wr_cycle[10647] = 1'b0;  addr_rom[10647]='h00000a1c;  wr_data_rom[10647]='h00000000;
    rd_cycle[10648] = 1'b1;  wr_cycle[10648] = 1'b0;  addr_rom[10648]='h00000a20;  wr_data_rom[10648]='h00000000;
    rd_cycle[10649] = 1'b1;  wr_cycle[10649] = 1'b0;  addr_rom[10649]='h00000a24;  wr_data_rom[10649]='h00000000;
    rd_cycle[10650] = 1'b1;  wr_cycle[10650] = 1'b0;  addr_rom[10650]='h00000a28;  wr_data_rom[10650]='h00000000;
    rd_cycle[10651] = 1'b1;  wr_cycle[10651] = 1'b0;  addr_rom[10651]='h00000a2c;  wr_data_rom[10651]='h00000000;
    rd_cycle[10652] = 1'b1;  wr_cycle[10652] = 1'b0;  addr_rom[10652]='h00000a30;  wr_data_rom[10652]='h00000000;
    rd_cycle[10653] = 1'b1;  wr_cycle[10653] = 1'b0;  addr_rom[10653]='h00000a34;  wr_data_rom[10653]='h00000000;
    rd_cycle[10654] = 1'b1;  wr_cycle[10654] = 1'b0;  addr_rom[10654]='h00000a38;  wr_data_rom[10654]='h00000000;
    rd_cycle[10655] = 1'b1;  wr_cycle[10655] = 1'b0;  addr_rom[10655]='h00000a3c;  wr_data_rom[10655]='h00000000;
    rd_cycle[10656] = 1'b1;  wr_cycle[10656] = 1'b0;  addr_rom[10656]='h00000a40;  wr_data_rom[10656]='h00000000;
    rd_cycle[10657] = 1'b1;  wr_cycle[10657] = 1'b0;  addr_rom[10657]='h00000a44;  wr_data_rom[10657]='h00000000;
    rd_cycle[10658] = 1'b1;  wr_cycle[10658] = 1'b0;  addr_rom[10658]='h00000a48;  wr_data_rom[10658]='h00000000;
    rd_cycle[10659] = 1'b1;  wr_cycle[10659] = 1'b0;  addr_rom[10659]='h00000a4c;  wr_data_rom[10659]='h00000000;
    rd_cycle[10660] = 1'b1;  wr_cycle[10660] = 1'b0;  addr_rom[10660]='h00000a50;  wr_data_rom[10660]='h00000000;
    rd_cycle[10661] = 1'b1;  wr_cycle[10661] = 1'b0;  addr_rom[10661]='h00000a54;  wr_data_rom[10661]='h00000000;
    rd_cycle[10662] = 1'b1;  wr_cycle[10662] = 1'b0;  addr_rom[10662]='h00000a58;  wr_data_rom[10662]='h00000000;
    rd_cycle[10663] = 1'b1;  wr_cycle[10663] = 1'b0;  addr_rom[10663]='h00000a5c;  wr_data_rom[10663]='h00000000;
    rd_cycle[10664] = 1'b1;  wr_cycle[10664] = 1'b0;  addr_rom[10664]='h00000a60;  wr_data_rom[10664]='h00000000;
    rd_cycle[10665] = 1'b1;  wr_cycle[10665] = 1'b0;  addr_rom[10665]='h00000a64;  wr_data_rom[10665]='h00000000;
    rd_cycle[10666] = 1'b1;  wr_cycle[10666] = 1'b0;  addr_rom[10666]='h00000a68;  wr_data_rom[10666]='h00000000;
    rd_cycle[10667] = 1'b1;  wr_cycle[10667] = 1'b0;  addr_rom[10667]='h00000a6c;  wr_data_rom[10667]='h00000000;
    rd_cycle[10668] = 1'b1;  wr_cycle[10668] = 1'b0;  addr_rom[10668]='h00000a70;  wr_data_rom[10668]='h00000000;
    rd_cycle[10669] = 1'b1;  wr_cycle[10669] = 1'b0;  addr_rom[10669]='h00000a74;  wr_data_rom[10669]='h00000000;
    rd_cycle[10670] = 1'b1;  wr_cycle[10670] = 1'b0;  addr_rom[10670]='h00000a78;  wr_data_rom[10670]='h00000000;
    rd_cycle[10671] = 1'b1;  wr_cycle[10671] = 1'b0;  addr_rom[10671]='h00000a7c;  wr_data_rom[10671]='h00000000;
    rd_cycle[10672] = 1'b1;  wr_cycle[10672] = 1'b0;  addr_rom[10672]='h00000a80;  wr_data_rom[10672]='h00000000;
    rd_cycle[10673] = 1'b1;  wr_cycle[10673] = 1'b0;  addr_rom[10673]='h00000a84;  wr_data_rom[10673]='h00000000;
    rd_cycle[10674] = 1'b1;  wr_cycle[10674] = 1'b0;  addr_rom[10674]='h00000a88;  wr_data_rom[10674]='h00000000;
    rd_cycle[10675] = 1'b1;  wr_cycle[10675] = 1'b0;  addr_rom[10675]='h00000a8c;  wr_data_rom[10675]='h00000000;
    rd_cycle[10676] = 1'b1;  wr_cycle[10676] = 1'b0;  addr_rom[10676]='h00000a90;  wr_data_rom[10676]='h00000000;
    rd_cycle[10677] = 1'b1;  wr_cycle[10677] = 1'b0;  addr_rom[10677]='h00000a94;  wr_data_rom[10677]='h00000000;
    rd_cycle[10678] = 1'b1;  wr_cycle[10678] = 1'b0;  addr_rom[10678]='h00000a98;  wr_data_rom[10678]='h00000000;
    rd_cycle[10679] = 1'b1;  wr_cycle[10679] = 1'b0;  addr_rom[10679]='h00000a9c;  wr_data_rom[10679]='h00000000;
    rd_cycle[10680] = 1'b1;  wr_cycle[10680] = 1'b0;  addr_rom[10680]='h00000aa0;  wr_data_rom[10680]='h00000000;
    rd_cycle[10681] = 1'b1;  wr_cycle[10681] = 1'b0;  addr_rom[10681]='h00000aa4;  wr_data_rom[10681]='h00000000;
    rd_cycle[10682] = 1'b1;  wr_cycle[10682] = 1'b0;  addr_rom[10682]='h00000aa8;  wr_data_rom[10682]='h00000000;
    rd_cycle[10683] = 1'b1;  wr_cycle[10683] = 1'b0;  addr_rom[10683]='h00000aac;  wr_data_rom[10683]='h00000000;
    rd_cycle[10684] = 1'b1;  wr_cycle[10684] = 1'b0;  addr_rom[10684]='h00000ab0;  wr_data_rom[10684]='h00000000;
    rd_cycle[10685] = 1'b1;  wr_cycle[10685] = 1'b0;  addr_rom[10685]='h00000ab4;  wr_data_rom[10685]='h00000000;
    rd_cycle[10686] = 1'b1;  wr_cycle[10686] = 1'b0;  addr_rom[10686]='h00000ab8;  wr_data_rom[10686]='h00000000;
    rd_cycle[10687] = 1'b1;  wr_cycle[10687] = 1'b0;  addr_rom[10687]='h00000abc;  wr_data_rom[10687]='h00000000;
    rd_cycle[10688] = 1'b1;  wr_cycle[10688] = 1'b0;  addr_rom[10688]='h00000ac0;  wr_data_rom[10688]='h00000000;
    rd_cycle[10689] = 1'b1;  wr_cycle[10689] = 1'b0;  addr_rom[10689]='h00000ac4;  wr_data_rom[10689]='h00000000;
    rd_cycle[10690] = 1'b1;  wr_cycle[10690] = 1'b0;  addr_rom[10690]='h00000ac8;  wr_data_rom[10690]='h00000000;
    rd_cycle[10691] = 1'b1;  wr_cycle[10691] = 1'b0;  addr_rom[10691]='h00000acc;  wr_data_rom[10691]='h00000000;
    rd_cycle[10692] = 1'b1;  wr_cycle[10692] = 1'b0;  addr_rom[10692]='h00000ad0;  wr_data_rom[10692]='h00000000;
    rd_cycle[10693] = 1'b1;  wr_cycle[10693] = 1'b0;  addr_rom[10693]='h00000ad4;  wr_data_rom[10693]='h00000000;
    rd_cycle[10694] = 1'b1;  wr_cycle[10694] = 1'b0;  addr_rom[10694]='h00000ad8;  wr_data_rom[10694]='h00000000;
    rd_cycle[10695] = 1'b1;  wr_cycle[10695] = 1'b0;  addr_rom[10695]='h00000adc;  wr_data_rom[10695]='h00000000;
    rd_cycle[10696] = 1'b1;  wr_cycle[10696] = 1'b0;  addr_rom[10696]='h00000ae0;  wr_data_rom[10696]='h00000000;
    rd_cycle[10697] = 1'b1;  wr_cycle[10697] = 1'b0;  addr_rom[10697]='h00000ae4;  wr_data_rom[10697]='h00000000;
    rd_cycle[10698] = 1'b1;  wr_cycle[10698] = 1'b0;  addr_rom[10698]='h00000ae8;  wr_data_rom[10698]='h00000000;
    rd_cycle[10699] = 1'b1;  wr_cycle[10699] = 1'b0;  addr_rom[10699]='h00000aec;  wr_data_rom[10699]='h00000000;
    rd_cycle[10700] = 1'b1;  wr_cycle[10700] = 1'b0;  addr_rom[10700]='h00000af0;  wr_data_rom[10700]='h00000000;
    rd_cycle[10701] = 1'b1;  wr_cycle[10701] = 1'b0;  addr_rom[10701]='h00000af4;  wr_data_rom[10701]='h00000000;
    rd_cycle[10702] = 1'b1;  wr_cycle[10702] = 1'b0;  addr_rom[10702]='h00000af8;  wr_data_rom[10702]='h00000000;
    rd_cycle[10703] = 1'b1;  wr_cycle[10703] = 1'b0;  addr_rom[10703]='h00000afc;  wr_data_rom[10703]='h00000000;
    rd_cycle[10704] = 1'b1;  wr_cycle[10704] = 1'b0;  addr_rom[10704]='h00000b00;  wr_data_rom[10704]='h00000000;
    rd_cycle[10705] = 1'b1;  wr_cycle[10705] = 1'b0;  addr_rom[10705]='h00000b04;  wr_data_rom[10705]='h00000000;
    rd_cycle[10706] = 1'b1;  wr_cycle[10706] = 1'b0;  addr_rom[10706]='h00000b08;  wr_data_rom[10706]='h00000000;
    rd_cycle[10707] = 1'b1;  wr_cycle[10707] = 1'b0;  addr_rom[10707]='h00000b0c;  wr_data_rom[10707]='h00000000;
    rd_cycle[10708] = 1'b1;  wr_cycle[10708] = 1'b0;  addr_rom[10708]='h00000b10;  wr_data_rom[10708]='h00000000;
    rd_cycle[10709] = 1'b1;  wr_cycle[10709] = 1'b0;  addr_rom[10709]='h00000b14;  wr_data_rom[10709]='h00000000;
    rd_cycle[10710] = 1'b1;  wr_cycle[10710] = 1'b0;  addr_rom[10710]='h00000b18;  wr_data_rom[10710]='h00000000;
    rd_cycle[10711] = 1'b1;  wr_cycle[10711] = 1'b0;  addr_rom[10711]='h00000b1c;  wr_data_rom[10711]='h00000000;
    rd_cycle[10712] = 1'b1;  wr_cycle[10712] = 1'b0;  addr_rom[10712]='h00000b20;  wr_data_rom[10712]='h00000000;
    rd_cycle[10713] = 1'b1;  wr_cycle[10713] = 1'b0;  addr_rom[10713]='h00000b24;  wr_data_rom[10713]='h00000000;
    rd_cycle[10714] = 1'b1;  wr_cycle[10714] = 1'b0;  addr_rom[10714]='h00000b28;  wr_data_rom[10714]='h00000000;
    rd_cycle[10715] = 1'b1;  wr_cycle[10715] = 1'b0;  addr_rom[10715]='h00000b2c;  wr_data_rom[10715]='h00000000;
    rd_cycle[10716] = 1'b1;  wr_cycle[10716] = 1'b0;  addr_rom[10716]='h00000b30;  wr_data_rom[10716]='h00000000;
    rd_cycle[10717] = 1'b1;  wr_cycle[10717] = 1'b0;  addr_rom[10717]='h00000b34;  wr_data_rom[10717]='h00000000;
    rd_cycle[10718] = 1'b1;  wr_cycle[10718] = 1'b0;  addr_rom[10718]='h00000b38;  wr_data_rom[10718]='h00000000;
    rd_cycle[10719] = 1'b1;  wr_cycle[10719] = 1'b0;  addr_rom[10719]='h00000b3c;  wr_data_rom[10719]='h00000000;
    rd_cycle[10720] = 1'b1;  wr_cycle[10720] = 1'b0;  addr_rom[10720]='h00000b40;  wr_data_rom[10720]='h00000000;
    rd_cycle[10721] = 1'b1;  wr_cycle[10721] = 1'b0;  addr_rom[10721]='h00000b44;  wr_data_rom[10721]='h00000000;
    rd_cycle[10722] = 1'b1;  wr_cycle[10722] = 1'b0;  addr_rom[10722]='h00000b48;  wr_data_rom[10722]='h00000000;
    rd_cycle[10723] = 1'b1;  wr_cycle[10723] = 1'b0;  addr_rom[10723]='h00000b4c;  wr_data_rom[10723]='h00000000;
    rd_cycle[10724] = 1'b1;  wr_cycle[10724] = 1'b0;  addr_rom[10724]='h00000b50;  wr_data_rom[10724]='h00000000;
    rd_cycle[10725] = 1'b1;  wr_cycle[10725] = 1'b0;  addr_rom[10725]='h00000b54;  wr_data_rom[10725]='h00000000;
    rd_cycle[10726] = 1'b1;  wr_cycle[10726] = 1'b0;  addr_rom[10726]='h00000b58;  wr_data_rom[10726]='h00000000;
    rd_cycle[10727] = 1'b1;  wr_cycle[10727] = 1'b0;  addr_rom[10727]='h00000b5c;  wr_data_rom[10727]='h00000000;
    rd_cycle[10728] = 1'b1;  wr_cycle[10728] = 1'b0;  addr_rom[10728]='h00000b60;  wr_data_rom[10728]='h00000000;
    rd_cycle[10729] = 1'b1;  wr_cycle[10729] = 1'b0;  addr_rom[10729]='h00000b64;  wr_data_rom[10729]='h00000000;
    rd_cycle[10730] = 1'b1;  wr_cycle[10730] = 1'b0;  addr_rom[10730]='h00000b68;  wr_data_rom[10730]='h00000000;
    rd_cycle[10731] = 1'b1;  wr_cycle[10731] = 1'b0;  addr_rom[10731]='h00000b6c;  wr_data_rom[10731]='h00000000;
    rd_cycle[10732] = 1'b1;  wr_cycle[10732] = 1'b0;  addr_rom[10732]='h00000b70;  wr_data_rom[10732]='h00000000;
    rd_cycle[10733] = 1'b1;  wr_cycle[10733] = 1'b0;  addr_rom[10733]='h00000b74;  wr_data_rom[10733]='h00000000;
    rd_cycle[10734] = 1'b1;  wr_cycle[10734] = 1'b0;  addr_rom[10734]='h00000b78;  wr_data_rom[10734]='h00000000;
    rd_cycle[10735] = 1'b1;  wr_cycle[10735] = 1'b0;  addr_rom[10735]='h00000b7c;  wr_data_rom[10735]='h00000000;
    rd_cycle[10736] = 1'b1;  wr_cycle[10736] = 1'b0;  addr_rom[10736]='h00000b80;  wr_data_rom[10736]='h00000000;
    rd_cycle[10737] = 1'b1;  wr_cycle[10737] = 1'b0;  addr_rom[10737]='h00000b84;  wr_data_rom[10737]='h00000000;
    rd_cycle[10738] = 1'b1;  wr_cycle[10738] = 1'b0;  addr_rom[10738]='h00000b88;  wr_data_rom[10738]='h00000000;
    rd_cycle[10739] = 1'b1;  wr_cycle[10739] = 1'b0;  addr_rom[10739]='h00000b8c;  wr_data_rom[10739]='h00000000;
    rd_cycle[10740] = 1'b1;  wr_cycle[10740] = 1'b0;  addr_rom[10740]='h00000b90;  wr_data_rom[10740]='h00000000;
    rd_cycle[10741] = 1'b1;  wr_cycle[10741] = 1'b0;  addr_rom[10741]='h00000b94;  wr_data_rom[10741]='h00000000;
    rd_cycle[10742] = 1'b1;  wr_cycle[10742] = 1'b0;  addr_rom[10742]='h00000b98;  wr_data_rom[10742]='h00000000;
    rd_cycle[10743] = 1'b1;  wr_cycle[10743] = 1'b0;  addr_rom[10743]='h00000b9c;  wr_data_rom[10743]='h00000000;
    rd_cycle[10744] = 1'b1;  wr_cycle[10744] = 1'b0;  addr_rom[10744]='h00000ba0;  wr_data_rom[10744]='h00000000;
    rd_cycle[10745] = 1'b1;  wr_cycle[10745] = 1'b0;  addr_rom[10745]='h00000ba4;  wr_data_rom[10745]='h00000000;
    rd_cycle[10746] = 1'b1;  wr_cycle[10746] = 1'b0;  addr_rom[10746]='h00000ba8;  wr_data_rom[10746]='h00000000;
    rd_cycle[10747] = 1'b1;  wr_cycle[10747] = 1'b0;  addr_rom[10747]='h00000bac;  wr_data_rom[10747]='h00000000;
    rd_cycle[10748] = 1'b1;  wr_cycle[10748] = 1'b0;  addr_rom[10748]='h00000bb0;  wr_data_rom[10748]='h00000000;
    rd_cycle[10749] = 1'b1;  wr_cycle[10749] = 1'b0;  addr_rom[10749]='h00000bb4;  wr_data_rom[10749]='h00000000;
    rd_cycle[10750] = 1'b1;  wr_cycle[10750] = 1'b0;  addr_rom[10750]='h00000bb8;  wr_data_rom[10750]='h00000000;
    rd_cycle[10751] = 1'b1;  wr_cycle[10751] = 1'b0;  addr_rom[10751]='h00000bbc;  wr_data_rom[10751]='h00000000;
    rd_cycle[10752] = 1'b1;  wr_cycle[10752] = 1'b0;  addr_rom[10752]='h00000bc0;  wr_data_rom[10752]='h00000000;
    rd_cycle[10753] = 1'b1;  wr_cycle[10753] = 1'b0;  addr_rom[10753]='h00000bc4;  wr_data_rom[10753]='h00000000;
    rd_cycle[10754] = 1'b1;  wr_cycle[10754] = 1'b0;  addr_rom[10754]='h00000bc8;  wr_data_rom[10754]='h00000000;
    rd_cycle[10755] = 1'b1;  wr_cycle[10755] = 1'b0;  addr_rom[10755]='h00000bcc;  wr_data_rom[10755]='h00000000;
    rd_cycle[10756] = 1'b1;  wr_cycle[10756] = 1'b0;  addr_rom[10756]='h00000bd0;  wr_data_rom[10756]='h00000000;
    rd_cycle[10757] = 1'b1;  wr_cycle[10757] = 1'b0;  addr_rom[10757]='h00000bd4;  wr_data_rom[10757]='h00000000;
    rd_cycle[10758] = 1'b1;  wr_cycle[10758] = 1'b0;  addr_rom[10758]='h00000bd8;  wr_data_rom[10758]='h00000000;
    rd_cycle[10759] = 1'b1;  wr_cycle[10759] = 1'b0;  addr_rom[10759]='h00000bdc;  wr_data_rom[10759]='h00000000;
    rd_cycle[10760] = 1'b1;  wr_cycle[10760] = 1'b0;  addr_rom[10760]='h00000be0;  wr_data_rom[10760]='h00000000;
    rd_cycle[10761] = 1'b1;  wr_cycle[10761] = 1'b0;  addr_rom[10761]='h00000be4;  wr_data_rom[10761]='h00000000;
    rd_cycle[10762] = 1'b1;  wr_cycle[10762] = 1'b0;  addr_rom[10762]='h00000be8;  wr_data_rom[10762]='h00000000;
    rd_cycle[10763] = 1'b1;  wr_cycle[10763] = 1'b0;  addr_rom[10763]='h00000bec;  wr_data_rom[10763]='h00000000;
    rd_cycle[10764] = 1'b1;  wr_cycle[10764] = 1'b0;  addr_rom[10764]='h00000bf0;  wr_data_rom[10764]='h00000000;
    rd_cycle[10765] = 1'b1;  wr_cycle[10765] = 1'b0;  addr_rom[10765]='h00000bf4;  wr_data_rom[10765]='h00000000;
    rd_cycle[10766] = 1'b1;  wr_cycle[10766] = 1'b0;  addr_rom[10766]='h00000bf8;  wr_data_rom[10766]='h00000000;
    rd_cycle[10767] = 1'b1;  wr_cycle[10767] = 1'b0;  addr_rom[10767]='h00000bfc;  wr_data_rom[10767]='h00000000;
    rd_cycle[10768] = 1'b1;  wr_cycle[10768] = 1'b0;  addr_rom[10768]='h00000c00;  wr_data_rom[10768]='h00000000;
    rd_cycle[10769] = 1'b1;  wr_cycle[10769] = 1'b0;  addr_rom[10769]='h00000c04;  wr_data_rom[10769]='h00000000;
    rd_cycle[10770] = 1'b1;  wr_cycle[10770] = 1'b0;  addr_rom[10770]='h00000c08;  wr_data_rom[10770]='h00000000;
    rd_cycle[10771] = 1'b1;  wr_cycle[10771] = 1'b0;  addr_rom[10771]='h00000c0c;  wr_data_rom[10771]='h00000000;
    rd_cycle[10772] = 1'b1;  wr_cycle[10772] = 1'b0;  addr_rom[10772]='h00000c10;  wr_data_rom[10772]='h00000000;
    rd_cycle[10773] = 1'b1;  wr_cycle[10773] = 1'b0;  addr_rom[10773]='h00000c14;  wr_data_rom[10773]='h00000000;
    rd_cycle[10774] = 1'b1;  wr_cycle[10774] = 1'b0;  addr_rom[10774]='h00000c18;  wr_data_rom[10774]='h00000000;
    rd_cycle[10775] = 1'b1;  wr_cycle[10775] = 1'b0;  addr_rom[10775]='h00000c1c;  wr_data_rom[10775]='h00000000;
    rd_cycle[10776] = 1'b1;  wr_cycle[10776] = 1'b0;  addr_rom[10776]='h00000c20;  wr_data_rom[10776]='h00000000;
    rd_cycle[10777] = 1'b1;  wr_cycle[10777] = 1'b0;  addr_rom[10777]='h00000c24;  wr_data_rom[10777]='h00000000;
    rd_cycle[10778] = 1'b1;  wr_cycle[10778] = 1'b0;  addr_rom[10778]='h00000c28;  wr_data_rom[10778]='h00000000;
    rd_cycle[10779] = 1'b1;  wr_cycle[10779] = 1'b0;  addr_rom[10779]='h00000c2c;  wr_data_rom[10779]='h00000000;
    rd_cycle[10780] = 1'b1;  wr_cycle[10780] = 1'b0;  addr_rom[10780]='h00000c30;  wr_data_rom[10780]='h00000000;
    rd_cycle[10781] = 1'b1;  wr_cycle[10781] = 1'b0;  addr_rom[10781]='h00000c34;  wr_data_rom[10781]='h00000000;
    rd_cycle[10782] = 1'b1;  wr_cycle[10782] = 1'b0;  addr_rom[10782]='h00000c38;  wr_data_rom[10782]='h00000000;
    rd_cycle[10783] = 1'b1;  wr_cycle[10783] = 1'b0;  addr_rom[10783]='h00000c3c;  wr_data_rom[10783]='h00000000;
    rd_cycle[10784] = 1'b1;  wr_cycle[10784] = 1'b0;  addr_rom[10784]='h00000c40;  wr_data_rom[10784]='h00000000;
    rd_cycle[10785] = 1'b1;  wr_cycle[10785] = 1'b0;  addr_rom[10785]='h00000c44;  wr_data_rom[10785]='h00000000;
    rd_cycle[10786] = 1'b1;  wr_cycle[10786] = 1'b0;  addr_rom[10786]='h00000c48;  wr_data_rom[10786]='h00000000;
    rd_cycle[10787] = 1'b1;  wr_cycle[10787] = 1'b0;  addr_rom[10787]='h00000c4c;  wr_data_rom[10787]='h00000000;
    rd_cycle[10788] = 1'b1;  wr_cycle[10788] = 1'b0;  addr_rom[10788]='h00000c50;  wr_data_rom[10788]='h00000000;
    rd_cycle[10789] = 1'b1;  wr_cycle[10789] = 1'b0;  addr_rom[10789]='h00000c54;  wr_data_rom[10789]='h00000000;
    rd_cycle[10790] = 1'b1;  wr_cycle[10790] = 1'b0;  addr_rom[10790]='h00000c58;  wr_data_rom[10790]='h00000000;
    rd_cycle[10791] = 1'b1;  wr_cycle[10791] = 1'b0;  addr_rom[10791]='h00000c5c;  wr_data_rom[10791]='h00000000;
    rd_cycle[10792] = 1'b1;  wr_cycle[10792] = 1'b0;  addr_rom[10792]='h00000c60;  wr_data_rom[10792]='h00000000;
    rd_cycle[10793] = 1'b1;  wr_cycle[10793] = 1'b0;  addr_rom[10793]='h00000c64;  wr_data_rom[10793]='h00000000;
    rd_cycle[10794] = 1'b1;  wr_cycle[10794] = 1'b0;  addr_rom[10794]='h00000c68;  wr_data_rom[10794]='h00000000;
    rd_cycle[10795] = 1'b1;  wr_cycle[10795] = 1'b0;  addr_rom[10795]='h00000c6c;  wr_data_rom[10795]='h00000000;
    rd_cycle[10796] = 1'b1;  wr_cycle[10796] = 1'b0;  addr_rom[10796]='h00000c70;  wr_data_rom[10796]='h00000000;
    rd_cycle[10797] = 1'b1;  wr_cycle[10797] = 1'b0;  addr_rom[10797]='h00000c74;  wr_data_rom[10797]='h00000000;
    rd_cycle[10798] = 1'b1;  wr_cycle[10798] = 1'b0;  addr_rom[10798]='h00000c78;  wr_data_rom[10798]='h00000000;
    rd_cycle[10799] = 1'b1;  wr_cycle[10799] = 1'b0;  addr_rom[10799]='h00000c7c;  wr_data_rom[10799]='h00000000;
    rd_cycle[10800] = 1'b1;  wr_cycle[10800] = 1'b0;  addr_rom[10800]='h00000c80;  wr_data_rom[10800]='h00000000;
    rd_cycle[10801] = 1'b1;  wr_cycle[10801] = 1'b0;  addr_rom[10801]='h00000c84;  wr_data_rom[10801]='h00000000;
    rd_cycle[10802] = 1'b1;  wr_cycle[10802] = 1'b0;  addr_rom[10802]='h00000c88;  wr_data_rom[10802]='h00000000;
    rd_cycle[10803] = 1'b1;  wr_cycle[10803] = 1'b0;  addr_rom[10803]='h00000c8c;  wr_data_rom[10803]='h00000000;
    rd_cycle[10804] = 1'b1;  wr_cycle[10804] = 1'b0;  addr_rom[10804]='h00000c90;  wr_data_rom[10804]='h00000000;
    rd_cycle[10805] = 1'b1;  wr_cycle[10805] = 1'b0;  addr_rom[10805]='h00000c94;  wr_data_rom[10805]='h00000000;
    rd_cycle[10806] = 1'b1;  wr_cycle[10806] = 1'b0;  addr_rom[10806]='h00000c98;  wr_data_rom[10806]='h00000000;
    rd_cycle[10807] = 1'b1;  wr_cycle[10807] = 1'b0;  addr_rom[10807]='h00000c9c;  wr_data_rom[10807]='h00000000;
    rd_cycle[10808] = 1'b1;  wr_cycle[10808] = 1'b0;  addr_rom[10808]='h00000ca0;  wr_data_rom[10808]='h00000000;
    rd_cycle[10809] = 1'b1;  wr_cycle[10809] = 1'b0;  addr_rom[10809]='h00000ca4;  wr_data_rom[10809]='h00000000;
    rd_cycle[10810] = 1'b1;  wr_cycle[10810] = 1'b0;  addr_rom[10810]='h00000ca8;  wr_data_rom[10810]='h00000000;
    rd_cycle[10811] = 1'b1;  wr_cycle[10811] = 1'b0;  addr_rom[10811]='h00000cac;  wr_data_rom[10811]='h00000000;
    rd_cycle[10812] = 1'b1;  wr_cycle[10812] = 1'b0;  addr_rom[10812]='h00000cb0;  wr_data_rom[10812]='h00000000;
    rd_cycle[10813] = 1'b1;  wr_cycle[10813] = 1'b0;  addr_rom[10813]='h00000cb4;  wr_data_rom[10813]='h00000000;
    rd_cycle[10814] = 1'b1;  wr_cycle[10814] = 1'b0;  addr_rom[10814]='h00000cb8;  wr_data_rom[10814]='h00000000;
    rd_cycle[10815] = 1'b1;  wr_cycle[10815] = 1'b0;  addr_rom[10815]='h00000cbc;  wr_data_rom[10815]='h00000000;
    rd_cycle[10816] = 1'b1;  wr_cycle[10816] = 1'b0;  addr_rom[10816]='h00000cc0;  wr_data_rom[10816]='h00000000;
    rd_cycle[10817] = 1'b1;  wr_cycle[10817] = 1'b0;  addr_rom[10817]='h00000cc4;  wr_data_rom[10817]='h00000000;
    rd_cycle[10818] = 1'b1;  wr_cycle[10818] = 1'b0;  addr_rom[10818]='h00000cc8;  wr_data_rom[10818]='h00000000;
    rd_cycle[10819] = 1'b1;  wr_cycle[10819] = 1'b0;  addr_rom[10819]='h00000ccc;  wr_data_rom[10819]='h00000000;
    rd_cycle[10820] = 1'b1;  wr_cycle[10820] = 1'b0;  addr_rom[10820]='h00000cd0;  wr_data_rom[10820]='h00000000;
    rd_cycle[10821] = 1'b1;  wr_cycle[10821] = 1'b0;  addr_rom[10821]='h00000cd4;  wr_data_rom[10821]='h00000000;
    rd_cycle[10822] = 1'b1;  wr_cycle[10822] = 1'b0;  addr_rom[10822]='h00000cd8;  wr_data_rom[10822]='h00000000;
    rd_cycle[10823] = 1'b1;  wr_cycle[10823] = 1'b0;  addr_rom[10823]='h00000cdc;  wr_data_rom[10823]='h00000000;
    rd_cycle[10824] = 1'b1;  wr_cycle[10824] = 1'b0;  addr_rom[10824]='h00000ce0;  wr_data_rom[10824]='h00000000;
    rd_cycle[10825] = 1'b1;  wr_cycle[10825] = 1'b0;  addr_rom[10825]='h00000ce4;  wr_data_rom[10825]='h00000000;
    rd_cycle[10826] = 1'b1;  wr_cycle[10826] = 1'b0;  addr_rom[10826]='h00000ce8;  wr_data_rom[10826]='h00000000;
    rd_cycle[10827] = 1'b1;  wr_cycle[10827] = 1'b0;  addr_rom[10827]='h00000cec;  wr_data_rom[10827]='h00000000;
    rd_cycle[10828] = 1'b1;  wr_cycle[10828] = 1'b0;  addr_rom[10828]='h00000cf0;  wr_data_rom[10828]='h00000000;
    rd_cycle[10829] = 1'b1;  wr_cycle[10829] = 1'b0;  addr_rom[10829]='h00000cf4;  wr_data_rom[10829]='h00000000;
    rd_cycle[10830] = 1'b1;  wr_cycle[10830] = 1'b0;  addr_rom[10830]='h00000cf8;  wr_data_rom[10830]='h00000000;
    rd_cycle[10831] = 1'b1;  wr_cycle[10831] = 1'b0;  addr_rom[10831]='h00000cfc;  wr_data_rom[10831]='h00000000;
    rd_cycle[10832] = 1'b1;  wr_cycle[10832] = 1'b0;  addr_rom[10832]='h00000d00;  wr_data_rom[10832]='h00000000;
    rd_cycle[10833] = 1'b1;  wr_cycle[10833] = 1'b0;  addr_rom[10833]='h00000d04;  wr_data_rom[10833]='h00000000;
    rd_cycle[10834] = 1'b1;  wr_cycle[10834] = 1'b0;  addr_rom[10834]='h00000d08;  wr_data_rom[10834]='h00000000;
    rd_cycle[10835] = 1'b1;  wr_cycle[10835] = 1'b0;  addr_rom[10835]='h00000d0c;  wr_data_rom[10835]='h00000000;
    rd_cycle[10836] = 1'b1;  wr_cycle[10836] = 1'b0;  addr_rom[10836]='h00000d10;  wr_data_rom[10836]='h00000000;
    rd_cycle[10837] = 1'b1;  wr_cycle[10837] = 1'b0;  addr_rom[10837]='h00000d14;  wr_data_rom[10837]='h00000000;
    rd_cycle[10838] = 1'b1;  wr_cycle[10838] = 1'b0;  addr_rom[10838]='h00000d18;  wr_data_rom[10838]='h00000000;
    rd_cycle[10839] = 1'b1;  wr_cycle[10839] = 1'b0;  addr_rom[10839]='h00000d1c;  wr_data_rom[10839]='h00000000;
    rd_cycle[10840] = 1'b1;  wr_cycle[10840] = 1'b0;  addr_rom[10840]='h00000d20;  wr_data_rom[10840]='h00000000;
    rd_cycle[10841] = 1'b1;  wr_cycle[10841] = 1'b0;  addr_rom[10841]='h00000d24;  wr_data_rom[10841]='h00000000;
    rd_cycle[10842] = 1'b1;  wr_cycle[10842] = 1'b0;  addr_rom[10842]='h00000d28;  wr_data_rom[10842]='h00000000;
    rd_cycle[10843] = 1'b1;  wr_cycle[10843] = 1'b0;  addr_rom[10843]='h00000d2c;  wr_data_rom[10843]='h00000000;
    rd_cycle[10844] = 1'b1;  wr_cycle[10844] = 1'b0;  addr_rom[10844]='h00000d30;  wr_data_rom[10844]='h00000000;
    rd_cycle[10845] = 1'b1;  wr_cycle[10845] = 1'b0;  addr_rom[10845]='h00000d34;  wr_data_rom[10845]='h00000000;
    rd_cycle[10846] = 1'b1;  wr_cycle[10846] = 1'b0;  addr_rom[10846]='h00000d38;  wr_data_rom[10846]='h00000000;
    rd_cycle[10847] = 1'b1;  wr_cycle[10847] = 1'b0;  addr_rom[10847]='h00000d3c;  wr_data_rom[10847]='h00000000;
    rd_cycle[10848] = 1'b1;  wr_cycle[10848] = 1'b0;  addr_rom[10848]='h00000d40;  wr_data_rom[10848]='h00000000;
    rd_cycle[10849] = 1'b1;  wr_cycle[10849] = 1'b0;  addr_rom[10849]='h00000d44;  wr_data_rom[10849]='h00000000;
    rd_cycle[10850] = 1'b1;  wr_cycle[10850] = 1'b0;  addr_rom[10850]='h00000d48;  wr_data_rom[10850]='h00000000;
    rd_cycle[10851] = 1'b1;  wr_cycle[10851] = 1'b0;  addr_rom[10851]='h00000d4c;  wr_data_rom[10851]='h00000000;
    rd_cycle[10852] = 1'b1;  wr_cycle[10852] = 1'b0;  addr_rom[10852]='h00000d50;  wr_data_rom[10852]='h00000000;
    rd_cycle[10853] = 1'b1;  wr_cycle[10853] = 1'b0;  addr_rom[10853]='h00000d54;  wr_data_rom[10853]='h00000000;
    rd_cycle[10854] = 1'b1;  wr_cycle[10854] = 1'b0;  addr_rom[10854]='h00000d58;  wr_data_rom[10854]='h00000000;
    rd_cycle[10855] = 1'b1;  wr_cycle[10855] = 1'b0;  addr_rom[10855]='h00000d5c;  wr_data_rom[10855]='h00000000;
    rd_cycle[10856] = 1'b1;  wr_cycle[10856] = 1'b0;  addr_rom[10856]='h00000d60;  wr_data_rom[10856]='h00000000;
    rd_cycle[10857] = 1'b1;  wr_cycle[10857] = 1'b0;  addr_rom[10857]='h00000d64;  wr_data_rom[10857]='h00000000;
    rd_cycle[10858] = 1'b1;  wr_cycle[10858] = 1'b0;  addr_rom[10858]='h00000d68;  wr_data_rom[10858]='h00000000;
    rd_cycle[10859] = 1'b1;  wr_cycle[10859] = 1'b0;  addr_rom[10859]='h00000d6c;  wr_data_rom[10859]='h00000000;
    rd_cycle[10860] = 1'b1;  wr_cycle[10860] = 1'b0;  addr_rom[10860]='h00000d70;  wr_data_rom[10860]='h00000000;
    rd_cycle[10861] = 1'b1;  wr_cycle[10861] = 1'b0;  addr_rom[10861]='h00000d74;  wr_data_rom[10861]='h00000000;
    rd_cycle[10862] = 1'b1;  wr_cycle[10862] = 1'b0;  addr_rom[10862]='h00000d78;  wr_data_rom[10862]='h00000000;
    rd_cycle[10863] = 1'b1;  wr_cycle[10863] = 1'b0;  addr_rom[10863]='h00000d7c;  wr_data_rom[10863]='h00000000;
    rd_cycle[10864] = 1'b1;  wr_cycle[10864] = 1'b0;  addr_rom[10864]='h00000d80;  wr_data_rom[10864]='h00000000;
    rd_cycle[10865] = 1'b1;  wr_cycle[10865] = 1'b0;  addr_rom[10865]='h00000d84;  wr_data_rom[10865]='h00000000;
    rd_cycle[10866] = 1'b1;  wr_cycle[10866] = 1'b0;  addr_rom[10866]='h00000d88;  wr_data_rom[10866]='h00000000;
    rd_cycle[10867] = 1'b1;  wr_cycle[10867] = 1'b0;  addr_rom[10867]='h00000d8c;  wr_data_rom[10867]='h00000000;
    rd_cycle[10868] = 1'b1;  wr_cycle[10868] = 1'b0;  addr_rom[10868]='h00000d90;  wr_data_rom[10868]='h00000000;
    rd_cycle[10869] = 1'b1;  wr_cycle[10869] = 1'b0;  addr_rom[10869]='h00000d94;  wr_data_rom[10869]='h00000000;
    rd_cycle[10870] = 1'b1;  wr_cycle[10870] = 1'b0;  addr_rom[10870]='h00000d98;  wr_data_rom[10870]='h00000000;
    rd_cycle[10871] = 1'b1;  wr_cycle[10871] = 1'b0;  addr_rom[10871]='h00000d9c;  wr_data_rom[10871]='h00000000;
    rd_cycle[10872] = 1'b1;  wr_cycle[10872] = 1'b0;  addr_rom[10872]='h00000da0;  wr_data_rom[10872]='h00000000;
    rd_cycle[10873] = 1'b1;  wr_cycle[10873] = 1'b0;  addr_rom[10873]='h00000da4;  wr_data_rom[10873]='h00000000;
    rd_cycle[10874] = 1'b1;  wr_cycle[10874] = 1'b0;  addr_rom[10874]='h00000da8;  wr_data_rom[10874]='h00000000;
    rd_cycle[10875] = 1'b1;  wr_cycle[10875] = 1'b0;  addr_rom[10875]='h00000dac;  wr_data_rom[10875]='h00000000;
    rd_cycle[10876] = 1'b1;  wr_cycle[10876] = 1'b0;  addr_rom[10876]='h00000db0;  wr_data_rom[10876]='h00000000;
    rd_cycle[10877] = 1'b1;  wr_cycle[10877] = 1'b0;  addr_rom[10877]='h00000db4;  wr_data_rom[10877]='h00000000;
    rd_cycle[10878] = 1'b1;  wr_cycle[10878] = 1'b0;  addr_rom[10878]='h00000db8;  wr_data_rom[10878]='h00000000;
    rd_cycle[10879] = 1'b1;  wr_cycle[10879] = 1'b0;  addr_rom[10879]='h00000dbc;  wr_data_rom[10879]='h00000000;
    rd_cycle[10880] = 1'b1;  wr_cycle[10880] = 1'b0;  addr_rom[10880]='h00000dc0;  wr_data_rom[10880]='h00000000;
    rd_cycle[10881] = 1'b1;  wr_cycle[10881] = 1'b0;  addr_rom[10881]='h00000dc4;  wr_data_rom[10881]='h00000000;
    rd_cycle[10882] = 1'b1;  wr_cycle[10882] = 1'b0;  addr_rom[10882]='h00000dc8;  wr_data_rom[10882]='h00000000;
    rd_cycle[10883] = 1'b1;  wr_cycle[10883] = 1'b0;  addr_rom[10883]='h00000dcc;  wr_data_rom[10883]='h00000000;
    rd_cycle[10884] = 1'b1;  wr_cycle[10884] = 1'b0;  addr_rom[10884]='h00000dd0;  wr_data_rom[10884]='h00000000;
    rd_cycle[10885] = 1'b1;  wr_cycle[10885] = 1'b0;  addr_rom[10885]='h00000dd4;  wr_data_rom[10885]='h00000000;
    rd_cycle[10886] = 1'b1;  wr_cycle[10886] = 1'b0;  addr_rom[10886]='h00000dd8;  wr_data_rom[10886]='h00000000;
    rd_cycle[10887] = 1'b1;  wr_cycle[10887] = 1'b0;  addr_rom[10887]='h00000ddc;  wr_data_rom[10887]='h00000000;
    rd_cycle[10888] = 1'b1;  wr_cycle[10888] = 1'b0;  addr_rom[10888]='h00000de0;  wr_data_rom[10888]='h00000000;
    rd_cycle[10889] = 1'b1;  wr_cycle[10889] = 1'b0;  addr_rom[10889]='h00000de4;  wr_data_rom[10889]='h00000000;
    rd_cycle[10890] = 1'b1;  wr_cycle[10890] = 1'b0;  addr_rom[10890]='h00000de8;  wr_data_rom[10890]='h00000000;
    rd_cycle[10891] = 1'b1;  wr_cycle[10891] = 1'b0;  addr_rom[10891]='h00000dec;  wr_data_rom[10891]='h00000000;
    rd_cycle[10892] = 1'b1;  wr_cycle[10892] = 1'b0;  addr_rom[10892]='h00000df0;  wr_data_rom[10892]='h00000000;
    rd_cycle[10893] = 1'b1;  wr_cycle[10893] = 1'b0;  addr_rom[10893]='h00000df4;  wr_data_rom[10893]='h00000000;
    rd_cycle[10894] = 1'b1;  wr_cycle[10894] = 1'b0;  addr_rom[10894]='h00000df8;  wr_data_rom[10894]='h00000000;
    rd_cycle[10895] = 1'b1;  wr_cycle[10895] = 1'b0;  addr_rom[10895]='h00000dfc;  wr_data_rom[10895]='h00000000;
    rd_cycle[10896] = 1'b1;  wr_cycle[10896] = 1'b0;  addr_rom[10896]='h00000e00;  wr_data_rom[10896]='h00000000;
    rd_cycle[10897] = 1'b1;  wr_cycle[10897] = 1'b0;  addr_rom[10897]='h00000e04;  wr_data_rom[10897]='h00000000;
    rd_cycle[10898] = 1'b1;  wr_cycle[10898] = 1'b0;  addr_rom[10898]='h00000e08;  wr_data_rom[10898]='h00000000;
    rd_cycle[10899] = 1'b1;  wr_cycle[10899] = 1'b0;  addr_rom[10899]='h00000e0c;  wr_data_rom[10899]='h00000000;
    rd_cycle[10900] = 1'b1;  wr_cycle[10900] = 1'b0;  addr_rom[10900]='h00000e10;  wr_data_rom[10900]='h00000000;
    rd_cycle[10901] = 1'b1;  wr_cycle[10901] = 1'b0;  addr_rom[10901]='h00000e14;  wr_data_rom[10901]='h00000000;
    rd_cycle[10902] = 1'b1;  wr_cycle[10902] = 1'b0;  addr_rom[10902]='h00000e18;  wr_data_rom[10902]='h00000000;
    rd_cycle[10903] = 1'b1;  wr_cycle[10903] = 1'b0;  addr_rom[10903]='h00000e1c;  wr_data_rom[10903]='h00000000;
    rd_cycle[10904] = 1'b1;  wr_cycle[10904] = 1'b0;  addr_rom[10904]='h00000e20;  wr_data_rom[10904]='h00000000;
    rd_cycle[10905] = 1'b1;  wr_cycle[10905] = 1'b0;  addr_rom[10905]='h00000e24;  wr_data_rom[10905]='h00000000;
    rd_cycle[10906] = 1'b1;  wr_cycle[10906] = 1'b0;  addr_rom[10906]='h00000e28;  wr_data_rom[10906]='h00000000;
    rd_cycle[10907] = 1'b1;  wr_cycle[10907] = 1'b0;  addr_rom[10907]='h00000e2c;  wr_data_rom[10907]='h00000000;
    rd_cycle[10908] = 1'b1;  wr_cycle[10908] = 1'b0;  addr_rom[10908]='h00000e30;  wr_data_rom[10908]='h00000000;
    rd_cycle[10909] = 1'b1;  wr_cycle[10909] = 1'b0;  addr_rom[10909]='h00000e34;  wr_data_rom[10909]='h00000000;
    rd_cycle[10910] = 1'b1;  wr_cycle[10910] = 1'b0;  addr_rom[10910]='h00000e38;  wr_data_rom[10910]='h00000000;
    rd_cycle[10911] = 1'b1;  wr_cycle[10911] = 1'b0;  addr_rom[10911]='h00000e3c;  wr_data_rom[10911]='h00000000;
    rd_cycle[10912] = 1'b1;  wr_cycle[10912] = 1'b0;  addr_rom[10912]='h00000e40;  wr_data_rom[10912]='h00000000;
    rd_cycle[10913] = 1'b1;  wr_cycle[10913] = 1'b0;  addr_rom[10913]='h00000e44;  wr_data_rom[10913]='h00000000;
    rd_cycle[10914] = 1'b1;  wr_cycle[10914] = 1'b0;  addr_rom[10914]='h00000e48;  wr_data_rom[10914]='h00000000;
    rd_cycle[10915] = 1'b1;  wr_cycle[10915] = 1'b0;  addr_rom[10915]='h00000e4c;  wr_data_rom[10915]='h00000000;
    rd_cycle[10916] = 1'b1;  wr_cycle[10916] = 1'b0;  addr_rom[10916]='h00000e50;  wr_data_rom[10916]='h00000000;
    rd_cycle[10917] = 1'b1;  wr_cycle[10917] = 1'b0;  addr_rom[10917]='h00000e54;  wr_data_rom[10917]='h00000000;
    rd_cycle[10918] = 1'b1;  wr_cycle[10918] = 1'b0;  addr_rom[10918]='h00000e58;  wr_data_rom[10918]='h00000000;
    rd_cycle[10919] = 1'b1;  wr_cycle[10919] = 1'b0;  addr_rom[10919]='h00000e5c;  wr_data_rom[10919]='h00000000;
    rd_cycle[10920] = 1'b1;  wr_cycle[10920] = 1'b0;  addr_rom[10920]='h00000e60;  wr_data_rom[10920]='h00000000;
    rd_cycle[10921] = 1'b1;  wr_cycle[10921] = 1'b0;  addr_rom[10921]='h00000e64;  wr_data_rom[10921]='h00000000;
    rd_cycle[10922] = 1'b1;  wr_cycle[10922] = 1'b0;  addr_rom[10922]='h00000e68;  wr_data_rom[10922]='h00000000;
    rd_cycle[10923] = 1'b1;  wr_cycle[10923] = 1'b0;  addr_rom[10923]='h00000e6c;  wr_data_rom[10923]='h00000000;
    rd_cycle[10924] = 1'b1;  wr_cycle[10924] = 1'b0;  addr_rom[10924]='h00000e70;  wr_data_rom[10924]='h00000000;
    rd_cycle[10925] = 1'b1;  wr_cycle[10925] = 1'b0;  addr_rom[10925]='h00000e74;  wr_data_rom[10925]='h00000000;
    rd_cycle[10926] = 1'b1;  wr_cycle[10926] = 1'b0;  addr_rom[10926]='h00000e78;  wr_data_rom[10926]='h00000000;
    rd_cycle[10927] = 1'b1;  wr_cycle[10927] = 1'b0;  addr_rom[10927]='h00000e7c;  wr_data_rom[10927]='h00000000;
    rd_cycle[10928] = 1'b1;  wr_cycle[10928] = 1'b0;  addr_rom[10928]='h00000e80;  wr_data_rom[10928]='h00000000;
    rd_cycle[10929] = 1'b1;  wr_cycle[10929] = 1'b0;  addr_rom[10929]='h00000e84;  wr_data_rom[10929]='h00000000;
    rd_cycle[10930] = 1'b1;  wr_cycle[10930] = 1'b0;  addr_rom[10930]='h00000e88;  wr_data_rom[10930]='h00000000;
    rd_cycle[10931] = 1'b1;  wr_cycle[10931] = 1'b0;  addr_rom[10931]='h00000e8c;  wr_data_rom[10931]='h00000000;
    rd_cycle[10932] = 1'b1;  wr_cycle[10932] = 1'b0;  addr_rom[10932]='h00000e90;  wr_data_rom[10932]='h00000000;
    rd_cycle[10933] = 1'b1;  wr_cycle[10933] = 1'b0;  addr_rom[10933]='h00000e94;  wr_data_rom[10933]='h00000000;
    rd_cycle[10934] = 1'b1;  wr_cycle[10934] = 1'b0;  addr_rom[10934]='h00000e98;  wr_data_rom[10934]='h00000000;
    rd_cycle[10935] = 1'b1;  wr_cycle[10935] = 1'b0;  addr_rom[10935]='h00000e9c;  wr_data_rom[10935]='h00000000;
    rd_cycle[10936] = 1'b1;  wr_cycle[10936] = 1'b0;  addr_rom[10936]='h00000ea0;  wr_data_rom[10936]='h00000000;
    rd_cycle[10937] = 1'b1;  wr_cycle[10937] = 1'b0;  addr_rom[10937]='h00000ea4;  wr_data_rom[10937]='h00000000;
    rd_cycle[10938] = 1'b1;  wr_cycle[10938] = 1'b0;  addr_rom[10938]='h00000ea8;  wr_data_rom[10938]='h00000000;
    rd_cycle[10939] = 1'b1;  wr_cycle[10939] = 1'b0;  addr_rom[10939]='h00000eac;  wr_data_rom[10939]='h00000000;
    rd_cycle[10940] = 1'b1;  wr_cycle[10940] = 1'b0;  addr_rom[10940]='h00000eb0;  wr_data_rom[10940]='h00000000;
    rd_cycle[10941] = 1'b1;  wr_cycle[10941] = 1'b0;  addr_rom[10941]='h00000eb4;  wr_data_rom[10941]='h00000000;
    rd_cycle[10942] = 1'b1;  wr_cycle[10942] = 1'b0;  addr_rom[10942]='h00000eb8;  wr_data_rom[10942]='h00000000;
    rd_cycle[10943] = 1'b1;  wr_cycle[10943] = 1'b0;  addr_rom[10943]='h00000ebc;  wr_data_rom[10943]='h00000000;
    rd_cycle[10944] = 1'b1;  wr_cycle[10944] = 1'b0;  addr_rom[10944]='h00000ec0;  wr_data_rom[10944]='h00000000;
    rd_cycle[10945] = 1'b1;  wr_cycle[10945] = 1'b0;  addr_rom[10945]='h00000ec4;  wr_data_rom[10945]='h00000000;
    rd_cycle[10946] = 1'b1;  wr_cycle[10946] = 1'b0;  addr_rom[10946]='h00000ec8;  wr_data_rom[10946]='h00000000;
    rd_cycle[10947] = 1'b1;  wr_cycle[10947] = 1'b0;  addr_rom[10947]='h00000ecc;  wr_data_rom[10947]='h00000000;
    rd_cycle[10948] = 1'b1;  wr_cycle[10948] = 1'b0;  addr_rom[10948]='h00000ed0;  wr_data_rom[10948]='h00000000;
    rd_cycle[10949] = 1'b1;  wr_cycle[10949] = 1'b0;  addr_rom[10949]='h00000ed4;  wr_data_rom[10949]='h00000000;
    rd_cycle[10950] = 1'b1;  wr_cycle[10950] = 1'b0;  addr_rom[10950]='h00000ed8;  wr_data_rom[10950]='h00000000;
    rd_cycle[10951] = 1'b1;  wr_cycle[10951] = 1'b0;  addr_rom[10951]='h00000edc;  wr_data_rom[10951]='h00000000;
    rd_cycle[10952] = 1'b1;  wr_cycle[10952] = 1'b0;  addr_rom[10952]='h00000ee0;  wr_data_rom[10952]='h00000000;
    rd_cycle[10953] = 1'b1;  wr_cycle[10953] = 1'b0;  addr_rom[10953]='h00000ee4;  wr_data_rom[10953]='h00000000;
    rd_cycle[10954] = 1'b1;  wr_cycle[10954] = 1'b0;  addr_rom[10954]='h00000ee8;  wr_data_rom[10954]='h00000000;
    rd_cycle[10955] = 1'b1;  wr_cycle[10955] = 1'b0;  addr_rom[10955]='h00000eec;  wr_data_rom[10955]='h00000000;
    rd_cycle[10956] = 1'b1;  wr_cycle[10956] = 1'b0;  addr_rom[10956]='h00000ef0;  wr_data_rom[10956]='h00000000;
    rd_cycle[10957] = 1'b1;  wr_cycle[10957] = 1'b0;  addr_rom[10957]='h00000ef4;  wr_data_rom[10957]='h00000000;
    rd_cycle[10958] = 1'b1;  wr_cycle[10958] = 1'b0;  addr_rom[10958]='h00000ef8;  wr_data_rom[10958]='h00000000;
    rd_cycle[10959] = 1'b1;  wr_cycle[10959] = 1'b0;  addr_rom[10959]='h00000efc;  wr_data_rom[10959]='h00000000;
    rd_cycle[10960] = 1'b1;  wr_cycle[10960] = 1'b0;  addr_rom[10960]='h00000f00;  wr_data_rom[10960]='h00000000;
    rd_cycle[10961] = 1'b1;  wr_cycle[10961] = 1'b0;  addr_rom[10961]='h00000f04;  wr_data_rom[10961]='h00000000;
    rd_cycle[10962] = 1'b1;  wr_cycle[10962] = 1'b0;  addr_rom[10962]='h00000f08;  wr_data_rom[10962]='h00000000;
    rd_cycle[10963] = 1'b1;  wr_cycle[10963] = 1'b0;  addr_rom[10963]='h00000f0c;  wr_data_rom[10963]='h00000000;
    rd_cycle[10964] = 1'b1;  wr_cycle[10964] = 1'b0;  addr_rom[10964]='h00000f10;  wr_data_rom[10964]='h00000000;
    rd_cycle[10965] = 1'b1;  wr_cycle[10965] = 1'b0;  addr_rom[10965]='h00000f14;  wr_data_rom[10965]='h00000000;
    rd_cycle[10966] = 1'b1;  wr_cycle[10966] = 1'b0;  addr_rom[10966]='h00000f18;  wr_data_rom[10966]='h00000000;
    rd_cycle[10967] = 1'b1;  wr_cycle[10967] = 1'b0;  addr_rom[10967]='h00000f1c;  wr_data_rom[10967]='h00000000;
    rd_cycle[10968] = 1'b1;  wr_cycle[10968] = 1'b0;  addr_rom[10968]='h00000f20;  wr_data_rom[10968]='h00000000;
    rd_cycle[10969] = 1'b1;  wr_cycle[10969] = 1'b0;  addr_rom[10969]='h00000f24;  wr_data_rom[10969]='h00000000;
    rd_cycle[10970] = 1'b1;  wr_cycle[10970] = 1'b0;  addr_rom[10970]='h00000f28;  wr_data_rom[10970]='h00000000;
    rd_cycle[10971] = 1'b1;  wr_cycle[10971] = 1'b0;  addr_rom[10971]='h00000f2c;  wr_data_rom[10971]='h00000000;
    rd_cycle[10972] = 1'b1;  wr_cycle[10972] = 1'b0;  addr_rom[10972]='h00000f30;  wr_data_rom[10972]='h00000000;
    rd_cycle[10973] = 1'b1;  wr_cycle[10973] = 1'b0;  addr_rom[10973]='h00000f34;  wr_data_rom[10973]='h00000000;
    rd_cycle[10974] = 1'b1;  wr_cycle[10974] = 1'b0;  addr_rom[10974]='h00000f38;  wr_data_rom[10974]='h00000000;
    rd_cycle[10975] = 1'b1;  wr_cycle[10975] = 1'b0;  addr_rom[10975]='h00000f3c;  wr_data_rom[10975]='h00000000;
    rd_cycle[10976] = 1'b1;  wr_cycle[10976] = 1'b0;  addr_rom[10976]='h00000f40;  wr_data_rom[10976]='h00000000;
    rd_cycle[10977] = 1'b1;  wr_cycle[10977] = 1'b0;  addr_rom[10977]='h00000f44;  wr_data_rom[10977]='h00000000;
    rd_cycle[10978] = 1'b1;  wr_cycle[10978] = 1'b0;  addr_rom[10978]='h00000f48;  wr_data_rom[10978]='h00000000;
    rd_cycle[10979] = 1'b1;  wr_cycle[10979] = 1'b0;  addr_rom[10979]='h00000f4c;  wr_data_rom[10979]='h00000000;
    rd_cycle[10980] = 1'b1;  wr_cycle[10980] = 1'b0;  addr_rom[10980]='h00000f50;  wr_data_rom[10980]='h00000000;
    rd_cycle[10981] = 1'b1;  wr_cycle[10981] = 1'b0;  addr_rom[10981]='h00000f54;  wr_data_rom[10981]='h00000000;
    rd_cycle[10982] = 1'b1;  wr_cycle[10982] = 1'b0;  addr_rom[10982]='h00000f58;  wr_data_rom[10982]='h00000000;
    rd_cycle[10983] = 1'b1;  wr_cycle[10983] = 1'b0;  addr_rom[10983]='h00000f5c;  wr_data_rom[10983]='h00000000;
    rd_cycle[10984] = 1'b1;  wr_cycle[10984] = 1'b0;  addr_rom[10984]='h00000f60;  wr_data_rom[10984]='h00000000;
    rd_cycle[10985] = 1'b1;  wr_cycle[10985] = 1'b0;  addr_rom[10985]='h00000f64;  wr_data_rom[10985]='h00000000;
    rd_cycle[10986] = 1'b1;  wr_cycle[10986] = 1'b0;  addr_rom[10986]='h00000f68;  wr_data_rom[10986]='h00000000;
    rd_cycle[10987] = 1'b1;  wr_cycle[10987] = 1'b0;  addr_rom[10987]='h00000f6c;  wr_data_rom[10987]='h00000000;
    rd_cycle[10988] = 1'b1;  wr_cycle[10988] = 1'b0;  addr_rom[10988]='h00000f70;  wr_data_rom[10988]='h00000000;
    rd_cycle[10989] = 1'b1;  wr_cycle[10989] = 1'b0;  addr_rom[10989]='h00000f74;  wr_data_rom[10989]='h00000000;
    rd_cycle[10990] = 1'b1;  wr_cycle[10990] = 1'b0;  addr_rom[10990]='h00000f78;  wr_data_rom[10990]='h00000000;
    rd_cycle[10991] = 1'b1;  wr_cycle[10991] = 1'b0;  addr_rom[10991]='h00000f7c;  wr_data_rom[10991]='h00000000;
    rd_cycle[10992] = 1'b1;  wr_cycle[10992] = 1'b0;  addr_rom[10992]='h00000f80;  wr_data_rom[10992]='h00000000;
    rd_cycle[10993] = 1'b1;  wr_cycle[10993] = 1'b0;  addr_rom[10993]='h00000f84;  wr_data_rom[10993]='h00000000;
    rd_cycle[10994] = 1'b1;  wr_cycle[10994] = 1'b0;  addr_rom[10994]='h00000f88;  wr_data_rom[10994]='h00000000;
    rd_cycle[10995] = 1'b1;  wr_cycle[10995] = 1'b0;  addr_rom[10995]='h00000f8c;  wr_data_rom[10995]='h00000000;
    rd_cycle[10996] = 1'b1;  wr_cycle[10996] = 1'b0;  addr_rom[10996]='h00000f90;  wr_data_rom[10996]='h00000000;
    rd_cycle[10997] = 1'b1;  wr_cycle[10997] = 1'b0;  addr_rom[10997]='h00000f94;  wr_data_rom[10997]='h00000000;
    rd_cycle[10998] = 1'b1;  wr_cycle[10998] = 1'b0;  addr_rom[10998]='h00000f98;  wr_data_rom[10998]='h00000000;
    rd_cycle[10999] = 1'b1;  wr_cycle[10999] = 1'b0;  addr_rom[10999]='h00000f9c;  wr_data_rom[10999]='h00000000;
    rd_cycle[11000] = 1'b1;  wr_cycle[11000] = 1'b0;  addr_rom[11000]='h00000fa0;  wr_data_rom[11000]='h00000000;
    rd_cycle[11001] = 1'b1;  wr_cycle[11001] = 1'b0;  addr_rom[11001]='h00000fa4;  wr_data_rom[11001]='h00000000;
    rd_cycle[11002] = 1'b1;  wr_cycle[11002] = 1'b0;  addr_rom[11002]='h00000fa8;  wr_data_rom[11002]='h00000000;
    rd_cycle[11003] = 1'b1;  wr_cycle[11003] = 1'b0;  addr_rom[11003]='h00000fac;  wr_data_rom[11003]='h00000000;
    rd_cycle[11004] = 1'b1;  wr_cycle[11004] = 1'b0;  addr_rom[11004]='h00000fb0;  wr_data_rom[11004]='h00000000;
    rd_cycle[11005] = 1'b1;  wr_cycle[11005] = 1'b0;  addr_rom[11005]='h00000fb4;  wr_data_rom[11005]='h00000000;
    rd_cycle[11006] = 1'b1;  wr_cycle[11006] = 1'b0;  addr_rom[11006]='h00000fb8;  wr_data_rom[11006]='h00000000;
    rd_cycle[11007] = 1'b1;  wr_cycle[11007] = 1'b0;  addr_rom[11007]='h00000fbc;  wr_data_rom[11007]='h00000000;
    rd_cycle[11008] = 1'b1;  wr_cycle[11008] = 1'b0;  addr_rom[11008]='h00000fc0;  wr_data_rom[11008]='h00000000;
    rd_cycle[11009] = 1'b1;  wr_cycle[11009] = 1'b0;  addr_rom[11009]='h00000fc4;  wr_data_rom[11009]='h00000000;
    rd_cycle[11010] = 1'b1;  wr_cycle[11010] = 1'b0;  addr_rom[11010]='h00000fc8;  wr_data_rom[11010]='h00000000;
    rd_cycle[11011] = 1'b1;  wr_cycle[11011] = 1'b0;  addr_rom[11011]='h00000fcc;  wr_data_rom[11011]='h00000000;
    rd_cycle[11012] = 1'b1;  wr_cycle[11012] = 1'b0;  addr_rom[11012]='h00000fd0;  wr_data_rom[11012]='h00000000;
    rd_cycle[11013] = 1'b1;  wr_cycle[11013] = 1'b0;  addr_rom[11013]='h00000fd4;  wr_data_rom[11013]='h00000000;
    rd_cycle[11014] = 1'b1;  wr_cycle[11014] = 1'b0;  addr_rom[11014]='h00000fd8;  wr_data_rom[11014]='h00000000;
    rd_cycle[11015] = 1'b1;  wr_cycle[11015] = 1'b0;  addr_rom[11015]='h00000fdc;  wr_data_rom[11015]='h00000000;
    rd_cycle[11016] = 1'b1;  wr_cycle[11016] = 1'b0;  addr_rom[11016]='h00000fe0;  wr_data_rom[11016]='h00000000;
    rd_cycle[11017] = 1'b1;  wr_cycle[11017] = 1'b0;  addr_rom[11017]='h00000fe4;  wr_data_rom[11017]='h00000000;
    rd_cycle[11018] = 1'b1;  wr_cycle[11018] = 1'b0;  addr_rom[11018]='h00000fe8;  wr_data_rom[11018]='h00000000;
    rd_cycle[11019] = 1'b1;  wr_cycle[11019] = 1'b0;  addr_rom[11019]='h00000fec;  wr_data_rom[11019]='h00000000;
    rd_cycle[11020] = 1'b1;  wr_cycle[11020] = 1'b0;  addr_rom[11020]='h00000ff0;  wr_data_rom[11020]='h00000000;
    rd_cycle[11021] = 1'b1;  wr_cycle[11021] = 1'b0;  addr_rom[11021]='h00000ff4;  wr_data_rom[11021]='h00000000;
    rd_cycle[11022] = 1'b1;  wr_cycle[11022] = 1'b0;  addr_rom[11022]='h00000ff8;  wr_data_rom[11022]='h00000000;
    rd_cycle[11023] = 1'b1;  wr_cycle[11023] = 1'b0;  addr_rom[11023]='h00000ffc;  wr_data_rom[11023]='h00000000;
    rd_cycle[11024] = 1'b1;  wr_cycle[11024] = 1'b0;  addr_rom[11024]='h00001000;  wr_data_rom[11024]='h00000000;
    rd_cycle[11025] = 1'b1;  wr_cycle[11025] = 1'b0;  addr_rom[11025]='h00001004;  wr_data_rom[11025]='h00000000;
    rd_cycle[11026] = 1'b1;  wr_cycle[11026] = 1'b0;  addr_rom[11026]='h00001008;  wr_data_rom[11026]='h00000000;
    rd_cycle[11027] = 1'b1;  wr_cycle[11027] = 1'b0;  addr_rom[11027]='h0000100c;  wr_data_rom[11027]='h00000000;
    rd_cycle[11028] = 1'b1;  wr_cycle[11028] = 1'b0;  addr_rom[11028]='h00001010;  wr_data_rom[11028]='h00000000;
    rd_cycle[11029] = 1'b1;  wr_cycle[11029] = 1'b0;  addr_rom[11029]='h00001014;  wr_data_rom[11029]='h00000000;
    rd_cycle[11030] = 1'b1;  wr_cycle[11030] = 1'b0;  addr_rom[11030]='h00001018;  wr_data_rom[11030]='h00000000;
    rd_cycle[11031] = 1'b1;  wr_cycle[11031] = 1'b0;  addr_rom[11031]='h0000101c;  wr_data_rom[11031]='h00000000;
    rd_cycle[11032] = 1'b1;  wr_cycle[11032] = 1'b0;  addr_rom[11032]='h00001020;  wr_data_rom[11032]='h00000000;
    rd_cycle[11033] = 1'b1;  wr_cycle[11033] = 1'b0;  addr_rom[11033]='h00001024;  wr_data_rom[11033]='h00000000;
    rd_cycle[11034] = 1'b1;  wr_cycle[11034] = 1'b0;  addr_rom[11034]='h00001028;  wr_data_rom[11034]='h00000000;
    rd_cycle[11035] = 1'b1;  wr_cycle[11035] = 1'b0;  addr_rom[11035]='h0000102c;  wr_data_rom[11035]='h00000000;
    rd_cycle[11036] = 1'b1;  wr_cycle[11036] = 1'b0;  addr_rom[11036]='h00001030;  wr_data_rom[11036]='h00000000;
    rd_cycle[11037] = 1'b1;  wr_cycle[11037] = 1'b0;  addr_rom[11037]='h00001034;  wr_data_rom[11037]='h00000000;
    rd_cycle[11038] = 1'b1;  wr_cycle[11038] = 1'b0;  addr_rom[11038]='h00001038;  wr_data_rom[11038]='h00000000;
    rd_cycle[11039] = 1'b1;  wr_cycle[11039] = 1'b0;  addr_rom[11039]='h0000103c;  wr_data_rom[11039]='h00000000;
    rd_cycle[11040] = 1'b1;  wr_cycle[11040] = 1'b0;  addr_rom[11040]='h00001040;  wr_data_rom[11040]='h00000000;
    rd_cycle[11041] = 1'b1;  wr_cycle[11041] = 1'b0;  addr_rom[11041]='h00001044;  wr_data_rom[11041]='h00000000;
    rd_cycle[11042] = 1'b1;  wr_cycle[11042] = 1'b0;  addr_rom[11042]='h00001048;  wr_data_rom[11042]='h00000000;
    rd_cycle[11043] = 1'b1;  wr_cycle[11043] = 1'b0;  addr_rom[11043]='h0000104c;  wr_data_rom[11043]='h00000000;
    rd_cycle[11044] = 1'b1;  wr_cycle[11044] = 1'b0;  addr_rom[11044]='h00001050;  wr_data_rom[11044]='h00000000;
    rd_cycle[11045] = 1'b1;  wr_cycle[11045] = 1'b0;  addr_rom[11045]='h00001054;  wr_data_rom[11045]='h00000000;
    rd_cycle[11046] = 1'b1;  wr_cycle[11046] = 1'b0;  addr_rom[11046]='h00001058;  wr_data_rom[11046]='h00000000;
    rd_cycle[11047] = 1'b1;  wr_cycle[11047] = 1'b0;  addr_rom[11047]='h0000105c;  wr_data_rom[11047]='h00000000;
    rd_cycle[11048] = 1'b1;  wr_cycle[11048] = 1'b0;  addr_rom[11048]='h00001060;  wr_data_rom[11048]='h00000000;
    rd_cycle[11049] = 1'b1;  wr_cycle[11049] = 1'b0;  addr_rom[11049]='h00001064;  wr_data_rom[11049]='h00000000;
    rd_cycle[11050] = 1'b1;  wr_cycle[11050] = 1'b0;  addr_rom[11050]='h00001068;  wr_data_rom[11050]='h00000000;
    rd_cycle[11051] = 1'b1;  wr_cycle[11051] = 1'b0;  addr_rom[11051]='h0000106c;  wr_data_rom[11051]='h00000000;
    rd_cycle[11052] = 1'b1;  wr_cycle[11052] = 1'b0;  addr_rom[11052]='h00001070;  wr_data_rom[11052]='h00000000;
    rd_cycle[11053] = 1'b1;  wr_cycle[11053] = 1'b0;  addr_rom[11053]='h00001074;  wr_data_rom[11053]='h00000000;
    rd_cycle[11054] = 1'b1;  wr_cycle[11054] = 1'b0;  addr_rom[11054]='h00001078;  wr_data_rom[11054]='h00000000;
    rd_cycle[11055] = 1'b1;  wr_cycle[11055] = 1'b0;  addr_rom[11055]='h0000107c;  wr_data_rom[11055]='h00000000;
    rd_cycle[11056] = 1'b1;  wr_cycle[11056] = 1'b0;  addr_rom[11056]='h00001080;  wr_data_rom[11056]='h00000000;
    rd_cycle[11057] = 1'b1;  wr_cycle[11057] = 1'b0;  addr_rom[11057]='h00001084;  wr_data_rom[11057]='h00000000;
    rd_cycle[11058] = 1'b1;  wr_cycle[11058] = 1'b0;  addr_rom[11058]='h00001088;  wr_data_rom[11058]='h00000000;
    rd_cycle[11059] = 1'b1;  wr_cycle[11059] = 1'b0;  addr_rom[11059]='h0000108c;  wr_data_rom[11059]='h00000000;
    rd_cycle[11060] = 1'b1;  wr_cycle[11060] = 1'b0;  addr_rom[11060]='h00001090;  wr_data_rom[11060]='h00000000;
    rd_cycle[11061] = 1'b1;  wr_cycle[11061] = 1'b0;  addr_rom[11061]='h00001094;  wr_data_rom[11061]='h00000000;
    rd_cycle[11062] = 1'b1;  wr_cycle[11062] = 1'b0;  addr_rom[11062]='h00001098;  wr_data_rom[11062]='h00000000;
    rd_cycle[11063] = 1'b1;  wr_cycle[11063] = 1'b0;  addr_rom[11063]='h0000109c;  wr_data_rom[11063]='h00000000;
    rd_cycle[11064] = 1'b1;  wr_cycle[11064] = 1'b0;  addr_rom[11064]='h000010a0;  wr_data_rom[11064]='h00000000;
    rd_cycle[11065] = 1'b1;  wr_cycle[11065] = 1'b0;  addr_rom[11065]='h000010a4;  wr_data_rom[11065]='h00000000;
    rd_cycle[11066] = 1'b1;  wr_cycle[11066] = 1'b0;  addr_rom[11066]='h000010a8;  wr_data_rom[11066]='h00000000;
    rd_cycle[11067] = 1'b1;  wr_cycle[11067] = 1'b0;  addr_rom[11067]='h000010ac;  wr_data_rom[11067]='h00000000;
    rd_cycle[11068] = 1'b1;  wr_cycle[11068] = 1'b0;  addr_rom[11068]='h000010b0;  wr_data_rom[11068]='h00000000;
    rd_cycle[11069] = 1'b1;  wr_cycle[11069] = 1'b0;  addr_rom[11069]='h000010b4;  wr_data_rom[11069]='h00000000;
    rd_cycle[11070] = 1'b1;  wr_cycle[11070] = 1'b0;  addr_rom[11070]='h000010b8;  wr_data_rom[11070]='h00000000;
    rd_cycle[11071] = 1'b1;  wr_cycle[11071] = 1'b0;  addr_rom[11071]='h000010bc;  wr_data_rom[11071]='h00000000;
    rd_cycle[11072] = 1'b1;  wr_cycle[11072] = 1'b0;  addr_rom[11072]='h000010c0;  wr_data_rom[11072]='h00000000;
    rd_cycle[11073] = 1'b1;  wr_cycle[11073] = 1'b0;  addr_rom[11073]='h000010c4;  wr_data_rom[11073]='h00000000;
    rd_cycle[11074] = 1'b1;  wr_cycle[11074] = 1'b0;  addr_rom[11074]='h000010c8;  wr_data_rom[11074]='h00000000;
    rd_cycle[11075] = 1'b1;  wr_cycle[11075] = 1'b0;  addr_rom[11075]='h000010cc;  wr_data_rom[11075]='h00000000;
    rd_cycle[11076] = 1'b1;  wr_cycle[11076] = 1'b0;  addr_rom[11076]='h000010d0;  wr_data_rom[11076]='h00000000;
    rd_cycle[11077] = 1'b1;  wr_cycle[11077] = 1'b0;  addr_rom[11077]='h000010d4;  wr_data_rom[11077]='h00000000;
    rd_cycle[11078] = 1'b1;  wr_cycle[11078] = 1'b0;  addr_rom[11078]='h000010d8;  wr_data_rom[11078]='h00000000;
    rd_cycle[11079] = 1'b1;  wr_cycle[11079] = 1'b0;  addr_rom[11079]='h000010dc;  wr_data_rom[11079]='h00000000;
    rd_cycle[11080] = 1'b1;  wr_cycle[11080] = 1'b0;  addr_rom[11080]='h000010e0;  wr_data_rom[11080]='h00000000;
    rd_cycle[11081] = 1'b1;  wr_cycle[11081] = 1'b0;  addr_rom[11081]='h000010e4;  wr_data_rom[11081]='h00000000;
    rd_cycle[11082] = 1'b1;  wr_cycle[11082] = 1'b0;  addr_rom[11082]='h000010e8;  wr_data_rom[11082]='h00000000;
    rd_cycle[11083] = 1'b1;  wr_cycle[11083] = 1'b0;  addr_rom[11083]='h000010ec;  wr_data_rom[11083]='h00000000;
    rd_cycle[11084] = 1'b1;  wr_cycle[11084] = 1'b0;  addr_rom[11084]='h000010f0;  wr_data_rom[11084]='h00000000;
    rd_cycle[11085] = 1'b1;  wr_cycle[11085] = 1'b0;  addr_rom[11085]='h000010f4;  wr_data_rom[11085]='h00000000;
    rd_cycle[11086] = 1'b1;  wr_cycle[11086] = 1'b0;  addr_rom[11086]='h000010f8;  wr_data_rom[11086]='h00000000;
    rd_cycle[11087] = 1'b1;  wr_cycle[11087] = 1'b0;  addr_rom[11087]='h000010fc;  wr_data_rom[11087]='h00000000;
    rd_cycle[11088] = 1'b1;  wr_cycle[11088] = 1'b0;  addr_rom[11088]='h00001100;  wr_data_rom[11088]='h00000000;
    rd_cycle[11089] = 1'b1;  wr_cycle[11089] = 1'b0;  addr_rom[11089]='h00001104;  wr_data_rom[11089]='h00000000;
    rd_cycle[11090] = 1'b1;  wr_cycle[11090] = 1'b0;  addr_rom[11090]='h00001108;  wr_data_rom[11090]='h00000000;
    rd_cycle[11091] = 1'b1;  wr_cycle[11091] = 1'b0;  addr_rom[11091]='h0000110c;  wr_data_rom[11091]='h00000000;
    rd_cycle[11092] = 1'b1;  wr_cycle[11092] = 1'b0;  addr_rom[11092]='h00001110;  wr_data_rom[11092]='h00000000;
    rd_cycle[11093] = 1'b1;  wr_cycle[11093] = 1'b0;  addr_rom[11093]='h00001114;  wr_data_rom[11093]='h00000000;
    rd_cycle[11094] = 1'b1;  wr_cycle[11094] = 1'b0;  addr_rom[11094]='h00001118;  wr_data_rom[11094]='h00000000;
    rd_cycle[11095] = 1'b1;  wr_cycle[11095] = 1'b0;  addr_rom[11095]='h0000111c;  wr_data_rom[11095]='h00000000;
    rd_cycle[11096] = 1'b1;  wr_cycle[11096] = 1'b0;  addr_rom[11096]='h00001120;  wr_data_rom[11096]='h00000000;
    rd_cycle[11097] = 1'b1;  wr_cycle[11097] = 1'b0;  addr_rom[11097]='h00001124;  wr_data_rom[11097]='h00000000;
    rd_cycle[11098] = 1'b1;  wr_cycle[11098] = 1'b0;  addr_rom[11098]='h00001128;  wr_data_rom[11098]='h00000000;
    rd_cycle[11099] = 1'b1;  wr_cycle[11099] = 1'b0;  addr_rom[11099]='h0000112c;  wr_data_rom[11099]='h00000000;
    rd_cycle[11100] = 1'b1;  wr_cycle[11100] = 1'b0;  addr_rom[11100]='h00001130;  wr_data_rom[11100]='h00000000;
    rd_cycle[11101] = 1'b1;  wr_cycle[11101] = 1'b0;  addr_rom[11101]='h00001134;  wr_data_rom[11101]='h00000000;
    rd_cycle[11102] = 1'b1;  wr_cycle[11102] = 1'b0;  addr_rom[11102]='h00001138;  wr_data_rom[11102]='h00000000;
    rd_cycle[11103] = 1'b1;  wr_cycle[11103] = 1'b0;  addr_rom[11103]='h0000113c;  wr_data_rom[11103]='h00000000;
    rd_cycle[11104] = 1'b1;  wr_cycle[11104] = 1'b0;  addr_rom[11104]='h00001140;  wr_data_rom[11104]='h00000000;
    rd_cycle[11105] = 1'b1;  wr_cycle[11105] = 1'b0;  addr_rom[11105]='h00001144;  wr_data_rom[11105]='h00000000;
    rd_cycle[11106] = 1'b1;  wr_cycle[11106] = 1'b0;  addr_rom[11106]='h00001148;  wr_data_rom[11106]='h00000000;
    rd_cycle[11107] = 1'b1;  wr_cycle[11107] = 1'b0;  addr_rom[11107]='h0000114c;  wr_data_rom[11107]='h00000000;
    rd_cycle[11108] = 1'b1;  wr_cycle[11108] = 1'b0;  addr_rom[11108]='h00001150;  wr_data_rom[11108]='h00000000;
    rd_cycle[11109] = 1'b1;  wr_cycle[11109] = 1'b0;  addr_rom[11109]='h00001154;  wr_data_rom[11109]='h00000000;
    rd_cycle[11110] = 1'b1;  wr_cycle[11110] = 1'b0;  addr_rom[11110]='h00001158;  wr_data_rom[11110]='h00000000;
    rd_cycle[11111] = 1'b1;  wr_cycle[11111] = 1'b0;  addr_rom[11111]='h0000115c;  wr_data_rom[11111]='h00000000;
    rd_cycle[11112] = 1'b1;  wr_cycle[11112] = 1'b0;  addr_rom[11112]='h00001160;  wr_data_rom[11112]='h00000000;
    rd_cycle[11113] = 1'b1;  wr_cycle[11113] = 1'b0;  addr_rom[11113]='h00001164;  wr_data_rom[11113]='h00000000;
    rd_cycle[11114] = 1'b1;  wr_cycle[11114] = 1'b0;  addr_rom[11114]='h00001168;  wr_data_rom[11114]='h00000000;
    rd_cycle[11115] = 1'b1;  wr_cycle[11115] = 1'b0;  addr_rom[11115]='h0000116c;  wr_data_rom[11115]='h00000000;
    rd_cycle[11116] = 1'b1;  wr_cycle[11116] = 1'b0;  addr_rom[11116]='h00001170;  wr_data_rom[11116]='h00000000;
    rd_cycle[11117] = 1'b1;  wr_cycle[11117] = 1'b0;  addr_rom[11117]='h00001174;  wr_data_rom[11117]='h00000000;
    rd_cycle[11118] = 1'b1;  wr_cycle[11118] = 1'b0;  addr_rom[11118]='h00001178;  wr_data_rom[11118]='h00000000;
    rd_cycle[11119] = 1'b1;  wr_cycle[11119] = 1'b0;  addr_rom[11119]='h0000117c;  wr_data_rom[11119]='h00000000;
    rd_cycle[11120] = 1'b1;  wr_cycle[11120] = 1'b0;  addr_rom[11120]='h00001180;  wr_data_rom[11120]='h00000000;
    rd_cycle[11121] = 1'b1;  wr_cycle[11121] = 1'b0;  addr_rom[11121]='h00001184;  wr_data_rom[11121]='h00000000;
    rd_cycle[11122] = 1'b1;  wr_cycle[11122] = 1'b0;  addr_rom[11122]='h00001188;  wr_data_rom[11122]='h00000000;
    rd_cycle[11123] = 1'b1;  wr_cycle[11123] = 1'b0;  addr_rom[11123]='h0000118c;  wr_data_rom[11123]='h00000000;
    rd_cycle[11124] = 1'b1;  wr_cycle[11124] = 1'b0;  addr_rom[11124]='h00001190;  wr_data_rom[11124]='h00000000;
    rd_cycle[11125] = 1'b1;  wr_cycle[11125] = 1'b0;  addr_rom[11125]='h00001194;  wr_data_rom[11125]='h00000000;
    rd_cycle[11126] = 1'b1;  wr_cycle[11126] = 1'b0;  addr_rom[11126]='h00001198;  wr_data_rom[11126]='h00000000;
    rd_cycle[11127] = 1'b1;  wr_cycle[11127] = 1'b0;  addr_rom[11127]='h0000119c;  wr_data_rom[11127]='h00000000;
    rd_cycle[11128] = 1'b1;  wr_cycle[11128] = 1'b0;  addr_rom[11128]='h000011a0;  wr_data_rom[11128]='h00000000;
    rd_cycle[11129] = 1'b1;  wr_cycle[11129] = 1'b0;  addr_rom[11129]='h000011a4;  wr_data_rom[11129]='h00000000;
    rd_cycle[11130] = 1'b1;  wr_cycle[11130] = 1'b0;  addr_rom[11130]='h000011a8;  wr_data_rom[11130]='h00000000;
    rd_cycle[11131] = 1'b1;  wr_cycle[11131] = 1'b0;  addr_rom[11131]='h000011ac;  wr_data_rom[11131]='h00000000;
    rd_cycle[11132] = 1'b1;  wr_cycle[11132] = 1'b0;  addr_rom[11132]='h000011b0;  wr_data_rom[11132]='h00000000;
    rd_cycle[11133] = 1'b1;  wr_cycle[11133] = 1'b0;  addr_rom[11133]='h000011b4;  wr_data_rom[11133]='h00000000;
    rd_cycle[11134] = 1'b1;  wr_cycle[11134] = 1'b0;  addr_rom[11134]='h000011b8;  wr_data_rom[11134]='h00000000;
    rd_cycle[11135] = 1'b1;  wr_cycle[11135] = 1'b0;  addr_rom[11135]='h000011bc;  wr_data_rom[11135]='h00000000;
    rd_cycle[11136] = 1'b1;  wr_cycle[11136] = 1'b0;  addr_rom[11136]='h000011c0;  wr_data_rom[11136]='h00000000;
    rd_cycle[11137] = 1'b1;  wr_cycle[11137] = 1'b0;  addr_rom[11137]='h000011c4;  wr_data_rom[11137]='h00000000;
    rd_cycle[11138] = 1'b1;  wr_cycle[11138] = 1'b0;  addr_rom[11138]='h000011c8;  wr_data_rom[11138]='h00000000;
    rd_cycle[11139] = 1'b1;  wr_cycle[11139] = 1'b0;  addr_rom[11139]='h000011cc;  wr_data_rom[11139]='h00000000;
    rd_cycle[11140] = 1'b1;  wr_cycle[11140] = 1'b0;  addr_rom[11140]='h000011d0;  wr_data_rom[11140]='h00000000;
    rd_cycle[11141] = 1'b1;  wr_cycle[11141] = 1'b0;  addr_rom[11141]='h000011d4;  wr_data_rom[11141]='h00000000;
    rd_cycle[11142] = 1'b1;  wr_cycle[11142] = 1'b0;  addr_rom[11142]='h000011d8;  wr_data_rom[11142]='h00000000;
    rd_cycle[11143] = 1'b1;  wr_cycle[11143] = 1'b0;  addr_rom[11143]='h000011dc;  wr_data_rom[11143]='h00000000;
    rd_cycle[11144] = 1'b1;  wr_cycle[11144] = 1'b0;  addr_rom[11144]='h000011e0;  wr_data_rom[11144]='h00000000;
    rd_cycle[11145] = 1'b1;  wr_cycle[11145] = 1'b0;  addr_rom[11145]='h000011e4;  wr_data_rom[11145]='h00000000;
    rd_cycle[11146] = 1'b1;  wr_cycle[11146] = 1'b0;  addr_rom[11146]='h000011e8;  wr_data_rom[11146]='h00000000;
    rd_cycle[11147] = 1'b1;  wr_cycle[11147] = 1'b0;  addr_rom[11147]='h000011ec;  wr_data_rom[11147]='h00000000;
    rd_cycle[11148] = 1'b1;  wr_cycle[11148] = 1'b0;  addr_rom[11148]='h000011f0;  wr_data_rom[11148]='h00000000;
    rd_cycle[11149] = 1'b1;  wr_cycle[11149] = 1'b0;  addr_rom[11149]='h000011f4;  wr_data_rom[11149]='h00000000;
    rd_cycle[11150] = 1'b1;  wr_cycle[11150] = 1'b0;  addr_rom[11150]='h000011f8;  wr_data_rom[11150]='h00000000;
    rd_cycle[11151] = 1'b1;  wr_cycle[11151] = 1'b0;  addr_rom[11151]='h000011fc;  wr_data_rom[11151]='h00000000;
    rd_cycle[11152] = 1'b1;  wr_cycle[11152] = 1'b0;  addr_rom[11152]='h00001200;  wr_data_rom[11152]='h00000000;
    rd_cycle[11153] = 1'b1;  wr_cycle[11153] = 1'b0;  addr_rom[11153]='h00001204;  wr_data_rom[11153]='h00000000;
    rd_cycle[11154] = 1'b1;  wr_cycle[11154] = 1'b0;  addr_rom[11154]='h00001208;  wr_data_rom[11154]='h00000000;
    rd_cycle[11155] = 1'b1;  wr_cycle[11155] = 1'b0;  addr_rom[11155]='h0000120c;  wr_data_rom[11155]='h00000000;
    rd_cycle[11156] = 1'b1;  wr_cycle[11156] = 1'b0;  addr_rom[11156]='h00001210;  wr_data_rom[11156]='h00000000;
    rd_cycle[11157] = 1'b1;  wr_cycle[11157] = 1'b0;  addr_rom[11157]='h00001214;  wr_data_rom[11157]='h00000000;
    rd_cycle[11158] = 1'b1;  wr_cycle[11158] = 1'b0;  addr_rom[11158]='h00001218;  wr_data_rom[11158]='h00000000;
    rd_cycle[11159] = 1'b1;  wr_cycle[11159] = 1'b0;  addr_rom[11159]='h0000121c;  wr_data_rom[11159]='h00000000;
    rd_cycle[11160] = 1'b1;  wr_cycle[11160] = 1'b0;  addr_rom[11160]='h00001220;  wr_data_rom[11160]='h00000000;
    rd_cycle[11161] = 1'b1;  wr_cycle[11161] = 1'b0;  addr_rom[11161]='h00001224;  wr_data_rom[11161]='h00000000;
    rd_cycle[11162] = 1'b1;  wr_cycle[11162] = 1'b0;  addr_rom[11162]='h00001228;  wr_data_rom[11162]='h00000000;
    rd_cycle[11163] = 1'b1;  wr_cycle[11163] = 1'b0;  addr_rom[11163]='h0000122c;  wr_data_rom[11163]='h00000000;
    rd_cycle[11164] = 1'b1;  wr_cycle[11164] = 1'b0;  addr_rom[11164]='h00001230;  wr_data_rom[11164]='h00000000;
    rd_cycle[11165] = 1'b1;  wr_cycle[11165] = 1'b0;  addr_rom[11165]='h00001234;  wr_data_rom[11165]='h00000000;
    rd_cycle[11166] = 1'b1;  wr_cycle[11166] = 1'b0;  addr_rom[11166]='h00001238;  wr_data_rom[11166]='h00000000;
    rd_cycle[11167] = 1'b1;  wr_cycle[11167] = 1'b0;  addr_rom[11167]='h0000123c;  wr_data_rom[11167]='h00000000;
    rd_cycle[11168] = 1'b1;  wr_cycle[11168] = 1'b0;  addr_rom[11168]='h00001240;  wr_data_rom[11168]='h00000000;
    rd_cycle[11169] = 1'b1;  wr_cycle[11169] = 1'b0;  addr_rom[11169]='h00001244;  wr_data_rom[11169]='h00000000;
    rd_cycle[11170] = 1'b1;  wr_cycle[11170] = 1'b0;  addr_rom[11170]='h00001248;  wr_data_rom[11170]='h00000000;
    rd_cycle[11171] = 1'b1;  wr_cycle[11171] = 1'b0;  addr_rom[11171]='h0000124c;  wr_data_rom[11171]='h00000000;
    rd_cycle[11172] = 1'b1;  wr_cycle[11172] = 1'b0;  addr_rom[11172]='h00001250;  wr_data_rom[11172]='h00000000;
    rd_cycle[11173] = 1'b1;  wr_cycle[11173] = 1'b0;  addr_rom[11173]='h00001254;  wr_data_rom[11173]='h00000000;
    rd_cycle[11174] = 1'b1;  wr_cycle[11174] = 1'b0;  addr_rom[11174]='h00001258;  wr_data_rom[11174]='h00000000;
    rd_cycle[11175] = 1'b1;  wr_cycle[11175] = 1'b0;  addr_rom[11175]='h0000125c;  wr_data_rom[11175]='h00000000;
    rd_cycle[11176] = 1'b1;  wr_cycle[11176] = 1'b0;  addr_rom[11176]='h00001260;  wr_data_rom[11176]='h00000000;
    rd_cycle[11177] = 1'b1;  wr_cycle[11177] = 1'b0;  addr_rom[11177]='h00001264;  wr_data_rom[11177]='h00000000;
    rd_cycle[11178] = 1'b1;  wr_cycle[11178] = 1'b0;  addr_rom[11178]='h00001268;  wr_data_rom[11178]='h00000000;
    rd_cycle[11179] = 1'b1;  wr_cycle[11179] = 1'b0;  addr_rom[11179]='h0000126c;  wr_data_rom[11179]='h00000000;
    rd_cycle[11180] = 1'b1;  wr_cycle[11180] = 1'b0;  addr_rom[11180]='h00001270;  wr_data_rom[11180]='h00000000;
    rd_cycle[11181] = 1'b1;  wr_cycle[11181] = 1'b0;  addr_rom[11181]='h00001274;  wr_data_rom[11181]='h00000000;
    rd_cycle[11182] = 1'b1;  wr_cycle[11182] = 1'b0;  addr_rom[11182]='h00001278;  wr_data_rom[11182]='h00000000;
    rd_cycle[11183] = 1'b1;  wr_cycle[11183] = 1'b0;  addr_rom[11183]='h0000127c;  wr_data_rom[11183]='h00000000;
    rd_cycle[11184] = 1'b1;  wr_cycle[11184] = 1'b0;  addr_rom[11184]='h00001280;  wr_data_rom[11184]='h00000000;
    rd_cycle[11185] = 1'b1;  wr_cycle[11185] = 1'b0;  addr_rom[11185]='h00001284;  wr_data_rom[11185]='h00000000;
    rd_cycle[11186] = 1'b1;  wr_cycle[11186] = 1'b0;  addr_rom[11186]='h00001288;  wr_data_rom[11186]='h00000000;
    rd_cycle[11187] = 1'b1;  wr_cycle[11187] = 1'b0;  addr_rom[11187]='h0000128c;  wr_data_rom[11187]='h00000000;
    rd_cycle[11188] = 1'b1;  wr_cycle[11188] = 1'b0;  addr_rom[11188]='h00001290;  wr_data_rom[11188]='h00000000;
    rd_cycle[11189] = 1'b1;  wr_cycle[11189] = 1'b0;  addr_rom[11189]='h00001294;  wr_data_rom[11189]='h00000000;
    rd_cycle[11190] = 1'b1;  wr_cycle[11190] = 1'b0;  addr_rom[11190]='h00001298;  wr_data_rom[11190]='h00000000;
    rd_cycle[11191] = 1'b1;  wr_cycle[11191] = 1'b0;  addr_rom[11191]='h0000129c;  wr_data_rom[11191]='h00000000;
    rd_cycle[11192] = 1'b1;  wr_cycle[11192] = 1'b0;  addr_rom[11192]='h000012a0;  wr_data_rom[11192]='h00000000;
    rd_cycle[11193] = 1'b1;  wr_cycle[11193] = 1'b0;  addr_rom[11193]='h000012a4;  wr_data_rom[11193]='h00000000;
    rd_cycle[11194] = 1'b1;  wr_cycle[11194] = 1'b0;  addr_rom[11194]='h000012a8;  wr_data_rom[11194]='h00000000;
    rd_cycle[11195] = 1'b1;  wr_cycle[11195] = 1'b0;  addr_rom[11195]='h000012ac;  wr_data_rom[11195]='h00000000;
    rd_cycle[11196] = 1'b1;  wr_cycle[11196] = 1'b0;  addr_rom[11196]='h000012b0;  wr_data_rom[11196]='h00000000;
    rd_cycle[11197] = 1'b1;  wr_cycle[11197] = 1'b0;  addr_rom[11197]='h000012b4;  wr_data_rom[11197]='h00000000;
    rd_cycle[11198] = 1'b1;  wr_cycle[11198] = 1'b0;  addr_rom[11198]='h000012b8;  wr_data_rom[11198]='h00000000;
    rd_cycle[11199] = 1'b1;  wr_cycle[11199] = 1'b0;  addr_rom[11199]='h000012bc;  wr_data_rom[11199]='h00000000;
    rd_cycle[11200] = 1'b1;  wr_cycle[11200] = 1'b0;  addr_rom[11200]='h000012c0;  wr_data_rom[11200]='h00000000;
    rd_cycle[11201] = 1'b1;  wr_cycle[11201] = 1'b0;  addr_rom[11201]='h000012c4;  wr_data_rom[11201]='h00000000;
    rd_cycle[11202] = 1'b1;  wr_cycle[11202] = 1'b0;  addr_rom[11202]='h000012c8;  wr_data_rom[11202]='h00000000;
    rd_cycle[11203] = 1'b1;  wr_cycle[11203] = 1'b0;  addr_rom[11203]='h000012cc;  wr_data_rom[11203]='h00000000;
    rd_cycle[11204] = 1'b1;  wr_cycle[11204] = 1'b0;  addr_rom[11204]='h000012d0;  wr_data_rom[11204]='h00000000;
    rd_cycle[11205] = 1'b1;  wr_cycle[11205] = 1'b0;  addr_rom[11205]='h000012d4;  wr_data_rom[11205]='h00000000;
    rd_cycle[11206] = 1'b1;  wr_cycle[11206] = 1'b0;  addr_rom[11206]='h000012d8;  wr_data_rom[11206]='h00000000;
    rd_cycle[11207] = 1'b1;  wr_cycle[11207] = 1'b0;  addr_rom[11207]='h000012dc;  wr_data_rom[11207]='h00000000;
    rd_cycle[11208] = 1'b1;  wr_cycle[11208] = 1'b0;  addr_rom[11208]='h000012e0;  wr_data_rom[11208]='h00000000;
    rd_cycle[11209] = 1'b1;  wr_cycle[11209] = 1'b0;  addr_rom[11209]='h000012e4;  wr_data_rom[11209]='h00000000;
    rd_cycle[11210] = 1'b1;  wr_cycle[11210] = 1'b0;  addr_rom[11210]='h000012e8;  wr_data_rom[11210]='h00000000;
    rd_cycle[11211] = 1'b1;  wr_cycle[11211] = 1'b0;  addr_rom[11211]='h000012ec;  wr_data_rom[11211]='h00000000;
    rd_cycle[11212] = 1'b1;  wr_cycle[11212] = 1'b0;  addr_rom[11212]='h000012f0;  wr_data_rom[11212]='h00000000;
    rd_cycle[11213] = 1'b1;  wr_cycle[11213] = 1'b0;  addr_rom[11213]='h000012f4;  wr_data_rom[11213]='h00000000;
    rd_cycle[11214] = 1'b1;  wr_cycle[11214] = 1'b0;  addr_rom[11214]='h000012f8;  wr_data_rom[11214]='h00000000;
    rd_cycle[11215] = 1'b1;  wr_cycle[11215] = 1'b0;  addr_rom[11215]='h000012fc;  wr_data_rom[11215]='h00000000;
    rd_cycle[11216] = 1'b1;  wr_cycle[11216] = 1'b0;  addr_rom[11216]='h00001300;  wr_data_rom[11216]='h00000000;
    rd_cycle[11217] = 1'b1;  wr_cycle[11217] = 1'b0;  addr_rom[11217]='h00001304;  wr_data_rom[11217]='h00000000;
    rd_cycle[11218] = 1'b1;  wr_cycle[11218] = 1'b0;  addr_rom[11218]='h00001308;  wr_data_rom[11218]='h00000000;
    rd_cycle[11219] = 1'b1;  wr_cycle[11219] = 1'b0;  addr_rom[11219]='h0000130c;  wr_data_rom[11219]='h00000000;
    rd_cycle[11220] = 1'b1;  wr_cycle[11220] = 1'b0;  addr_rom[11220]='h00001310;  wr_data_rom[11220]='h00000000;
    rd_cycle[11221] = 1'b1;  wr_cycle[11221] = 1'b0;  addr_rom[11221]='h00001314;  wr_data_rom[11221]='h00000000;
    rd_cycle[11222] = 1'b1;  wr_cycle[11222] = 1'b0;  addr_rom[11222]='h00001318;  wr_data_rom[11222]='h00000000;
    rd_cycle[11223] = 1'b1;  wr_cycle[11223] = 1'b0;  addr_rom[11223]='h0000131c;  wr_data_rom[11223]='h00000000;
    rd_cycle[11224] = 1'b1;  wr_cycle[11224] = 1'b0;  addr_rom[11224]='h00001320;  wr_data_rom[11224]='h00000000;
    rd_cycle[11225] = 1'b1;  wr_cycle[11225] = 1'b0;  addr_rom[11225]='h00001324;  wr_data_rom[11225]='h00000000;
    rd_cycle[11226] = 1'b1;  wr_cycle[11226] = 1'b0;  addr_rom[11226]='h00001328;  wr_data_rom[11226]='h00000000;
    rd_cycle[11227] = 1'b1;  wr_cycle[11227] = 1'b0;  addr_rom[11227]='h0000132c;  wr_data_rom[11227]='h00000000;
    rd_cycle[11228] = 1'b1;  wr_cycle[11228] = 1'b0;  addr_rom[11228]='h00001330;  wr_data_rom[11228]='h00000000;
    rd_cycle[11229] = 1'b1;  wr_cycle[11229] = 1'b0;  addr_rom[11229]='h00001334;  wr_data_rom[11229]='h00000000;
    rd_cycle[11230] = 1'b1;  wr_cycle[11230] = 1'b0;  addr_rom[11230]='h00001338;  wr_data_rom[11230]='h00000000;
    rd_cycle[11231] = 1'b1;  wr_cycle[11231] = 1'b0;  addr_rom[11231]='h0000133c;  wr_data_rom[11231]='h00000000;
    rd_cycle[11232] = 1'b1;  wr_cycle[11232] = 1'b0;  addr_rom[11232]='h00001340;  wr_data_rom[11232]='h00000000;
    rd_cycle[11233] = 1'b1;  wr_cycle[11233] = 1'b0;  addr_rom[11233]='h00001344;  wr_data_rom[11233]='h00000000;
    rd_cycle[11234] = 1'b1;  wr_cycle[11234] = 1'b0;  addr_rom[11234]='h00001348;  wr_data_rom[11234]='h00000000;
    rd_cycle[11235] = 1'b1;  wr_cycle[11235] = 1'b0;  addr_rom[11235]='h0000134c;  wr_data_rom[11235]='h00000000;
    rd_cycle[11236] = 1'b1;  wr_cycle[11236] = 1'b0;  addr_rom[11236]='h00001350;  wr_data_rom[11236]='h00000000;
    rd_cycle[11237] = 1'b1;  wr_cycle[11237] = 1'b0;  addr_rom[11237]='h00001354;  wr_data_rom[11237]='h00000000;
    rd_cycle[11238] = 1'b1;  wr_cycle[11238] = 1'b0;  addr_rom[11238]='h00001358;  wr_data_rom[11238]='h00000000;
    rd_cycle[11239] = 1'b1;  wr_cycle[11239] = 1'b0;  addr_rom[11239]='h0000135c;  wr_data_rom[11239]='h00000000;
    rd_cycle[11240] = 1'b1;  wr_cycle[11240] = 1'b0;  addr_rom[11240]='h00001360;  wr_data_rom[11240]='h00000000;
    rd_cycle[11241] = 1'b1;  wr_cycle[11241] = 1'b0;  addr_rom[11241]='h00001364;  wr_data_rom[11241]='h00000000;
    rd_cycle[11242] = 1'b1;  wr_cycle[11242] = 1'b0;  addr_rom[11242]='h00001368;  wr_data_rom[11242]='h00000000;
    rd_cycle[11243] = 1'b1;  wr_cycle[11243] = 1'b0;  addr_rom[11243]='h0000136c;  wr_data_rom[11243]='h00000000;
    rd_cycle[11244] = 1'b1;  wr_cycle[11244] = 1'b0;  addr_rom[11244]='h00001370;  wr_data_rom[11244]='h00000000;
    rd_cycle[11245] = 1'b1;  wr_cycle[11245] = 1'b0;  addr_rom[11245]='h00001374;  wr_data_rom[11245]='h00000000;
    rd_cycle[11246] = 1'b1;  wr_cycle[11246] = 1'b0;  addr_rom[11246]='h00001378;  wr_data_rom[11246]='h00000000;
    rd_cycle[11247] = 1'b1;  wr_cycle[11247] = 1'b0;  addr_rom[11247]='h0000137c;  wr_data_rom[11247]='h00000000;
    rd_cycle[11248] = 1'b1;  wr_cycle[11248] = 1'b0;  addr_rom[11248]='h00001380;  wr_data_rom[11248]='h00000000;
    rd_cycle[11249] = 1'b1;  wr_cycle[11249] = 1'b0;  addr_rom[11249]='h00001384;  wr_data_rom[11249]='h00000000;
    rd_cycle[11250] = 1'b1;  wr_cycle[11250] = 1'b0;  addr_rom[11250]='h00001388;  wr_data_rom[11250]='h00000000;
    rd_cycle[11251] = 1'b1;  wr_cycle[11251] = 1'b0;  addr_rom[11251]='h0000138c;  wr_data_rom[11251]='h00000000;
    rd_cycle[11252] = 1'b1;  wr_cycle[11252] = 1'b0;  addr_rom[11252]='h00001390;  wr_data_rom[11252]='h00000000;
    rd_cycle[11253] = 1'b1;  wr_cycle[11253] = 1'b0;  addr_rom[11253]='h00001394;  wr_data_rom[11253]='h00000000;
    rd_cycle[11254] = 1'b1;  wr_cycle[11254] = 1'b0;  addr_rom[11254]='h00001398;  wr_data_rom[11254]='h00000000;
    rd_cycle[11255] = 1'b1;  wr_cycle[11255] = 1'b0;  addr_rom[11255]='h0000139c;  wr_data_rom[11255]='h00000000;
    rd_cycle[11256] = 1'b1;  wr_cycle[11256] = 1'b0;  addr_rom[11256]='h000013a0;  wr_data_rom[11256]='h00000000;
    rd_cycle[11257] = 1'b1;  wr_cycle[11257] = 1'b0;  addr_rom[11257]='h000013a4;  wr_data_rom[11257]='h00000000;
    rd_cycle[11258] = 1'b1;  wr_cycle[11258] = 1'b0;  addr_rom[11258]='h000013a8;  wr_data_rom[11258]='h00000000;
    rd_cycle[11259] = 1'b1;  wr_cycle[11259] = 1'b0;  addr_rom[11259]='h000013ac;  wr_data_rom[11259]='h00000000;
    rd_cycle[11260] = 1'b1;  wr_cycle[11260] = 1'b0;  addr_rom[11260]='h000013b0;  wr_data_rom[11260]='h00000000;
    rd_cycle[11261] = 1'b1;  wr_cycle[11261] = 1'b0;  addr_rom[11261]='h000013b4;  wr_data_rom[11261]='h00000000;
    rd_cycle[11262] = 1'b1;  wr_cycle[11262] = 1'b0;  addr_rom[11262]='h000013b8;  wr_data_rom[11262]='h00000000;
    rd_cycle[11263] = 1'b1;  wr_cycle[11263] = 1'b0;  addr_rom[11263]='h000013bc;  wr_data_rom[11263]='h00000000;
    rd_cycle[11264] = 1'b1;  wr_cycle[11264] = 1'b0;  addr_rom[11264]='h000013c0;  wr_data_rom[11264]='h00000000;
    rd_cycle[11265] = 1'b1;  wr_cycle[11265] = 1'b0;  addr_rom[11265]='h000013c4;  wr_data_rom[11265]='h00000000;
    rd_cycle[11266] = 1'b1;  wr_cycle[11266] = 1'b0;  addr_rom[11266]='h000013c8;  wr_data_rom[11266]='h00000000;
    rd_cycle[11267] = 1'b1;  wr_cycle[11267] = 1'b0;  addr_rom[11267]='h000013cc;  wr_data_rom[11267]='h00000000;
    rd_cycle[11268] = 1'b1;  wr_cycle[11268] = 1'b0;  addr_rom[11268]='h000013d0;  wr_data_rom[11268]='h00000000;
    rd_cycle[11269] = 1'b1;  wr_cycle[11269] = 1'b0;  addr_rom[11269]='h000013d4;  wr_data_rom[11269]='h00000000;
    rd_cycle[11270] = 1'b1;  wr_cycle[11270] = 1'b0;  addr_rom[11270]='h000013d8;  wr_data_rom[11270]='h00000000;
    rd_cycle[11271] = 1'b1;  wr_cycle[11271] = 1'b0;  addr_rom[11271]='h000013dc;  wr_data_rom[11271]='h00000000;
    rd_cycle[11272] = 1'b1;  wr_cycle[11272] = 1'b0;  addr_rom[11272]='h000013e0;  wr_data_rom[11272]='h00000000;
    rd_cycle[11273] = 1'b1;  wr_cycle[11273] = 1'b0;  addr_rom[11273]='h000013e4;  wr_data_rom[11273]='h00000000;
    rd_cycle[11274] = 1'b1;  wr_cycle[11274] = 1'b0;  addr_rom[11274]='h000013e8;  wr_data_rom[11274]='h00000000;
    rd_cycle[11275] = 1'b1;  wr_cycle[11275] = 1'b0;  addr_rom[11275]='h000013ec;  wr_data_rom[11275]='h00000000;
    rd_cycle[11276] = 1'b1;  wr_cycle[11276] = 1'b0;  addr_rom[11276]='h000013f0;  wr_data_rom[11276]='h00000000;
    rd_cycle[11277] = 1'b1;  wr_cycle[11277] = 1'b0;  addr_rom[11277]='h000013f4;  wr_data_rom[11277]='h00000000;
    rd_cycle[11278] = 1'b1;  wr_cycle[11278] = 1'b0;  addr_rom[11278]='h000013f8;  wr_data_rom[11278]='h00000000;
    rd_cycle[11279] = 1'b1;  wr_cycle[11279] = 1'b0;  addr_rom[11279]='h000013fc;  wr_data_rom[11279]='h00000000;
    rd_cycle[11280] = 1'b1;  wr_cycle[11280] = 1'b0;  addr_rom[11280]='h00001400;  wr_data_rom[11280]='h00000000;
    rd_cycle[11281] = 1'b1;  wr_cycle[11281] = 1'b0;  addr_rom[11281]='h00001404;  wr_data_rom[11281]='h00000000;
    rd_cycle[11282] = 1'b1;  wr_cycle[11282] = 1'b0;  addr_rom[11282]='h00001408;  wr_data_rom[11282]='h00000000;
    rd_cycle[11283] = 1'b1;  wr_cycle[11283] = 1'b0;  addr_rom[11283]='h0000140c;  wr_data_rom[11283]='h00000000;
    rd_cycle[11284] = 1'b1;  wr_cycle[11284] = 1'b0;  addr_rom[11284]='h00001410;  wr_data_rom[11284]='h00000000;
    rd_cycle[11285] = 1'b1;  wr_cycle[11285] = 1'b0;  addr_rom[11285]='h00001414;  wr_data_rom[11285]='h00000000;
    rd_cycle[11286] = 1'b1;  wr_cycle[11286] = 1'b0;  addr_rom[11286]='h00001418;  wr_data_rom[11286]='h00000000;
    rd_cycle[11287] = 1'b1;  wr_cycle[11287] = 1'b0;  addr_rom[11287]='h0000141c;  wr_data_rom[11287]='h00000000;
    rd_cycle[11288] = 1'b1;  wr_cycle[11288] = 1'b0;  addr_rom[11288]='h00001420;  wr_data_rom[11288]='h00000000;
    rd_cycle[11289] = 1'b1;  wr_cycle[11289] = 1'b0;  addr_rom[11289]='h00001424;  wr_data_rom[11289]='h00000000;
    rd_cycle[11290] = 1'b1;  wr_cycle[11290] = 1'b0;  addr_rom[11290]='h00001428;  wr_data_rom[11290]='h00000000;
    rd_cycle[11291] = 1'b1;  wr_cycle[11291] = 1'b0;  addr_rom[11291]='h0000142c;  wr_data_rom[11291]='h00000000;
    rd_cycle[11292] = 1'b1;  wr_cycle[11292] = 1'b0;  addr_rom[11292]='h00001430;  wr_data_rom[11292]='h00000000;
    rd_cycle[11293] = 1'b1;  wr_cycle[11293] = 1'b0;  addr_rom[11293]='h00001434;  wr_data_rom[11293]='h00000000;
    rd_cycle[11294] = 1'b1;  wr_cycle[11294] = 1'b0;  addr_rom[11294]='h00001438;  wr_data_rom[11294]='h00000000;
    rd_cycle[11295] = 1'b1;  wr_cycle[11295] = 1'b0;  addr_rom[11295]='h0000143c;  wr_data_rom[11295]='h00000000;
    rd_cycle[11296] = 1'b1;  wr_cycle[11296] = 1'b0;  addr_rom[11296]='h00001440;  wr_data_rom[11296]='h00000000;
    rd_cycle[11297] = 1'b1;  wr_cycle[11297] = 1'b0;  addr_rom[11297]='h00001444;  wr_data_rom[11297]='h00000000;
    rd_cycle[11298] = 1'b1;  wr_cycle[11298] = 1'b0;  addr_rom[11298]='h00001448;  wr_data_rom[11298]='h00000000;
    rd_cycle[11299] = 1'b1;  wr_cycle[11299] = 1'b0;  addr_rom[11299]='h0000144c;  wr_data_rom[11299]='h00000000;
    rd_cycle[11300] = 1'b1;  wr_cycle[11300] = 1'b0;  addr_rom[11300]='h00001450;  wr_data_rom[11300]='h00000000;
    rd_cycle[11301] = 1'b1;  wr_cycle[11301] = 1'b0;  addr_rom[11301]='h00001454;  wr_data_rom[11301]='h00000000;
    rd_cycle[11302] = 1'b1;  wr_cycle[11302] = 1'b0;  addr_rom[11302]='h00001458;  wr_data_rom[11302]='h00000000;
    rd_cycle[11303] = 1'b1;  wr_cycle[11303] = 1'b0;  addr_rom[11303]='h0000145c;  wr_data_rom[11303]='h00000000;
    rd_cycle[11304] = 1'b1;  wr_cycle[11304] = 1'b0;  addr_rom[11304]='h00001460;  wr_data_rom[11304]='h00000000;
    rd_cycle[11305] = 1'b1;  wr_cycle[11305] = 1'b0;  addr_rom[11305]='h00001464;  wr_data_rom[11305]='h00000000;
    rd_cycle[11306] = 1'b1;  wr_cycle[11306] = 1'b0;  addr_rom[11306]='h00001468;  wr_data_rom[11306]='h00000000;
    rd_cycle[11307] = 1'b1;  wr_cycle[11307] = 1'b0;  addr_rom[11307]='h0000146c;  wr_data_rom[11307]='h00000000;
    rd_cycle[11308] = 1'b1;  wr_cycle[11308] = 1'b0;  addr_rom[11308]='h00001470;  wr_data_rom[11308]='h00000000;
    rd_cycle[11309] = 1'b1;  wr_cycle[11309] = 1'b0;  addr_rom[11309]='h00001474;  wr_data_rom[11309]='h00000000;
    rd_cycle[11310] = 1'b1;  wr_cycle[11310] = 1'b0;  addr_rom[11310]='h00001478;  wr_data_rom[11310]='h00000000;
    rd_cycle[11311] = 1'b1;  wr_cycle[11311] = 1'b0;  addr_rom[11311]='h0000147c;  wr_data_rom[11311]='h00000000;
    rd_cycle[11312] = 1'b1;  wr_cycle[11312] = 1'b0;  addr_rom[11312]='h00001480;  wr_data_rom[11312]='h00000000;
    rd_cycle[11313] = 1'b1;  wr_cycle[11313] = 1'b0;  addr_rom[11313]='h00001484;  wr_data_rom[11313]='h00000000;
    rd_cycle[11314] = 1'b1;  wr_cycle[11314] = 1'b0;  addr_rom[11314]='h00001488;  wr_data_rom[11314]='h00000000;
    rd_cycle[11315] = 1'b1;  wr_cycle[11315] = 1'b0;  addr_rom[11315]='h0000148c;  wr_data_rom[11315]='h00000000;
    rd_cycle[11316] = 1'b1;  wr_cycle[11316] = 1'b0;  addr_rom[11316]='h00001490;  wr_data_rom[11316]='h00000000;
    rd_cycle[11317] = 1'b1;  wr_cycle[11317] = 1'b0;  addr_rom[11317]='h00001494;  wr_data_rom[11317]='h00000000;
    rd_cycle[11318] = 1'b1;  wr_cycle[11318] = 1'b0;  addr_rom[11318]='h00001498;  wr_data_rom[11318]='h00000000;
    rd_cycle[11319] = 1'b1;  wr_cycle[11319] = 1'b0;  addr_rom[11319]='h0000149c;  wr_data_rom[11319]='h00000000;
    rd_cycle[11320] = 1'b1;  wr_cycle[11320] = 1'b0;  addr_rom[11320]='h000014a0;  wr_data_rom[11320]='h00000000;
    rd_cycle[11321] = 1'b1;  wr_cycle[11321] = 1'b0;  addr_rom[11321]='h000014a4;  wr_data_rom[11321]='h00000000;
    rd_cycle[11322] = 1'b1;  wr_cycle[11322] = 1'b0;  addr_rom[11322]='h000014a8;  wr_data_rom[11322]='h00000000;
    rd_cycle[11323] = 1'b1;  wr_cycle[11323] = 1'b0;  addr_rom[11323]='h000014ac;  wr_data_rom[11323]='h00000000;
    rd_cycle[11324] = 1'b1;  wr_cycle[11324] = 1'b0;  addr_rom[11324]='h000014b0;  wr_data_rom[11324]='h00000000;
    rd_cycle[11325] = 1'b1;  wr_cycle[11325] = 1'b0;  addr_rom[11325]='h000014b4;  wr_data_rom[11325]='h00000000;
    rd_cycle[11326] = 1'b1;  wr_cycle[11326] = 1'b0;  addr_rom[11326]='h000014b8;  wr_data_rom[11326]='h00000000;
    rd_cycle[11327] = 1'b1;  wr_cycle[11327] = 1'b0;  addr_rom[11327]='h000014bc;  wr_data_rom[11327]='h00000000;
    rd_cycle[11328] = 1'b1;  wr_cycle[11328] = 1'b0;  addr_rom[11328]='h000014c0;  wr_data_rom[11328]='h00000000;
    rd_cycle[11329] = 1'b1;  wr_cycle[11329] = 1'b0;  addr_rom[11329]='h000014c4;  wr_data_rom[11329]='h00000000;
    rd_cycle[11330] = 1'b1;  wr_cycle[11330] = 1'b0;  addr_rom[11330]='h000014c8;  wr_data_rom[11330]='h00000000;
    rd_cycle[11331] = 1'b1;  wr_cycle[11331] = 1'b0;  addr_rom[11331]='h000014cc;  wr_data_rom[11331]='h00000000;
    rd_cycle[11332] = 1'b1;  wr_cycle[11332] = 1'b0;  addr_rom[11332]='h000014d0;  wr_data_rom[11332]='h00000000;
    rd_cycle[11333] = 1'b1;  wr_cycle[11333] = 1'b0;  addr_rom[11333]='h000014d4;  wr_data_rom[11333]='h00000000;
    rd_cycle[11334] = 1'b1;  wr_cycle[11334] = 1'b0;  addr_rom[11334]='h000014d8;  wr_data_rom[11334]='h00000000;
    rd_cycle[11335] = 1'b1;  wr_cycle[11335] = 1'b0;  addr_rom[11335]='h000014dc;  wr_data_rom[11335]='h00000000;
    rd_cycle[11336] = 1'b1;  wr_cycle[11336] = 1'b0;  addr_rom[11336]='h000014e0;  wr_data_rom[11336]='h00000000;
    rd_cycle[11337] = 1'b1;  wr_cycle[11337] = 1'b0;  addr_rom[11337]='h000014e4;  wr_data_rom[11337]='h00000000;
    rd_cycle[11338] = 1'b1;  wr_cycle[11338] = 1'b0;  addr_rom[11338]='h000014e8;  wr_data_rom[11338]='h00000000;
    rd_cycle[11339] = 1'b1;  wr_cycle[11339] = 1'b0;  addr_rom[11339]='h000014ec;  wr_data_rom[11339]='h00000000;
    rd_cycle[11340] = 1'b1;  wr_cycle[11340] = 1'b0;  addr_rom[11340]='h000014f0;  wr_data_rom[11340]='h00000000;
    rd_cycle[11341] = 1'b1;  wr_cycle[11341] = 1'b0;  addr_rom[11341]='h000014f4;  wr_data_rom[11341]='h00000000;
    rd_cycle[11342] = 1'b1;  wr_cycle[11342] = 1'b0;  addr_rom[11342]='h000014f8;  wr_data_rom[11342]='h00000000;
    rd_cycle[11343] = 1'b1;  wr_cycle[11343] = 1'b0;  addr_rom[11343]='h000014fc;  wr_data_rom[11343]='h00000000;
    rd_cycle[11344] = 1'b1;  wr_cycle[11344] = 1'b0;  addr_rom[11344]='h00001500;  wr_data_rom[11344]='h00000000;
    rd_cycle[11345] = 1'b1;  wr_cycle[11345] = 1'b0;  addr_rom[11345]='h00001504;  wr_data_rom[11345]='h00000000;
    rd_cycle[11346] = 1'b1;  wr_cycle[11346] = 1'b0;  addr_rom[11346]='h00001508;  wr_data_rom[11346]='h00000000;
    rd_cycle[11347] = 1'b1;  wr_cycle[11347] = 1'b0;  addr_rom[11347]='h0000150c;  wr_data_rom[11347]='h00000000;
    rd_cycle[11348] = 1'b1;  wr_cycle[11348] = 1'b0;  addr_rom[11348]='h00001510;  wr_data_rom[11348]='h00000000;
    rd_cycle[11349] = 1'b1;  wr_cycle[11349] = 1'b0;  addr_rom[11349]='h00001514;  wr_data_rom[11349]='h00000000;
    rd_cycle[11350] = 1'b1;  wr_cycle[11350] = 1'b0;  addr_rom[11350]='h00001518;  wr_data_rom[11350]='h00000000;
    rd_cycle[11351] = 1'b1;  wr_cycle[11351] = 1'b0;  addr_rom[11351]='h0000151c;  wr_data_rom[11351]='h00000000;
    rd_cycle[11352] = 1'b1;  wr_cycle[11352] = 1'b0;  addr_rom[11352]='h00001520;  wr_data_rom[11352]='h00000000;
    rd_cycle[11353] = 1'b1;  wr_cycle[11353] = 1'b0;  addr_rom[11353]='h00001524;  wr_data_rom[11353]='h00000000;
    rd_cycle[11354] = 1'b1;  wr_cycle[11354] = 1'b0;  addr_rom[11354]='h00001528;  wr_data_rom[11354]='h00000000;
    rd_cycle[11355] = 1'b1;  wr_cycle[11355] = 1'b0;  addr_rom[11355]='h0000152c;  wr_data_rom[11355]='h00000000;
    rd_cycle[11356] = 1'b1;  wr_cycle[11356] = 1'b0;  addr_rom[11356]='h00001530;  wr_data_rom[11356]='h00000000;
    rd_cycle[11357] = 1'b1;  wr_cycle[11357] = 1'b0;  addr_rom[11357]='h00001534;  wr_data_rom[11357]='h00000000;
    rd_cycle[11358] = 1'b1;  wr_cycle[11358] = 1'b0;  addr_rom[11358]='h00001538;  wr_data_rom[11358]='h00000000;
    rd_cycle[11359] = 1'b1;  wr_cycle[11359] = 1'b0;  addr_rom[11359]='h0000153c;  wr_data_rom[11359]='h00000000;
    rd_cycle[11360] = 1'b1;  wr_cycle[11360] = 1'b0;  addr_rom[11360]='h00001540;  wr_data_rom[11360]='h00000000;
    rd_cycle[11361] = 1'b1;  wr_cycle[11361] = 1'b0;  addr_rom[11361]='h00001544;  wr_data_rom[11361]='h00000000;
    rd_cycle[11362] = 1'b1;  wr_cycle[11362] = 1'b0;  addr_rom[11362]='h00001548;  wr_data_rom[11362]='h00000000;
    rd_cycle[11363] = 1'b1;  wr_cycle[11363] = 1'b0;  addr_rom[11363]='h0000154c;  wr_data_rom[11363]='h00000000;
    rd_cycle[11364] = 1'b1;  wr_cycle[11364] = 1'b0;  addr_rom[11364]='h00001550;  wr_data_rom[11364]='h00000000;
    rd_cycle[11365] = 1'b1;  wr_cycle[11365] = 1'b0;  addr_rom[11365]='h00001554;  wr_data_rom[11365]='h00000000;
    rd_cycle[11366] = 1'b1;  wr_cycle[11366] = 1'b0;  addr_rom[11366]='h00001558;  wr_data_rom[11366]='h00000000;
    rd_cycle[11367] = 1'b1;  wr_cycle[11367] = 1'b0;  addr_rom[11367]='h0000155c;  wr_data_rom[11367]='h00000000;
    rd_cycle[11368] = 1'b1;  wr_cycle[11368] = 1'b0;  addr_rom[11368]='h00001560;  wr_data_rom[11368]='h00000000;
    rd_cycle[11369] = 1'b1;  wr_cycle[11369] = 1'b0;  addr_rom[11369]='h00001564;  wr_data_rom[11369]='h00000000;
    rd_cycle[11370] = 1'b1;  wr_cycle[11370] = 1'b0;  addr_rom[11370]='h00001568;  wr_data_rom[11370]='h00000000;
    rd_cycle[11371] = 1'b1;  wr_cycle[11371] = 1'b0;  addr_rom[11371]='h0000156c;  wr_data_rom[11371]='h00000000;
    rd_cycle[11372] = 1'b1;  wr_cycle[11372] = 1'b0;  addr_rom[11372]='h00001570;  wr_data_rom[11372]='h00000000;
    rd_cycle[11373] = 1'b1;  wr_cycle[11373] = 1'b0;  addr_rom[11373]='h00001574;  wr_data_rom[11373]='h00000000;
    rd_cycle[11374] = 1'b1;  wr_cycle[11374] = 1'b0;  addr_rom[11374]='h00001578;  wr_data_rom[11374]='h00000000;
    rd_cycle[11375] = 1'b1;  wr_cycle[11375] = 1'b0;  addr_rom[11375]='h0000157c;  wr_data_rom[11375]='h00000000;
    rd_cycle[11376] = 1'b1;  wr_cycle[11376] = 1'b0;  addr_rom[11376]='h00001580;  wr_data_rom[11376]='h00000000;
    rd_cycle[11377] = 1'b1;  wr_cycle[11377] = 1'b0;  addr_rom[11377]='h00001584;  wr_data_rom[11377]='h00000000;
    rd_cycle[11378] = 1'b1;  wr_cycle[11378] = 1'b0;  addr_rom[11378]='h00001588;  wr_data_rom[11378]='h00000000;
    rd_cycle[11379] = 1'b1;  wr_cycle[11379] = 1'b0;  addr_rom[11379]='h0000158c;  wr_data_rom[11379]='h00000000;
    rd_cycle[11380] = 1'b1;  wr_cycle[11380] = 1'b0;  addr_rom[11380]='h00001590;  wr_data_rom[11380]='h00000000;
    rd_cycle[11381] = 1'b1;  wr_cycle[11381] = 1'b0;  addr_rom[11381]='h00001594;  wr_data_rom[11381]='h00000000;
    rd_cycle[11382] = 1'b1;  wr_cycle[11382] = 1'b0;  addr_rom[11382]='h00001598;  wr_data_rom[11382]='h00000000;
    rd_cycle[11383] = 1'b1;  wr_cycle[11383] = 1'b0;  addr_rom[11383]='h0000159c;  wr_data_rom[11383]='h00000000;
    rd_cycle[11384] = 1'b1;  wr_cycle[11384] = 1'b0;  addr_rom[11384]='h000015a0;  wr_data_rom[11384]='h00000000;
    rd_cycle[11385] = 1'b1;  wr_cycle[11385] = 1'b0;  addr_rom[11385]='h000015a4;  wr_data_rom[11385]='h00000000;
    rd_cycle[11386] = 1'b1;  wr_cycle[11386] = 1'b0;  addr_rom[11386]='h000015a8;  wr_data_rom[11386]='h00000000;
    rd_cycle[11387] = 1'b1;  wr_cycle[11387] = 1'b0;  addr_rom[11387]='h000015ac;  wr_data_rom[11387]='h00000000;
    rd_cycle[11388] = 1'b1;  wr_cycle[11388] = 1'b0;  addr_rom[11388]='h000015b0;  wr_data_rom[11388]='h00000000;
    rd_cycle[11389] = 1'b1;  wr_cycle[11389] = 1'b0;  addr_rom[11389]='h000015b4;  wr_data_rom[11389]='h00000000;
    rd_cycle[11390] = 1'b1;  wr_cycle[11390] = 1'b0;  addr_rom[11390]='h000015b8;  wr_data_rom[11390]='h00000000;
    rd_cycle[11391] = 1'b1;  wr_cycle[11391] = 1'b0;  addr_rom[11391]='h000015bc;  wr_data_rom[11391]='h00000000;
    rd_cycle[11392] = 1'b1;  wr_cycle[11392] = 1'b0;  addr_rom[11392]='h000015c0;  wr_data_rom[11392]='h00000000;
    rd_cycle[11393] = 1'b1;  wr_cycle[11393] = 1'b0;  addr_rom[11393]='h000015c4;  wr_data_rom[11393]='h00000000;
    rd_cycle[11394] = 1'b1;  wr_cycle[11394] = 1'b0;  addr_rom[11394]='h000015c8;  wr_data_rom[11394]='h00000000;
    rd_cycle[11395] = 1'b1;  wr_cycle[11395] = 1'b0;  addr_rom[11395]='h000015cc;  wr_data_rom[11395]='h00000000;
    rd_cycle[11396] = 1'b1;  wr_cycle[11396] = 1'b0;  addr_rom[11396]='h000015d0;  wr_data_rom[11396]='h00000000;
    rd_cycle[11397] = 1'b1;  wr_cycle[11397] = 1'b0;  addr_rom[11397]='h000015d4;  wr_data_rom[11397]='h00000000;
    rd_cycle[11398] = 1'b1;  wr_cycle[11398] = 1'b0;  addr_rom[11398]='h000015d8;  wr_data_rom[11398]='h00000000;
    rd_cycle[11399] = 1'b1;  wr_cycle[11399] = 1'b0;  addr_rom[11399]='h000015dc;  wr_data_rom[11399]='h00000000;
    rd_cycle[11400] = 1'b1;  wr_cycle[11400] = 1'b0;  addr_rom[11400]='h000015e0;  wr_data_rom[11400]='h00000000;
    rd_cycle[11401] = 1'b1;  wr_cycle[11401] = 1'b0;  addr_rom[11401]='h000015e4;  wr_data_rom[11401]='h00000000;
    rd_cycle[11402] = 1'b1;  wr_cycle[11402] = 1'b0;  addr_rom[11402]='h000015e8;  wr_data_rom[11402]='h00000000;
    rd_cycle[11403] = 1'b1;  wr_cycle[11403] = 1'b0;  addr_rom[11403]='h000015ec;  wr_data_rom[11403]='h00000000;
    rd_cycle[11404] = 1'b1;  wr_cycle[11404] = 1'b0;  addr_rom[11404]='h000015f0;  wr_data_rom[11404]='h00000000;
    rd_cycle[11405] = 1'b1;  wr_cycle[11405] = 1'b0;  addr_rom[11405]='h000015f4;  wr_data_rom[11405]='h00000000;
    rd_cycle[11406] = 1'b1;  wr_cycle[11406] = 1'b0;  addr_rom[11406]='h000015f8;  wr_data_rom[11406]='h00000000;
    rd_cycle[11407] = 1'b1;  wr_cycle[11407] = 1'b0;  addr_rom[11407]='h000015fc;  wr_data_rom[11407]='h00000000;
    rd_cycle[11408] = 1'b1;  wr_cycle[11408] = 1'b0;  addr_rom[11408]='h00001600;  wr_data_rom[11408]='h00000000;
    rd_cycle[11409] = 1'b1;  wr_cycle[11409] = 1'b0;  addr_rom[11409]='h00001604;  wr_data_rom[11409]='h00000000;
    rd_cycle[11410] = 1'b1;  wr_cycle[11410] = 1'b0;  addr_rom[11410]='h00001608;  wr_data_rom[11410]='h00000000;
    rd_cycle[11411] = 1'b1;  wr_cycle[11411] = 1'b0;  addr_rom[11411]='h0000160c;  wr_data_rom[11411]='h00000000;
    rd_cycle[11412] = 1'b1;  wr_cycle[11412] = 1'b0;  addr_rom[11412]='h00001610;  wr_data_rom[11412]='h00000000;
    rd_cycle[11413] = 1'b1;  wr_cycle[11413] = 1'b0;  addr_rom[11413]='h00001614;  wr_data_rom[11413]='h00000000;
    rd_cycle[11414] = 1'b1;  wr_cycle[11414] = 1'b0;  addr_rom[11414]='h00001618;  wr_data_rom[11414]='h00000000;
    rd_cycle[11415] = 1'b1;  wr_cycle[11415] = 1'b0;  addr_rom[11415]='h0000161c;  wr_data_rom[11415]='h00000000;
    rd_cycle[11416] = 1'b1;  wr_cycle[11416] = 1'b0;  addr_rom[11416]='h00001620;  wr_data_rom[11416]='h00000000;
    rd_cycle[11417] = 1'b1;  wr_cycle[11417] = 1'b0;  addr_rom[11417]='h00001624;  wr_data_rom[11417]='h00000000;
    rd_cycle[11418] = 1'b1;  wr_cycle[11418] = 1'b0;  addr_rom[11418]='h00001628;  wr_data_rom[11418]='h00000000;
    rd_cycle[11419] = 1'b1;  wr_cycle[11419] = 1'b0;  addr_rom[11419]='h0000162c;  wr_data_rom[11419]='h00000000;
    rd_cycle[11420] = 1'b1;  wr_cycle[11420] = 1'b0;  addr_rom[11420]='h00001630;  wr_data_rom[11420]='h00000000;
    rd_cycle[11421] = 1'b1;  wr_cycle[11421] = 1'b0;  addr_rom[11421]='h00001634;  wr_data_rom[11421]='h00000000;
    rd_cycle[11422] = 1'b1;  wr_cycle[11422] = 1'b0;  addr_rom[11422]='h00001638;  wr_data_rom[11422]='h00000000;
    rd_cycle[11423] = 1'b1;  wr_cycle[11423] = 1'b0;  addr_rom[11423]='h0000163c;  wr_data_rom[11423]='h00000000;
    rd_cycle[11424] = 1'b1;  wr_cycle[11424] = 1'b0;  addr_rom[11424]='h00001640;  wr_data_rom[11424]='h00000000;
    rd_cycle[11425] = 1'b1;  wr_cycle[11425] = 1'b0;  addr_rom[11425]='h00001644;  wr_data_rom[11425]='h00000000;
    rd_cycle[11426] = 1'b1;  wr_cycle[11426] = 1'b0;  addr_rom[11426]='h00001648;  wr_data_rom[11426]='h00000000;
    rd_cycle[11427] = 1'b1;  wr_cycle[11427] = 1'b0;  addr_rom[11427]='h0000164c;  wr_data_rom[11427]='h00000000;
    rd_cycle[11428] = 1'b1;  wr_cycle[11428] = 1'b0;  addr_rom[11428]='h00001650;  wr_data_rom[11428]='h00000000;
    rd_cycle[11429] = 1'b1;  wr_cycle[11429] = 1'b0;  addr_rom[11429]='h00001654;  wr_data_rom[11429]='h00000000;
    rd_cycle[11430] = 1'b1;  wr_cycle[11430] = 1'b0;  addr_rom[11430]='h00001658;  wr_data_rom[11430]='h00000000;
    rd_cycle[11431] = 1'b1;  wr_cycle[11431] = 1'b0;  addr_rom[11431]='h0000165c;  wr_data_rom[11431]='h00000000;
    rd_cycle[11432] = 1'b1;  wr_cycle[11432] = 1'b0;  addr_rom[11432]='h00001660;  wr_data_rom[11432]='h00000000;
    rd_cycle[11433] = 1'b1;  wr_cycle[11433] = 1'b0;  addr_rom[11433]='h00001664;  wr_data_rom[11433]='h00000000;
    rd_cycle[11434] = 1'b1;  wr_cycle[11434] = 1'b0;  addr_rom[11434]='h00001668;  wr_data_rom[11434]='h00000000;
    rd_cycle[11435] = 1'b1;  wr_cycle[11435] = 1'b0;  addr_rom[11435]='h0000166c;  wr_data_rom[11435]='h00000000;
    rd_cycle[11436] = 1'b1;  wr_cycle[11436] = 1'b0;  addr_rom[11436]='h00001670;  wr_data_rom[11436]='h00000000;
    rd_cycle[11437] = 1'b1;  wr_cycle[11437] = 1'b0;  addr_rom[11437]='h00001674;  wr_data_rom[11437]='h00000000;
    rd_cycle[11438] = 1'b1;  wr_cycle[11438] = 1'b0;  addr_rom[11438]='h00001678;  wr_data_rom[11438]='h00000000;
    rd_cycle[11439] = 1'b1;  wr_cycle[11439] = 1'b0;  addr_rom[11439]='h0000167c;  wr_data_rom[11439]='h00000000;
    rd_cycle[11440] = 1'b1;  wr_cycle[11440] = 1'b0;  addr_rom[11440]='h00001680;  wr_data_rom[11440]='h00000000;
    rd_cycle[11441] = 1'b1;  wr_cycle[11441] = 1'b0;  addr_rom[11441]='h00001684;  wr_data_rom[11441]='h00000000;
    rd_cycle[11442] = 1'b1;  wr_cycle[11442] = 1'b0;  addr_rom[11442]='h00001688;  wr_data_rom[11442]='h00000000;
    rd_cycle[11443] = 1'b1;  wr_cycle[11443] = 1'b0;  addr_rom[11443]='h0000168c;  wr_data_rom[11443]='h00000000;
    rd_cycle[11444] = 1'b1;  wr_cycle[11444] = 1'b0;  addr_rom[11444]='h00001690;  wr_data_rom[11444]='h00000000;
    rd_cycle[11445] = 1'b1;  wr_cycle[11445] = 1'b0;  addr_rom[11445]='h00001694;  wr_data_rom[11445]='h00000000;
    rd_cycle[11446] = 1'b1;  wr_cycle[11446] = 1'b0;  addr_rom[11446]='h00001698;  wr_data_rom[11446]='h00000000;
    rd_cycle[11447] = 1'b1;  wr_cycle[11447] = 1'b0;  addr_rom[11447]='h0000169c;  wr_data_rom[11447]='h00000000;
    rd_cycle[11448] = 1'b1;  wr_cycle[11448] = 1'b0;  addr_rom[11448]='h000016a0;  wr_data_rom[11448]='h00000000;
    rd_cycle[11449] = 1'b1;  wr_cycle[11449] = 1'b0;  addr_rom[11449]='h000016a4;  wr_data_rom[11449]='h00000000;
    rd_cycle[11450] = 1'b1;  wr_cycle[11450] = 1'b0;  addr_rom[11450]='h000016a8;  wr_data_rom[11450]='h00000000;
    rd_cycle[11451] = 1'b1;  wr_cycle[11451] = 1'b0;  addr_rom[11451]='h000016ac;  wr_data_rom[11451]='h00000000;
    rd_cycle[11452] = 1'b1;  wr_cycle[11452] = 1'b0;  addr_rom[11452]='h000016b0;  wr_data_rom[11452]='h00000000;
    rd_cycle[11453] = 1'b1;  wr_cycle[11453] = 1'b0;  addr_rom[11453]='h000016b4;  wr_data_rom[11453]='h00000000;
    rd_cycle[11454] = 1'b1;  wr_cycle[11454] = 1'b0;  addr_rom[11454]='h000016b8;  wr_data_rom[11454]='h00000000;
    rd_cycle[11455] = 1'b1;  wr_cycle[11455] = 1'b0;  addr_rom[11455]='h000016bc;  wr_data_rom[11455]='h00000000;
    rd_cycle[11456] = 1'b1;  wr_cycle[11456] = 1'b0;  addr_rom[11456]='h000016c0;  wr_data_rom[11456]='h00000000;
    rd_cycle[11457] = 1'b1;  wr_cycle[11457] = 1'b0;  addr_rom[11457]='h000016c4;  wr_data_rom[11457]='h00000000;
    rd_cycle[11458] = 1'b1;  wr_cycle[11458] = 1'b0;  addr_rom[11458]='h000016c8;  wr_data_rom[11458]='h00000000;
    rd_cycle[11459] = 1'b1;  wr_cycle[11459] = 1'b0;  addr_rom[11459]='h000016cc;  wr_data_rom[11459]='h00000000;
    rd_cycle[11460] = 1'b1;  wr_cycle[11460] = 1'b0;  addr_rom[11460]='h000016d0;  wr_data_rom[11460]='h00000000;
    rd_cycle[11461] = 1'b1;  wr_cycle[11461] = 1'b0;  addr_rom[11461]='h000016d4;  wr_data_rom[11461]='h00000000;
    rd_cycle[11462] = 1'b1;  wr_cycle[11462] = 1'b0;  addr_rom[11462]='h000016d8;  wr_data_rom[11462]='h00000000;
    rd_cycle[11463] = 1'b1;  wr_cycle[11463] = 1'b0;  addr_rom[11463]='h000016dc;  wr_data_rom[11463]='h00000000;
    rd_cycle[11464] = 1'b1;  wr_cycle[11464] = 1'b0;  addr_rom[11464]='h000016e0;  wr_data_rom[11464]='h00000000;
    rd_cycle[11465] = 1'b1;  wr_cycle[11465] = 1'b0;  addr_rom[11465]='h000016e4;  wr_data_rom[11465]='h00000000;
    rd_cycle[11466] = 1'b1;  wr_cycle[11466] = 1'b0;  addr_rom[11466]='h000016e8;  wr_data_rom[11466]='h00000000;
    rd_cycle[11467] = 1'b1;  wr_cycle[11467] = 1'b0;  addr_rom[11467]='h000016ec;  wr_data_rom[11467]='h00000000;
    rd_cycle[11468] = 1'b1;  wr_cycle[11468] = 1'b0;  addr_rom[11468]='h000016f0;  wr_data_rom[11468]='h00000000;
    rd_cycle[11469] = 1'b1;  wr_cycle[11469] = 1'b0;  addr_rom[11469]='h000016f4;  wr_data_rom[11469]='h00000000;
    rd_cycle[11470] = 1'b1;  wr_cycle[11470] = 1'b0;  addr_rom[11470]='h000016f8;  wr_data_rom[11470]='h00000000;
    rd_cycle[11471] = 1'b1;  wr_cycle[11471] = 1'b0;  addr_rom[11471]='h000016fc;  wr_data_rom[11471]='h00000000;
    rd_cycle[11472] = 1'b1;  wr_cycle[11472] = 1'b0;  addr_rom[11472]='h00001700;  wr_data_rom[11472]='h00000000;
    rd_cycle[11473] = 1'b1;  wr_cycle[11473] = 1'b0;  addr_rom[11473]='h00001704;  wr_data_rom[11473]='h00000000;
    rd_cycle[11474] = 1'b1;  wr_cycle[11474] = 1'b0;  addr_rom[11474]='h00001708;  wr_data_rom[11474]='h00000000;
    rd_cycle[11475] = 1'b1;  wr_cycle[11475] = 1'b0;  addr_rom[11475]='h0000170c;  wr_data_rom[11475]='h00000000;
    rd_cycle[11476] = 1'b1;  wr_cycle[11476] = 1'b0;  addr_rom[11476]='h00001710;  wr_data_rom[11476]='h00000000;
    rd_cycle[11477] = 1'b1;  wr_cycle[11477] = 1'b0;  addr_rom[11477]='h00001714;  wr_data_rom[11477]='h00000000;
    rd_cycle[11478] = 1'b1;  wr_cycle[11478] = 1'b0;  addr_rom[11478]='h00001718;  wr_data_rom[11478]='h00000000;
    rd_cycle[11479] = 1'b1;  wr_cycle[11479] = 1'b0;  addr_rom[11479]='h0000171c;  wr_data_rom[11479]='h00000000;
    rd_cycle[11480] = 1'b1;  wr_cycle[11480] = 1'b0;  addr_rom[11480]='h00001720;  wr_data_rom[11480]='h00000000;
    rd_cycle[11481] = 1'b1;  wr_cycle[11481] = 1'b0;  addr_rom[11481]='h00001724;  wr_data_rom[11481]='h00000000;
    rd_cycle[11482] = 1'b1;  wr_cycle[11482] = 1'b0;  addr_rom[11482]='h00001728;  wr_data_rom[11482]='h00000000;
    rd_cycle[11483] = 1'b1;  wr_cycle[11483] = 1'b0;  addr_rom[11483]='h0000172c;  wr_data_rom[11483]='h00000000;
    rd_cycle[11484] = 1'b1;  wr_cycle[11484] = 1'b0;  addr_rom[11484]='h00001730;  wr_data_rom[11484]='h00000000;
    rd_cycle[11485] = 1'b1;  wr_cycle[11485] = 1'b0;  addr_rom[11485]='h00001734;  wr_data_rom[11485]='h00000000;
    rd_cycle[11486] = 1'b1;  wr_cycle[11486] = 1'b0;  addr_rom[11486]='h00001738;  wr_data_rom[11486]='h00000000;
    rd_cycle[11487] = 1'b1;  wr_cycle[11487] = 1'b0;  addr_rom[11487]='h0000173c;  wr_data_rom[11487]='h00000000;
    rd_cycle[11488] = 1'b1;  wr_cycle[11488] = 1'b0;  addr_rom[11488]='h00001740;  wr_data_rom[11488]='h00000000;
    rd_cycle[11489] = 1'b1;  wr_cycle[11489] = 1'b0;  addr_rom[11489]='h00001744;  wr_data_rom[11489]='h00000000;
    rd_cycle[11490] = 1'b1;  wr_cycle[11490] = 1'b0;  addr_rom[11490]='h00001748;  wr_data_rom[11490]='h00000000;
    rd_cycle[11491] = 1'b1;  wr_cycle[11491] = 1'b0;  addr_rom[11491]='h0000174c;  wr_data_rom[11491]='h00000000;
    rd_cycle[11492] = 1'b1;  wr_cycle[11492] = 1'b0;  addr_rom[11492]='h00001750;  wr_data_rom[11492]='h00000000;
    rd_cycle[11493] = 1'b1;  wr_cycle[11493] = 1'b0;  addr_rom[11493]='h00001754;  wr_data_rom[11493]='h00000000;
    rd_cycle[11494] = 1'b1;  wr_cycle[11494] = 1'b0;  addr_rom[11494]='h00001758;  wr_data_rom[11494]='h00000000;
    rd_cycle[11495] = 1'b1;  wr_cycle[11495] = 1'b0;  addr_rom[11495]='h0000175c;  wr_data_rom[11495]='h00000000;
    rd_cycle[11496] = 1'b1;  wr_cycle[11496] = 1'b0;  addr_rom[11496]='h00001760;  wr_data_rom[11496]='h00000000;
    rd_cycle[11497] = 1'b1;  wr_cycle[11497] = 1'b0;  addr_rom[11497]='h00001764;  wr_data_rom[11497]='h00000000;
    rd_cycle[11498] = 1'b1;  wr_cycle[11498] = 1'b0;  addr_rom[11498]='h00001768;  wr_data_rom[11498]='h00000000;
    rd_cycle[11499] = 1'b1;  wr_cycle[11499] = 1'b0;  addr_rom[11499]='h0000176c;  wr_data_rom[11499]='h00000000;
    rd_cycle[11500] = 1'b1;  wr_cycle[11500] = 1'b0;  addr_rom[11500]='h00001770;  wr_data_rom[11500]='h00000000;
    rd_cycle[11501] = 1'b1;  wr_cycle[11501] = 1'b0;  addr_rom[11501]='h00001774;  wr_data_rom[11501]='h00000000;
    rd_cycle[11502] = 1'b1;  wr_cycle[11502] = 1'b0;  addr_rom[11502]='h00001778;  wr_data_rom[11502]='h00000000;
    rd_cycle[11503] = 1'b1;  wr_cycle[11503] = 1'b0;  addr_rom[11503]='h0000177c;  wr_data_rom[11503]='h00000000;
    rd_cycle[11504] = 1'b1;  wr_cycle[11504] = 1'b0;  addr_rom[11504]='h00001780;  wr_data_rom[11504]='h00000000;
    rd_cycle[11505] = 1'b1;  wr_cycle[11505] = 1'b0;  addr_rom[11505]='h00001784;  wr_data_rom[11505]='h00000000;
    rd_cycle[11506] = 1'b1;  wr_cycle[11506] = 1'b0;  addr_rom[11506]='h00001788;  wr_data_rom[11506]='h00000000;
    rd_cycle[11507] = 1'b1;  wr_cycle[11507] = 1'b0;  addr_rom[11507]='h0000178c;  wr_data_rom[11507]='h00000000;
    rd_cycle[11508] = 1'b1;  wr_cycle[11508] = 1'b0;  addr_rom[11508]='h00001790;  wr_data_rom[11508]='h00000000;
    rd_cycle[11509] = 1'b1;  wr_cycle[11509] = 1'b0;  addr_rom[11509]='h00001794;  wr_data_rom[11509]='h00000000;
    rd_cycle[11510] = 1'b1;  wr_cycle[11510] = 1'b0;  addr_rom[11510]='h00001798;  wr_data_rom[11510]='h00000000;
    rd_cycle[11511] = 1'b1;  wr_cycle[11511] = 1'b0;  addr_rom[11511]='h0000179c;  wr_data_rom[11511]='h00000000;
    rd_cycle[11512] = 1'b1;  wr_cycle[11512] = 1'b0;  addr_rom[11512]='h000017a0;  wr_data_rom[11512]='h00000000;
    rd_cycle[11513] = 1'b1;  wr_cycle[11513] = 1'b0;  addr_rom[11513]='h000017a4;  wr_data_rom[11513]='h00000000;
    rd_cycle[11514] = 1'b1;  wr_cycle[11514] = 1'b0;  addr_rom[11514]='h000017a8;  wr_data_rom[11514]='h00000000;
    rd_cycle[11515] = 1'b1;  wr_cycle[11515] = 1'b0;  addr_rom[11515]='h000017ac;  wr_data_rom[11515]='h00000000;
    rd_cycle[11516] = 1'b1;  wr_cycle[11516] = 1'b0;  addr_rom[11516]='h000017b0;  wr_data_rom[11516]='h00000000;
    rd_cycle[11517] = 1'b1;  wr_cycle[11517] = 1'b0;  addr_rom[11517]='h000017b4;  wr_data_rom[11517]='h00000000;
    rd_cycle[11518] = 1'b1;  wr_cycle[11518] = 1'b0;  addr_rom[11518]='h000017b8;  wr_data_rom[11518]='h00000000;
    rd_cycle[11519] = 1'b1;  wr_cycle[11519] = 1'b0;  addr_rom[11519]='h000017bc;  wr_data_rom[11519]='h00000000;
    rd_cycle[11520] = 1'b1;  wr_cycle[11520] = 1'b0;  addr_rom[11520]='h000017c0;  wr_data_rom[11520]='h00000000;
    rd_cycle[11521] = 1'b1;  wr_cycle[11521] = 1'b0;  addr_rom[11521]='h000017c4;  wr_data_rom[11521]='h00000000;
    rd_cycle[11522] = 1'b1;  wr_cycle[11522] = 1'b0;  addr_rom[11522]='h000017c8;  wr_data_rom[11522]='h00000000;
    rd_cycle[11523] = 1'b1;  wr_cycle[11523] = 1'b0;  addr_rom[11523]='h000017cc;  wr_data_rom[11523]='h00000000;
    rd_cycle[11524] = 1'b1;  wr_cycle[11524] = 1'b0;  addr_rom[11524]='h000017d0;  wr_data_rom[11524]='h00000000;
    rd_cycle[11525] = 1'b1;  wr_cycle[11525] = 1'b0;  addr_rom[11525]='h000017d4;  wr_data_rom[11525]='h00000000;
    rd_cycle[11526] = 1'b1;  wr_cycle[11526] = 1'b0;  addr_rom[11526]='h000017d8;  wr_data_rom[11526]='h00000000;
    rd_cycle[11527] = 1'b1;  wr_cycle[11527] = 1'b0;  addr_rom[11527]='h000017dc;  wr_data_rom[11527]='h00000000;
    rd_cycle[11528] = 1'b1;  wr_cycle[11528] = 1'b0;  addr_rom[11528]='h000017e0;  wr_data_rom[11528]='h00000000;
    rd_cycle[11529] = 1'b1;  wr_cycle[11529] = 1'b0;  addr_rom[11529]='h000017e4;  wr_data_rom[11529]='h00000000;
    rd_cycle[11530] = 1'b1;  wr_cycle[11530] = 1'b0;  addr_rom[11530]='h000017e8;  wr_data_rom[11530]='h00000000;
    rd_cycle[11531] = 1'b1;  wr_cycle[11531] = 1'b0;  addr_rom[11531]='h000017ec;  wr_data_rom[11531]='h00000000;
    rd_cycle[11532] = 1'b1;  wr_cycle[11532] = 1'b0;  addr_rom[11532]='h000017f0;  wr_data_rom[11532]='h00000000;
    rd_cycle[11533] = 1'b1;  wr_cycle[11533] = 1'b0;  addr_rom[11533]='h000017f4;  wr_data_rom[11533]='h00000000;
    rd_cycle[11534] = 1'b1;  wr_cycle[11534] = 1'b0;  addr_rom[11534]='h000017f8;  wr_data_rom[11534]='h00000000;
    rd_cycle[11535] = 1'b1;  wr_cycle[11535] = 1'b0;  addr_rom[11535]='h000017fc;  wr_data_rom[11535]='h00000000;
    rd_cycle[11536] = 1'b1;  wr_cycle[11536] = 1'b0;  addr_rom[11536]='h00001800;  wr_data_rom[11536]='h00000000;
    rd_cycle[11537] = 1'b1;  wr_cycle[11537] = 1'b0;  addr_rom[11537]='h00001804;  wr_data_rom[11537]='h00000000;
    rd_cycle[11538] = 1'b1;  wr_cycle[11538] = 1'b0;  addr_rom[11538]='h00001808;  wr_data_rom[11538]='h00000000;
    rd_cycle[11539] = 1'b1;  wr_cycle[11539] = 1'b0;  addr_rom[11539]='h0000180c;  wr_data_rom[11539]='h00000000;
    rd_cycle[11540] = 1'b1;  wr_cycle[11540] = 1'b0;  addr_rom[11540]='h00001810;  wr_data_rom[11540]='h00000000;
    rd_cycle[11541] = 1'b1;  wr_cycle[11541] = 1'b0;  addr_rom[11541]='h00001814;  wr_data_rom[11541]='h00000000;
    rd_cycle[11542] = 1'b1;  wr_cycle[11542] = 1'b0;  addr_rom[11542]='h00001818;  wr_data_rom[11542]='h00000000;
    rd_cycle[11543] = 1'b1;  wr_cycle[11543] = 1'b0;  addr_rom[11543]='h0000181c;  wr_data_rom[11543]='h00000000;
    rd_cycle[11544] = 1'b1;  wr_cycle[11544] = 1'b0;  addr_rom[11544]='h00001820;  wr_data_rom[11544]='h00000000;
    rd_cycle[11545] = 1'b1;  wr_cycle[11545] = 1'b0;  addr_rom[11545]='h00001824;  wr_data_rom[11545]='h00000000;
    rd_cycle[11546] = 1'b1;  wr_cycle[11546] = 1'b0;  addr_rom[11546]='h00001828;  wr_data_rom[11546]='h00000000;
    rd_cycle[11547] = 1'b1;  wr_cycle[11547] = 1'b0;  addr_rom[11547]='h0000182c;  wr_data_rom[11547]='h00000000;
    rd_cycle[11548] = 1'b1;  wr_cycle[11548] = 1'b0;  addr_rom[11548]='h00001830;  wr_data_rom[11548]='h00000000;
    rd_cycle[11549] = 1'b1;  wr_cycle[11549] = 1'b0;  addr_rom[11549]='h00001834;  wr_data_rom[11549]='h00000000;
    rd_cycle[11550] = 1'b1;  wr_cycle[11550] = 1'b0;  addr_rom[11550]='h00001838;  wr_data_rom[11550]='h00000000;
    rd_cycle[11551] = 1'b1;  wr_cycle[11551] = 1'b0;  addr_rom[11551]='h0000183c;  wr_data_rom[11551]='h00000000;
    rd_cycle[11552] = 1'b1;  wr_cycle[11552] = 1'b0;  addr_rom[11552]='h00001840;  wr_data_rom[11552]='h00000000;
    rd_cycle[11553] = 1'b1;  wr_cycle[11553] = 1'b0;  addr_rom[11553]='h00001844;  wr_data_rom[11553]='h00000000;
    rd_cycle[11554] = 1'b1;  wr_cycle[11554] = 1'b0;  addr_rom[11554]='h00001848;  wr_data_rom[11554]='h00000000;
    rd_cycle[11555] = 1'b1;  wr_cycle[11555] = 1'b0;  addr_rom[11555]='h0000184c;  wr_data_rom[11555]='h00000000;
    rd_cycle[11556] = 1'b1;  wr_cycle[11556] = 1'b0;  addr_rom[11556]='h00001850;  wr_data_rom[11556]='h00000000;
    rd_cycle[11557] = 1'b1;  wr_cycle[11557] = 1'b0;  addr_rom[11557]='h00001854;  wr_data_rom[11557]='h00000000;
    rd_cycle[11558] = 1'b1;  wr_cycle[11558] = 1'b0;  addr_rom[11558]='h00001858;  wr_data_rom[11558]='h00000000;
    rd_cycle[11559] = 1'b1;  wr_cycle[11559] = 1'b0;  addr_rom[11559]='h0000185c;  wr_data_rom[11559]='h00000000;
    rd_cycle[11560] = 1'b1;  wr_cycle[11560] = 1'b0;  addr_rom[11560]='h00001860;  wr_data_rom[11560]='h00000000;
    rd_cycle[11561] = 1'b1;  wr_cycle[11561] = 1'b0;  addr_rom[11561]='h00001864;  wr_data_rom[11561]='h00000000;
    rd_cycle[11562] = 1'b1;  wr_cycle[11562] = 1'b0;  addr_rom[11562]='h00001868;  wr_data_rom[11562]='h00000000;
    rd_cycle[11563] = 1'b1;  wr_cycle[11563] = 1'b0;  addr_rom[11563]='h0000186c;  wr_data_rom[11563]='h00000000;
    rd_cycle[11564] = 1'b1;  wr_cycle[11564] = 1'b0;  addr_rom[11564]='h00001870;  wr_data_rom[11564]='h00000000;
    rd_cycle[11565] = 1'b1;  wr_cycle[11565] = 1'b0;  addr_rom[11565]='h00001874;  wr_data_rom[11565]='h00000000;
    rd_cycle[11566] = 1'b1;  wr_cycle[11566] = 1'b0;  addr_rom[11566]='h00001878;  wr_data_rom[11566]='h00000000;
    rd_cycle[11567] = 1'b1;  wr_cycle[11567] = 1'b0;  addr_rom[11567]='h0000187c;  wr_data_rom[11567]='h00000000;
    rd_cycle[11568] = 1'b1;  wr_cycle[11568] = 1'b0;  addr_rom[11568]='h00001880;  wr_data_rom[11568]='h00000000;
    rd_cycle[11569] = 1'b1;  wr_cycle[11569] = 1'b0;  addr_rom[11569]='h00001884;  wr_data_rom[11569]='h00000000;
    rd_cycle[11570] = 1'b1;  wr_cycle[11570] = 1'b0;  addr_rom[11570]='h00001888;  wr_data_rom[11570]='h00000000;
    rd_cycle[11571] = 1'b1;  wr_cycle[11571] = 1'b0;  addr_rom[11571]='h0000188c;  wr_data_rom[11571]='h00000000;
    rd_cycle[11572] = 1'b1;  wr_cycle[11572] = 1'b0;  addr_rom[11572]='h00001890;  wr_data_rom[11572]='h00000000;
    rd_cycle[11573] = 1'b1;  wr_cycle[11573] = 1'b0;  addr_rom[11573]='h00001894;  wr_data_rom[11573]='h00000000;
    rd_cycle[11574] = 1'b1;  wr_cycle[11574] = 1'b0;  addr_rom[11574]='h00001898;  wr_data_rom[11574]='h00000000;
    rd_cycle[11575] = 1'b1;  wr_cycle[11575] = 1'b0;  addr_rom[11575]='h0000189c;  wr_data_rom[11575]='h00000000;
    rd_cycle[11576] = 1'b1;  wr_cycle[11576] = 1'b0;  addr_rom[11576]='h000018a0;  wr_data_rom[11576]='h00000000;
    rd_cycle[11577] = 1'b1;  wr_cycle[11577] = 1'b0;  addr_rom[11577]='h000018a4;  wr_data_rom[11577]='h00000000;
    rd_cycle[11578] = 1'b1;  wr_cycle[11578] = 1'b0;  addr_rom[11578]='h000018a8;  wr_data_rom[11578]='h00000000;
    rd_cycle[11579] = 1'b1;  wr_cycle[11579] = 1'b0;  addr_rom[11579]='h000018ac;  wr_data_rom[11579]='h00000000;
    rd_cycle[11580] = 1'b1;  wr_cycle[11580] = 1'b0;  addr_rom[11580]='h000018b0;  wr_data_rom[11580]='h00000000;
    rd_cycle[11581] = 1'b1;  wr_cycle[11581] = 1'b0;  addr_rom[11581]='h000018b4;  wr_data_rom[11581]='h00000000;
    rd_cycle[11582] = 1'b1;  wr_cycle[11582] = 1'b0;  addr_rom[11582]='h000018b8;  wr_data_rom[11582]='h00000000;
    rd_cycle[11583] = 1'b1;  wr_cycle[11583] = 1'b0;  addr_rom[11583]='h000018bc;  wr_data_rom[11583]='h00000000;
    rd_cycle[11584] = 1'b1;  wr_cycle[11584] = 1'b0;  addr_rom[11584]='h000018c0;  wr_data_rom[11584]='h00000000;
    rd_cycle[11585] = 1'b1;  wr_cycle[11585] = 1'b0;  addr_rom[11585]='h000018c4;  wr_data_rom[11585]='h00000000;
    rd_cycle[11586] = 1'b1;  wr_cycle[11586] = 1'b0;  addr_rom[11586]='h000018c8;  wr_data_rom[11586]='h00000000;
    rd_cycle[11587] = 1'b1;  wr_cycle[11587] = 1'b0;  addr_rom[11587]='h000018cc;  wr_data_rom[11587]='h00000000;
    rd_cycle[11588] = 1'b1;  wr_cycle[11588] = 1'b0;  addr_rom[11588]='h000018d0;  wr_data_rom[11588]='h00000000;
    rd_cycle[11589] = 1'b1;  wr_cycle[11589] = 1'b0;  addr_rom[11589]='h000018d4;  wr_data_rom[11589]='h00000000;
    rd_cycle[11590] = 1'b1;  wr_cycle[11590] = 1'b0;  addr_rom[11590]='h000018d8;  wr_data_rom[11590]='h00000000;
    rd_cycle[11591] = 1'b1;  wr_cycle[11591] = 1'b0;  addr_rom[11591]='h000018dc;  wr_data_rom[11591]='h00000000;
    rd_cycle[11592] = 1'b1;  wr_cycle[11592] = 1'b0;  addr_rom[11592]='h000018e0;  wr_data_rom[11592]='h00000000;
    rd_cycle[11593] = 1'b1;  wr_cycle[11593] = 1'b0;  addr_rom[11593]='h000018e4;  wr_data_rom[11593]='h00000000;
    rd_cycle[11594] = 1'b1;  wr_cycle[11594] = 1'b0;  addr_rom[11594]='h000018e8;  wr_data_rom[11594]='h00000000;
    rd_cycle[11595] = 1'b1;  wr_cycle[11595] = 1'b0;  addr_rom[11595]='h000018ec;  wr_data_rom[11595]='h00000000;
    rd_cycle[11596] = 1'b1;  wr_cycle[11596] = 1'b0;  addr_rom[11596]='h000018f0;  wr_data_rom[11596]='h00000000;
    rd_cycle[11597] = 1'b1;  wr_cycle[11597] = 1'b0;  addr_rom[11597]='h000018f4;  wr_data_rom[11597]='h00000000;
    rd_cycle[11598] = 1'b1;  wr_cycle[11598] = 1'b0;  addr_rom[11598]='h000018f8;  wr_data_rom[11598]='h00000000;
    rd_cycle[11599] = 1'b1;  wr_cycle[11599] = 1'b0;  addr_rom[11599]='h000018fc;  wr_data_rom[11599]='h00000000;
    rd_cycle[11600] = 1'b1;  wr_cycle[11600] = 1'b0;  addr_rom[11600]='h00001900;  wr_data_rom[11600]='h00000000;
    rd_cycle[11601] = 1'b1;  wr_cycle[11601] = 1'b0;  addr_rom[11601]='h00001904;  wr_data_rom[11601]='h00000000;
    rd_cycle[11602] = 1'b1;  wr_cycle[11602] = 1'b0;  addr_rom[11602]='h00001908;  wr_data_rom[11602]='h00000000;
    rd_cycle[11603] = 1'b1;  wr_cycle[11603] = 1'b0;  addr_rom[11603]='h0000190c;  wr_data_rom[11603]='h00000000;
    rd_cycle[11604] = 1'b1;  wr_cycle[11604] = 1'b0;  addr_rom[11604]='h00001910;  wr_data_rom[11604]='h00000000;
    rd_cycle[11605] = 1'b1;  wr_cycle[11605] = 1'b0;  addr_rom[11605]='h00001914;  wr_data_rom[11605]='h00000000;
    rd_cycle[11606] = 1'b1;  wr_cycle[11606] = 1'b0;  addr_rom[11606]='h00001918;  wr_data_rom[11606]='h00000000;
    rd_cycle[11607] = 1'b1;  wr_cycle[11607] = 1'b0;  addr_rom[11607]='h0000191c;  wr_data_rom[11607]='h00000000;
    rd_cycle[11608] = 1'b1;  wr_cycle[11608] = 1'b0;  addr_rom[11608]='h00001920;  wr_data_rom[11608]='h00000000;
    rd_cycle[11609] = 1'b1;  wr_cycle[11609] = 1'b0;  addr_rom[11609]='h00001924;  wr_data_rom[11609]='h00000000;
    rd_cycle[11610] = 1'b1;  wr_cycle[11610] = 1'b0;  addr_rom[11610]='h00001928;  wr_data_rom[11610]='h00000000;
    rd_cycle[11611] = 1'b1;  wr_cycle[11611] = 1'b0;  addr_rom[11611]='h0000192c;  wr_data_rom[11611]='h00000000;
    rd_cycle[11612] = 1'b1;  wr_cycle[11612] = 1'b0;  addr_rom[11612]='h00001930;  wr_data_rom[11612]='h00000000;
    rd_cycle[11613] = 1'b1;  wr_cycle[11613] = 1'b0;  addr_rom[11613]='h00001934;  wr_data_rom[11613]='h00000000;
    rd_cycle[11614] = 1'b1;  wr_cycle[11614] = 1'b0;  addr_rom[11614]='h00001938;  wr_data_rom[11614]='h00000000;
    rd_cycle[11615] = 1'b1;  wr_cycle[11615] = 1'b0;  addr_rom[11615]='h0000193c;  wr_data_rom[11615]='h00000000;
    rd_cycle[11616] = 1'b1;  wr_cycle[11616] = 1'b0;  addr_rom[11616]='h00001940;  wr_data_rom[11616]='h00000000;
    rd_cycle[11617] = 1'b1;  wr_cycle[11617] = 1'b0;  addr_rom[11617]='h00001944;  wr_data_rom[11617]='h00000000;
    rd_cycle[11618] = 1'b1;  wr_cycle[11618] = 1'b0;  addr_rom[11618]='h00001948;  wr_data_rom[11618]='h00000000;
    rd_cycle[11619] = 1'b1;  wr_cycle[11619] = 1'b0;  addr_rom[11619]='h0000194c;  wr_data_rom[11619]='h00000000;
    rd_cycle[11620] = 1'b1;  wr_cycle[11620] = 1'b0;  addr_rom[11620]='h00001950;  wr_data_rom[11620]='h00000000;
    rd_cycle[11621] = 1'b1;  wr_cycle[11621] = 1'b0;  addr_rom[11621]='h00001954;  wr_data_rom[11621]='h00000000;
    rd_cycle[11622] = 1'b1;  wr_cycle[11622] = 1'b0;  addr_rom[11622]='h00001958;  wr_data_rom[11622]='h00000000;
    rd_cycle[11623] = 1'b1;  wr_cycle[11623] = 1'b0;  addr_rom[11623]='h0000195c;  wr_data_rom[11623]='h00000000;
    rd_cycle[11624] = 1'b1;  wr_cycle[11624] = 1'b0;  addr_rom[11624]='h00001960;  wr_data_rom[11624]='h00000000;
    rd_cycle[11625] = 1'b1;  wr_cycle[11625] = 1'b0;  addr_rom[11625]='h00001964;  wr_data_rom[11625]='h00000000;
    rd_cycle[11626] = 1'b1;  wr_cycle[11626] = 1'b0;  addr_rom[11626]='h00001968;  wr_data_rom[11626]='h00000000;
    rd_cycle[11627] = 1'b1;  wr_cycle[11627] = 1'b0;  addr_rom[11627]='h0000196c;  wr_data_rom[11627]='h00000000;
    rd_cycle[11628] = 1'b1;  wr_cycle[11628] = 1'b0;  addr_rom[11628]='h00001970;  wr_data_rom[11628]='h00000000;
    rd_cycle[11629] = 1'b1;  wr_cycle[11629] = 1'b0;  addr_rom[11629]='h00001974;  wr_data_rom[11629]='h00000000;
    rd_cycle[11630] = 1'b1;  wr_cycle[11630] = 1'b0;  addr_rom[11630]='h00001978;  wr_data_rom[11630]='h00000000;
    rd_cycle[11631] = 1'b1;  wr_cycle[11631] = 1'b0;  addr_rom[11631]='h0000197c;  wr_data_rom[11631]='h00000000;
    rd_cycle[11632] = 1'b1;  wr_cycle[11632] = 1'b0;  addr_rom[11632]='h00001980;  wr_data_rom[11632]='h00000000;
    rd_cycle[11633] = 1'b1;  wr_cycle[11633] = 1'b0;  addr_rom[11633]='h00001984;  wr_data_rom[11633]='h00000000;
    rd_cycle[11634] = 1'b1;  wr_cycle[11634] = 1'b0;  addr_rom[11634]='h00001988;  wr_data_rom[11634]='h00000000;
    rd_cycle[11635] = 1'b1;  wr_cycle[11635] = 1'b0;  addr_rom[11635]='h0000198c;  wr_data_rom[11635]='h00000000;
    rd_cycle[11636] = 1'b1;  wr_cycle[11636] = 1'b0;  addr_rom[11636]='h00001990;  wr_data_rom[11636]='h00000000;
    rd_cycle[11637] = 1'b1;  wr_cycle[11637] = 1'b0;  addr_rom[11637]='h00001994;  wr_data_rom[11637]='h00000000;
    rd_cycle[11638] = 1'b1;  wr_cycle[11638] = 1'b0;  addr_rom[11638]='h00001998;  wr_data_rom[11638]='h00000000;
    rd_cycle[11639] = 1'b1;  wr_cycle[11639] = 1'b0;  addr_rom[11639]='h0000199c;  wr_data_rom[11639]='h00000000;
    rd_cycle[11640] = 1'b1;  wr_cycle[11640] = 1'b0;  addr_rom[11640]='h000019a0;  wr_data_rom[11640]='h00000000;
    rd_cycle[11641] = 1'b1;  wr_cycle[11641] = 1'b0;  addr_rom[11641]='h000019a4;  wr_data_rom[11641]='h00000000;
    rd_cycle[11642] = 1'b1;  wr_cycle[11642] = 1'b0;  addr_rom[11642]='h000019a8;  wr_data_rom[11642]='h00000000;
    rd_cycle[11643] = 1'b1;  wr_cycle[11643] = 1'b0;  addr_rom[11643]='h000019ac;  wr_data_rom[11643]='h00000000;
    rd_cycle[11644] = 1'b1;  wr_cycle[11644] = 1'b0;  addr_rom[11644]='h000019b0;  wr_data_rom[11644]='h00000000;
    rd_cycle[11645] = 1'b1;  wr_cycle[11645] = 1'b0;  addr_rom[11645]='h000019b4;  wr_data_rom[11645]='h00000000;
    rd_cycle[11646] = 1'b1;  wr_cycle[11646] = 1'b0;  addr_rom[11646]='h000019b8;  wr_data_rom[11646]='h00000000;
    rd_cycle[11647] = 1'b1;  wr_cycle[11647] = 1'b0;  addr_rom[11647]='h000019bc;  wr_data_rom[11647]='h00000000;
    rd_cycle[11648] = 1'b1;  wr_cycle[11648] = 1'b0;  addr_rom[11648]='h000019c0;  wr_data_rom[11648]='h00000000;
    rd_cycle[11649] = 1'b1;  wr_cycle[11649] = 1'b0;  addr_rom[11649]='h000019c4;  wr_data_rom[11649]='h00000000;
    rd_cycle[11650] = 1'b1;  wr_cycle[11650] = 1'b0;  addr_rom[11650]='h000019c8;  wr_data_rom[11650]='h00000000;
    rd_cycle[11651] = 1'b1;  wr_cycle[11651] = 1'b0;  addr_rom[11651]='h000019cc;  wr_data_rom[11651]='h00000000;
    rd_cycle[11652] = 1'b1;  wr_cycle[11652] = 1'b0;  addr_rom[11652]='h000019d0;  wr_data_rom[11652]='h00000000;
    rd_cycle[11653] = 1'b1;  wr_cycle[11653] = 1'b0;  addr_rom[11653]='h000019d4;  wr_data_rom[11653]='h00000000;
    rd_cycle[11654] = 1'b1;  wr_cycle[11654] = 1'b0;  addr_rom[11654]='h000019d8;  wr_data_rom[11654]='h00000000;
    rd_cycle[11655] = 1'b1;  wr_cycle[11655] = 1'b0;  addr_rom[11655]='h000019dc;  wr_data_rom[11655]='h00000000;
    rd_cycle[11656] = 1'b1;  wr_cycle[11656] = 1'b0;  addr_rom[11656]='h000019e0;  wr_data_rom[11656]='h00000000;
    rd_cycle[11657] = 1'b1;  wr_cycle[11657] = 1'b0;  addr_rom[11657]='h000019e4;  wr_data_rom[11657]='h00000000;
    rd_cycle[11658] = 1'b1;  wr_cycle[11658] = 1'b0;  addr_rom[11658]='h000019e8;  wr_data_rom[11658]='h00000000;
    rd_cycle[11659] = 1'b1;  wr_cycle[11659] = 1'b0;  addr_rom[11659]='h000019ec;  wr_data_rom[11659]='h00000000;
    rd_cycle[11660] = 1'b1;  wr_cycle[11660] = 1'b0;  addr_rom[11660]='h000019f0;  wr_data_rom[11660]='h00000000;
    rd_cycle[11661] = 1'b1;  wr_cycle[11661] = 1'b0;  addr_rom[11661]='h000019f4;  wr_data_rom[11661]='h00000000;
    rd_cycle[11662] = 1'b1;  wr_cycle[11662] = 1'b0;  addr_rom[11662]='h000019f8;  wr_data_rom[11662]='h00000000;
    rd_cycle[11663] = 1'b1;  wr_cycle[11663] = 1'b0;  addr_rom[11663]='h000019fc;  wr_data_rom[11663]='h00000000;
    rd_cycle[11664] = 1'b1;  wr_cycle[11664] = 1'b0;  addr_rom[11664]='h00001a00;  wr_data_rom[11664]='h00000000;
    rd_cycle[11665] = 1'b1;  wr_cycle[11665] = 1'b0;  addr_rom[11665]='h00001a04;  wr_data_rom[11665]='h00000000;
    rd_cycle[11666] = 1'b1;  wr_cycle[11666] = 1'b0;  addr_rom[11666]='h00001a08;  wr_data_rom[11666]='h00000000;
    rd_cycle[11667] = 1'b1;  wr_cycle[11667] = 1'b0;  addr_rom[11667]='h00001a0c;  wr_data_rom[11667]='h00000000;
    rd_cycle[11668] = 1'b1;  wr_cycle[11668] = 1'b0;  addr_rom[11668]='h00001a10;  wr_data_rom[11668]='h00000000;
    rd_cycle[11669] = 1'b1;  wr_cycle[11669] = 1'b0;  addr_rom[11669]='h00001a14;  wr_data_rom[11669]='h00000000;
    rd_cycle[11670] = 1'b1;  wr_cycle[11670] = 1'b0;  addr_rom[11670]='h00001a18;  wr_data_rom[11670]='h00000000;
    rd_cycle[11671] = 1'b1;  wr_cycle[11671] = 1'b0;  addr_rom[11671]='h00001a1c;  wr_data_rom[11671]='h00000000;
    rd_cycle[11672] = 1'b1;  wr_cycle[11672] = 1'b0;  addr_rom[11672]='h00001a20;  wr_data_rom[11672]='h00000000;
    rd_cycle[11673] = 1'b1;  wr_cycle[11673] = 1'b0;  addr_rom[11673]='h00001a24;  wr_data_rom[11673]='h00000000;
    rd_cycle[11674] = 1'b1;  wr_cycle[11674] = 1'b0;  addr_rom[11674]='h00001a28;  wr_data_rom[11674]='h00000000;
    rd_cycle[11675] = 1'b1;  wr_cycle[11675] = 1'b0;  addr_rom[11675]='h00001a2c;  wr_data_rom[11675]='h00000000;
    rd_cycle[11676] = 1'b1;  wr_cycle[11676] = 1'b0;  addr_rom[11676]='h00001a30;  wr_data_rom[11676]='h00000000;
    rd_cycle[11677] = 1'b1;  wr_cycle[11677] = 1'b0;  addr_rom[11677]='h00001a34;  wr_data_rom[11677]='h00000000;
    rd_cycle[11678] = 1'b1;  wr_cycle[11678] = 1'b0;  addr_rom[11678]='h00001a38;  wr_data_rom[11678]='h00000000;
    rd_cycle[11679] = 1'b1;  wr_cycle[11679] = 1'b0;  addr_rom[11679]='h00001a3c;  wr_data_rom[11679]='h00000000;
    rd_cycle[11680] = 1'b1;  wr_cycle[11680] = 1'b0;  addr_rom[11680]='h00001a40;  wr_data_rom[11680]='h00000000;
    rd_cycle[11681] = 1'b1;  wr_cycle[11681] = 1'b0;  addr_rom[11681]='h00001a44;  wr_data_rom[11681]='h00000000;
    rd_cycle[11682] = 1'b1;  wr_cycle[11682] = 1'b0;  addr_rom[11682]='h00001a48;  wr_data_rom[11682]='h00000000;
    rd_cycle[11683] = 1'b1;  wr_cycle[11683] = 1'b0;  addr_rom[11683]='h00001a4c;  wr_data_rom[11683]='h00000000;
    rd_cycle[11684] = 1'b1;  wr_cycle[11684] = 1'b0;  addr_rom[11684]='h00001a50;  wr_data_rom[11684]='h00000000;
    rd_cycle[11685] = 1'b1;  wr_cycle[11685] = 1'b0;  addr_rom[11685]='h00001a54;  wr_data_rom[11685]='h00000000;
    rd_cycle[11686] = 1'b1;  wr_cycle[11686] = 1'b0;  addr_rom[11686]='h00001a58;  wr_data_rom[11686]='h00000000;
    rd_cycle[11687] = 1'b1;  wr_cycle[11687] = 1'b0;  addr_rom[11687]='h00001a5c;  wr_data_rom[11687]='h00000000;
    rd_cycle[11688] = 1'b1;  wr_cycle[11688] = 1'b0;  addr_rom[11688]='h00001a60;  wr_data_rom[11688]='h00000000;
    rd_cycle[11689] = 1'b1;  wr_cycle[11689] = 1'b0;  addr_rom[11689]='h00001a64;  wr_data_rom[11689]='h00000000;
    rd_cycle[11690] = 1'b1;  wr_cycle[11690] = 1'b0;  addr_rom[11690]='h00001a68;  wr_data_rom[11690]='h00000000;
    rd_cycle[11691] = 1'b1;  wr_cycle[11691] = 1'b0;  addr_rom[11691]='h00001a6c;  wr_data_rom[11691]='h00000000;
    rd_cycle[11692] = 1'b1;  wr_cycle[11692] = 1'b0;  addr_rom[11692]='h00001a70;  wr_data_rom[11692]='h00000000;
    rd_cycle[11693] = 1'b1;  wr_cycle[11693] = 1'b0;  addr_rom[11693]='h00001a74;  wr_data_rom[11693]='h00000000;
    rd_cycle[11694] = 1'b1;  wr_cycle[11694] = 1'b0;  addr_rom[11694]='h00001a78;  wr_data_rom[11694]='h00000000;
    rd_cycle[11695] = 1'b1;  wr_cycle[11695] = 1'b0;  addr_rom[11695]='h00001a7c;  wr_data_rom[11695]='h00000000;
    rd_cycle[11696] = 1'b1;  wr_cycle[11696] = 1'b0;  addr_rom[11696]='h00001a80;  wr_data_rom[11696]='h00000000;
    rd_cycle[11697] = 1'b1;  wr_cycle[11697] = 1'b0;  addr_rom[11697]='h00001a84;  wr_data_rom[11697]='h00000000;
    rd_cycle[11698] = 1'b1;  wr_cycle[11698] = 1'b0;  addr_rom[11698]='h00001a88;  wr_data_rom[11698]='h00000000;
    rd_cycle[11699] = 1'b1;  wr_cycle[11699] = 1'b0;  addr_rom[11699]='h00001a8c;  wr_data_rom[11699]='h00000000;
    rd_cycle[11700] = 1'b1;  wr_cycle[11700] = 1'b0;  addr_rom[11700]='h00001a90;  wr_data_rom[11700]='h00000000;
    rd_cycle[11701] = 1'b1;  wr_cycle[11701] = 1'b0;  addr_rom[11701]='h00001a94;  wr_data_rom[11701]='h00000000;
    rd_cycle[11702] = 1'b1;  wr_cycle[11702] = 1'b0;  addr_rom[11702]='h00001a98;  wr_data_rom[11702]='h00000000;
    rd_cycle[11703] = 1'b1;  wr_cycle[11703] = 1'b0;  addr_rom[11703]='h00001a9c;  wr_data_rom[11703]='h00000000;
    rd_cycle[11704] = 1'b1;  wr_cycle[11704] = 1'b0;  addr_rom[11704]='h00001aa0;  wr_data_rom[11704]='h00000000;
    rd_cycle[11705] = 1'b1;  wr_cycle[11705] = 1'b0;  addr_rom[11705]='h00001aa4;  wr_data_rom[11705]='h00000000;
    rd_cycle[11706] = 1'b1;  wr_cycle[11706] = 1'b0;  addr_rom[11706]='h00001aa8;  wr_data_rom[11706]='h00000000;
    rd_cycle[11707] = 1'b1;  wr_cycle[11707] = 1'b0;  addr_rom[11707]='h00001aac;  wr_data_rom[11707]='h00000000;
    rd_cycle[11708] = 1'b1;  wr_cycle[11708] = 1'b0;  addr_rom[11708]='h00001ab0;  wr_data_rom[11708]='h00000000;
    rd_cycle[11709] = 1'b1;  wr_cycle[11709] = 1'b0;  addr_rom[11709]='h00001ab4;  wr_data_rom[11709]='h00000000;
    rd_cycle[11710] = 1'b1;  wr_cycle[11710] = 1'b0;  addr_rom[11710]='h00001ab8;  wr_data_rom[11710]='h00000000;
    rd_cycle[11711] = 1'b1;  wr_cycle[11711] = 1'b0;  addr_rom[11711]='h00001abc;  wr_data_rom[11711]='h00000000;
    rd_cycle[11712] = 1'b1;  wr_cycle[11712] = 1'b0;  addr_rom[11712]='h00001ac0;  wr_data_rom[11712]='h00000000;
    rd_cycle[11713] = 1'b1;  wr_cycle[11713] = 1'b0;  addr_rom[11713]='h00001ac4;  wr_data_rom[11713]='h00000000;
    rd_cycle[11714] = 1'b1;  wr_cycle[11714] = 1'b0;  addr_rom[11714]='h00001ac8;  wr_data_rom[11714]='h00000000;
    rd_cycle[11715] = 1'b1;  wr_cycle[11715] = 1'b0;  addr_rom[11715]='h00001acc;  wr_data_rom[11715]='h00000000;
    rd_cycle[11716] = 1'b1;  wr_cycle[11716] = 1'b0;  addr_rom[11716]='h00001ad0;  wr_data_rom[11716]='h00000000;
    rd_cycle[11717] = 1'b1;  wr_cycle[11717] = 1'b0;  addr_rom[11717]='h00001ad4;  wr_data_rom[11717]='h00000000;
    rd_cycle[11718] = 1'b1;  wr_cycle[11718] = 1'b0;  addr_rom[11718]='h00001ad8;  wr_data_rom[11718]='h00000000;
    rd_cycle[11719] = 1'b1;  wr_cycle[11719] = 1'b0;  addr_rom[11719]='h00001adc;  wr_data_rom[11719]='h00000000;
    rd_cycle[11720] = 1'b1;  wr_cycle[11720] = 1'b0;  addr_rom[11720]='h00001ae0;  wr_data_rom[11720]='h00000000;
    rd_cycle[11721] = 1'b1;  wr_cycle[11721] = 1'b0;  addr_rom[11721]='h00001ae4;  wr_data_rom[11721]='h00000000;
    rd_cycle[11722] = 1'b1;  wr_cycle[11722] = 1'b0;  addr_rom[11722]='h00001ae8;  wr_data_rom[11722]='h00000000;
    rd_cycle[11723] = 1'b1;  wr_cycle[11723] = 1'b0;  addr_rom[11723]='h00001aec;  wr_data_rom[11723]='h00000000;
    rd_cycle[11724] = 1'b1;  wr_cycle[11724] = 1'b0;  addr_rom[11724]='h00001af0;  wr_data_rom[11724]='h00000000;
    rd_cycle[11725] = 1'b1;  wr_cycle[11725] = 1'b0;  addr_rom[11725]='h00001af4;  wr_data_rom[11725]='h00000000;
    rd_cycle[11726] = 1'b1;  wr_cycle[11726] = 1'b0;  addr_rom[11726]='h00001af8;  wr_data_rom[11726]='h00000000;
    rd_cycle[11727] = 1'b1;  wr_cycle[11727] = 1'b0;  addr_rom[11727]='h00001afc;  wr_data_rom[11727]='h00000000;
    rd_cycle[11728] = 1'b1;  wr_cycle[11728] = 1'b0;  addr_rom[11728]='h00001b00;  wr_data_rom[11728]='h00000000;
    rd_cycle[11729] = 1'b1;  wr_cycle[11729] = 1'b0;  addr_rom[11729]='h00001b04;  wr_data_rom[11729]='h00000000;
    rd_cycle[11730] = 1'b1;  wr_cycle[11730] = 1'b0;  addr_rom[11730]='h00001b08;  wr_data_rom[11730]='h00000000;
    rd_cycle[11731] = 1'b1;  wr_cycle[11731] = 1'b0;  addr_rom[11731]='h00001b0c;  wr_data_rom[11731]='h00000000;
    rd_cycle[11732] = 1'b1;  wr_cycle[11732] = 1'b0;  addr_rom[11732]='h00001b10;  wr_data_rom[11732]='h00000000;
    rd_cycle[11733] = 1'b1;  wr_cycle[11733] = 1'b0;  addr_rom[11733]='h00001b14;  wr_data_rom[11733]='h00000000;
    rd_cycle[11734] = 1'b1;  wr_cycle[11734] = 1'b0;  addr_rom[11734]='h00001b18;  wr_data_rom[11734]='h00000000;
    rd_cycle[11735] = 1'b1;  wr_cycle[11735] = 1'b0;  addr_rom[11735]='h00001b1c;  wr_data_rom[11735]='h00000000;
    rd_cycle[11736] = 1'b1;  wr_cycle[11736] = 1'b0;  addr_rom[11736]='h00001b20;  wr_data_rom[11736]='h00000000;
    rd_cycle[11737] = 1'b1;  wr_cycle[11737] = 1'b0;  addr_rom[11737]='h00001b24;  wr_data_rom[11737]='h00000000;
    rd_cycle[11738] = 1'b1;  wr_cycle[11738] = 1'b0;  addr_rom[11738]='h00001b28;  wr_data_rom[11738]='h00000000;
    rd_cycle[11739] = 1'b1;  wr_cycle[11739] = 1'b0;  addr_rom[11739]='h00001b2c;  wr_data_rom[11739]='h00000000;
    rd_cycle[11740] = 1'b1;  wr_cycle[11740] = 1'b0;  addr_rom[11740]='h00001b30;  wr_data_rom[11740]='h00000000;
    rd_cycle[11741] = 1'b1;  wr_cycle[11741] = 1'b0;  addr_rom[11741]='h00001b34;  wr_data_rom[11741]='h00000000;
    rd_cycle[11742] = 1'b1;  wr_cycle[11742] = 1'b0;  addr_rom[11742]='h00001b38;  wr_data_rom[11742]='h00000000;
    rd_cycle[11743] = 1'b1;  wr_cycle[11743] = 1'b0;  addr_rom[11743]='h00001b3c;  wr_data_rom[11743]='h00000000;
    rd_cycle[11744] = 1'b1;  wr_cycle[11744] = 1'b0;  addr_rom[11744]='h00001b40;  wr_data_rom[11744]='h00000000;
    rd_cycle[11745] = 1'b1;  wr_cycle[11745] = 1'b0;  addr_rom[11745]='h00001b44;  wr_data_rom[11745]='h00000000;
    rd_cycle[11746] = 1'b1;  wr_cycle[11746] = 1'b0;  addr_rom[11746]='h00001b48;  wr_data_rom[11746]='h00000000;
    rd_cycle[11747] = 1'b1;  wr_cycle[11747] = 1'b0;  addr_rom[11747]='h00001b4c;  wr_data_rom[11747]='h00000000;
    rd_cycle[11748] = 1'b1;  wr_cycle[11748] = 1'b0;  addr_rom[11748]='h00001b50;  wr_data_rom[11748]='h00000000;
    rd_cycle[11749] = 1'b1;  wr_cycle[11749] = 1'b0;  addr_rom[11749]='h00001b54;  wr_data_rom[11749]='h00000000;
    rd_cycle[11750] = 1'b1;  wr_cycle[11750] = 1'b0;  addr_rom[11750]='h00001b58;  wr_data_rom[11750]='h00000000;
    rd_cycle[11751] = 1'b1;  wr_cycle[11751] = 1'b0;  addr_rom[11751]='h00001b5c;  wr_data_rom[11751]='h00000000;
    rd_cycle[11752] = 1'b1;  wr_cycle[11752] = 1'b0;  addr_rom[11752]='h00001b60;  wr_data_rom[11752]='h00000000;
    rd_cycle[11753] = 1'b1;  wr_cycle[11753] = 1'b0;  addr_rom[11753]='h00001b64;  wr_data_rom[11753]='h00000000;
    rd_cycle[11754] = 1'b1;  wr_cycle[11754] = 1'b0;  addr_rom[11754]='h00001b68;  wr_data_rom[11754]='h00000000;
    rd_cycle[11755] = 1'b1;  wr_cycle[11755] = 1'b0;  addr_rom[11755]='h00001b6c;  wr_data_rom[11755]='h00000000;
    rd_cycle[11756] = 1'b1;  wr_cycle[11756] = 1'b0;  addr_rom[11756]='h00001b70;  wr_data_rom[11756]='h00000000;
    rd_cycle[11757] = 1'b1;  wr_cycle[11757] = 1'b0;  addr_rom[11757]='h00001b74;  wr_data_rom[11757]='h00000000;
    rd_cycle[11758] = 1'b1;  wr_cycle[11758] = 1'b0;  addr_rom[11758]='h00001b78;  wr_data_rom[11758]='h00000000;
    rd_cycle[11759] = 1'b1;  wr_cycle[11759] = 1'b0;  addr_rom[11759]='h00001b7c;  wr_data_rom[11759]='h00000000;
    rd_cycle[11760] = 1'b1;  wr_cycle[11760] = 1'b0;  addr_rom[11760]='h00001b80;  wr_data_rom[11760]='h00000000;
    rd_cycle[11761] = 1'b1;  wr_cycle[11761] = 1'b0;  addr_rom[11761]='h00001b84;  wr_data_rom[11761]='h00000000;
    rd_cycle[11762] = 1'b1;  wr_cycle[11762] = 1'b0;  addr_rom[11762]='h00001b88;  wr_data_rom[11762]='h00000000;
    rd_cycle[11763] = 1'b1;  wr_cycle[11763] = 1'b0;  addr_rom[11763]='h00001b8c;  wr_data_rom[11763]='h00000000;
    rd_cycle[11764] = 1'b1;  wr_cycle[11764] = 1'b0;  addr_rom[11764]='h00001b90;  wr_data_rom[11764]='h00000000;
    rd_cycle[11765] = 1'b1;  wr_cycle[11765] = 1'b0;  addr_rom[11765]='h00001b94;  wr_data_rom[11765]='h00000000;
    rd_cycle[11766] = 1'b1;  wr_cycle[11766] = 1'b0;  addr_rom[11766]='h00001b98;  wr_data_rom[11766]='h00000000;
    rd_cycle[11767] = 1'b1;  wr_cycle[11767] = 1'b0;  addr_rom[11767]='h00001b9c;  wr_data_rom[11767]='h00000000;
    rd_cycle[11768] = 1'b1;  wr_cycle[11768] = 1'b0;  addr_rom[11768]='h00001ba0;  wr_data_rom[11768]='h00000000;
    rd_cycle[11769] = 1'b1;  wr_cycle[11769] = 1'b0;  addr_rom[11769]='h00001ba4;  wr_data_rom[11769]='h00000000;
    rd_cycle[11770] = 1'b1;  wr_cycle[11770] = 1'b0;  addr_rom[11770]='h00001ba8;  wr_data_rom[11770]='h00000000;
    rd_cycle[11771] = 1'b1;  wr_cycle[11771] = 1'b0;  addr_rom[11771]='h00001bac;  wr_data_rom[11771]='h00000000;
    rd_cycle[11772] = 1'b1;  wr_cycle[11772] = 1'b0;  addr_rom[11772]='h00001bb0;  wr_data_rom[11772]='h00000000;
    rd_cycle[11773] = 1'b1;  wr_cycle[11773] = 1'b0;  addr_rom[11773]='h00001bb4;  wr_data_rom[11773]='h00000000;
    rd_cycle[11774] = 1'b1;  wr_cycle[11774] = 1'b0;  addr_rom[11774]='h00001bb8;  wr_data_rom[11774]='h00000000;
    rd_cycle[11775] = 1'b1;  wr_cycle[11775] = 1'b0;  addr_rom[11775]='h00001bbc;  wr_data_rom[11775]='h00000000;
    rd_cycle[11776] = 1'b1;  wr_cycle[11776] = 1'b0;  addr_rom[11776]='h00001bc0;  wr_data_rom[11776]='h00000000;
    rd_cycle[11777] = 1'b1;  wr_cycle[11777] = 1'b0;  addr_rom[11777]='h00001bc4;  wr_data_rom[11777]='h00000000;
    rd_cycle[11778] = 1'b1;  wr_cycle[11778] = 1'b0;  addr_rom[11778]='h00001bc8;  wr_data_rom[11778]='h00000000;
    rd_cycle[11779] = 1'b1;  wr_cycle[11779] = 1'b0;  addr_rom[11779]='h00001bcc;  wr_data_rom[11779]='h00000000;
    rd_cycle[11780] = 1'b1;  wr_cycle[11780] = 1'b0;  addr_rom[11780]='h00001bd0;  wr_data_rom[11780]='h00000000;
    rd_cycle[11781] = 1'b1;  wr_cycle[11781] = 1'b0;  addr_rom[11781]='h00001bd4;  wr_data_rom[11781]='h00000000;
    rd_cycle[11782] = 1'b1;  wr_cycle[11782] = 1'b0;  addr_rom[11782]='h00001bd8;  wr_data_rom[11782]='h00000000;
    rd_cycle[11783] = 1'b1;  wr_cycle[11783] = 1'b0;  addr_rom[11783]='h00001bdc;  wr_data_rom[11783]='h00000000;
    rd_cycle[11784] = 1'b1;  wr_cycle[11784] = 1'b0;  addr_rom[11784]='h00001be0;  wr_data_rom[11784]='h00000000;
    rd_cycle[11785] = 1'b1;  wr_cycle[11785] = 1'b0;  addr_rom[11785]='h00001be4;  wr_data_rom[11785]='h00000000;
    rd_cycle[11786] = 1'b1;  wr_cycle[11786] = 1'b0;  addr_rom[11786]='h00001be8;  wr_data_rom[11786]='h00000000;
    rd_cycle[11787] = 1'b1;  wr_cycle[11787] = 1'b0;  addr_rom[11787]='h00001bec;  wr_data_rom[11787]='h00000000;
    rd_cycle[11788] = 1'b1;  wr_cycle[11788] = 1'b0;  addr_rom[11788]='h00001bf0;  wr_data_rom[11788]='h00000000;
    rd_cycle[11789] = 1'b1;  wr_cycle[11789] = 1'b0;  addr_rom[11789]='h00001bf4;  wr_data_rom[11789]='h00000000;
    rd_cycle[11790] = 1'b1;  wr_cycle[11790] = 1'b0;  addr_rom[11790]='h00001bf8;  wr_data_rom[11790]='h00000000;
    rd_cycle[11791] = 1'b1;  wr_cycle[11791] = 1'b0;  addr_rom[11791]='h00001bfc;  wr_data_rom[11791]='h00000000;
    rd_cycle[11792] = 1'b1;  wr_cycle[11792] = 1'b0;  addr_rom[11792]='h00001c00;  wr_data_rom[11792]='h00000000;
    rd_cycle[11793] = 1'b1;  wr_cycle[11793] = 1'b0;  addr_rom[11793]='h00001c04;  wr_data_rom[11793]='h00000000;
    rd_cycle[11794] = 1'b1;  wr_cycle[11794] = 1'b0;  addr_rom[11794]='h00001c08;  wr_data_rom[11794]='h00000000;
    rd_cycle[11795] = 1'b1;  wr_cycle[11795] = 1'b0;  addr_rom[11795]='h00001c0c;  wr_data_rom[11795]='h00000000;
    rd_cycle[11796] = 1'b1;  wr_cycle[11796] = 1'b0;  addr_rom[11796]='h00001c10;  wr_data_rom[11796]='h00000000;
    rd_cycle[11797] = 1'b1;  wr_cycle[11797] = 1'b0;  addr_rom[11797]='h00001c14;  wr_data_rom[11797]='h00000000;
    rd_cycle[11798] = 1'b1;  wr_cycle[11798] = 1'b0;  addr_rom[11798]='h00001c18;  wr_data_rom[11798]='h00000000;
    rd_cycle[11799] = 1'b1;  wr_cycle[11799] = 1'b0;  addr_rom[11799]='h00001c1c;  wr_data_rom[11799]='h00000000;
    rd_cycle[11800] = 1'b1;  wr_cycle[11800] = 1'b0;  addr_rom[11800]='h00001c20;  wr_data_rom[11800]='h00000000;
    rd_cycle[11801] = 1'b1;  wr_cycle[11801] = 1'b0;  addr_rom[11801]='h00001c24;  wr_data_rom[11801]='h00000000;
    rd_cycle[11802] = 1'b1;  wr_cycle[11802] = 1'b0;  addr_rom[11802]='h00001c28;  wr_data_rom[11802]='h00000000;
    rd_cycle[11803] = 1'b1;  wr_cycle[11803] = 1'b0;  addr_rom[11803]='h00001c2c;  wr_data_rom[11803]='h00000000;
    rd_cycle[11804] = 1'b1;  wr_cycle[11804] = 1'b0;  addr_rom[11804]='h00001c30;  wr_data_rom[11804]='h00000000;
    rd_cycle[11805] = 1'b1;  wr_cycle[11805] = 1'b0;  addr_rom[11805]='h00001c34;  wr_data_rom[11805]='h00000000;
    rd_cycle[11806] = 1'b1;  wr_cycle[11806] = 1'b0;  addr_rom[11806]='h00001c38;  wr_data_rom[11806]='h00000000;
    rd_cycle[11807] = 1'b1;  wr_cycle[11807] = 1'b0;  addr_rom[11807]='h00001c3c;  wr_data_rom[11807]='h00000000;
    rd_cycle[11808] = 1'b1;  wr_cycle[11808] = 1'b0;  addr_rom[11808]='h00001c40;  wr_data_rom[11808]='h00000000;
    rd_cycle[11809] = 1'b1;  wr_cycle[11809] = 1'b0;  addr_rom[11809]='h00001c44;  wr_data_rom[11809]='h00000000;
    rd_cycle[11810] = 1'b1;  wr_cycle[11810] = 1'b0;  addr_rom[11810]='h00001c48;  wr_data_rom[11810]='h00000000;
    rd_cycle[11811] = 1'b1;  wr_cycle[11811] = 1'b0;  addr_rom[11811]='h00001c4c;  wr_data_rom[11811]='h00000000;
    rd_cycle[11812] = 1'b1;  wr_cycle[11812] = 1'b0;  addr_rom[11812]='h00001c50;  wr_data_rom[11812]='h00000000;
    rd_cycle[11813] = 1'b1;  wr_cycle[11813] = 1'b0;  addr_rom[11813]='h00001c54;  wr_data_rom[11813]='h00000000;
    rd_cycle[11814] = 1'b1;  wr_cycle[11814] = 1'b0;  addr_rom[11814]='h00001c58;  wr_data_rom[11814]='h00000000;
    rd_cycle[11815] = 1'b1;  wr_cycle[11815] = 1'b0;  addr_rom[11815]='h00001c5c;  wr_data_rom[11815]='h00000000;
    rd_cycle[11816] = 1'b1;  wr_cycle[11816] = 1'b0;  addr_rom[11816]='h00001c60;  wr_data_rom[11816]='h00000000;
    rd_cycle[11817] = 1'b1;  wr_cycle[11817] = 1'b0;  addr_rom[11817]='h00001c64;  wr_data_rom[11817]='h00000000;
    rd_cycle[11818] = 1'b1;  wr_cycle[11818] = 1'b0;  addr_rom[11818]='h00001c68;  wr_data_rom[11818]='h00000000;
    rd_cycle[11819] = 1'b1;  wr_cycle[11819] = 1'b0;  addr_rom[11819]='h00001c6c;  wr_data_rom[11819]='h00000000;
    rd_cycle[11820] = 1'b1;  wr_cycle[11820] = 1'b0;  addr_rom[11820]='h00001c70;  wr_data_rom[11820]='h00000000;
    rd_cycle[11821] = 1'b1;  wr_cycle[11821] = 1'b0;  addr_rom[11821]='h00001c74;  wr_data_rom[11821]='h00000000;
    rd_cycle[11822] = 1'b1;  wr_cycle[11822] = 1'b0;  addr_rom[11822]='h00001c78;  wr_data_rom[11822]='h00000000;
    rd_cycle[11823] = 1'b1;  wr_cycle[11823] = 1'b0;  addr_rom[11823]='h00001c7c;  wr_data_rom[11823]='h00000000;
    rd_cycle[11824] = 1'b1;  wr_cycle[11824] = 1'b0;  addr_rom[11824]='h00001c80;  wr_data_rom[11824]='h00000000;
    rd_cycle[11825] = 1'b1;  wr_cycle[11825] = 1'b0;  addr_rom[11825]='h00001c84;  wr_data_rom[11825]='h00000000;
    rd_cycle[11826] = 1'b1;  wr_cycle[11826] = 1'b0;  addr_rom[11826]='h00001c88;  wr_data_rom[11826]='h00000000;
    rd_cycle[11827] = 1'b1;  wr_cycle[11827] = 1'b0;  addr_rom[11827]='h00001c8c;  wr_data_rom[11827]='h00000000;
    rd_cycle[11828] = 1'b1;  wr_cycle[11828] = 1'b0;  addr_rom[11828]='h00001c90;  wr_data_rom[11828]='h00000000;
    rd_cycle[11829] = 1'b1;  wr_cycle[11829] = 1'b0;  addr_rom[11829]='h00001c94;  wr_data_rom[11829]='h00000000;
    rd_cycle[11830] = 1'b1;  wr_cycle[11830] = 1'b0;  addr_rom[11830]='h00001c98;  wr_data_rom[11830]='h00000000;
    rd_cycle[11831] = 1'b1;  wr_cycle[11831] = 1'b0;  addr_rom[11831]='h00001c9c;  wr_data_rom[11831]='h00000000;
    rd_cycle[11832] = 1'b1;  wr_cycle[11832] = 1'b0;  addr_rom[11832]='h00001ca0;  wr_data_rom[11832]='h00000000;
    rd_cycle[11833] = 1'b1;  wr_cycle[11833] = 1'b0;  addr_rom[11833]='h00001ca4;  wr_data_rom[11833]='h00000000;
    rd_cycle[11834] = 1'b1;  wr_cycle[11834] = 1'b0;  addr_rom[11834]='h00001ca8;  wr_data_rom[11834]='h00000000;
    rd_cycle[11835] = 1'b1;  wr_cycle[11835] = 1'b0;  addr_rom[11835]='h00001cac;  wr_data_rom[11835]='h00000000;
    rd_cycle[11836] = 1'b1;  wr_cycle[11836] = 1'b0;  addr_rom[11836]='h00001cb0;  wr_data_rom[11836]='h00000000;
    rd_cycle[11837] = 1'b1;  wr_cycle[11837] = 1'b0;  addr_rom[11837]='h00001cb4;  wr_data_rom[11837]='h00000000;
    rd_cycle[11838] = 1'b1;  wr_cycle[11838] = 1'b0;  addr_rom[11838]='h00001cb8;  wr_data_rom[11838]='h00000000;
    rd_cycle[11839] = 1'b1;  wr_cycle[11839] = 1'b0;  addr_rom[11839]='h00001cbc;  wr_data_rom[11839]='h00000000;
    rd_cycle[11840] = 1'b1;  wr_cycle[11840] = 1'b0;  addr_rom[11840]='h00001cc0;  wr_data_rom[11840]='h00000000;
    rd_cycle[11841] = 1'b1;  wr_cycle[11841] = 1'b0;  addr_rom[11841]='h00001cc4;  wr_data_rom[11841]='h00000000;
    rd_cycle[11842] = 1'b1;  wr_cycle[11842] = 1'b0;  addr_rom[11842]='h00001cc8;  wr_data_rom[11842]='h00000000;
    rd_cycle[11843] = 1'b1;  wr_cycle[11843] = 1'b0;  addr_rom[11843]='h00001ccc;  wr_data_rom[11843]='h00000000;
    rd_cycle[11844] = 1'b1;  wr_cycle[11844] = 1'b0;  addr_rom[11844]='h00001cd0;  wr_data_rom[11844]='h00000000;
    rd_cycle[11845] = 1'b1;  wr_cycle[11845] = 1'b0;  addr_rom[11845]='h00001cd4;  wr_data_rom[11845]='h00000000;
    rd_cycle[11846] = 1'b1;  wr_cycle[11846] = 1'b0;  addr_rom[11846]='h00001cd8;  wr_data_rom[11846]='h00000000;
    rd_cycle[11847] = 1'b1;  wr_cycle[11847] = 1'b0;  addr_rom[11847]='h00001cdc;  wr_data_rom[11847]='h00000000;
    rd_cycle[11848] = 1'b1;  wr_cycle[11848] = 1'b0;  addr_rom[11848]='h00001ce0;  wr_data_rom[11848]='h00000000;
    rd_cycle[11849] = 1'b1;  wr_cycle[11849] = 1'b0;  addr_rom[11849]='h00001ce4;  wr_data_rom[11849]='h00000000;
    rd_cycle[11850] = 1'b1;  wr_cycle[11850] = 1'b0;  addr_rom[11850]='h00001ce8;  wr_data_rom[11850]='h00000000;
    rd_cycle[11851] = 1'b1;  wr_cycle[11851] = 1'b0;  addr_rom[11851]='h00001cec;  wr_data_rom[11851]='h00000000;
    rd_cycle[11852] = 1'b1;  wr_cycle[11852] = 1'b0;  addr_rom[11852]='h00001cf0;  wr_data_rom[11852]='h00000000;
    rd_cycle[11853] = 1'b1;  wr_cycle[11853] = 1'b0;  addr_rom[11853]='h00001cf4;  wr_data_rom[11853]='h00000000;
    rd_cycle[11854] = 1'b1;  wr_cycle[11854] = 1'b0;  addr_rom[11854]='h00001cf8;  wr_data_rom[11854]='h00000000;
    rd_cycle[11855] = 1'b1;  wr_cycle[11855] = 1'b0;  addr_rom[11855]='h00001cfc;  wr_data_rom[11855]='h00000000;
    rd_cycle[11856] = 1'b1;  wr_cycle[11856] = 1'b0;  addr_rom[11856]='h00001d00;  wr_data_rom[11856]='h00000000;
    rd_cycle[11857] = 1'b1;  wr_cycle[11857] = 1'b0;  addr_rom[11857]='h00001d04;  wr_data_rom[11857]='h00000000;
    rd_cycle[11858] = 1'b1;  wr_cycle[11858] = 1'b0;  addr_rom[11858]='h00001d08;  wr_data_rom[11858]='h00000000;
    rd_cycle[11859] = 1'b1;  wr_cycle[11859] = 1'b0;  addr_rom[11859]='h00001d0c;  wr_data_rom[11859]='h00000000;
    rd_cycle[11860] = 1'b1;  wr_cycle[11860] = 1'b0;  addr_rom[11860]='h00001d10;  wr_data_rom[11860]='h00000000;
    rd_cycle[11861] = 1'b1;  wr_cycle[11861] = 1'b0;  addr_rom[11861]='h00001d14;  wr_data_rom[11861]='h00000000;
    rd_cycle[11862] = 1'b1;  wr_cycle[11862] = 1'b0;  addr_rom[11862]='h00001d18;  wr_data_rom[11862]='h00000000;
    rd_cycle[11863] = 1'b1;  wr_cycle[11863] = 1'b0;  addr_rom[11863]='h00001d1c;  wr_data_rom[11863]='h00000000;
    rd_cycle[11864] = 1'b1;  wr_cycle[11864] = 1'b0;  addr_rom[11864]='h00001d20;  wr_data_rom[11864]='h00000000;
    rd_cycle[11865] = 1'b1;  wr_cycle[11865] = 1'b0;  addr_rom[11865]='h00001d24;  wr_data_rom[11865]='h00000000;
    rd_cycle[11866] = 1'b1;  wr_cycle[11866] = 1'b0;  addr_rom[11866]='h00001d28;  wr_data_rom[11866]='h00000000;
    rd_cycle[11867] = 1'b1;  wr_cycle[11867] = 1'b0;  addr_rom[11867]='h00001d2c;  wr_data_rom[11867]='h00000000;
    rd_cycle[11868] = 1'b1;  wr_cycle[11868] = 1'b0;  addr_rom[11868]='h00001d30;  wr_data_rom[11868]='h00000000;
    rd_cycle[11869] = 1'b1;  wr_cycle[11869] = 1'b0;  addr_rom[11869]='h00001d34;  wr_data_rom[11869]='h00000000;
    rd_cycle[11870] = 1'b1;  wr_cycle[11870] = 1'b0;  addr_rom[11870]='h00001d38;  wr_data_rom[11870]='h00000000;
    rd_cycle[11871] = 1'b1;  wr_cycle[11871] = 1'b0;  addr_rom[11871]='h00001d3c;  wr_data_rom[11871]='h00000000;
    rd_cycle[11872] = 1'b1;  wr_cycle[11872] = 1'b0;  addr_rom[11872]='h00001d40;  wr_data_rom[11872]='h00000000;
    rd_cycle[11873] = 1'b1;  wr_cycle[11873] = 1'b0;  addr_rom[11873]='h00001d44;  wr_data_rom[11873]='h00000000;
    rd_cycle[11874] = 1'b1;  wr_cycle[11874] = 1'b0;  addr_rom[11874]='h00001d48;  wr_data_rom[11874]='h00000000;
    rd_cycle[11875] = 1'b1;  wr_cycle[11875] = 1'b0;  addr_rom[11875]='h00001d4c;  wr_data_rom[11875]='h00000000;
    rd_cycle[11876] = 1'b1;  wr_cycle[11876] = 1'b0;  addr_rom[11876]='h00001d50;  wr_data_rom[11876]='h00000000;
    rd_cycle[11877] = 1'b1;  wr_cycle[11877] = 1'b0;  addr_rom[11877]='h00001d54;  wr_data_rom[11877]='h00000000;
    rd_cycle[11878] = 1'b1;  wr_cycle[11878] = 1'b0;  addr_rom[11878]='h00001d58;  wr_data_rom[11878]='h00000000;
    rd_cycle[11879] = 1'b1;  wr_cycle[11879] = 1'b0;  addr_rom[11879]='h00001d5c;  wr_data_rom[11879]='h00000000;
    rd_cycle[11880] = 1'b1;  wr_cycle[11880] = 1'b0;  addr_rom[11880]='h00001d60;  wr_data_rom[11880]='h00000000;
    rd_cycle[11881] = 1'b1;  wr_cycle[11881] = 1'b0;  addr_rom[11881]='h00001d64;  wr_data_rom[11881]='h00000000;
    rd_cycle[11882] = 1'b1;  wr_cycle[11882] = 1'b0;  addr_rom[11882]='h00001d68;  wr_data_rom[11882]='h00000000;
    rd_cycle[11883] = 1'b1;  wr_cycle[11883] = 1'b0;  addr_rom[11883]='h00001d6c;  wr_data_rom[11883]='h00000000;
    rd_cycle[11884] = 1'b1;  wr_cycle[11884] = 1'b0;  addr_rom[11884]='h00001d70;  wr_data_rom[11884]='h00000000;
    rd_cycle[11885] = 1'b1;  wr_cycle[11885] = 1'b0;  addr_rom[11885]='h00001d74;  wr_data_rom[11885]='h00000000;
    rd_cycle[11886] = 1'b1;  wr_cycle[11886] = 1'b0;  addr_rom[11886]='h00001d78;  wr_data_rom[11886]='h00000000;
    rd_cycle[11887] = 1'b1;  wr_cycle[11887] = 1'b0;  addr_rom[11887]='h00001d7c;  wr_data_rom[11887]='h00000000;
    rd_cycle[11888] = 1'b1;  wr_cycle[11888] = 1'b0;  addr_rom[11888]='h00001d80;  wr_data_rom[11888]='h00000000;
    rd_cycle[11889] = 1'b1;  wr_cycle[11889] = 1'b0;  addr_rom[11889]='h00001d84;  wr_data_rom[11889]='h00000000;
    rd_cycle[11890] = 1'b1;  wr_cycle[11890] = 1'b0;  addr_rom[11890]='h00001d88;  wr_data_rom[11890]='h00000000;
    rd_cycle[11891] = 1'b1;  wr_cycle[11891] = 1'b0;  addr_rom[11891]='h00001d8c;  wr_data_rom[11891]='h00000000;
    rd_cycle[11892] = 1'b1;  wr_cycle[11892] = 1'b0;  addr_rom[11892]='h00001d90;  wr_data_rom[11892]='h00000000;
    rd_cycle[11893] = 1'b1;  wr_cycle[11893] = 1'b0;  addr_rom[11893]='h00001d94;  wr_data_rom[11893]='h00000000;
    rd_cycle[11894] = 1'b1;  wr_cycle[11894] = 1'b0;  addr_rom[11894]='h00001d98;  wr_data_rom[11894]='h00000000;
    rd_cycle[11895] = 1'b1;  wr_cycle[11895] = 1'b0;  addr_rom[11895]='h00001d9c;  wr_data_rom[11895]='h00000000;
    rd_cycle[11896] = 1'b1;  wr_cycle[11896] = 1'b0;  addr_rom[11896]='h00001da0;  wr_data_rom[11896]='h00000000;
    rd_cycle[11897] = 1'b1;  wr_cycle[11897] = 1'b0;  addr_rom[11897]='h00001da4;  wr_data_rom[11897]='h00000000;
    rd_cycle[11898] = 1'b1;  wr_cycle[11898] = 1'b0;  addr_rom[11898]='h00001da8;  wr_data_rom[11898]='h00000000;
    rd_cycle[11899] = 1'b1;  wr_cycle[11899] = 1'b0;  addr_rom[11899]='h00001dac;  wr_data_rom[11899]='h00000000;
    rd_cycle[11900] = 1'b1;  wr_cycle[11900] = 1'b0;  addr_rom[11900]='h00001db0;  wr_data_rom[11900]='h00000000;
    rd_cycle[11901] = 1'b1;  wr_cycle[11901] = 1'b0;  addr_rom[11901]='h00001db4;  wr_data_rom[11901]='h00000000;
    rd_cycle[11902] = 1'b1;  wr_cycle[11902] = 1'b0;  addr_rom[11902]='h00001db8;  wr_data_rom[11902]='h00000000;
    rd_cycle[11903] = 1'b1;  wr_cycle[11903] = 1'b0;  addr_rom[11903]='h00001dbc;  wr_data_rom[11903]='h00000000;
    rd_cycle[11904] = 1'b1;  wr_cycle[11904] = 1'b0;  addr_rom[11904]='h00001dc0;  wr_data_rom[11904]='h00000000;
    rd_cycle[11905] = 1'b1;  wr_cycle[11905] = 1'b0;  addr_rom[11905]='h00001dc4;  wr_data_rom[11905]='h00000000;
    rd_cycle[11906] = 1'b1;  wr_cycle[11906] = 1'b0;  addr_rom[11906]='h00001dc8;  wr_data_rom[11906]='h00000000;
    rd_cycle[11907] = 1'b1;  wr_cycle[11907] = 1'b0;  addr_rom[11907]='h00001dcc;  wr_data_rom[11907]='h00000000;
    rd_cycle[11908] = 1'b1;  wr_cycle[11908] = 1'b0;  addr_rom[11908]='h00001dd0;  wr_data_rom[11908]='h00000000;
    rd_cycle[11909] = 1'b1;  wr_cycle[11909] = 1'b0;  addr_rom[11909]='h00001dd4;  wr_data_rom[11909]='h00000000;
    rd_cycle[11910] = 1'b1;  wr_cycle[11910] = 1'b0;  addr_rom[11910]='h00001dd8;  wr_data_rom[11910]='h00000000;
    rd_cycle[11911] = 1'b1;  wr_cycle[11911] = 1'b0;  addr_rom[11911]='h00001ddc;  wr_data_rom[11911]='h00000000;
    rd_cycle[11912] = 1'b1;  wr_cycle[11912] = 1'b0;  addr_rom[11912]='h00001de0;  wr_data_rom[11912]='h00000000;
    rd_cycle[11913] = 1'b1;  wr_cycle[11913] = 1'b0;  addr_rom[11913]='h00001de4;  wr_data_rom[11913]='h00000000;
    rd_cycle[11914] = 1'b1;  wr_cycle[11914] = 1'b0;  addr_rom[11914]='h00001de8;  wr_data_rom[11914]='h00000000;
    rd_cycle[11915] = 1'b1;  wr_cycle[11915] = 1'b0;  addr_rom[11915]='h00001dec;  wr_data_rom[11915]='h00000000;
    rd_cycle[11916] = 1'b1;  wr_cycle[11916] = 1'b0;  addr_rom[11916]='h00001df0;  wr_data_rom[11916]='h00000000;
    rd_cycle[11917] = 1'b1;  wr_cycle[11917] = 1'b0;  addr_rom[11917]='h00001df4;  wr_data_rom[11917]='h00000000;
    rd_cycle[11918] = 1'b1;  wr_cycle[11918] = 1'b0;  addr_rom[11918]='h00001df8;  wr_data_rom[11918]='h00000000;
    rd_cycle[11919] = 1'b1;  wr_cycle[11919] = 1'b0;  addr_rom[11919]='h00001dfc;  wr_data_rom[11919]='h00000000;
    rd_cycle[11920] = 1'b1;  wr_cycle[11920] = 1'b0;  addr_rom[11920]='h00001e00;  wr_data_rom[11920]='h00000000;
    rd_cycle[11921] = 1'b1;  wr_cycle[11921] = 1'b0;  addr_rom[11921]='h00001e04;  wr_data_rom[11921]='h00000000;
    rd_cycle[11922] = 1'b1;  wr_cycle[11922] = 1'b0;  addr_rom[11922]='h00001e08;  wr_data_rom[11922]='h00000000;
    rd_cycle[11923] = 1'b1;  wr_cycle[11923] = 1'b0;  addr_rom[11923]='h00001e0c;  wr_data_rom[11923]='h00000000;
    rd_cycle[11924] = 1'b1;  wr_cycle[11924] = 1'b0;  addr_rom[11924]='h00001e10;  wr_data_rom[11924]='h00000000;
    rd_cycle[11925] = 1'b1;  wr_cycle[11925] = 1'b0;  addr_rom[11925]='h00001e14;  wr_data_rom[11925]='h00000000;
    rd_cycle[11926] = 1'b1;  wr_cycle[11926] = 1'b0;  addr_rom[11926]='h00001e18;  wr_data_rom[11926]='h00000000;
    rd_cycle[11927] = 1'b1;  wr_cycle[11927] = 1'b0;  addr_rom[11927]='h00001e1c;  wr_data_rom[11927]='h00000000;
    rd_cycle[11928] = 1'b1;  wr_cycle[11928] = 1'b0;  addr_rom[11928]='h00001e20;  wr_data_rom[11928]='h00000000;
    rd_cycle[11929] = 1'b1;  wr_cycle[11929] = 1'b0;  addr_rom[11929]='h00001e24;  wr_data_rom[11929]='h00000000;
    rd_cycle[11930] = 1'b1;  wr_cycle[11930] = 1'b0;  addr_rom[11930]='h00001e28;  wr_data_rom[11930]='h00000000;
    rd_cycle[11931] = 1'b1;  wr_cycle[11931] = 1'b0;  addr_rom[11931]='h00001e2c;  wr_data_rom[11931]='h00000000;
    rd_cycle[11932] = 1'b1;  wr_cycle[11932] = 1'b0;  addr_rom[11932]='h00001e30;  wr_data_rom[11932]='h00000000;
    rd_cycle[11933] = 1'b1;  wr_cycle[11933] = 1'b0;  addr_rom[11933]='h00001e34;  wr_data_rom[11933]='h00000000;
    rd_cycle[11934] = 1'b1;  wr_cycle[11934] = 1'b0;  addr_rom[11934]='h00001e38;  wr_data_rom[11934]='h00000000;
    rd_cycle[11935] = 1'b1;  wr_cycle[11935] = 1'b0;  addr_rom[11935]='h00001e3c;  wr_data_rom[11935]='h00000000;
    rd_cycle[11936] = 1'b1;  wr_cycle[11936] = 1'b0;  addr_rom[11936]='h00001e40;  wr_data_rom[11936]='h00000000;
    rd_cycle[11937] = 1'b1;  wr_cycle[11937] = 1'b0;  addr_rom[11937]='h00001e44;  wr_data_rom[11937]='h00000000;
    rd_cycle[11938] = 1'b1;  wr_cycle[11938] = 1'b0;  addr_rom[11938]='h00001e48;  wr_data_rom[11938]='h00000000;
    rd_cycle[11939] = 1'b1;  wr_cycle[11939] = 1'b0;  addr_rom[11939]='h00001e4c;  wr_data_rom[11939]='h00000000;
    rd_cycle[11940] = 1'b1;  wr_cycle[11940] = 1'b0;  addr_rom[11940]='h00001e50;  wr_data_rom[11940]='h00000000;
    rd_cycle[11941] = 1'b1;  wr_cycle[11941] = 1'b0;  addr_rom[11941]='h00001e54;  wr_data_rom[11941]='h00000000;
    rd_cycle[11942] = 1'b1;  wr_cycle[11942] = 1'b0;  addr_rom[11942]='h00001e58;  wr_data_rom[11942]='h00000000;
    rd_cycle[11943] = 1'b1;  wr_cycle[11943] = 1'b0;  addr_rom[11943]='h00001e5c;  wr_data_rom[11943]='h00000000;
    rd_cycle[11944] = 1'b1;  wr_cycle[11944] = 1'b0;  addr_rom[11944]='h00001e60;  wr_data_rom[11944]='h00000000;
    rd_cycle[11945] = 1'b1;  wr_cycle[11945] = 1'b0;  addr_rom[11945]='h00001e64;  wr_data_rom[11945]='h00000000;
    rd_cycle[11946] = 1'b1;  wr_cycle[11946] = 1'b0;  addr_rom[11946]='h00001e68;  wr_data_rom[11946]='h00000000;
    rd_cycle[11947] = 1'b1;  wr_cycle[11947] = 1'b0;  addr_rom[11947]='h00001e6c;  wr_data_rom[11947]='h00000000;
    rd_cycle[11948] = 1'b1;  wr_cycle[11948] = 1'b0;  addr_rom[11948]='h00001e70;  wr_data_rom[11948]='h00000000;
    rd_cycle[11949] = 1'b1;  wr_cycle[11949] = 1'b0;  addr_rom[11949]='h00001e74;  wr_data_rom[11949]='h00000000;
    rd_cycle[11950] = 1'b1;  wr_cycle[11950] = 1'b0;  addr_rom[11950]='h00001e78;  wr_data_rom[11950]='h00000000;
    rd_cycle[11951] = 1'b1;  wr_cycle[11951] = 1'b0;  addr_rom[11951]='h00001e7c;  wr_data_rom[11951]='h00000000;
    rd_cycle[11952] = 1'b1;  wr_cycle[11952] = 1'b0;  addr_rom[11952]='h00001e80;  wr_data_rom[11952]='h00000000;
    rd_cycle[11953] = 1'b1;  wr_cycle[11953] = 1'b0;  addr_rom[11953]='h00001e84;  wr_data_rom[11953]='h00000000;
    rd_cycle[11954] = 1'b1;  wr_cycle[11954] = 1'b0;  addr_rom[11954]='h00001e88;  wr_data_rom[11954]='h00000000;
    rd_cycle[11955] = 1'b1;  wr_cycle[11955] = 1'b0;  addr_rom[11955]='h00001e8c;  wr_data_rom[11955]='h00000000;
    rd_cycle[11956] = 1'b1;  wr_cycle[11956] = 1'b0;  addr_rom[11956]='h00001e90;  wr_data_rom[11956]='h00000000;
    rd_cycle[11957] = 1'b1;  wr_cycle[11957] = 1'b0;  addr_rom[11957]='h00001e94;  wr_data_rom[11957]='h00000000;
    rd_cycle[11958] = 1'b1;  wr_cycle[11958] = 1'b0;  addr_rom[11958]='h00001e98;  wr_data_rom[11958]='h00000000;
    rd_cycle[11959] = 1'b1;  wr_cycle[11959] = 1'b0;  addr_rom[11959]='h00001e9c;  wr_data_rom[11959]='h00000000;
    rd_cycle[11960] = 1'b1;  wr_cycle[11960] = 1'b0;  addr_rom[11960]='h00001ea0;  wr_data_rom[11960]='h00000000;
    rd_cycle[11961] = 1'b1;  wr_cycle[11961] = 1'b0;  addr_rom[11961]='h00001ea4;  wr_data_rom[11961]='h00000000;
    rd_cycle[11962] = 1'b1;  wr_cycle[11962] = 1'b0;  addr_rom[11962]='h00001ea8;  wr_data_rom[11962]='h00000000;
    rd_cycle[11963] = 1'b1;  wr_cycle[11963] = 1'b0;  addr_rom[11963]='h00001eac;  wr_data_rom[11963]='h00000000;
    rd_cycle[11964] = 1'b1;  wr_cycle[11964] = 1'b0;  addr_rom[11964]='h00001eb0;  wr_data_rom[11964]='h00000000;
    rd_cycle[11965] = 1'b1;  wr_cycle[11965] = 1'b0;  addr_rom[11965]='h00001eb4;  wr_data_rom[11965]='h00000000;
    rd_cycle[11966] = 1'b1;  wr_cycle[11966] = 1'b0;  addr_rom[11966]='h00001eb8;  wr_data_rom[11966]='h00000000;
    rd_cycle[11967] = 1'b1;  wr_cycle[11967] = 1'b0;  addr_rom[11967]='h00001ebc;  wr_data_rom[11967]='h00000000;
    rd_cycle[11968] = 1'b1;  wr_cycle[11968] = 1'b0;  addr_rom[11968]='h00001ec0;  wr_data_rom[11968]='h00000000;
    rd_cycle[11969] = 1'b1;  wr_cycle[11969] = 1'b0;  addr_rom[11969]='h00001ec4;  wr_data_rom[11969]='h00000000;
    rd_cycle[11970] = 1'b1;  wr_cycle[11970] = 1'b0;  addr_rom[11970]='h00001ec8;  wr_data_rom[11970]='h00000000;
    rd_cycle[11971] = 1'b1;  wr_cycle[11971] = 1'b0;  addr_rom[11971]='h00001ecc;  wr_data_rom[11971]='h00000000;
    rd_cycle[11972] = 1'b1;  wr_cycle[11972] = 1'b0;  addr_rom[11972]='h00001ed0;  wr_data_rom[11972]='h00000000;
    rd_cycle[11973] = 1'b1;  wr_cycle[11973] = 1'b0;  addr_rom[11973]='h00001ed4;  wr_data_rom[11973]='h00000000;
    rd_cycle[11974] = 1'b1;  wr_cycle[11974] = 1'b0;  addr_rom[11974]='h00001ed8;  wr_data_rom[11974]='h00000000;
    rd_cycle[11975] = 1'b1;  wr_cycle[11975] = 1'b0;  addr_rom[11975]='h00001edc;  wr_data_rom[11975]='h00000000;
    rd_cycle[11976] = 1'b1;  wr_cycle[11976] = 1'b0;  addr_rom[11976]='h00001ee0;  wr_data_rom[11976]='h00000000;
    rd_cycle[11977] = 1'b1;  wr_cycle[11977] = 1'b0;  addr_rom[11977]='h00001ee4;  wr_data_rom[11977]='h00000000;
    rd_cycle[11978] = 1'b1;  wr_cycle[11978] = 1'b0;  addr_rom[11978]='h00001ee8;  wr_data_rom[11978]='h00000000;
    rd_cycle[11979] = 1'b1;  wr_cycle[11979] = 1'b0;  addr_rom[11979]='h00001eec;  wr_data_rom[11979]='h00000000;
    rd_cycle[11980] = 1'b1;  wr_cycle[11980] = 1'b0;  addr_rom[11980]='h00001ef0;  wr_data_rom[11980]='h00000000;
    rd_cycle[11981] = 1'b1;  wr_cycle[11981] = 1'b0;  addr_rom[11981]='h00001ef4;  wr_data_rom[11981]='h00000000;
    rd_cycle[11982] = 1'b1;  wr_cycle[11982] = 1'b0;  addr_rom[11982]='h00001ef8;  wr_data_rom[11982]='h00000000;
    rd_cycle[11983] = 1'b1;  wr_cycle[11983] = 1'b0;  addr_rom[11983]='h00001efc;  wr_data_rom[11983]='h00000000;
    rd_cycle[11984] = 1'b1;  wr_cycle[11984] = 1'b0;  addr_rom[11984]='h00001f00;  wr_data_rom[11984]='h00000000;
    rd_cycle[11985] = 1'b1;  wr_cycle[11985] = 1'b0;  addr_rom[11985]='h00001f04;  wr_data_rom[11985]='h00000000;
    rd_cycle[11986] = 1'b1;  wr_cycle[11986] = 1'b0;  addr_rom[11986]='h00001f08;  wr_data_rom[11986]='h00000000;
    rd_cycle[11987] = 1'b1;  wr_cycle[11987] = 1'b0;  addr_rom[11987]='h00001f0c;  wr_data_rom[11987]='h00000000;
    rd_cycle[11988] = 1'b1;  wr_cycle[11988] = 1'b0;  addr_rom[11988]='h00001f10;  wr_data_rom[11988]='h00000000;
    rd_cycle[11989] = 1'b1;  wr_cycle[11989] = 1'b0;  addr_rom[11989]='h00001f14;  wr_data_rom[11989]='h00000000;
    rd_cycle[11990] = 1'b1;  wr_cycle[11990] = 1'b0;  addr_rom[11990]='h00001f18;  wr_data_rom[11990]='h00000000;
    rd_cycle[11991] = 1'b1;  wr_cycle[11991] = 1'b0;  addr_rom[11991]='h00001f1c;  wr_data_rom[11991]='h00000000;
    rd_cycle[11992] = 1'b1;  wr_cycle[11992] = 1'b0;  addr_rom[11992]='h00001f20;  wr_data_rom[11992]='h00000000;
    rd_cycle[11993] = 1'b1;  wr_cycle[11993] = 1'b0;  addr_rom[11993]='h00001f24;  wr_data_rom[11993]='h00000000;
    rd_cycle[11994] = 1'b1;  wr_cycle[11994] = 1'b0;  addr_rom[11994]='h00001f28;  wr_data_rom[11994]='h00000000;
    rd_cycle[11995] = 1'b1;  wr_cycle[11995] = 1'b0;  addr_rom[11995]='h00001f2c;  wr_data_rom[11995]='h00000000;
    rd_cycle[11996] = 1'b1;  wr_cycle[11996] = 1'b0;  addr_rom[11996]='h00001f30;  wr_data_rom[11996]='h00000000;
    rd_cycle[11997] = 1'b1;  wr_cycle[11997] = 1'b0;  addr_rom[11997]='h00001f34;  wr_data_rom[11997]='h00000000;
    rd_cycle[11998] = 1'b1;  wr_cycle[11998] = 1'b0;  addr_rom[11998]='h00001f38;  wr_data_rom[11998]='h00000000;
    rd_cycle[11999] = 1'b1;  wr_cycle[11999] = 1'b0;  addr_rom[11999]='h00001f3c;  wr_data_rom[11999]='h00000000;
end

initial begin
    validation_data[    0] = 'h00000042; 
    validation_data[    1] = 'h0000161a; 
    validation_data[    2] = 'h0000142c; 
    validation_data[    3] = 'h00000c3c; 
    validation_data[    4] = 'h00000c86; 
    validation_data[    5] = 'h000004fb; 
    validation_data[    6] = 'h00001064; 
    validation_data[    7] = 'h00000f20; 
    validation_data[    8] = 'h000001a3; 
    validation_data[    9] = 'h000004ef; 
    validation_data[   10] = 'h000019eb; 
    validation_data[   11] = 'h0000086f; 
    validation_data[   12] = 'h00001f14; 
    validation_data[   13] = 'h00001b9b; 
    validation_data[   14] = 'h00000e73; 
    validation_data[   15] = 'h00000e13; 
    validation_data[   16] = 'h00000c17; 
    validation_data[   17] = 'h00001570; 
    validation_data[   18] = 'h0000011e; 
    validation_data[   19] = 'h00000512; 
    validation_data[   20] = 'h00000b8a; 
    validation_data[   21] = 'h000008b8; 
    validation_data[   22] = 'h00000858; 
    validation_data[   23] = 'h000004d1; 
    validation_data[   24] = 'h00001082; 
    validation_data[   25] = 'h0000156c; 
    validation_data[   26] = 'h00000665; 
    validation_data[   27] = 'h00000979; 
    validation_data[   28] = 'h000019d3; 
    validation_data[   29] = 'h00000967; 
    validation_data[   30] = 'h0000127b; 
    validation_data[   31] = 'h00001f06; 
    validation_data[   32] = 'h00001f25; 
    validation_data[   33] = 'h00001766; 
    validation_data[   34] = 'h00000c2a; 
    validation_data[   35] = 'h000010f4; 
    validation_data[   36] = 'h0000078a; 
    validation_data[   37] = 'h00000ae5; 
    validation_data[   38] = 'h000016db; 
    validation_data[   39] = 'h0000131c; 
    validation_data[   40] = 'h000010db; 
    validation_data[   41] = 'h0000127e; 
    validation_data[   42] = 'h000017d8; 
    validation_data[   43] = 'h000011c7; 
    validation_data[   44] = 'h00001219; 
    validation_data[   45] = 'h00000ede; 
    validation_data[   46] = 'h00001842; 
    validation_data[   47] = 'h00001c84; 
    validation_data[   48] = 'h0000107a; 
    validation_data[   49] = 'h00001474; 
    validation_data[   50] = 'h0000197f; 
    validation_data[   51] = 'h00000f15; 
    validation_data[   52] = 'h00000cf0; 
    validation_data[   53] = 'h00001e4e; 
    validation_data[   54] = 'h00001b60; 
    validation_data[   55] = 'h00000107; 
    validation_data[   56] = 'h00001449; 
    validation_data[   57] = 'h00001147; 
    validation_data[   58] = 'h00000997; 
    validation_data[   59] = 'h00000008; 
    validation_data[   60] = 'h000012de; 
    validation_data[   61] = 'h00001e74; 
    validation_data[   62] = 'h00000f07; 
    validation_data[   63] = 'h000005a1; 
    validation_data[   64] = 'h0000069f; 
    validation_data[   65] = 'h00000d73; 
    validation_data[   66] = 'h00001cab; 
    validation_data[   67] = 'h00001002; 
    validation_data[   68] = 'h0000140c; 
    validation_data[   69] = 'h00001e3d; 
    validation_data[   70] = 'h000011eb; 
    validation_data[   71] = 'h00001126; 
    validation_data[   72] = 'h00001d92; 
    validation_data[   73] = 'h000019bc; 
    validation_data[   74] = 'h00001a2e; 
    validation_data[   75] = 'h00000b99; 
    validation_data[   76] = 'h00001a60; 
    validation_data[   77] = 'h000018eb; 
    validation_data[   78] = 'h0000179d; 
    validation_data[   79] = 'h00001969; 
    validation_data[   80] = 'h00000ce7; 
    validation_data[   81] = 'h000000a3; 
    validation_data[   82] = 'h00001724; 
    validation_data[   83] = 'h00000453; 
    validation_data[   84] = 'h00001d70; 
    validation_data[   85] = 'h00000315; 
    validation_data[   86] = 'h00000cd9; 
    validation_data[   87] = 'h00001516; 
    validation_data[   88] = 'h000006ae; 
    validation_data[   89] = 'h000007c2; 
    validation_data[   90] = 'h00000618; 
    validation_data[   91] = 'h00000ac7; 
    validation_data[   92] = 'h0000062f; 
    validation_data[   93] = 'h00000600; 
    validation_data[   94] = 'h000016d9; 
    validation_data[   95] = 'h00001881; 
    validation_data[   96] = 'h00000a68; 
    validation_data[   97] = 'h0000187f; 
    validation_data[   98] = 'h00000902; 
    validation_data[   99] = 'h0000143d; 
    validation_data[  100] = 'h00001590; 
    validation_data[  101] = 'h00000746; 
    validation_data[  102] = 'h00000616; 
    validation_data[  103] = 'h00001220; 
    validation_data[  104] = 'h00001783; 
    validation_data[  105] = 'h000018e4; 
    validation_data[  106] = 'h000017e0; 
    validation_data[  107] = 'h0000050f; 
    validation_data[  108] = 'h000007bc; 
    validation_data[  109] = 'h00000f69; 
    validation_data[  110] = 'h00000ae3; 
    validation_data[  111] = 'h0000023d; 
    validation_data[  112] = 'h000009ec; 
    validation_data[  113] = 'h00000e08; 
    validation_data[  114] = 'h00000cdb; 
    validation_data[  115] = 'h00001dd3; 
    validation_data[  116] = 'h00001eac; 
    validation_data[  117] = 'h00001aa8; 
    validation_data[  118] = 'h00001088; 
    validation_data[  119] = 'h00001aca; 
    validation_data[  120] = 'h000001d1; 
    validation_data[  121] = 'h000011f3; 
    validation_data[  122] = 'h000004eb; 
    validation_data[  123] = 'h0000180b; 
    validation_data[  124] = 'h00000dd4; 
    validation_data[  125] = 'h00000760; 
    validation_data[  126] = 'h00001f2e; 
    validation_data[  127] = 'h000007d7; 
    validation_data[  128] = 'h00000176; 
    validation_data[  129] = 'h000004a1; 
    validation_data[  130] = 'h0000185e; 
    validation_data[  131] = 'h00000326; 
    validation_data[  132] = 'h00000e3b; 
    validation_data[  133] = 'h00000551; 
    validation_data[  134] = 'h00000de0; 
    validation_data[  135] = 'h000017cd; 
    validation_data[  136] = 'h000009b8; 
    validation_data[  137] = 'h00000f51; 
    validation_data[  138] = 'h00000bc1; 
    validation_data[  139] = 'h00001632; 
    validation_data[  140] = 'h00000579; 
    validation_data[  141] = 'h00001b0f; 
    validation_data[  142] = 'h0000134c; 
    validation_data[  143] = 'h00001d37; 
    validation_data[  144] = 'h00000243; 
    validation_data[  145] = 'h00001631; 
    validation_data[  146] = 'h000019e8; 
    validation_data[  147] = 'h000018cc; 
    validation_data[  148] = 'h00000bc1; 
    validation_data[  149] = 'h00001352; 
    validation_data[  150] = 'h00000c51; 
    validation_data[  151] = 'h00000e23; 
    validation_data[  152] = 'h0000118f; 
    validation_data[  153] = 'h0000009c; 
    validation_data[  154] = 'h00000070; 
    validation_data[  155] = 'h00000d92; 
    validation_data[  156] = 'h00001629; 
    validation_data[  157] = 'h000002bc; 
    validation_data[  158] = 'h00001777; 
    validation_data[  159] = 'h00001098; 
    validation_data[  160] = 'h00001da0; 
    validation_data[  161] = 'h00001326; 
    validation_data[  162] = 'h00000de2; 
    validation_data[  163] = 'h0000066a; 
    validation_data[  164] = 'h00001648; 
    validation_data[  165] = 'h00000405; 
    validation_data[  166] = 'h00000325; 
    validation_data[  167] = 'h00000fb7; 
    validation_data[  168] = 'h00000ac4; 
    validation_data[  169] = 'h0000107f; 
    validation_data[  170] = 'h00000261; 
    validation_data[  171] = 'h00000e39; 
    validation_data[  172] = 'h000001f8; 
    validation_data[  173] = 'h00001884; 
    validation_data[  174] = 'h00000261; 
    validation_data[  175] = 'h00000aa4; 
    validation_data[  176] = 'h00000e4a; 
    validation_data[  177] = 'h00000ef3; 
    validation_data[  178] = 'h00000902; 
    validation_data[  179] = 'h00000885; 
    validation_data[  180] = 'h00000fde; 
    validation_data[  181] = 'h00001f2c; 
    validation_data[  182] = 'h00001035; 
    validation_data[  183] = 'h000004d5; 
    validation_data[  184] = 'h0000140c; 
    validation_data[  185] = 'h00000dc8; 
    validation_data[  186] = 'h000015e4; 
    validation_data[  187] = 'h00001350; 
    validation_data[  188] = 'h000009c0; 
    validation_data[  189] = 'h000011a4; 
    validation_data[  190] = 'h00000d91; 
    validation_data[  191] = 'h00001ab1; 
    validation_data[  192] = 'h000007a0; 
    validation_data[  193] = 'h0000188e; 
    validation_data[  194] = 'h000008f9; 
    validation_data[  195] = 'h00000aff; 
    validation_data[  196] = 'h0000019b; 
    validation_data[  197] = 'h00000c12; 
    validation_data[  198] = 'h00001aa0; 
    validation_data[  199] = 'h00000fd7; 
    validation_data[  200] = 'h00000327; 
    validation_data[  201] = 'h00001cf3; 
    validation_data[  202] = 'h000017f8; 
    validation_data[  203] = 'h00001e03; 
    validation_data[  204] = 'h000012e7; 
    validation_data[  205] = 'h000009d0; 
    validation_data[  206] = 'h00000654; 
    validation_data[  207] = 'h000000fe; 
    validation_data[  208] = 'h000010d0; 
    validation_data[  209] = 'h00001e0f; 
    validation_data[  210] = 'h00001c18; 
    validation_data[  211] = 'h00000000; 
    validation_data[  212] = 'h00001b42; 
    validation_data[  213] = 'h00001b70; 
    validation_data[  214] = 'h0000016d; 
    validation_data[  215] = 'h000013d4; 
    validation_data[  216] = 'h00000462; 
    validation_data[  217] = 'h00000872; 
    validation_data[  218] = 'h00001d6f; 
    validation_data[  219] = 'h00000c0a; 
    validation_data[  220] = 'h00000cb6; 
    validation_data[  221] = 'h000019a4; 
    validation_data[  222] = 'h00001aa0; 
    validation_data[  223] = 'h00000f7b; 
    validation_data[  224] = 'h00000ca4; 
    validation_data[  225] = 'h00000eaa; 
    validation_data[  226] = 'h000010aa; 
    validation_data[  227] = 'h000007c1; 
    validation_data[  228] = 'h00001c15; 
    validation_data[  229] = 'h000012fb; 
    validation_data[  230] = 'h00000212; 
    validation_data[  231] = 'h00000238; 
    validation_data[  232] = 'h00000c98; 
    validation_data[  233] = 'h00001a43; 
    validation_data[  234] = 'h000009ef; 
    validation_data[  235] = 'h0000023d; 
    validation_data[  236] = 'h000008d8; 
    validation_data[  237] = 'h00001216; 
    validation_data[  238] = 'h00001924; 
    validation_data[  239] = 'h0000137d; 
    validation_data[  240] = 'h00001b29; 
    validation_data[  241] = 'h00000279; 
    validation_data[  242] = 'h00000462; 
    validation_data[  243] = 'h00001b38; 
    validation_data[  244] = 'h00000041; 
    validation_data[  245] = 'h00001247; 
    validation_data[  246] = 'h00000e78; 
    validation_data[  247] = 'h00001689; 
    validation_data[  248] = 'h00000578; 
    validation_data[  249] = 'h000019aa; 
    validation_data[  250] = 'h00000488; 
    validation_data[  251] = 'h00000f56; 
    validation_data[  252] = 'h000002c5; 
    validation_data[  253] = 'h00001902; 
    validation_data[  254] = 'h0000013a; 
    validation_data[  255] = 'h00000fe8; 
    validation_data[  256] = 'h00001ccb; 
    validation_data[  257] = 'h00001c2a; 
    validation_data[  258] = 'h000017d3; 
    validation_data[  259] = 'h0000170f; 
    validation_data[  260] = 'h000004ab; 
    validation_data[  261] = 'h00000c48; 
    validation_data[  262] = 'h000003b3; 
    validation_data[  263] = 'h000019ce; 
    validation_data[  264] = 'h00001ebf; 
    validation_data[  265] = 'h00000f8d; 
    validation_data[  266] = 'h00001f0d; 
    validation_data[  267] = 'h000014f8; 
    validation_data[  268] = 'h00001bfe; 
    validation_data[  269] = 'h000015cb; 
    validation_data[  270] = 'h00001abd; 
    validation_data[  271] = 'h0000145f; 
    validation_data[  272] = 'h00001502; 
    validation_data[  273] = 'h00000a55; 
    validation_data[  274] = 'h00001095; 
    validation_data[  275] = 'h0000058f; 
    validation_data[  276] = 'h00000096; 
    validation_data[  277] = 'h00000eb3; 
    validation_data[  278] = 'h000015ff; 
    validation_data[  279] = 'h00001be4; 
    validation_data[  280] = 'h0000136d; 
    validation_data[  281] = 'h000015e8; 
    validation_data[  282] = 'h0000014e; 
    validation_data[  283] = 'h00000656; 
    validation_data[  284] = 'h00000e71; 
    validation_data[  285] = 'h0000159e; 
    validation_data[  286] = 'h00000f1c; 
    validation_data[  287] = 'h00001be4; 
    validation_data[  288] = 'h0000172a; 
    validation_data[  289] = 'h00001d12; 
    validation_data[  290] = 'h00000de2; 
    validation_data[  291] = 'h0000055d; 
    validation_data[  292] = 'h00001285; 
    validation_data[  293] = 'h0000075e; 
    validation_data[  294] = 'h00000e25; 
    validation_data[  295] = 'h000010a4; 
    validation_data[  296] = 'h00000541; 
    validation_data[  297] = 'h00000635; 
    validation_data[  298] = 'h00001b11; 
    validation_data[  299] = 'h00000dad; 
    validation_data[  300] = 'h00001d05; 
    validation_data[  301] = 'h00000cff; 
    validation_data[  302] = 'h00000dfc; 
    validation_data[  303] = 'h0000063c; 
    validation_data[  304] = 'h00000f02; 
    validation_data[  305] = 'h00000416; 
    validation_data[  306] = 'h0000193a; 
    validation_data[  307] = 'h00001b6b; 
    validation_data[  308] = 'h00001ce1; 
    validation_data[  309] = 'h000013b0; 
    validation_data[  310] = 'h00000bc3; 
    validation_data[  311] = 'h00001aa7; 
    validation_data[  312] = 'h00001847; 
    validation_data[  313] = 'h00001dbb; 
    validation_data[  314] = 'h00000769; 
    validation_data[  315] = 'h00001c24; 
    validation_data[  316] = 'h000017d3; 
    validation_data[  317] = 'h000008f6; 
    validation_data[  318] = 'h00000662; 
    validation_data[  319] = 'h0000039b; 
    validation_data[  320] = 'h0000042a; 
    validation_data[  321] = 'h000007f6; 
    validation_data[  322] = 'h000004dd; 
    validation_data[  323] = 'h00001173; 
    validation_data[  324] = 'h00000020; 
    validation_data[  325] = 'h00001b15; 
    validation_data[  326] = 'h000000e4; 
    validation_data[  327] = 'h00001a7a; 
    validation_data[  328] = 'h00000d53; 
    validation_data[  329] = 'h0000144a; 
    validation_data[  330] = 'h000017c3; 
    validation_data[  331] = 'h0000173c; 
    validation_data[  332] = 'h000008bc; 
    validation_data[  333] = 'h00000c2e; 
    validation_data[  334] = 'h00001377; 
    validation_data[  335] = 'h00001169; 
    validation_data[  336] = 'h00001092; 
    validation_data[  337] = 'h00000a68; 
    validation_data[  338] = 'h00000510; 
    validation_data[  339] = 'h00001838; 
    validation_data[  340] = 'h000013f7; 
    validation_data[  341] = 'h00001bd2; 
    validation_data[  342] = 'h00001b43; 
    validation_data[  343] = 'h0000124f; 
    validation_data[  344] = 'h0000016f; 
    validation_data[  345] = 'h0000104e; 
    validation_data[  346] = 'h000002c0; 
    validation_data[  347] = 'h00000db7; 
    validation_data[  348] = 'h00001e3e; 
    validation_data[  349] = 'h00001a77; 
    validation_data[  350] = 'h00000e41; 
    validation_data[  351] = 'h00001581; 
    validation_data[  352] = 'h00000246; 
    validation_data[  353] = 'h00001053; 
    validation_data[  354] = 'h00000b0f; 
    validation_data[  355] = 'h00000cc4; 
    validation_data[  356] = 'h00000ad5; 
    validation_data[  357] = 'h00001783; 
    validation_data[  358] = 'h000009c9; 
    validation_data[  359] = 'h00000ab0; 
    validation_data[  360] = 'h00000964; 
    validation_data[  361] = 'h00000c53; 
    validation_data[  362] = 'h000017a9; 
    validation_data[  363] = 'h00000ee6; 
    validation_data[  364] = 'h0000103a; 
    validation_data[  365] = 'h000016c6; 
    validation_data[  366] = 'h00001979; 
    validation_data[  367] = 'h00001e01; 
    validation_data[  368] = 'h000011f5; 
    validation_data[  369] = 'h00000d8f; 
    validation_data[  370] = 'h000010ff; 
    validation_data[  371] = 'h00000f53; 
    validation_data[  372] = 'h0000146e; 
    validation_data[  373] = 'h00000ee4; 
    validation_data[  374] = 'h00000009; 
    validation_data[  375] = 'h0000149c; 
    validation_data[  376] = 'h00000682; 
    validation_data[  377] = 'h000007c9; 
    validation_data[  378] = 'h00000115; 
    validation_data[  379] = 'h00000609; 
    validation_data[  380] = 'h00001b14; 
    validation_data[  381] = 'h000005d3; 
    validation_data[  382] = 'h00000692; 
    validation_data[  383] = 'h000002e6; 
    validation_data[  384] = 'h000005e8; 
    validation_data[  385] = 'h0000194a; 
    validation_data[  386] = 'h000010e3; 
    validation_data[  387] = 'h0000039b; 
    validation_data[  388] = 'h00001cc8; 
    validation_data[  389] = 'h00001c8b; 
    validation_data[  390] = 'h00000591; 
    validation_data[  391] = 'h00000765; 
    validation_data[  392] = 'h00000dda; 
    validation_data[  393] = 'h000002cf; 
    validation_data[  394] = 'h00001227; 
    validation_data[  395] = 'h00000b94; 
    validation_data[  396] = 'h00001861; 
    validation_data[  397] = 'h00000cce; 
    validation_data[  398] = 'h0000057b; 
    validation_data[  399] = 'h0000110e; 
    validation_data[  400] = 'h000008c8; 
    validation_data[  401] = 'h00001278; 
    validation_data[  402] = 'h00000d4b; 
    validation_data[  403] = 'h000007c8; 
    validation_data[  404] = 'h000000d2; 
    validation_data[  405] = 'h000001ec; 
    validation_data[  406] = 'h00001d2a; 
    validation_data[  407] = 'h00001957; 
    validation_data[  408] = 'h00001510; 
    validation_data[  409] = 'h000009f6; 
    validation_data[  410] = 'h000019c8; 
    validation_data[  411] = 'h0000125e; 
    validation_data[  412] = 'h000004a8; 
    validation_data[  413] = 'h00000eba; 
    validation_data[  414] = 'h000015dc; 
    validation_data[  415] = 'h00000c42; 
    validation_data[  416] = 'h0000111d; 
    validation_data[  417] = 'h00000e2b; 
    validation_data[  418] = 'h0000153d; 
    validation_data[  419] = 'h00000b0d; 
    validation_data[  420] = 'h00001c73; 
    validation_data[  421] = 'h000012cf; 
    validation_data[  422] = 'h000007ac; 
    validation_data[  423] = 'h00001d43; 
    validation_data[  424] = 'h00001595; 
    validation_data[  425] = 'h00000d29; 
    validation_data[  426] = 'h00001979; 
    validation_data[  427] = 'h000013fe; 
    validation_data[  428] = 'h00001119; 
    validation_data[  429] = 'h00001ad3; 
    validation_data[  430] = 'h00000472; 
    validation_data[  431] = 'h000016fe; 
    validation_data[  432] = 'h00001783; 
    validation_data[  433] = 'h00001bd3; 
    validation_data[  434] = 'h000004df; 
    validation_data[  435] = 'h00001507; 
    validation_data[  436] = 'h00000266; 
    validation_data[  437] = 'h000002dd; 
    validation_data[  438] = 'h00000afc; 
    validation_data[  439] = 'h00000dfc; 
    validation_data[  440] = 'h00000e5c; 
    validation_data[  441] = 'h000018e0; 
    validation_data[  442] = 'h00001609; 
    validation_data[  443] = 'h00001c28; 
    validation_data[  444] = 'h00000afd; 
    validation_data[  445] = 'h0000154e; 
    validation_data[  446] = 'h00001146; 
    validation_data[  447] = 'h00001d89; 
    validation_data[  448] = 'h00001dbd; 
    validation_data[  449] = 'h00001177; 
    validation_data[  450] = 'h00000b7c; 
    validation_data[  451] = 'h000011e9; 
    validation_data[  452] = 'h0000190e; 
    validation_data[  453] = 'h00001cd2; 
    validation_data[  454] = 'h0000022c; 
    validation_data[  455] = 'h00000dfe; 
    validation_data[  456] = 'h000010ad; 
    validation_data[  457] = 'h00000509; 
    validation_data[  458] = 'h00001bf3; 
    validation_data[  459] = 'h0000146e; 
    validation_data[  460] = 'h00001e69; 
    validation_data[  461] = 'h00001cf5; 
    validation_data[  462] = 'h00001d52; 
    validation_data[  463] = 'h000002ad; 
    validation_data[  464] = 'h000001a2; 
    validation_data[  465] = 'h000001a7; 
    validation_data[  466] = 'h0000132d; 
    validation_data[  467] = 'h00001dd4; 
    validation_data[  468] = 'h00000ea4; 
    validation_data[  469] = 'h00001188; 
    validation_data[  470] = 'h00001820; 
    validation_data[  471] = 'h0000101a; 
    validation_data[  472] = 'h000007ef; 
    validation_data[  473] = 'h00001646; 
    validation_data[  474] = 'h00001aa1; 
    validation_data[  475] = 'h0000158b; 
    validation_data[  476] = 'h0000185e; 
    validation_data[  477] = 'h000006c5; 
    validation_data[  478] = 'h000013d7; 
    validation_data[  479] = 'h00001a48; 
    validation_data[  480] = 'h00000d39; 
    validation_data[  481] = 'h000000b1; 
    validation_data[  482] = 'h000006a9; 
    validation_data[  483] = 'h00000ac5; 
    validation_data[  484] = 'h00000877; 
    validation_data[  485] = 'h00000532; 
    validation_data[  486] = 'h00001d5d; 
    validation_data[  487] = 'h000012a9; 
    validation_data[  488] = 'h00001020; 
    validation_data[  489] = 'h00000d22; 
    validation_data[  490] = 'h00000934; 
    validation_data[  491] = 'h00000171; 
    validation_data[  492] = 'h000003fc; 
    validation_data[  493] = 'h00001c31; 
    validation_data[  494] = 'h00001154; 
    validation_data[  495] = 'h00001c9a; 
    validation_data[  496] = 'h000003a5; 
    validation_data[  497] = 'h00001dbd; 
    validation_data[  498] = 'h00001065; 
    validation_data[  499] = 'h00001f27; 
    validation_data[  500] = 'h000003bf; 
    validation_data[  501] = 'h0000072b; 
    validation_data[  502] = 'h0000062c; 
    validation_data[  503] = 'h00000f80; 
    validation_data[  504] = 'h0000156b; 
    validation_data[  505] = 'h00001d2d; 
    validation_data[  506] = 'h000001c4; 
    validation_data[  507] = 'h00000785; 
    validation_data[  508] = 'h00000133; 
    validation_data[  509] = 'h0000095d; 
    validation_data[  510] = 'h000000f3; 
    validation_data[  511] = 'h00001327; 
    validation_data[  512] = 'h00000d56; 
    validation_data[  513] = 'h00000cad; 
    validation_data[  514] = 'h000015f5; 
    validation_data[  515] = 'h00000256; 
    validation_data[  516] = 'h000004cc; 
    validation_data[  517] = 'h00000e5b; 
    validation_data[  518] = 'h000019be; 
    validation_data[  519] = 'h00000320; 
    validation_data[  520] = 'h000011ae; 
    validation_data[  521] = 'h000003cf; 
    validation_data[  522] = 'h000017cd; 
    validation_data[  523] = 'h00000ef4; 
    validation_data[  524] = 'h0000035c; 
    validation_data[  525] = 'h00000902; 
    validation_data[  526] = 'h00000b92; 
    validation_data[  527] = 'h000010f9; 
    validation_data[  528] = 'h00001693; 
    validation_data[  529] = 'h0000134c; 
    validation_data[  530] = 'h00000355; 
    validation_data[  531] = 'h00000748; 
    validation_data[  532] = 'h000008b9; 
    validation_data[  533] = 'h00000fd7; 
    validation_data[  534] = 'h000013fa; 
    validation_data[  535] = 'h00000eb8; 
    validation_data[  536] = 'h00000051; 
    validation_data[  537] = 'h00001b75; 
    validation_data[  538] = 'h000003cd; 
    validation_data[  539] = 'h0000038a; 
    validation_data[  540] = 'h00001731; 
    validation_data[  541] = 'h00001b85; 
    validation_data[  542] = 'h00001bac; 
    validation_data[  543] = 'h00000e2b; 
    validation_data[  544] = 'h00000491; 
    validation_data[  545] = 'h000009b9; 
    validation_data[  546] = 'h00000249; 
    validation_data[  547] = 'h00001d9a; 
    validation_data[  548] = 'h000005c2; 
    validation_data[  549] = 'h00000226; 
    validation_data[  550] = 'h00001cbf; 
    validation_data[  551] = 'h00001e8d; 
    validation_data[  552] = 'h00001b33; 
    validation_data[  553] = 'h000015ac; 
    validation_data[  554] = 'h000016cc; 
    validation_data[  555] = 'h00001a47; 
    validation_data[  556] = 'h00001463; 
    validation_data[  557] = 'h0000046b; 
    validation_data[  558] = 'h00000013; 
    validation_data[  559] = 'h00001a9e; 
    validation_data[  560] = 'h000009e7; 
    validation_data[  561] = 'h00001483; 
    validation_data[  562] = 'h00001bbc; 
    validation_data[  563] = 'h000014e2; 
    validation_data[  564] = 'h00000a59; 
    validation_data[  565] = 'h000014fe; 
    validation_data[  566] = 'h00001df3; 
    validation_data[  567] = 'h0000150d; 
    validation_data[  568] = 'h000004c0; 
    validation_data[  569] = 'h00001e72; 
    validation_data[  570] = 'h0000056e; 
    validation_data[  571] = 'h0000164f; 
    validation_data[  572] = 'h000016ca; 
    validation_data[  573] = 'h000019f9; 
    validation_data[  574] = 'h00000e89; 
    validation_data[  575] = 'h00000fa4; 
    validation_data[  576] = 'h00000165; 
    validation_data[  577] = 'h00001558; 
    validation_data[  578] = 'h000011e1; 
    validation_data[  579] = 'h00001800; 
    validation_data[  580] = 'h000016ac; 
    validation_data[  581] = 'h00000418; 
    validation_data[  582] = 'h00001d61; 
    validation_data[  583] = 'h00000ce2; 
    validation_data[  584] = 'h00000d21; 
    validation_data[  585] = 'h0000070a; 
    validation_data[  586] = 'h00001b3d; 
    validation_data[  587] = 'h00000fa5; 
    validation_data[  588] = 'h00000f0f; 
    validation_data[  589] = 'h00001ef0; 
    validation_data[  590] = 'h00001c11; 
    validation_data[  591] = 'h000003af; 
    validation_data[  592] = 'h00000279; 
    validation_data[  593] = 'h000015d0; 
    validation_data[  594] = 'h00001851; 
    validation_data[  595] = 'h00001c3b; 
    validation_data[  596] = 'h000002ee; 
    validation_data[  597] = 'h00001c14; 
    validation_data[  598] = 'h00000217; 
    validation_data[  599] = 'h000014d9; 
    validation_data[  600] = 'h00001c64; 
    validation_data[  601] = 'h00000379; 
    validation_data[  602] = 'h000019b5; 
    validation_data[  603] = 'h000014e4; 
    validation_data[  604] = 'h00000f0a; 
    validation_data[  605] = 'h00000dc9; 
    validation_data[  606] = 'h00001ba0; 
    validation_data[  607] = 'h00000e3d; 
    validation_data[  608] = 'h000018d2; 
    validation_data[  609] = 'h00001872; 
    validation_data[  610] = 'h00001d77; 
    validation_data[  611] = 'h00001171; 
    validation_data[  612] = 'h00001bd2; 
    validation_data[  613] = 'h0000076f; 
    validation_data[  614] = 'h0000057b; 
    validation_data[  615] = 'h00000fc0; 
    validation_data[  616] = 'h00000293; 
    validation_data[  617] = 'h00000fef; 
    validation_data[  618] = 'h0000030e; 
    validation_data[  619] = 'h00001bf8; 
    validation_data[  620] = 'h00001506; 
    validation_data[  621] = 'h0000119b; 
    validation_data[  622] = 'h00001866; 
    validation_data[  623] = 'h000001be; 
    validation_data[  624] = 'h00000d7e; 
    validation_data[  625] = 'h00000444; 
    validation_data[  626] = 'h00001aa5; 
    validation_data[  627] = 'h00001970; 
    validation_data[  628] = 'h00001030; 
    validation_data[  629] = 'h00000a68; 
    validation_data[  630] = 'h00000cf2; 
    validation_data[  631] = 'h00001284; 
    validation_data[  632] = 'h0000045b; 
    validation_data[  633] = 'h0000148f; 
    validation_data[  634] = 'h00000b4d; 
    validation_data[  635] = 'h000008c6; 
    validation_data[  636] = 'h00000e4f; 
    validation_data[  637] = 'h00001e50; 
    validation_data[  638] = 'h00001ca3; 
    validation_data[  639] = 'h000006d0; 
    validation_data[  640] = 'h000001d6; 
    validation_data[  641] = 'h00000aee; 
    validation_data[  642] = 'h00001c95; 
    validation_data[  643] = 'h000009b1; 
    validation_data[  644] = 'h00001526; 
    validation_data[  645] = 'h0000113f; 
    validation_data[  646] = 'h000011b3; 
    validation_data[  647] = 'h0000125d; 
    validation_data[  648] = 'h00000497; 
    validation_data[  649] = 'h000009b5; 
    validation_data[  650] = 'h000014d8; 
    validation_data[  651] = 'h0000173c; 
    validation_data[  652] = 'h0000143d; 
    validation_data[  653] = 'h00000ff9; 
    validation_data[  654] = 'h0000197c; 
    validation_data[  655] = 'h00001cda; 
    validation_data[  656] = 'h0000077a; 
    validation_data[  657] = 'h000015ad; 
    validation_data[  658] = 'h0000013e; 
    validation_data[  659] = 'h0000163a; 
    validation_data[  660] = 'h00001183; 
    validation_data[  661] = 'h00001340; 
    validation_data[  662] = 'h0000166f; 
    validation_data[  663] = 'h000001f9; 
    validation_data[  664] = 'h000003e1; 
    validation_data[  665] = 'h00000ba2; 
    validation_data[  666] = 'h00000bc9; 
    validation_data[  667] = 'h00001758; 
    validation_data[  668] = 'h00001619; 
    validation_data[  669] = 'h00000b7f; 
    validation_data[  670] = 'h000013af; 
    validation_data[  671] = 'h00000cac; 
    validation_data[  672] = 'h00001755; 
    validation_data[  673] = 'h00000022; 
    validation_data[  674] = 'h00001c8a; 
    validation_data[  675] = 'h0000090f; 
    validation_data[  676] = 'h00000aa7; 
    validation_data[  677] = 'h00000a1d; 
    validation_data[  678] = 'h00000755; 
    validation_data[  679] = 'h000012d0; 
    validation_data[  680] = 'h00000090; 
    validation_data[  681] = 'h00001675; 
    validation_data[  682] = 'h000014cc; 
    validation_data[  683] = 'h00000ddc; 
    validation_data[  684] = 'h0000110c; 
    validation_data[  685] = 'h00000513; 
    validation_data[  686] = 'h00000b76; 
    validation_data[  687] = 'h000003f7; 
    validation_data[  688] = 'h00000a02; 
    validation_data[  689] = 'h00001eb6; 
    validation_data[  690] = 'h00001640; 
    validation_data[  691] = 'h00001ccd; 
    validation_data[  692] = 'h00001c8f; 
    validation_data[  693] = 'h000001b3; 
    validation_data[  694] = 'h000010a7; 
    validation_data[  695] = 'h00001d4a; 
    validation_data[  696] = 'h00001932; 
    validation_data[  697] = 'h000007f7; 
    validation_data[  698] = 'h000009b1; 
    validation_data[  699] = 'h0000028f; 
    validation_data[  700] = 'h000019e8; 
    validation_data[  701] = 'h00000f66; 
    validation_data[  702] = 'h0000141e; 
    validation_data[  703] = 'h00000a9d; 
    validation_data[  704] = 'h0000140c; 
    validation_data[  705] = 'h0000177b; 
    validation_data[  706] = 'h00001e5c; 
    validation_data[  707] = 'h00000dd6; 
    validation_data[  708] = 'h00000a29; 
    validation_data[  709] = 'h00000ceb; 
    validation_data[  710] = 'h00000805; 
    validation_data[  711] = 'h00001c3d; 
    validation_data[  712] = 'h00001ae8; 
    validation_data[  713] = 'h000001b2; 
    validation_data[  714] = 'h0000064f; 
    validation_data[  715] = 'h000014a7; 
    validation_data[  716] = 'h000015d6; 
    validation_data[  717] = 'h00000d88; 
    validation_data[  718] = 'h00001946; 
    validation_data[  719] = 'h000000ff; 
    validation_data[  720] = 'h000003f1; 
    validation_data[  721] = 'h00001441; 
    validation_data[  722] = 'h00001047; 
    validation_data[  723] = 'h00000631; 
    validation_data[  724] = 'h0000076c; 
    validation_data[  725] = 'h00001464; 
    validation_data[  726] = 'h00000b45; 
    validation_data[  727] = 'h0000141d; 
    validation_data[  728] = 'h00000e66; 
    validation_data[  729] = 'h0000012b; 
    validation_data[  730] = 'h000008dc; 
    validation_data[  731] = 'h00001403; 
    validation_data[  732] = 'h00000b59; 
    validation_data[  733] = 'h00001ae9; 
    validation_data[  734] = 'h0000147e; 
    validation_data[  735] = 'h000012e3; 
    validation_data[  736] = 'h00001dde; 
    validation_data[  737] = 'h00000092; 
    validation_data[  738] = 'h000012d3; 
    validation_data[  739] = 'h00001e38; 
    validation_data[  740] = 'h0000127e; 
    validation_data[  741] = 'h00000dde; 
    validation_data[  742] = 'h0000011d; 
    validation_data[  743] = 'h00000f01; 
    validation_data[  744] = 'h00000887; 
    validation_data[  745] = 'h0000014b; 
    validation_data[  746] = 'h00001df2; 
    validation_data[  747] = 'h000017b5; 
    validation_data[  748] = 'h00001ba1; 
    validation_data[  749] = 'h00001393; 
    validation_data[  750] = 'h000009b0; 
    validation_data[  751] = 'h00000c2c; 
    validation_data[  752] = 'h00000846; 
    validation_data[  753] = 'h00001b78; 
    validation_data[  754] = 'h00001dcd; 
    validation_data[  755] = 'h00000bc6; 
    validation_data[  756] = 'h00001b24; 
    validation_data[  757] = 'h00000a8f; 
    validation_data[  758] = 'h00000da3; 
    validation_data[  759] = 'h0000145d; 
    validation_data[  760] = 'h0000142c; 
    validation_data[  761] = 'h000018ad; 
    validation_data[  762] = 'h00001828; 
    validation_data[  763] = 'h0000163f; 
    validation_data[  764] = 'h00000a6a; 
    validation_data[  765] = 'h000007dc; 
    validation_data[  766] = 'h00001d45; 
    validation_data[  767] = 'h00000634; 
    validation_data[  768] = 'h00001913; 
    validation_data[  769] = 'h00000fa9; 
    validation_data[  770] = 'h000014fa; 
    validation_data[  771] = 'h00001cec; 
    validation_data[  772] = 'h0000016a; 
    validation_data[  773] = 'h0000044c; 
    validation_data[  774] = 'h000001d0; 
    validation_data[  775] = 'h000012fe; 
    validation_data[  776] = 'h00000663; 
    validation_data[  777] = 'h000004b4; 
    validation_data[  778] = 'h00000af9; 
    validation_data[  779] = 'h00001e05; 
    validation_data[  780] = 'h000015dc; 
    validation_data[  781] = 'h00001a24; 
    validation_data[  782] = 'h00001a2f; 
    validation_data[  783] = 'h00001b06; 
    validation_data[  784] = 'h00001c5b; 
    validation_data[  785] = 'h00001217; 
    validation_data[  786] = 'h00001813; 
    validation_data[  787] = 'h000011b4; 
    validation_data[  788] = 'h00001eb3; 
    validation_data[  789] = 'h00000d1d; 
    validation_data[  790] = 'h00000c83; 
    validation_data[  791] = 'h00001bcc; 
    validation_data[  792] = 'h00000c61; 
    validation_data[  793] = 'h000008c3; 
    validation_data[  794] = 'h0000173e; 
    validation_data[  795] = 'h0000132b; 
    validation_data[  796] = 'h0000015d; 
    validation_data[  797] = 'h0000196b; 
    validation_data[  798] = 'h000007af; 
    validation_data[  799] = 'h00000817; 
    validation_data[  800] = 'h00001307; 
    validation_data[  801] = 'h000007fc; 
    validation_data[  802] = 'h0000137b; 
    validation_data[  803] = 'h0000071b; 
    validation_data[  804] = 'h00000dab; 
    validation_data[  805] = 'h000013ea; 
    validation_data[  806] = 'h000016e8; 
    validation_data[  807] = 'h00000077; 
    validation_data[  808] = 'h00000aad; 
    validation_data[  809] = 'h00001dc1; 
    validation_data[  810] = 'h00001577; 
    validation_data[  811] = 'h00000e9b; 
    validation_data[  812] = 'h00001d92; 
    validation_data[  813] = 'h00000405; 
    validation_data[  814] = 'h0000122c; 
    validation_data[  815] = 'h00000eca; 
    validation_data[  816] = 'h000011cd; 
    validation_data[  817] = 'h0000088c; 
    validation_data[  818] = 'h00000c31; 
    validation_data[  819] = 'h00001e6f; 
    validation_data[  820] = 'h000002ee; 
    validation_data[  821] = 'h00000173; 
    validation_data[  822] = 'h00000b14; 
    validation_data[  823] = 'h0000078f; 
    validation_data[  824] = 'h00001c37; 
    validation_data[  825] = 'h000012c9; 
    validation_data[  826] = 'h00001c5f; 
    validation_data[  827] = 'h00000abb; 
    validation_data[  828] = 'h00001acc; 
    validation_data[  829] = 'h00000e58; 
    validation_data[  830] = 'h00001da1; 
    validation_data[  831] = 'h00000075; 
    validation_data[  832] = 'h00001de4; 
    validation_data[  833] = 'h00000d52; 
    validation_data[  834] = 'h00000dd8; 
    validation_data[  835] = 'h00000197; 
    validation_data[  836] = 'h00001b3c; 
    validation_data[  837] = 'h000010fb; 
    validation_data[  838] = 'h00000baf; 
    validation_data[  839] = 'h000014f2; 
    validation_data[  840] = 'h0000084d; 
    validation_data[  841] = 'h00000ae8; 
    validation_data[  842] = 'h00000206; 
    validation_data[  843] = 'h0000181a; 
    validation_data[  844] = 'h0000126a; 
    validation_data[  845] = 'h000019fa; 
    validation_data[  846] = 'h00000b7f; 
    validation_data[  847] = 'h00001b4d; 
    validation_data[  848] = 'h000002ec; 
    validation_data[  849] = 'h00000d2b; 
    validation_data[  850] = 'h00000851; 
    validation_data[  851] = 'h000015bd; 
    validation_data[  852] = 'h00000750; 
    validation_data[  853] = 'h00000c25; 
    validation_data[  854] = 'h00001abe; 
    validation_data[  855] = 'h00001c5a; 
    validation_data[  856] = 'h00001445; 
    validation_data[  857] = 'h00001ecf; 
    validation_data[  858] = 'h000012ef; 
    validation_data[  859] = 'h000000e6; 
    validation_data[  860] = 'h00001426; 
    validation_data[  861] = 'h00000186; 
    validation_data[  862] = 'h00000dd6; 
    validation_data[  863] = 'h00000a6c; 
    validation_data[  864] = 'h0000020b; 
    validation_data[  865] = 'h00000e79; 
    validation_data[  866] = 'h00000f1b; 
    validation_data[  867] = 'h00001e5a; 
    validation_data[  868] = 'h00000fb2; 
    validation_data[  869] = 'h00000786; 
    validation_data[  870] = 'h00000f07; 
    validation_data[  871] = 'h0000074f; 
    validation_data[  872] = 'h00001dcb; 
    validation_data[  873] = 'h0000137d; 
    validation_data[  874] = 'h00000979; 
    validation_data[  875] = 'h00000182; 
    validation_data[  876] = 'h00001a11; 
    validation_data[  877] = 'h00000b0a; 
    validation_data[  878] = 'h00000291; 
    validation_data[  879] = 'h0000021a; 
    validation_data[  880] = 'h000003a9; 
    validation_data[  881] = 'h000017f6; 
    validation_data[  882] = 'h0000044a; 
    validation_data[  883] = 'h00000b43; 
    validation_data[  884] = 'h00000200; 
    validation_data[  885] = 'h000008ec; 
    validation_data[  886] = 'h00001017; 
    validation_data[  887] = 'h00001ed1; 
    validation_data[  888] = 'h00000175; 
    validation_data[  889] = 'h00001a9a; 
    validation_data[  890] = 'h00001592; 
    validation_data[  891] = 'h00000ffd; 
    validation_data[  892] = 'h00000356; 
    validation_data[  893] = 'h00000b73; 
    validation_data[  894] = 'h00000c62; 
    validation_data[  895] = 'h00001245; 
    validation_data[  896] = 'h000009b6; 
    validation_data[  897] = 'h00001ae3; 
    validation_data[  898] = 'h0000075f; 
    validation_data[  899] = 'h00000385; 
    validation_data[  900] = 'h000011f4; 
    validation_data[  901] = 'h0000029a; 
    validation_data[  902] = 'h000012c4; 
    validation_data[  903] = 'h0000170c; 
    validation_data[  904] = 'h00000f95; 
    validation_data[  905] = 'h00001e76; 
    validation_data[  906] = 'h000012b5; 
    validation_data[  907] = 'h000016ce; 
    validation_data[  908] = 'h00001322; 
    validation_data[  909] = 'h000014b2; 
    validation_data[  910] = 'h00000b64; 
    validation_data[  911] = 'h0000004f; 
    validation_data[  912] = 'h000007fa; 
    validation_data[  913] = 'h00001974; 
    validation_data[  914] = 'h00001267; 
    validation_data[  915] = 'h00001271; 
    validation_data[  916] = 'h000005e6; 
    validation_data[  917] = 'h00000c47; 
    validation_data[  918] = 'h00001677; 
    validation_data[  919] = 'h000002a1; 
    validation_data[  920] = 'h00001700; 
    validation_data[  921] = 'h000015e8; 
    validation_data[  922] = 'h00001864; 
    validation_data[  923] = 'h00000ac6; 
    validation_data[  924] = 'h000007ea; 
    validation_data[  925] = 'h00001359; 
    validation_data[  926] = 'h000001a4; 
    validation_data[  927] = 'h00000536; 
    validation_data[  928] = 'h000010a6; 
    validation_data[  929] = 'h00001294; 
    validation_data[  930] = 'h00000173; 
    validation_data[  931] = 'h00000ed7; 
    validation_data[  932] = 'h00000e42; 
    validation_data[  933] = 'h00000a7a; 
    validation_data[  934] = 'h00000e8a; 
    validation_data[  935] = 'h0000057e; 
    validation_data[  936] = 'h000005ec; 
    validation_data[  937] = 'h00001391; 
    validation_data[  938] = 'h000013d1; 
    validation_data[  939] = 'h0000128a; 
    validation_data[  940] = 'h00000bda; 
    validation_data[  941] = 'h0000048e; 
    validation_data[  942] = 'h0000138e; 
    validation_data[  943] = 'h0000047a; 
    validation_data[  944] = 'h00001bea; 
    validation_data[  945] = 'h0000040d; 
    validation_data[  946] = 'h00001437; 
    validation_data[  947] = 'h0000018b; 
    validation_data[  948] = 'h00000f8e; 
    validation_data[  949] = 'h000011af; 
    validation_data[  950] = 'h000001d5; 
    validation_data[  951] = 'h0000109b; 
    validation_data[  952] = 'h00001a90; 
    validation_data[  953] = 'h000009b6; 
    validation_data[  954] = 'h00001f1c; 
    validation_data[  955] = 'h0000082a; 
    validation_data[  956] = 'h000011b9; 
    validation_data[  957] = 'h000009dd; 
    validation_data[  958] = 'h000006df; 
    validation_data[  959] = 'h000001b5; 
    validation_data[  960] = 'h0000113e; 
    validation_data[  961] = 'h00000d0f; 
    validation_data[  962] = 'h00000c40; 
    validation_data[  963] = 'h000002e3; 
    validation_data[  964] = 'h000003e3; 
    validation_data[  965] = 'h00000f7b; 
    validation_data[  966] = 'h00000c9c; 
    validation_data[  967] = 'h0000017f; 
    validation_data[  968] = 'h00000345; 
    validation_data[  969] = 'h00001c59; 
    validation_data[  970] = 'h00001460; 
    validation_data[  971] = 'h00001725; 
    validation_data[  972] = 'h0000037a; 
    validation_data[  973] = 'h000010a5; 
    validation_data[  974] = 'h00000edb; 
    validation_data[  975] = 'h00000923; 
    validation_data[  976] = 'h00001254; 
    validation_data[  977] = 'h00000748; 
    validation_data[  978] = 'h000019dc; 
    validation_data[  979] = 'h00001cae; 
    validation_data[  980] = 'h00000dec; 
    validation_data[  981] = 'h0000072d; 
    validation_data[  982] = 'h00000491; 
    validation_data[  983] = 'h00000fa1; 
    validation_data[  984] = 'h00001358; 
    validation_data[  985] = 'h0000156f; 
    validation_data[  986] = 'h00000ea5; 
    validation_data[  987] = 'h000007ab; 
    validation_data[  988] = 'h00001893; 
    validation_data[  989] = 'h00000bc1; 
    validation_data[  990] = 'h00000b08; 
    validation_data[  991] = 'h0000011b; 
    validation_data[  992] = 'h00000187; 
    validation_data[  993] = 'h000016ea; 
    validation_data[  994] = 'h00000b93; 
    validation_data[  995] = 'h0000132a; 
    validation_data[  996] = 'h00001d99; 
    validation_data[  997] = 'h0000157f; 
    validation_data[  998] = 'h0000104b; 
    validation_data[  999] = 'h000017de; 
    validation_data[ 1000] = 'h0000196a; 
    validation_data[ 1001] = 'h000000c9; 
    validation_data[ 1002] = 'h00000f42; 
    validation_data[ 1003] = 'h00000298; 
    validation_data[ 1004] = 'h00000f91; 
    validation_data[ 1005] = 'h00001604; 
    validation_data[ 1006] = 'h00001ad7; 
    validation_data[ 1007] = 'h00000984; 
    validation_data[ 1008] = 'h00000a99; 
    validation_data[ 1009] = 'h00001af7; 
    validation_data[ 1010] = 'h00001f3a; 
    validation_data[ 1011] = 'h000006a5; 
    validation_data[ 1012] = 'h0000105c; 
    validation_data[ 1013] = 'h000019e5; 
    validation_data[ 1014] = 'h00000c31; 
    validation_data[ 1015] = 'h00001f03; 
    validation_data[ 1016] = 'h00000fd5; 
    validation_data[ 1017] = 'h000017f0; 
    validation_data[ 1018] = 'h00001df1; 
    validation_data[ 1019] = 'h00001a75; 
    validation_data[ 1020] = 'h00000bfc; 
    validation_data[ 1021] = 'h00000f4f; 
    validation_data[ 1022] = 'h00000df4; 
    validation_data[ 1023] = 'h000004a1; 
    validation_data[ 1024] = 'h00000f40; 
    validation_data[ 1025] = 'h000009f3; 
    validation_data[ 1026] = 'h00001e2f; 
    validation_data[ 1027] = 'h00000183; 
    validation_data[ 1028] = 'h000010f8; 
    validation_data[ 1029] = 'h00001a5a; 
    validation_data[ 1030] = 'h00000537; 
    validation_data[ 1031] = 'h00001bfc; 
    validation_data[ 1032] = 'h00000779; 
    validation_data[ 1033] = 'h00001df6; 
    validation_data[ 1034] = 'h000013aa; 
    validation_data[ 1035] = 'h00000075; 
    validation_data[ 1036] = 'h0000098c; 
    validation_data[ 1037] = 'h00001c38; 
    validation_data[ 1038] = 'h000018ee; 
    validation_data[ 1039] = 'h0000166e; 
    validation_data[ 1040] = 'h0000126f; 
    validation_data[ 1041] = 'h00000620; 
    validation_data[ 1042] = 'h00000839; 
    validation_data[ 1043] = 'h000014f1; 
    validation_data[ 1044] = 'h0000128c; 
    validation_data[ 1045] = 'h00000af6; 
    validation_data[ 1046] = 'h000011f3; 
    validation_data[ 1047] = 'h00001d31; 
    validation_data[ 1048] = 'h000018de; 
    validation_data[ 1049] = 'h00000ff7; 
    validation_data[ 1050] = 'h0000064b; 
    validation_data[ 1051] = 'h0000036f; 
    validation_data[ 1052] = 'h00000556; 
    validation_data[ 1053] = 'h00001ce6; 
    validation_data[ 1054] = 'h0000041c; 
    validation_data[ 1055] = 'h00000668; 
    validation_data[ 1056] = 'h00000616; 
    validation_data[ 1057] = 'h0000130c; 
    validation_data[ 1058] = 'h00001304; 
    validation_data[ 1059] = 'h000019f9; 
    validation_data[ 1060] = 'h00001559; 
    validation_data[ 1061] = 'h00000675; 
    validation_data[ 1062] = 'h00000956; 
    validation_data[ 1063] = 'h00001d67; 
    validation_data[ 1064] = 'h000001fa; 
    validation_data[ 1065] = 'h00001139; 
    validation_data[ 1066] = 'h00001edd; 
    validation_data[ 1067] = 'h0000006a; 
    validation_data[ 1068] = 'h00001d69; 
    validation_data[ 1069] = 'h00001ac6; 
    validation_data[ 1070] = 'h00001783; 
    validation_data[ 1071] = 'h00001b0e; 
    validation_data[ 1072] = 'h00000b66; 
    validation_data[ 1073] = 'h00001991; 
    validation_data[ 1074] = 'h000001e7; 
    validation_data[ 1075] = 'h0000186b; 
    validation_data[ 1076] = 'h00000a79; 
    validation_data[ 1077] = 'h00001ccd; 
    validation_data[ 1078] = 'h00001b59; 
    validation_data[ 1079] = 'h0000128b; 
    validation_data[ 1080] = 'h00001380; 
    validation_data[ 1081] = 'h0000157e; 
    validation_data[ 1082] = 'h0000036e; 
    validation_data[ 1083] = 'h000007cc; 
    validation_data[ 1084] = 'h0000121b; 
    validation_data[ 1085] = 'h000015c9; 
    validation_data[ 1086] = 'h000004b3; 
    validation_data[ 1087] = 'h00001852; 
    validation_data[ 1088] = 'h0000003c; 
    validation_data[ 1089] = 'h00000077; 
    validation_data[ 1090] = 'h000000dd; 
    validation_data[ 1091] = 'h00000bd2; 
    validation_data[ 1092] = 'h00000440; 
    validation_data[ 1093] = 'h0000098d; 
    validation_data[ 1094] = 'h000015fb; 
    validation_data[ 1095] = 'h000008d2; 
    validation_data[ 1096] = 'h00000984; 
    validation_data[ 1097] = 'h00000a00; 
    validation_data[ 1098] = 'h00000fdf; 
    validation_data[ 1099] = 'h00001b52; 
    validation_data[ 1100] = 'h000001df; 
    validation_data[ 1101] = 'h00000834; 
    validation_data[ 1102] = 'h00001457; 
    validation_data[ 1103] = 'h00000159; 
    validation_data[ 1104] = 'h00001a85; 
    validation_data[ 1105] = 'h00001c6a; 
    validation_data[ 1106] = 'h00000e61; 
    validation_data[ 1107] = 'h000004ee; 
    validation_data[ 1108] = 'h00001635; 
    validation_data[ 1109] = 'h00000c96; 
    validation_data[ 1110] = 'h0000156d; 
    validation_data[ 1111] = 'h00000078; 
    validation_data[ 1112] = 'h00000a39; 
    validation_data[ 1113] = 'h00000fc6; 
    validation_data[ 1114] = 'h000013d3; 
    validation_data[ 1115] = 'h00001b1f; 
    validation_data[ 1116] = 'h000014f0; 
    validation_data[ 1117] = 'h00000db6; 
    validation_data[ 1118] = 'h0000151f; 
    validation_data[ 1119] = 'h0000095b; 
    validation_data[ 1120] = 'h000000a2; 
    validation_data[ 1121] = 'h00000116; 
    validation_data[ 1122] = 'h00001ad4; 
    validation_data[ 1123] = 'h00001e77; 
    validation_data[ 1124] = 'h00001935; 
    validation_data[ 1125] = 'h000005ac; 
    validation_data[ 1126] = 'h00001d78; 
    validation_data[ 1127] = 'h00001269; 
    validation_data[ 1128] = 'h0000131e; 
    validation_data[ 1129] = 'h000009b3; 
    validation_data[ 1130] = 'h00000dbc; 
    validation_data[ 1131] = 'h00000926; 
    validation_data[ 1132] = 'h0000081c; 
    validation_data[ 1133] = 'h00001c84; 
    validation_data[ 1134] = 'h00000e52; 
    validation_data[ 1135] = 'h00000a95; 
    validation_data[ 1136] = 'h000009f1; 
    validation_data[ 1137] = 'h00000a25; 
    validation_data[ 1138] = 'h00000979; 
    validation_data[ 1139] = 'h00001b9a; 
    validation_data[ 1140] = 'h00000ccf; 
    validation_data[ 1141] = 'h0000110b; 
    validation_data[ 1142] = 'h00000862; 
    validation_data[ 1143] = 'h00000561; 
    validation_data[ 1144] = 'h0000184a; 
    validation_data[ 1145] = 'h00000303; 
    validation_data[ 1146] = 'h00001c07; 
    validation_data[ 1147] = 'h00001e87; 
    validation_data[ 1148] = 'h000013a8; 
    validation_data[ 1149] = 'h00001d3b; 
    validation_data[ 1150] = 'h0000184e; 
    validation_data[ 1151] = 'h00001068; 
    validation_data[ 1152] = 'h000013ed; 
    validation_data[ 1153] = 'h00000061; 
    validation_data[ 1154] = 'h00001033; 
    validation_data[ 1155] = 'h000010e1; 
    validation_data[ 1156] = 'h000019c6; 
    validation_data[ 1157] = 'h0000048b; 
    validation_data[ 1158] = 'h00000acc; 
    validation_data[ 1159] = 'h00001eef; 
    validation_data[ 1160] = 'h000016de; 
    validation_data[ 1161] = 'h000009c0; 
    validation_data[ 1162] = 'h00001d9f; 
    validation_data[ 1163] = 'h00000be6; 
    validation_data[ 1164] = 'h00000589; 
    validation_data[ 1165] = 'h00001b92; 
    validation_data[ 1166] = 'h000005c8; 
    validation_data[ 1167] = 'h0000084a; 
    validation_data[ 1168] = 'h00000fd2; 
    validation_data[ 1169] = 'h00000c72; 
    validation_data[ 1170] = 'h00000ce3; 
    validation_data[ 1171] = 'h00000bdb; 
    validation_data[ 1172] = 'h00001b1c; 
    validation_data[ 1173] = 'h0000166f; 
    validation_data[ 1174] = 'h00000905; 
    validation_data[ 1175] = 'h0000171d; 
    validation_data[ 1176] = 'h0000068b; 
    validation_data[ 1177] = 'h00000171; 
    validation_data[ 1178] = 'h00000449; 
    validation_data[ 1179] = 'h00000a7b; 
    validation_data[ 1180] = 'h0000192e; 
    validation_data[ 1181] = 'h000017db; 
    validation_data[ 1182] = 'h00000b20; 
    validation_data[ 1183] = 'h00001ee5; 
    validation_data[ 1184] = 'h000001de; 
    validation_data[ 1185] = 'h00000d05; 
    validation_data[ 1186] = 'h000004a5; 
    validation_data[ 1187] = 'h00001345; 
    validation_data[ 1188] = 'h00000864; 
    validation_data[ 1189] = 'h0000059a; 
    validation_data[ 1190] = 'h00001537; 
    validation_data[ 1191] = 'h00001dd3; 
    validation_data[ 1192] = 'h00001143; 
    validation_data[ 1193] = 'h00000639; 
    validation_data[ 1194] = 'h000004e4; 
    validation_data[ 1195] = 'h0000156e; 
    validation_data[ 1196] = 'h000002f6; 
    validation_data[ 1197] = 'h00001e20; 
    validation_data[ 1198] = 'h00001f0d; 
    validation_data[ 1199] = 'h00000ceb; 
    validation_data[ 1200] = 'h00000853; 
    validation_data[ 1201] = 'h00000466; 
    validation_data[ 1202] = 'h00000abf; 
    validation_data[ 1203] = 'h00001834; 
    validation_data[ 1204] = 'h00001e5c; 
    validation_data[ 1205] = 'h0000059e; 
    validation_data[ 1206] = 'h000014e0; 
    validation_data[ 1207] = 'h00001d7c; 
    validation_data[ 1208] = 'h0000162d; 
    validation_data[ 1209] = 'h0000132b; 
    validation_data[ 1210] = 'h0000159b; 
    validation_data[ 1211] = 'h000009d0; 
    validation_data[ 1212] = 'h000000bc; 
    validation_data[ 1213] = 'h00000cff; 
    validation_data[ 1214] = 'h00000581; 
    validation_data[ 1215] = 'h00000732; 
    validation_data[ 1216] = 'h000010c2; 
    validation_data[ 1217] = 'h000006c0; 
    validation_data[ 1218] = 'h0000188f; 
    validation_data[ 1219] = 'h0000115f; 
    validation_data[ 1220] = 'h0000016b; 
    validation_data[ 1221] = 'h00000f82; 
    validation_data[ 1222] = 'h000003ea; 
    validation_data[ 1223] = 'h00001df2; 
    validation_data[ 1224] = 'h00001e10; 
    validation_data[ 1225] = 'h00001cd1; 
    validation_data[ 1226] = 'h00000a79; 
    validation_data[ 1227] = 'h00000cc5; 
    validation_data[ 1228] = 'h000001b1; 
    validation_data[ 1229] = 'h000019a5; 
    validation_data[ 1230] = 'h00001c32; 
    validation_data[ 1231] = 'h00000389; 
    validation_data[ 1232] = 'h00001b61; 
    validation_data[ 1233] = 'h000019a2; 
    validation_data[ 1234] = 'h0000169d; 
    validation_data[ 1235] = 'h00000a2c; 
    validation_data[ 1236] = 'h00000fc8; 
    validation_data[ 1237] = 'h0000021a; 
    validation_data[ 1238] = 'h00000108; 
    validation_data[ 1239] = 'h00000dfc; 
    validation_data[ 1240] = 'h00001748; 
    validation_data[ 1241] = 'h00000b94; 
    validation_data[ 1242] = 'h000011e2; 
    validation_data[ 1243] = 'h00000613; 
    validation_data[ 1244] = 'h00001838; 
    validation_data[ 1245] = 'h000014e3; 
    validation_data[ 1246] = 'h0000166f; 
    validation_data[ 1247] = 'h000010ed; 
    validation_data[ 1248] = 'h0000044e; 
    validation_data[ 1249] = 'h000007fe; 
    validation_data[ 1250] = 'h000012c5; 
    validation_data[ 1251] = 'h0000071c; 
    validation_data[ 1252] = 'h0000144e; 
    validation_data[ 1253] = 'h000000eb; 
    validation_data[ 1254] = 'h000010db; 
    validation_data[ 1255] = 'h0000066d; 
    validation_data[ 1256] = 'h00001edc; 
    validation_data[ 1257] = 'h00001ca8; 
    validation_data[ 1258] = 'h00001b39; 
    validation_data[ 1259] = 'h00001bd1; 
    validation_data[ 1260] = 'h00001579; 
    validation_data[ 1261] = 'h0000070d; 
    validation_data[ 1262] = 'h00000f47; 
    validation_data[ 1263] = 'h000000b7; 
    validation_data[ 1264] = 'h00000655; 
    validation_data[ 1265] = 'h00000320; 
    validation_data[ 1266] = 'h000013d6; 
    validation_data[ 1267] = 'h000017cf; 
    validation_data[ 1268] = 'h000012d4; 
    validation_data[ 1269] = 'h00001549; 
    validation_data[ 1270] = 'h00000204; 
    validation_data[ 1271] = 'h0000152f; 
    validation_data[ 1272] = 'h000004c7; 
    validation_data[ 1273] = 'h00000d45; 
    validation_data[ 1274] = 'h00000b9b; 
    validation_data[ 1275] = 'h0000174d; 
    validation_data[ 1276] = 'h00000400; 
    validation_data[ 1277] = 'h000012e2; 
    validation_data[ 1278] = 'h00001c23; 
    validation_data[ 1279] = 'h0000133f; 
    validation_data[ 1280] = 'h00001ddd; 
    validation_data[ 1281] = 'h0000001f; 
    validation_data[ 1282] = 'h000002a7; 
    validation_data[ 1283] = 'h000008e3; 
    validation_data[ 1284] = 'h00000484; 
    validation_data[ 1285] = 'h00000c4a; 
    validation_data[ 1286] = 'h00000e51; 
    validation_data[ 1287] = 'h00000012; 
    validation_data[ 1288] = 'h00000e6c; 
    validation_data[ 1289] = 'h000009dc; 
    validation_data[ 1290] = 'h00001864; 
    validation_data[ 1291] = 'h000017f9; 
    validation_data[ 1292] = 'h00001b32; 
    validation_data[ 1293] = 'h00000260; 
    validation_data[ 1294] = 'h00001784; 
    validation_data[ 1295] = 'h00001c7f; 
    validation_data[ 1296] = 'h00001698; 
    validation_data[ 1297] = 'h00001905; 
    validation_data[ 1298] = 'h000012b0; 
    validation_data[ 1299] = 'h000014c5; 
    validation_data[ 1300] = 'h00001def; 
    validation_data[ 1301] = 'h00001588; 
    validation_data[ 1302] = 'h00000b84; 
    validation_data[ 1303] = 'h000000af; 
    validation_data[ 1304] = 'h00000192; 
    validation_data[ 1305] = 'h00001d89; 
    validation_data[ 1306] = 'h00000a01; 
    validation_data[ 1307] = 'h000002c4; 
    validation_data[ 1308] = 'h00001a01; 
    validation_data[ 1309] = 'h00001f1e; 
    validation_data[ 1310] = 'h00001c91; 
    validation_data[ 1311] = 'h00000d53; 
    validation_data[ 1312] = 'h0000158f; 
    validation_data[ 1313] = 'h00000536; 
    validation_data[ 1314] = 'h00001985; 
    validation_data[ 1315] = 'h00001db0; 
    validation_data[ 1316] = 'h0000089d; 
    validation_data[ 1317] = 'h00001215; 
    validation_data[ 1318] = 'h000009b5; 
    validation_data[ 1319] = 'h00000310; 
    validation_data[ 1320] = 'h0000111e; 
    validation_data[ 1321] = 'h00001474; 
    validation_data[ 1322] = 'h00001323; 
    validation_data[ 1323] = 'h00000954; 
    validation_data[ 1324] = 'h00001036; 
    validation_data[ 1325] = 'h00001b34; 
    validation_data[ 1326] = 'h00001d88; 
    validation_data[ 1327] = 'h00001bcb; 
    validation_data[ 1328] = 'h000010bb; 
    validation_data[ 1329] = 'h000004ad; 
    validation_data[ 1330] = 'h0000047f; 
    validation_data[ 1331] = 'h000014d6; 
    validation_data[ 1332] = 'h00000983; 
    validation_data[ 1333] = 'h000016bc; 
    validation_data[ 1334] = 'h00000a3e; 
    validation_data[ 1335] = 'h00001004; 
    validation_data[ 1336] = 'h00001d2c; 
    validation_data[ 1337] = 'h00001015; 
    validation_data[ 1338] = 'h00000eee; 
    validation_data[ 1339] = 'h000002f1; 
    validation_data[ 1340] = 'h0000132b; 
    validation_data[ 1341] = 'h00001083; 
    validation_data[ 1342] = 'h000009fa; 
    validation_data[ 1343] = 'h00000a1f; 
    validation_data[ 1344] = 'h00001ca7; 
    validation_data[ 1345] = 'h000009e0; 
    validation_data[ 1346] = 'h00001355; 
    validation_data[ 1347] = 'h0000133f; 
    validation_data[ 1348] = 'h000003ed; 
    validation_data[ 1349] = 'h0000053d; 
    validation_data[ 1350] = 'h00000fca; 
    validation_data[ 1351] = 'h00000bf6; 
    validation_data[ 1352] = 'h00001605; 
    validation_data[ 1353] = 'h000006ea; 
    validation_data[ 1354] = 'h000007a8; 
    validation_data[ 1355] = 'h00001b39; 
    validation_data[ 1356] = 'h00000d7a; 
    validation_data[ 1357] = 'h00001732; 
    validation_data[ 1358] = 'h00000b6f; 
    validation_data[ 1359] = 'h0000038d; 
    validation_data[ 1360] = 'h000013e5; 
    validation_data[ 1361] = 'h0000192d; 
    validation_data[ 1362] = 'h00000015; 
    validation_data[ 1363] = 'h000007ea; 
    validation_data[ 1364] = 'h00000efa; 
    validation_data[ 1365] = 'h00001ec1; 
    validation_data[ 1366] = 'h00000fad; 
    validation_data[ 1367] = 'h00000a30; 
    validation_data[ 1368] = 'h00001548; 
    validation_data[ 1369] = 'h00001102; 
    validation_data[ 1370] = 'h000005bf; 
    validation_data[ 1371] = 'h00001b72; 
    validation_data[ 1372] = 'h00000b55; 
    validation_data[ 1373] = 'h00000247; 
    validation_data[ 1374] = 'h000004bf; 
    validation_data[ 1375] = 'h00001631; 
    validation_data[ 1376] = 'h00001815; 
    validation_data[ 1377] = 'h000004fb; 
    validation_data[ 1378] = 'h00001841; 
    validation_data[ 1379] = 'h00000ae8; 
    validation_data[ 1380] = 'h000005c7; 
    validation_data[ 1381] = 'h0000008a; 
    validation_data[ 1382] = 'h000018e5; 
    validation_data[ 1383] = 'h00001e70; 
    validation_data[ 1384] = 'h000000dc; 
    validation_data[ 1385] = 'h00001c81; 
    validation_data[ 1386] = 'h00000de4; 
    validation_data[ 1387] = 'h000001be; 
    validation_data[ 1388] = 'h00000054; 
    validation_data[ 1389] = 'h00001349; 
    validation_data[ 1390] = 'h000008d5; 
    validation_data[ 1391] = 'h0000175e; 
    validation_data[ 1392] = 'h00001890; 
    validation_data[ 1393] = 'h0000139c; 
    validation_data[ 1394] = 'h00001437; 
    validation_data[ 1395] = 'h00000008; 
    validation_data[ 1396] = 'h0000109d; 
    validation_data[ 1397] = 'h0000097e; 
    validation_data[ 1398] = 'h00000411; 
    validation_data[ 1399] = 'h00001cad; 
    validation_data[ 1400] = 'h000009e4; 
    validation_data[ 1401] = 'h000013c6; 
    validation_data[ 1402] = 'h0000188e; 
    validation_data[ 1403] = 'h00001068; 
    validation_data[ 1404] = 'h0000178d; 
    validation_data[ 1405] = 'h00001e06; 
    validation_data[ 1406] = 'h0000061a; 
    validation_data[ 1407] = 'h00001d2e; 
    validation_data[ 1408] = 'h000010ac; 
    validation_data[ 1409] = 'h000005ae; 
    validation_data[ 1410] = 'h00000dbc; 
    validation_data[ 1411] = 'h00000339; 
    validation_data[ 1412] = 'h000002ee; 
    validation_data[ 1413] = 'h00001db6; 
    validation_data[ 1414] = 'h00000755; 
    validation_data[ 1415] = 'h000000d5; 
    validation_data[ 1416] = 'h00000acb; 
    validation_data[ 1417] = 'h000007e0; 
    validation_data[ 1418] = 'h00001a47; 
    validation_data[ 1419] = 'h00001404; 
    validation_data[ 1420] = 'h00001878; 
    validation_data[ 1421] = 'h0000005a; 
    validation_data[ 1422] = 'h0000080b; 
    validation_data[ 1423] = 'h0000084b; 
    validation_data[ 1424] = 'h00001e30; 
    validation_data[ 1425] = 'h00001450; 
    validation_data[ 1426] = 'h00000533; 
    validation_data[ 1427] = 'h00001760; 
    validation_data[ 1428] = 'h00001f3b; 
    validation_data[ 1429] = 'h000014f4; 
    validation_data[ 1430] = 'h00000926; 
    validation_data[ 1431] = 'h00000180; 
    validation_data[ 1432] = 'h00000e8b; 
    validation_data[ 1433] = 'h00001a1e; 
    validation_data[ 1434] = 'h00001442; 
    validation_data[ 1435] = 'h00000691; 
    validation_data[ 1436] = 'h00000cee; 
    validation_data[ 1437] = 'h00000dbf; 
    validation_data[ 1438] = 'h000017ed; 
    validation_data[ 1439] = 'h00001826; 
    validation_data[ 1440] = 'h000002e3; 
    validation_data[ 1441] = 'h00001515; 
    validation_data[ 1442] = 'h0000101a; 
    validation_data[ 1443] = 'h00001ac0; 
    validation_data[ 1444] = 'h0000162a; 
    validation_data[ 1445] = 'h00000f1f; 
    validation_data[ 1446] = 'h00001898; 
    validation_data[ 1447] = 'h00000f19; 
    validation_data[ 1448] = 'h000018e8; 
    validation_data[ 1449] = 'h00001d8f; 
    validation_data[ 1450] = 'h00000ae2; 
    validation_data[ 1451] = 'h00001eaf; 
    validation_data[ 1452] = 'h00001c94; 
    validation_data[ 1453] = 'h00001918; 
    validation_data[ 1454] = 'h00000847; 
    validation_data[ 1455] = 'h00000bd6; 
    validation_data[ 1456] = 'h0000111b; 
    validation_data[ 1457] = 'h0000009e; 
    validation_data[ 1458] = 'h00001aa3; 
    validation_data[ 1459] = 'h0000117a; 
    validation_data[ 1460] = 'h000015aa; 
    validation_data[ 1461] = 'h0000012b; 
    validation_data[ 1462] = 'h00001d1e; 
    validation_data[ 1463] = 'h00001a5b; 
    validation_data[ 1464] = 'h00001d57; 
    validation_data[ 1465] = 'h0000039f; 
    validation_data[ 1466] = 'h000005be; 
    validation_data[ 1467] = 'h00001dc8; 
    validation_data[ 1468] = 'h00000754; 
    validation_data[ 1469] = 'h000013e8; 
    validation_data[ 1470] = 'h000000a0; 
    validation_data[ 1471] = 'h00001859; 
    validation_data[ 1472] = 'h0000095f; 
    validation_data[ 1473] = 'h00001a1d; 
    validation_data[ 1474] = 'h000011cd; 
    validation_data[ 1475] = 'h00000cda; 
    validation_data[ 1476] = 'h00001d93; 
    validation_data[ 1477] = 'h00000cf1; 
    validation_data[ 1478] = 'h000004e0; 
    validation_data[ 1479] = 'h00000a23; 
    validation_data[ 1480] = 'h00000cee; 
    validation_data[ 1481] = 'h0000004f; 
    validation_data[ 1482] = 'h00001270; 
    validation_data[ 1483] = 'h00000ac8; 
    validation_data[ 1484] = 'h00000b79; 
    validation_data[ 1485] = 'h00000cfe; 
    validation_data[ 1486] = 'h000000ab; 
    validation_data[ 1487] = 'h000012ea; 
    validation_data[ 1488] = 'h000004e4; 
    validation_data[ 1489] = 'h00001559; 
    validation_data[ 1490] = 'h0000042c; 
    validation_data[ 1491] = 'h0000052f; 
    validation_data[ 1492] = 'h000019b0; 
    validation_data[ 1493] = 'h00000ac7; 
    validation_data[ 1494] = 'h00000f62; 
    validation_data[ 1495] = 'h000018e2; 
    validation_data[ 1496] = 'h000000b2; 
    validation_data[ 1497] = 'h0000172d; 
    validation_data[ 1498] = 'h000011d1; 
    validation_data[ 1499] = 'h00000c16; 
    validation_data[ 1500] = 'h00000d38; 
    validation_data[ 1501] = 'h00000f15; 
    validation_data[ 1502] = 'h00001da8; 
    validation_data[ 1503] = 'h00001d3a; 
    validation_data[ 1504] = 'h000010f7; 
    validation_data[ 1505] = 'h00001dbf; 
    validation_data[ 1506] = 'h00001871; 
    validation_data[ 1507] = 'h00000a68; 
    validation_data[ 1508] = 'h0000139d; 
    validation_data[ 1509] = 'h00001e89; 
    validation_data[ 1510] = 'h000011e3; 
    validation_data[ 1511] = 'h00001cc5; 
    validation_data[ 1512] = 'h000004a6; 
    validation_data[ 1513] = 'h00000baf; 
    validation_data[ 1514] = 'h000008a7; 
    validation_data[ 1515] = 'h000000f7; 
    validation_data[ 1516] = 'h000001ed; 
    validation_data[ 1517] = 'h00000abe; 
    validation_data[ 1518] = 'h00001314; 
    validation_data[ 1519] = 'h0000118d; 
    validation_data[ 1520] = 'h00000250; 
    validation_data[ 1521] = 'h0000062d; 
    validation_data[ 1522] = 'h000009f8; 
    validation_data[ 1523] = 'h000012c5; 
    validation_data[ 1524] = 'h0000116a; 
    validation_data[ 1525] = 'h00001713; 
    validation_data[ 1526] = 'h000011b0; 
    validation_data[ 1527] = 'h000003d5; 
    validation_data[ 1528] = 'h000015c5; 
    validation_data[ 1529] = 'h00000a69; 
    validation_data[ 1530] = 'h000012e3; 
    validation_data[ 1531] = 'h0000137b; 
    validation_data[ 1532] = 'h00001952; 
    validation_data[ 1533] = 'h000001b3; 
    validation_data[ 1534] = 'h000015f8; 
    validation_data[ 1535] = 'h0000046e; 
    validation_data[ 1536] = 'h000007eb; 
    validation_data[ 1537] = 'h0000061b; 
    validation_data[ 1538] = 'h00001bdc; 
    validation_data[ 1539] = 'h00000ab6; 
    validation_data[ 1540] = 'h0000012a; 
    validation_data[ 1541] = 'h00000196; 
    validation_data[ 1542] = 'h00000234; 
    validation_data[ 1543] = 'h00001b94; 
    validation_data[ 1544] = 'h00000557; 
    validation_data[ 1545] = 'h00001d81; 
    validation_data[ 1546] = 'h0000048c; 
    validation_data[ 1547] = 'h00001d36; 
    validation_data[ 1548] = 'h00001a6d; 
    validation_data[ 1549] = 'h0000108d; 
    validation_data[ 1550] = 'h00000446; 
    validation_data[ 1551] = 'h0000075f; 
    validation_data[ 1552] = 'h00000873; 
    validation_data[ 1553] = 'h00000797; 
    validation_data[ 1554] = 'h00001763; 
    validation_data[ 1555] = 'h00001b45; 
    validation_data[ 1556] = 'h00001879; 
    validation_data[ 1557] = 'h000014c7; 
    validation_data[ 1558] = 'h00000ec7; 
    validation_data[ 1559] = 'h00000845; 
    validation_data[ 1560] = 'h00000028; 
    validation_data[ 1561] = 'h0000142a; 
    validation_data[ 1562] = 'h00000df9; 
    validation_data[ 1563] = 'h000009b1; 
    validation_data[ 1564] = 'h00000ece; 
    validation_data[ 1565] = 'h00000bdb; 
    validation_data[ 1566] = 'h0000181b; 
    validation_data[ 1567] = 'h00001d33; 
    validation_data[ 1568] = 'h00001bda; 
    validation_data[ 1569] = 'h000000df; 
    validation_data[ 1570] = 'h000000a9; 
    validation_data[ 1571] = 'h00000501; 
    validation_data[ 1572] = 'h00001a99; 
    validation_data[ 1573] = 'h00001b27; 
    validation_data[ 1574] = 'h00001e00; 
    validation_data[ 1575] = 'h00000578; 
    validation_data[ 1576] = 'h000000ec; 
    validation_data[ 1577] = 'h00001e8d; 
    validation_data[ 1578] = 'h0000091f; 
    validation_data[ 1579] = 'h00001468; 
    validation_data[ 1580] = 'h0000078a; 
    validation_data[ 1581] = 'h0000062c; 
    validation_data[ 1582] = 'h00000052; 
    validation_data[ 1583] = 'h00000a95; 
    validation_data[ 1584] = 'h00000824; 
    validation_data[ 1585] = 'h000012bb; 
    validation_data[ 1586] = 'h000013d3; 
    validation_data[ 1587] = 'h00000ba7; 
    validation_data[ 1588] = 'h0000141e; 
    validation_data[ 1589] = 'h00001d2d; 
    validation_data[ 1590] = 'h000014eb; 
    validation_data[ 1591] = 'h0000093a; 
    validation_data[ 1592] = 'h00000d14; 
    validation_data[ 1593] = 'h0000087d; 
    validation_data[ 1594] = 'h00000a30; 
    validation_data[ 1595] = 'h000006ac; 
    validation_data[ 1596] = 'h00001ee8; 
    validation_data[ 1597] = 'h0000140e; 
    validation_data[ 1598] = 'h00000d99; 
    validation_data[ 1599] = 'h00000b6d; 
    validation_data[ 1600] = 'h0000076d; 
    validation_data[ 1601] = 'h00001bbd; 
    validation_data[ 1602] = 'h00001dcf; 
    validation_data[ 1603] = 'h0000013d; 
    validation_data[ 1604] = 'h00000926; 
    validation_data[ 1605] = 'h000010dc; 
    validation_data[ 1606] = 'h00000f0b; 
    validation_data[ 1607] = 'h00001d26; 
    validation_data[ 1608] = 'h00000871; 
    validation_data[ 1609] = 'h00001200; 
    validation_data[ 1610] = 'h00001349; 
    validation_data[ 1611] = 'h00001406; 
    validation_data[ 1612] = 'h00000114; 
    validation_data[ 1613] = 'h00000095; 
    validation_data[ 1614] = 'h00001436; 
    validation_data[ 1615] = 'h000019ba; 
    validation_data[ 1616] = 'h00001801; 
    validation_data[ 1617] = 'h00000cba; 
    validation_data[ 1618] = 'h0000137c; 
    validation_data[ 1619] = 'h00001abe; 
    validation_data[ 1620] = 'h00000254; 
    validation_data[ 1621] = 'h0000085f; 
    validation_data[ 1622] = 'h00000452; 
    validation_data[ 1623] = 'h00001cae; 
    validation_data[ 1624] = 'h0000068f; 
    validation_data[ 1625] = 'h0000090c; 
    validation_data[ 1626] = 'h0000057b; 
    validation_data[ 1627] = 'h000013a8; 
    validation_data[ 1628] = 'h00000319; 
    validation_data[ 1629] = 'h00001d95; 
    validation_data[ 1630] = 'h000019cb; 
    validation_data[ 1631] = 'h00000e4b; 
    validation_data[ 1632] = 'h00000694; 
    validation_data[ 1633] = 'h0000174e; 
    validation_data[ 1634] = 'h00001ee5; 
    validation_data[ 1635] = 'h000000fe; 
    validation_data[ 1636] = 'h00000271; 
    validation_data[ 1637] = 'h00000d2e; 
    validation_data[ 1638] = 'h00000ca3; 
    validation_data[ 1639] = 'h00000be7; 
    validation_data[ 1640] = 'h00000622; 
    validation_data[ 1641] = 'h000001df; 
    validation_data[ 1642] = 'h00000db8; 
    validation_data[ 1643] = 'h00001c5d; 
    validation_data[ 1644] = 'h00001f0c; 
    validation_data[ 1645] = 'h00001188; 
    validation_data[ 1646] = 'h00001908; 
    validation_data[ 1647] = 'h000010b9; 
    validation_data[ 1648] = 'h00000ba9; 
    validation_data[ 1649] = 'h000016c3; 
    validation_data[ 1650] = 'h000004ad; 
    validation_data[ 1651] = 'h00000681; 
    validation_data[ 1652] = 'h00001e90; 
    validation_data[ 1653] = 'h00001069; 
    validation_data[ 1654] = 'h000015b2; 
    validation_data[ 1655] = 'h00000456; 
    validation_data[ 1656] = 'h0000096e; 
    validation_data[ 1657] = 'h000010e8; 
    validation_data[ 1658] = 'h0000123e; 
    validation_data[ 1659] = 'h000018f3; 
    validation_data[ 1660] = 'h00001094; 
    validation_data[ 1661] = 'h0000006c; 
    validation_data[ 1662] = 'h00000a4a; 
    validation_data[ 1663] = 'h00000e5f; 
    validation_data[ 1664] = 'h00001878; 
    validation_data[ 1665] = 'h000001cd; 
    validation_data[ 1666] = 'h000015b6; 
    validation_data[ 1667] = 'h00001b72; 
    validation_data[ 1668] = 'h00000150; 
    validation_data[ 1669] = 'h00001a84; 
    validation_data[ 1670] = 'h00001f16; 
    validation_data[ 1671] = 'h00001044; 
    validation_data[ 1672] = 'h00000b64; 
    validation_data[ 1673] = 'h000012c5; 
    validation_data[ 1674] = 'h000006fc; 
    validation_data[ 1675] = 'h000007e2; 
    validation_data[ 1676] = 'h00000fe7; 
    validation_data[ 1677] = 'h00000da6; 
    validation_data[ 1678] = 'h00000b48; 
    validation_data[ 1679] = 'h0000011d; 
    validation_data[ 1680] = 'h00001776; 
    validation_data[ 1681] = 'h00000a54; 
    validation_data[ 1682] = 'h000013cd; 
    validation_data[ 1683] = 'h00001457; 
    validation_data[ 1684] = 'h0000176a; 
    validation_data[ 1685] = 'h00001054; 
    validation_data[ 1686] = 'h000000c6; 
    validation_data[ 1687] = 'h00000d4c; 
    validation_data[ 1688] = 'h00000f6b; 
    validation_data[ 1689] = 'h00001909; 
    validation_data[ 1690] = 'h00001d32; 
    validation_data[ 1691] = 'h00001705; 
    validation_data[ 1692] = 'h000008e4; 
    validation_data[ 1693] = 'h00001084; 
    validation_data[ 1694] = 'h00001dcd; 
    validation_data[ 1695] = 'h00000d8f; 
    validation_data[ 1696] = 'h0000047b; 
    validation_data[ 1697] = 'h00000987; 
    validation_data[ 1698] = 'h00000f8e; 
    validation_data[ 1699] = 'h000002cd; 
    validation_data[ 1700] = 'h000001e9; 
    validation_data[ 1701] = 'h00001933; 
    validation_data[ 1702] = 'h00001d2c; 
    validation_data[ 1703] = 'h00000778; 
    validation_data[ 1704] = 'h00001aab; 
    validation_data[ 1705] = 'h00001a41; 
    validation_data[ 1706] = 'h00000651; 
    validation_data[ 1707] = 'h00000d4b; 
    validation_data[ 1708] = 'h00001223; 
    validation_data[ 1709] = 'h000011e9; 
    validation_data[ 1710] = 'h000018a5; 
    validation_data[ 1711] = 'h00000456; 
    validation_data[ 1712] = 'h00001c0e; 
    validation_data[ 1713] = 'h0000123c; 
    validation_data[ 1714] = 'h00001e3b; 
    validation_data[ 1715] = 'h00000209; 
    validation_data[ 1716] = 'h0000013f; 
    validation_data[ 1717] = 'h000009f8; 
    validation_data[ 1718] = 'h00000889; 
    validation_data[ 1719] = 'h000014b8; 
    validation_data[ 1720] = 'h0000157c; 
    validation_data[ 1721] = 'h000017d3; 
    validation_data[ 1722] = 'h00001103; 
    validation_data[ 1723] = 'h00000abb; 
    validation_data[ 1724] = 'h000012a5; 
    validation_data[ 1725] = 'h000013fd; 
    validation_data[ 1726] = 'h00001c84; 
    validation_data[ 1727] = 'h000016f7; 
    validation_data[ 1728] = 'h00000257; 
    validation_data[ 1729] = 'h00001f05; 
    validation_data[ 1730] = 'h000001e7; 
    validation_data[ 1731] = 'h00001a0c; 
    validation_data[ 1732] = 'h0000020f; 
    validation_data[ 1733] = 'h00000777; 
    validation_data[ 1734] = 'h00000394; 
    validation_data[ 1735] = 'h00000254; 
    validation_data[ 1736] = 'h00000e43; 
    validation_data[ 1737] = 'h00001015; 
    validation_data[ 1738] = 'h00001ec3; 
    validation_data[ 1739] = 'h00000c57; 
    validation_data[ 1740] = 'h00001bba; 
    validation_data[ 1741] = 'h000008b2; 
    validation_data[ 1742] = 'h00001076; 
    validation_data[ 1743] = 'h00000a28; 
    validation_data[ 1744] = 'h000003bd; 
    validation_data[ 1745] = 'h00000027; 
    validation_data[ 1746] = 'h0000151c; 
    validation_data[ 1747] = 'h000016fa; 
    validation_data[ 1748] = 'h0000052f; 
    validation_data[ 1749] = 'h0000199f; 
    validation_data[ 1750] = 'h0000015e; 
    validation_data[ 1751] = 'h0000154d; 
    validation_data[ 1752] = 'h00001199; 
    validation_data[ 1753] = 'h00000843; 
    validation_data[ 1754] = 'h00000cab; 
    validation_data[ 1755] = 'h00001350; 
    validation_data[ 1756] = 'h000011d7; 
    validation_data[ 1757] = 'h00001ec3; 
    validation_data[ 1758] = 'h00000eab; 
    validation_data[ 1759] = 'h00001c92; 
    validation_data[ 1760] = 'h00001671; 
    validation_data[ 1761] = 'h0000096a; 
    validation_data[ 1762] = 'h000005ed; 
    validation_data[ 1763] = 'h000008ad; 
    validation_data[ 1764] = 'h00001dd5; 
    validation_data[ 1765] = 'h00001dc1; 
    validation_data[ 1766] = 'h000010d6; 
    validation_data[ 1767] = 'h00001cea; 
    validation_data[ 1768] = 'h00000848; 
    validation_data[ 1769] = 'h00001d5e; 
    validation_data[ 1770] = 'h00000e3e; 
    validation_data[ 1771] = 'h00000ada; 
    validation_data[ 1772] = 'h000006f3; 
    validation_data[ 1773] = 'h000011ca; 
    validation_data[ 1774] = 'h000002a7; 
    validation_data[ 1775] = 'h00001c6f; 
    validation_data[ 1776] = 'h00000eb5; 
    validation_data[ 1777] = 'h0000169c; 
    validation_data[ 1778] = 'h000009fb; 
    validation_data[ 1779] = 'h00000c83; 
    validation_data[ 1780] = 'h00001c8b; 
    validation_data[ 1781] = 'h00001928; 
    validation_data[ 1782] = 'h0000159c; 
    validation_data[ 1783] = 'h00000c15; 
    validation_data[ 1784] = 'h00000b12; 
    validation_data[ 1785] = 'h0000190d; 
    validation_data[ 1786] = 'h00000ac4; 
    validation_data[ 1787] = 'h000006c1; 
    validation_data[ 1788] = 'h000012bc; 
    validation_data[ 1789] = 'h00001338; 
    validation_data[ 1790] = 'h00000dc7; 
    validation_data[ 1791] = 'h0000093f; 
    validation_data[ 1792] = 'h000006db; 
    validation_data[ 1793] = 'h000018fe; 
    validation_data[ 1794] = 'h00001576; 
    validation_data[ 1795] = 'h00000efb; 
    validation_data[ 1796] = 'h00000cb6; 
    validation_data[ 1797] = 'h000004e4; 
    validation_data[ 1798] = 'h00001a19; 
    validation_data[ 1799] = 'h00000168; 
    validation_data[ 1800] = 'h00000bee; 
    validation_data[ 1801] = 'h00000068; 
    validation_data[ 1802] = 'h00000cc0; 
    validation_data[ 1803] = 'h0000155d; 
    validation_data[ 1804] = 'h000001cc; 
    validation_data[ 1805] = 'h00000053; 
    validation_data[ 1806] = 'h00000f17; 
    validation_data[ 1807] = 'h0000191a; 
    validation_data[ 1808] = 'h0000095d; 
    validation_data[ 1809] = 'h00000da1; 
    validation_data[ 1810] = 'h00001192; 
    validation_data[ 1811] = 'h00001b7d; 
    validation_data[ 1812] = 'h00000024; 
    validation_data[ 1813] = 'h000001f5; 
    validation_data[ 1814] = 'h000010d2; 
    validation_data[ 1815] = 'h00000b87; 
    validation_data[ 1816] = 'h00000670; 
    validation_data[ 1817] = 'h00001e60; 
    validation_data[ 1818] = 'h000008e4; 
    validation_data[ 1819] = 'h00001ec8; 
    validation_data[ 1820] = 'h000015e8; 
    validation_data[ 1821] = 'h00000429; 
    validation_data[ 1822] = 'h00000bd2; 
    validation_data[ 1823] = 'h000017c3; 
    validation_data[ 1824] = 'h00001d44; 
    validation_data[ 1825] = 'h00001994; 
    validation_data[ 1826] = 'h00000bae; 
    validation_data[ 1827] = 'h00000a69; 
    validation_data[ 1828] = 'h00000916; 
    validation_data[ 1829] = 'h00000b5f; 
    validation_data[ 1830] = 'h00001516; 
    validation_data[ 1831] = 'h00000c4b; 
    validation_data[ 1832] = 'h000009e0; 
    validation_data[ 1833] = 'h00000eb9; 
    validation_data[ 1834] = 'h00001f39; 
    validation_data[ 1835] = 'h000017d8; 
    validation_data[ 1836] = 'h00000e04; 
    validation_data[ 1837] = 'h00001664; 
    validation_data[ 1838] = 'h00000951; 
    validation_data[ 1839] = 'h00000cdb; 
    validation_data[ 1840] = 'h000009e7; 
    validation_data[ 1841] = 'h0000049f; 
    validation_data[ 1842] = 'h000011c0; 
    validation_data[ 1843] = 'h00001ac7; 
    validation_data[ 1844] = 'h00001734; 
    validation_data[ 1845] = 'h00001064; 
    validation_data[ 1846] = 'h00000a85; 
    validation_data[ 1847] = 'h00000d18; 
    validation_data[ 1848] = 'h000000f7; 
    validation_data[ 1849] = 'h00001040; 
    validation_data[ 1850] = 'h00000433; 
    validation_data[ 1851] = 'h00000406; 
    validation_data[ 1852] = 'h00001da2; 
    validation_data[ 1853] = 'h0000153f; 
    validation_data[ 1854] = 'h00001380; 
    validation_data[ 1855] = 'h000001b3; 
    validation_data[ 1856] = 'h00001a32; 
    validation_data[ 1857] = 'h00000a46; 
    validation_data[ 1858] = 'h00001c2b; 
    validation_data[ 1859] = 'h000017ab; 
    validation_data[ 1860] = 'h00000f0b; 
    validation_data[ 1861] = 'h0000130c; 
    validation_data[ 1862] = 'h00000052; 
    validation_data[ 1863] = 'h00001944; 
    validation_data[ 1864] = 'h000014da; 
    validation_data[ 1865] = 'h000011eb; 
    validation_data[ 1866] = 'h00000b8f; 
    validation_data[ 1867] = 'h000011e2; 
    validation_data[ 1868] = 'h00000932; 
    validation_data[ 1869] = 'h0000191a; 
    validation_data[ 1870] = 'h00001d2e; 
    validation_data[ 1871] = 'h00000529; 
    validation_data[ 1872] = 'h00000e9f; 
    validation_data[ 1873] = 'h00000e43; 
    validation_data[ 1874] = 'h0000178f; 
    validation_data[ 1875] = 'h000011a1; 
    validation_data[ 1876] = 'h000006af; 
    validation_data[ 1877] = 'h000012a2; 
    validation_data[ 1878] = 'h00001690; 
    validation_data[ 1879] = 'h00000b53; 
    validation_data[ 1880] = 'h00000620; 
    validation_data[ 1881] = 'h00001794; 
    validation_data[ 1882] = 'h00001900; 
    validation_data[ 1883] = 'h0000072c; 
    validation_data[ 1884] = 'h000016c6; 
    validation_data[ 1885] = 'h0000060b; 
    validation_data[ 1886] = 'h00000fa7; 
    validation_data[ 1887] = 'h000009d6; 
    validation_data[ 1888] = 'h00001712; 
    validation_data[ 1889] = 'h0000169c; 
    validation_data[ 1890] = 'h00001afb; 
    validation_data[ 1891] = 'h00001e75; 
    validation_data[ 1892] = 'h0000083d; 
    validation_data[ 1893] = 'h00001f11; 
    validation_data[ 1894] = 'h00001c11; 
    validation_data[ 1895] = 'h0000069b; 
    validation_data[ 1896] = 'h000013bd; 
    validation_data[ 1897] = 'h00000625; 
    validation_data[ 1898] = 'h00001172; 
    validation_data[ 1899] = 'h00000790; 
    validation_data[ 1900] = 'h00001574; 
    validation_data[ 1901] = 'h00000e4e; 
    validation_data[ 1902] = 'h000005bc; 
    validation_data[ 1903] = 'h0000124a; 
    validation_data[ 1904] = 'h00000654; 
    validation_data[ 1905] = 'h00000b7c; 
    validation_data[ 1906] = 'h00001a72; 
    validation_data[ 1907] = 'h00000a72; 
    validation_data[ 1908] = 'h000013fa; 
    validation_data[ 1909] = 'h0000084f; 
    validation_data[ 1910] = 'h0000037d; 
    validation_data[ 1911] = 'h000011ac; 
    validation_data[ 1912] = 'h000014c2; 
    validation_data[ 1913] = 'h000000e5; 
    validation_data[ 1914] = 'h00000083; 
    validation_data[ 1915] = 'h00000975; 
    validation_data[ 1916] = 'h00001934; 
    validation_data[ 1917] = 'h0000135b; 
    validation_data[ 1918] = 'h00001728; 
    validation_data[ 1919] = 'h0000012c; 
    validation_data[ 1920] = 'h000000d4; 
    validation_data[ 1921] = 'h000004ae; 
    validation_data[ 1922] = 'h00000d2d; 
    validation_data[ 1923] = 'h00001b54; 
    validation_data[ 1924] = 'h00000dd8; 
    validation_data[ 1925] = 'h000000d2; 
    validation_data[ 1926] = 'h00000f22; 
    validation_data[ 1927] = 'h00000b01; 
    validation_data[ 1928] = 'h000001ec; 
    validation_data[ 1929] = 'h00001a53; 
    validation_data[ 1930] = 'h00000b40; 
    validation_data[ 1931] = 'h000007b5; 
    validation_data[ 1932] = 'h00001d2e; 
    validation_data[ 1933] = 'h00000169; 
    validation_data[ 1934] = 'h00001d27; 
    validation_data[ 1935] = 'h00000eea; 
    validation_data[ 1936] = 'h00000254; 
    validation_data[ 1937] = 'h00000665; 
    validation_data[ 1938] = 'h0000177f; 
    validation_data[ 1939] = 'h00000411; 
    validation_data[ 1940] = 'h00001c70; 
    validation_data[ 1941] = 'h00000123; 
    validation_data[ 1942] = 'h00001de9; 
    validation_data[ 1943] = 'h00001bd6; 
    validation_data[ 1944] = 'h00001c18; 
    validation_data[ 1945] = 'h00001a9d; 
    validation_data[ 1946] = 'h00000f45; 
    validation_data[ 1947] = 'h000000eb; 
    validation_data[ 1948] = 'h0000151e; 
    validation_data[ 1949] = 'h000016a6; 
    validation_data[ 1950] = 'h000011cd; 
    validation_data[ 1951] = 'h00001285; 
    validation_data[ 1952] = 'h0000117c; 
    validation_data[ 1953] = 'h00001805; 
    validation_data[ 1954] = 'h00000131; 
    validation_data[ 1955] = 'h00000746; 
    validation_data[ 1956] = 'h00001b1e; 
    validation_data[ 1957] = 'h0000050c; 
    validation_data[ 1958] = 'h000013ee; 
    validation_data[ 1959] = 'h00000ca0; 
    validation_data[ 1960] = 'h00001a04; 
    validation_data[ 1961] = 'h00001ad0; 
    validation_data[ 1962] = 'h0000171c; 
    validation_data[ 1963] = 'h000002e1; 
    validation_data[ 1964] = 'h00000e3a; 
    validation_data[ 1965] = 'h00001d58; 
    validation_data[ 1966] = 'h00001770; 
    validation_data[ 1967] = 'h00000a2a; 
    validation_data[ 1968] = 'h00000e7d; 
    validation_data[ 1969] = 'h00001339; 
    validation_data[ 1970] = 'h00001488; 
    validation_data[ 1971] = 'h00001793; 
    validation_data[ 1972] = 'h0000108e; 
    validation_data[ 1973] = 'h00001661; 
    validation_data[ 1974] = 'h00000665; 
    validation_data[ 1975] = 'h000003c2; 
    validation_data[ 1976] = 'h00000785; 
    validation_data[ 1977] = 'h00001c91; 
    validation_data[ 1978] = 'h0000157a; 
    validation_data[ 1979] = 'h00001bf4; 
    validation_data[ 1980] = 'h00001c2c; 
    validation_data[ 1981] = 'h00001110; 
    validation_data[ 1982] = 'h00000e67; 
    validation_data[ 1983] = 'h000015d0; 
    validation_data[ 1984] = 'h00001a0e; 
    validation_data[ 1985] = 'h0000056a; 
    validation_data[ 1986] = 'h0000008d; 
    validation_data[ 1987] = 'h00001b6d; 
    validation_data[ 1988] = 'h00001629; 
    validation_data[ 1989] = 'h00000523; 
    validation_data[ 1990] = 'h00000b99; 
    validation_data[ 1991] = 'h0000067b; 
    validation_data[ 1992] = 'h00000496; 
    validation_data[ 1993] = 'h00000160; 
    validation_data[ 1994] = 'h00001810; 
    validation_data[ 1995] = 'h00001148; 
    validation_data[ 1996] = 'h0000045f; 
    validation_data[ 1997] = 'h0000017d; 
    validation_data[ 1998] = 'h0000054e; 
    validation_data[ 1999] = 'h00001427; 

end


reg clk = 1'b1, rst = 1'b1;
initial #4 rst = 1'b0;
always  #1 clk = ~clk;

wire  miss;
wire [31:0] rd_data;
reg  [31:0] index = 0, wr_data = 0, addr = 0;
reg  rd_req = 1'b0, wr_req = 1'b0;
reg rd_req_ff = 1'b0, miss_ff = 1'b0;
reg [31:0] validation_count = 0;

always @ (posedge clk or posedge rst)
    if(rst) begin
        rd_req_ff <= 1'b0;
        miss_ff   <= 1'b0;
    end else begin
        rd_req_ff <= rd_req;
        miss_ff   <= miss;
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        validation_count <= 0;
    end else begin
        if(validation_count>=`DATA_COUNT) begin
            validation_count <= 'hffffffff;
        end else if(rd_req_ff && (index>(4*`DATA_COUNT))) begin
            if(~miss_ff) begin
                if(validation_data[validation_count]==rd_data)
                    validation_count <= validation_count+1;
                else
                    validation_count <= 0;
            end
        end else begin
            validation_count <= 0;
        end
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        index   <= 0;
        wr_data <= 0;
        addr    <= 0;
        rd_req  <= 1'b0;
        wr_req  <= 1'b0;
    end else begin
        if(~miss) begin
            if(index<`RDWR_COUNT) begin
                if(wr_cycle[index]) begin
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b1;
                end else if(rd_cycle[index]) begin
                    wr_data <= 0;
                    rd_req  <= 1'b1;
                    wr_req  <= 1'b0;
                end else begin
                    wr_data <= 0;
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b0;
                end
                wr_data <= wr_data_rom[index];
                addr    <= addr_rom[index];
                index <= index + 1;
            end else begin
                wr_data <= 0;
                addr    <= 0;
                rd_req  <= 1'b0;
                wr_req  <= 1'b0;
            end
        end
    end

cache #(
    .LINE_ADDR_LEN  ( 3             ),
    .SET_ADDR_LEN   ( 2             ),
    .TAG_ADDR_LEN   ( 12            ),
    .WAY_CNT        ( 3             )
) cache_test_instance (
    .clk            ( clk           ),
    .rst            ( rst           ),
    .miss           ( miss          ),
    .addr           ( addr          ),
    .rd_req         ( rd_req        ),
    .rd_data        ( rd_data       ),
    .wr_req         ( wr_req        ),
    .wr_data        ( wr_data       )
);

endmodule

