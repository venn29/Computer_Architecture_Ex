`timescale 1ns/100ps
//correct read result:
// 00000cc5 00000421 00000221 00000a99 00000030 00000963 000004e5 000007c0 00000503 00000731 0000090a 00000b6e 00000645 0000088c 00000a7e 000008f5 0000031f 00000251 00000c3b 00000c1e 00000d8a 00000946 00000d40 00000e7a 000004bf 00000f34 00000907 0000011b 000008ce 000001c8 000008f1 00000f88 00000ddc 00000a22 00000a79 00000c68 00000cca 0000073d 00000bb1 00000e24 00000241 00000108 00000257 000009a3 00000bdc 000009bd 000004b8 000006d8 000007a0 00000472 000006b6 00000ddf 00000607 00000f70 0000058b 000006ce 0000039e 0000017f 000000de 00000b73 00000126 00000867 0000086d 000002c1 00000ee8 00000276 00000f21 00000bbb 00000831 000006d8 00000e89 00000e4b 00000cd5 000001a3 00000cd7 00000f99 00000d00 000000e1 00000e15 00000c17 0000094c 00000ed0 00000e88 00000267 00000411 00000aa9 00000eb7 0000031d 00000c5e 00000c7f 000003a2 00000358 000009d8 000005ac 0000004f 00000b42 000001c8 0000091f 00000d4a 000006ad 000007b1 0000062e 0000071b 00000b3f 000003dd 00000f3a 00000203 000008b7 000008f5 0000036e 00000763 0000028f 000009ad 00000611 000008c2 00000730 000001ad 000004b6 0000028c 00000628 00000c8d 000008f2 00000a1e 00000758 00000ba3 00000750 00000ea5 000003fc 00000884 0000082a 00000ad3 000007c8 00000f81 00000121 00000476 000005e5 000009db 000000d6 00000749 00000ef3 00000c25 00000158 0000044e 00000d23 000008db 0000085d 00000c99 00000f13 000007e0 00000057 00000670 00000376 00000443 00000e05 000006df 00000b54 00000604 000004d9 000003d4 00000f8a 00000829 00000ce3 0000094c 00000e7a 00000157 00000835 00000926 00000af4 00000918 000007e5 000009ce 00000a7a 000009d9 000007de 00000bd3 00000530 000009b7 00000ce5 00000a50 00000a4b 00000056 0000084d 00000c56 000002cf 0000080e 00000c79 00000c71 000007cf 0000093b 00000038 00000609 00000b83 000001d1 00000c6e 00000217 00000e3a 00000b94 0000065d 00000359 00000cdf 00000f3f 00000131 00000338 00000080 0000051c 000006e9 00000133 00000351 000004a6 0000027e 00000992 00000bf7 00000307 000003e8 00000317 000003c4 00000d9d 00000e56 00000117 00000719 00000d32 00000d7d 00000195 000003cc 00000233 00000212 00000124 00000b1f 00000f63 000007b2 00000447 00000b69 000001df 00000b7d 00000d12 00000b4a 000007f6 000008fc 00000289 00000080 00000f33 0000028d 00000d2c 000009f2 00000df5 000008b2 00000e76 00000653 0000011c 00000097 00000660 0000000e 000005c0 0000011d 00000489 00000431 0000012e 00000786 00000614 000006f8 000000d9 000005c3 00000e48 00000d52 00000118 000004a6 00000766 00000473 00000d6c 00000c13 00000ab0 00000e34 000006be 00000690 0000055f 00000017 00000f31 000001e2 00000439 000006c8 00000c9b 00000a93 00000e5d 00000549 000000c0 000000b6 00000017 000003c6 000004da 00000635 0000077a 00000973 000006d5 00000c15 00000a12 00000ad4 00000b12 0000065e 00000620 00000564 00000b43 00000457 000001b1 00000ae6 00000cc0 000005a1 00000959 0000068f 000006bf 00000563 00000edf 00000919 000008fd 00000f65 0000000a 000004b8 00000637 000003a0 00000e2b 00000f40 00000123 00000f2b 0000025f 00000e7b 00000d9d 00000d8e 000005de 000000c9 00000903 00000238 00000405 0000027f 000002fa 00000bdc 00000ed2 00000a61 0000061c 00000a7f 00000b44 000005c6 00000551 000007ab 000000f6 000004ca 00000228 000007a7 0000023f 000006a0 00000323 000007f0 00000bfb 00000e1b 00000554 00000add 0000056a 00000287 00000540 00000a9a 0000079e 000000f9 00000e8c 000008cd 00000af9 00000677 000006a1 00000a04 00000820 0000023a 00000cb8 00000128 0000055d 00000f79 000001c5 0000020c 00000552 00000659 0000070e 000005be 00000cec 0000063e 0000049b 00000f9b 000009ef 00000199 00000e07 00000839 000008e8 00000477 00000897 00000421 000009c1 00000ecc 0000008c 00000d0c 0000021f 00000a64 00000f93 00000513 000003f3 00000f3d 000005d7 00000c12 000005c7 0000042c 00000487 0000007f 00000309 00000f13 000008b0 00000a36 00000b7c 00000ef0 00000cf8 00000400 000006d7 00000a3c 00000899 000007f7 00000f1f 00000741 0000083c 000007e2 0000098b 000004c7 0000069f 00000a81 00000502 0000029f 00000f62 000004d1 00000f1d 00000d81 0000070c 000003b7 00000a62 00000036 00000e0d 0000064d 00000295 00000115 00000e81 00000c0a 00000421 00000347 000006db 00000568 00000c0a 00000011 00000b4e 00000197 000000e9 000000c1 0000056d 00000cad 00000080 00000b54 00000107 00000598 0000084f 0000016c 00000dc8 000007c7 00000af2 00000414 00000aad 000003bf 000007d4 00000d4c 00000571 00000ee4 00000eaf 00000f1d 00000aa0 00000911 00000945 00000c25 00000be4 00000e3e 00000bf4 00000352 00000704 000004cb 000004b1 00000f67 000003de 0000015a 00000e6b 00000a5e 00000994 00000738 0000017c 00000ad1 0000094b 000001c2 00000a99 000006fb 0000035b 00000ceb 00000ea2 00000709 00000559 00000264 00000ab1 00000495 000007c8 000005ad 00000086 000003f1 00000f7d 00000445 00000ad9 00000331 000005a3 000009fb 0000038d 00000969 00000877 00000782 0000004a 00000187 000002b9 00000a46 00000541 000000af 00000c3c 00000779 00000b4b 00000371 000004ec 00000ad6 00000e8a 00000d4f 00000a0d 00000b36 000001e7 0000045a 000004a0 00000e79 000002a1 00000180 000007a6 0000052d 000000c5 00000614 00000786 00000678 00000e65 0000096e 0000063f 00000bd6 00000748 000001e5 00000970 000002cd 00000dbd 000004c9 000005c5 0000084d 00000552 00000186 0000011c 00000708 00000875 000001a9 0000027b 000002f8 00000c42 00000a0a 00000438 0000048d 00000e5f 00000609 00000334 000006be 00000bec 000006f1 00000a61 00000461 0000065e 00000b0e 00000870 00000ef4 00000dcb 000001f7 0000052d 00000b03 00000685 00000f91 00000250 00000153 000008af 000007f5 00000c28 00000dd3 00000bf9 00000176 00000205 0000075c 00000113 00000f41 00000c9a 0000075c 000002c1 0000032d 00000e46 00000357 00000ae1 00000bab 00000ab8 0000071a 0000095e 0000077b 00000017 000003da 00000670 00000a1c 000007a9 00000565 00000233 00000c15 000009b5 00000990 00000a50 00000ed3 000009bd 00000524 00000543 00000e89 000008fc 000008aa 0000096b 000008f2 00000257 00000047 0000053b 000008d3 00000932 0000038b 00000774 00000751 00000c3c 00000a9a 00000a98 0000024f 0000078f 00000a51 000007db 00000d22 000003bd 00000b72 000007ec 0000030f 00000453 000004ec 00000870 00000a79 00000792 00000b90 00000686 00000a23 000002eb 00000d57 00000b5e 0000028a 000004cd 00000cc3 0000071f 00000d5b 00000e55 00000e20 0000096b 0000096f 00000194 00000959 00000401 00000edb 00000ee5 00000eb7 00000bcd 00000c4b 000000f2 0000008f 00000383 0000084c 00000570 0000077f 00000c41 000001f0 000001f9 00000d3e 00000160 00000f92 000000c6 00000836 00000bfd 00000ee7 00000d64 00000074 00000cb4 00000362 00000065 00000c50 00000d02 00000865 000003cd 00000a00 00000a70 00000a0c 000008ea 00000cab 00000edd 00000f7a 00000219 00000652 0000063b 00000d93 0000024e 00000f9f 00000350 0000000a 000008d5 000000e4 000003fc 00000cea 00000d49 00000dc6 00000aba 00000ae7 00000431 00000ce9 000009e8 000008e4 00000137 00000133 00000072 00000a1d 00000dc3 000004a8 00000563 00000862 00000f10 000007be 00000be0 00000082 00000383 00000882 000006a0 0000004f 000001f6 00000886 0000073b 00000b85 00000978 00000516 000009c2 0000069d 00000d51 00000f87 000005dc 00000c40 00000a31 0000003e 00000860 000009c9 00000b7d 00000f78 00000a30 00000a99 0000046a 000009f2 00000a3c 000008fb 00000f60 00000049 000009ad 000006db 000003da 00000579 00000549 000002f3 000008ea 00000418 00000734 00000269 00000867 00000253 00000711 00000cd7 000004e5 000004e2 0000019c 00000b5d 0000085f 000007c0 00000501 00000cc9 0000049f 00000e8a 00000d03 000007c3 00000439 00000657 00000401 0000084e 00000eec 000004bc 0000035b 000001ca 00000111 00000335 00000dd1 000003cd 00000c7a 00000c61 00000af5 00000878 00000384 00000ed4 00000296 000007b2 000009bf 00000cef 00000d95 00000c96 00000488 000008f9 00000926 00000a7c 000000f3 00000415 00000946 00000a24 0000095b 0000011e 00000f74 000002e4 00000eed 0000072c 00000f52 000007f4 000001b5 00000261 000005c4 00000276 000003f5 00000c44 00000a1d 00000306 00000448 00000c13 00000ea0 00000186 00000f93 00000d8a 00000d1e 0000007f 000008d0 00000eac 00000d6e 00000a57 0000097a 00000c5e 0000069a 00000c73 00000b0b 00000b6a 00000212 0000008e 00000a7c 00000118 00000f8c 00000338 000005a6 00000034 00000078 00000af4 000002dc 00000a85 00000f20 0000047c 00000065 00000d5c 00000051 00000419 000000f1 0000064f 00000eef 00000e27 00000ee6 00000102 000007f3 0000041f 00000cef 000003c0 00000ca7 00000623 000002f8 0000026d 000007f4 0000011e 00000312 000006bf 00000bcf 00000926 00000654 00000686 000008e5 000009b9 0000032b 00000d2e 00000186 00000823 00000266 0000098f 000005b0 00000b91 00000acc 000003bf 00000c0a 00000a96 00000d68 000009a4 00000cf3 000004b0 00000519 00000bb3 000001b3 00000069 00000884 0000099c 0000003b 00000f7f 00000294 000007e7 0000058f 00000b58 00000352 00000ba0 00000330 000000c1 0000060f 000009be 00000317 000001be 0000052e 0000023f 00000442 00000c5a 000005e8 000005a1 00000cc8 00000ef0 000008a3 000006b5 00000dfb 00000111 00000c51 00000f35 00000f7c 000006bc 000009a6 000006f3 0000012f 00000ace 00000b62 00000840 000005ea 00000236 00000e64 00000392 00000c19 0000062f 00000e92 00000623 0000062c 00000433 00000bcd 00000b7a 000001c0 00000133 0000058d 000008e6 00000802 000003f8 00000f6e 00000512 00000b8e 00000bc0 00000a23 0000099b 00000c84 00000e93 000005e8 0000049c 00000b8c 00000a0e 0000076f 00000609 0000076b 00000e29

module cache_tb();

`define DATA_COUNT (1000)
`define RDWR_COUNT (6*`DATA_COUNT)

reg wr_cycle           [`RDWR_COUNT];
reg rd_cycle           [`RDWR_COUNT];
reg [31:0] addr_rom    [`RDWR_COUNT];
reg [31:0] wr_data_rom [`RDWR_COUNT];
reg [31:0] validation_data [`DATA_COUNT];

initial begin
    // 1000 sequence write cycles
    rd_cycle[    0] = 1'b0;  wr_cycle[    0] = 1'b1;  addr_rom[    0]='h00000000;  wr_data_rom[    0]='h00000cc5;
    rd_cycle[    1] = 1'b0;  wr_cycle[    1] = 1'b1;  addr_rom[    1]='h00000004;  wr_data_rom[    1]='h00000421;
    rd_cycle[    2] = 1'b0;  wr_cycle[    2] = 1'b1;  addr_rom[    2]='h00000008;  wr_data_rom[    2]='h00000a58;
    rd_cycle[    3] = 1'b0;  wr_cycle[    3] = 1'b1;  addr_rom[    3]='h0000000c;  wr_data_rom[    3]='h00000a99;
    rd_cycle[    4] = 1'b0;  wr_cycle[    4] = 1'b1;  addr_rom[    4]='h00000010;  wr_data_rom[    4]='h00000030;
    rd_cycle[    5] = 1'b0;  wr_cycle[    5] = 1'b1;  addr_rom[    5]='h00000014;  wr_data_rom[    5]='h00000b7a;
    rd_cycle[    6] = 1'b0;  wr_cycle[    6] = 1'b1;  addr_rom[    6]='h00000018;  wr_data_rom[    6]='h000004e5;
    rd_cycle[    7] = 1'b0;  wr_cycle[    7] = 1'b1;  addr_rom[    7]='h0000001c;  wr_data_rom[    7]='h00000728;
    rd_cycle[    8] = 1'b0;  wr_cycle[    8] = 1'b1;  addr_rom[    8]='h00000020;  wr_data_rom[    8]='h00000ed9;
    rd_cycle[    9] = 1'b0;  wr_cycle[    9] = 1'b1;  addr_rom[    9]='h00000024;  wr_data_rom[    9]='h00000e11;
    rd_cycle[   10] = 1'b0;  wr_cycle[   10] = 1'b1;  addr_rom[   10]='h00000028;  wr_data_rom[   10]='h00000572;
    rd_cycle[   11] = 1'b0;  wr_cycle[   11] = 1'b1;  addr_rom[   11]='h0000002c;  wr_data_rom[   11]='h00000b6e;
    rd_cycle[   12] = 1'b0;  wr_cycle[   12] = 1'b1;  addr_rom[   12]='h00000030;  wr_data_rom[   12]='h00000645;
    rd_cycle[   13] = 1'b0;  wr_cycle[   13] = 1'b1;  addr_rom[   13]='h00000034;  wr_data_rom[   13]='h0000088c;
    rd_cycle[   14] = 1'b0;  wr_cycle[   14] = 1'b1;  addr_rom[   14]='h00000038;  wr_data_rom[   14]='h00000a7e;
    rd_cycle[   15] = 1'b0;  wr_cycle[   15] = 1'b1;  addr_rom[   15]='h0000003c;  wr_data_rom[   15]='h000008f5;
    rd_cycle[   16] = 1'b0;  wr_cycle[   16] = 1'b1;  addr_rom[   16]='h00000040;  wr_data_rom[   16]='h0000043e;
    rd_cycle[   17] = 1'b0;  wr_cycle[   17] = 1'b1;  addr_rom[   17]='h00000044;  wr_data_rom[   17]='h000007ca;
    rd_cycle[   18] = 1'b0;  wr_cycle[   18] = 1'b1;  addr_rom[   18]='h00000048;  wr_data_rom[   18]='h00000da3;
    rd_cycle[   19] = 1'b0;  wr_cycle[   19] = 1'b1;  addr_rom[   19]='h0000004c;  wr_data_rom[   19]='h00000638;
    rd_cycle[   20] = 1'b0;  wr_cycle[   20] = 1'b1;  addr_rom[   20]='h00000050;  wr_data_rom[   20]='h00000369;
    rd_cycle[   21] = 1'b0;  wr_cycle[   21] = 1'b1;  addr_rom[   21]='h00000054;  wr_data_rom[   21]='h00000d0f;
    rd_cycle[   22] = 1'b0;  wr_cycle[   22] = 1'b1;  addr_rom[   22]='h00000058;  wr_data_rom[   22]='h00000f6a;
    rd_cycle[   23] = 1'b0;  wr_cycle[   23] = 1'b1;  addr_rom[   23]='h0000005c;  wr_data_rom[   23]='h0000044d;
    rd_cycle[   24] = 1'b0;  wr_cycle[   24] = 1'b1;  addr_rom[   24]='h00000060;  wr_data_rom[   24]='h00000e3c;
    rd_cycle[   25] = 1'b0;  wr_cycle[   25] = 1'b1;  addr_rom[   25]='h00000064;  wr_data_rom[   25]='h00000d2d;
    rd_cycle[   26] = 1'b0;  wr_cycle[   26] = 1'b1;  addr_rom[   26]='h00000068;  wr_data_rom[   26]='h00000907;
    rd_cycle[   27] = 1'b0;  wr_cycle[   27] = 1'b1;  addr_rom[   27]='h0000006c;  wr_data_rom[   27]='h0000011b;
    rd_cycle[   28] = 1'b0;  wr_cycle[   28] = 1'b1;  addr_rom[   28]='h00000070;  wr_data_rom[   28]='h00000ecc;
    rd_cycle[   29] = 1'b0;  wr_cycle[   29] = 1'b1;  addr_rom[   29]='h00000074;  wr_data_rom[   29]='h000009d8;
    rd_cycle[   30] = 1'b0;  wr_cycle[   30] = 1'b1;  addr_rom[   30]='h00000078;  wr_data_rom[   30]='h00000f48;
    rd_cycle[   31] = 1'b0;  wr_cycle[   31] = 1'b1;  addr_rom[   31]='h0000007c;  wr_data_rom[   31]='h00000f88;
    rd_cycle[   32] = 1'b0;  wr_cycle[   32] = 1'b1;  addr_rom[   32]='h00000080;  wr_data_rom[   32]='h00000ddc;
    rd_cycle[   33] = 1'b0;  wr_cycle[   33] = 1'b1;  addr_rom[   33]='h00000084;  wr_data_rom[   33]='h00000a22;
    rd_cycle[   34] = 1'b0;  wr_cycle[   34] = 1'b1;  addr_rom[   34]='h00000088;  wr_data_rom[   34]='h00000c58;
    rd_cycle[   35] = 1'b0;  wr_cycle[   35] = 1'b1;  addr_rom[   35]='h0000008c;  wr_data_rom[   35]='h00000525;
    rd_cycle[   36] = 1'b0;  wr_cycle[   36] = 1'b1;  addr_rom[   36]='h00000090;  wr_data_rom[   36]='h000001ce;
    rd_cycle[   37] = 1'b0;  wr_cycle[   37] = 1'b1;  addr_rom[   37]='h00000094;  wr_data_rom[   37]='h00000609;
    rd_cycle[   38] = 1'b0;  wr_cycle[   38] = 1'b1;  addr_rom[   38]='h00000098;  wr_data_rom[   38]='h0000013b;
    rd_cycle[   39] = 1'b0;  wr_cycle[   39] = 1'b1;  addr_rom[   39]='h0000009c;  wr_data_rom[   39]='h000004c3;
    rd_cycle[   40] = 1'b0;  wr_cycle[   40] = 1'b1;  addr_rom[   40]='h000000a0;  wr_data_rom[   40]='h00000273;
    rd_cycle[   41] = 1'b0;  wr_cycle[   41] = 1'b1;  addr_rom[   41]='h000000a4;  wr_data_rom[   41]='h00000ee0;
    rd_cycle[   42] = 1'b0;  wr_cycle[   42] = 1'b1;  addr_rom[   42]='h000000a8;  wr_data_rom[   42]='h00000784;
    rd_cycle[   43] = 1'b0;  wr_cycle[   43] = 1'b1;  addr_rom[   43]='h000000ac;  wr_data_rom[   43]='h00000909;
    rd_cycle[   44] = 1'b0;  wr_cycle[   44] = 1'b1;  addr_rom[   44]='h000000b0;  wr_data_rom[   44]='h00000bdc;
    rd_cycle[   45] = 1'b0;  wr_cycle[   45] = 1'b1;  addr_rom[   45]='h000000b4;  wr_data_rom[   45]='h000009bd;
    rd_cycle[   46] = 1'b0;  wr_cycle[   46] = 1'b1;  addr_rom[   46]='h000000b8;  wr_data_rom[   46]='h0000005f;
    rd_cycle[   47] = 1'b0;  wr_cycle[   47] = 1'b1;  addr_rom[   47]='h000000bc;  wr_data_rom[   47]='h000006d8;
    rd_cycle[   48] = 1'b0;  wr_cycle[   48] = 1'b1;  addr_rom[   48]='h000000c0;  wr_data_rom[   48]='h00000799;
    rd_cycle[   49] = 1'b0;  wr_cycle[   49] = 1'b1;  addr_rom[   49]='h000000c4;  wr_data_rom[   49]='h00000079;
    rd_cycle[   50] = 1'b0;  wr_cycle[   50] = 1'b1;  addr_rom[   50]='h000000c8;  wr_data_rom[   50]='h00000125;
    rd_cycle[   51] = 1'b0;  wr_cycle[   51] = 1'b1;  addr_rom[   51]='h000000cc;  wr_data_rom[   51]='h00000ee0;
    rd_cycle[   52] = 1'b0;  wr_cycle[   52] = 1'b1;  addr_rom[   52]='h000000d0;  wr_data_rom[   52]='h00000d1e;
    rd_cycle[   53] = 1'b0;  wr_cycle[   53] = 1'b1;  addr_rom[   53]='h000000d4;  wr_data_rom[   53]='h00000dbd;
    rd_cycle[   54] = 1'b0;  wr_cycle[   54] = 1'b1;  addr_rom[   54]='h000000d8;  wr_data_rom[   54]='h00000ac1;
    rd_cycle[   55] = 1'b0;  wr_cycle[   55] = 1'b1;  addr_rom[   55]='h000000dc;  wr_data_rom[   55]='h000006ce;
    rd_cycle[   56] = 1'b0;  wr_cycle[   56] = 1'b1;  addr_rom[   56]='h000000e0;  wr_data_rom[   56]='h00000c88;
    rd_cycle[   57] = 1'b0;  wr_cycle[   57] = 1'b1;  addr_rom[   57]='h000000e4;  wr_data_rom[   57]='h0000017f;
    rd_cycle[   58] = 1'b0;  wr_cycle[   58] = 1'b1;  addr_rom[   58]='h000000e8;  wr_data_rom[   58]='h000007b1;
    rd_cycle[   59] = 1'b0;  wr_cycle[   59] = 1'b1;  addr_rom[   59]='h000000ec;  wr_data_rom[   59]='h00000b73;
    rd_cycle[   60] = 1'b0;  wr_cycle[   60] = 1'b1;  addr_rom[   60]='h000000f0;  wr_data_rom[   60]='h00000126;
    rd_cycle[   61] = 1'b0;  wr_cycle[   61] = 1'b1;  addr_rom[   61]='h000000f4;  wr_data_rom[   61]='h00000acd;
    rd_cycle[   62] = 1'b0;  wr_cycle[   62] = 1'b1;  addr_rom[   62]='h000000f8;  wr_data_rom[   62]='h00000c8d;
    rd_cycle[   63] = 1'b0;  wr_cycle[   63] = 1'b1;  addr_rom[   63]='h000000fc;  wr_data_rom[   63]='h00000de3;
    rd_cycle[   64] = 1'b0;  wr_cycle[   64] = 1'b1;  addr_rom[   64]='h00000100;  wr_data_rom[   64]='h000005cd;
    rd_cycle[   65] = 1'b0;  wr_cycle[   65] = 1'b1;  addr_rom[   65]='h00000104;  wr_data_rom[   65]='h000001b8;
    rd_cycle[   66] = 1'b0;  wr_cycle[   66] = 1'b1;  addr_rom[   66]='h00000108;  wr_data_rom[   66]='h00000f21;
    rd_cycle[   67] = 1'b0;  wr_cycle[   67] = 1'b1;  addr_rom[   67]='h0000010c;  wr_data_rom[   67]='h00000d75;
    rd_cycle[   68] = 1'b0;  wr_cycle[   68] = 1'b1;  addr_rom[   68]='h00000110;  wr_data_rom[   68]='h00000f67;
    rd_cycle[   69] = 1'b0;  wr_cycle[   69] = 1'b1;  addr_rom[   69]='h00000114;  wr_data_rom[   69]='h00000ef7;
    rd_cycle[   70] = 1'b0;  wr_cycle[   70] = 1'b1;  addr_rom[   70]='h00000118;  wr_data_rom[   70]='h00000e89;
    rd_cycle[   71] = 1'b0;  wr_cycle[   71] = 1'b1;  addr_rom[   71]='h0000011c;  wr_data_rom[   71]='h00000cd9;
    rd_cycle[   72] = 1'b0;  wr_cycle[   72] = 1'b1;  addr_rom[   72]='h00000120;  wr_data_rom[   72]='h0000041e;
    rd_cycle[   73] = 1'b0;  wr_cycle[   73] = 1'b1;  addr_rom[   73]='h00000124;  wr_data_rom[   73]='h000006b3;
    rd_cycle[   74] = 1'b0;  wr_cycle[   74] = 1'b1;  addr_rom[   74]='h00000128;  wr_data_rom[   74]='h000003c4;
    rd_cycle[   75] = 1'b0;  wr_cycle[   75] = 1'b1;  addr_rom[   75]='h0000012c;  wr_data_rom[   75]='h00000da3;
    rd_cycle[   76] = 1'b0;  wr_cycle[   76] = 1'b1;  addr_rom[   76]='h00000130;  wr_data_rom[   76]='h00000d00;
    rd_cycle[   77] = 1'b0;  wr_cycle[   77] = 1'b1;  addr_rom[   77]='h00000134;  wr_data_rom[   77]='h00000bfd;
    rd_cycle[   78] = 1'b0;  wr_cycle[   78] = 1'b1;  addr_rom[   78]='h00000138;  wr_data_rom[   78]='h000000d5;
    rd_cycle[   79] = 1'b0;  wr_cycle[   79] = 1'b1;  addr_rom[   79]='h0000013c;  wr_data_rom[   79]='h00000c17;
    rd_cycle[   80] = 1'b0;  wr_cycle[   80] = 1'b1;  addr_rom[   80]='h00000140;  wr_data_rom[   80]='h00000ea6;
    rd_cycle[   81] = 1'b0;  wr_cycle[   81] = 1'b1;  addr_rom[   81]='h00000144;  wr_data_rom[   81]='h000002ea;
    rd_cycle[   82] = 1'b0;  wr_cycle[   82] = 1'b1;  addr_rom[   82]='h00000148;  wr_data_rom[   82]='h000002cf;
    rd_cycle[   83] = 1'b0;  wr_cycle[   83] = 1'b1;  addr_rom[   83]='h0000014c;  wr_data_rom[   83]='h00000348;
    rd_cycle[   84] = 1'b0;  wr_cycle[   84] = 1'b1;  addr_rom[   84]='h00000150;  wr_data_rom[   84]='h0000076d;
    rd_cycle[   85] = 1'b0;  wr_cycle[   85] = 1'b1;  addr_rom[   85]='h00000154;  wr_data_rom[   85]='h00000aa9;
    rd_cycle[   86] = 1'b0;  wr_cycle[   86] = 1'b1;  addr_rom[   86]='h00000158;  wr_data_rom[   86]='h00000eb7;
    rd_cycle[   87] = 1'b0;  wr_cycle[   87] = 1'b1;  addr_rom[   87]='h0000015c;  wr_data_rom[   87]='h00000de7;
    rd_cycle[   88] = 1'b0;  wr_cycle[   88] = 1'b1;  addr_rom[   88]='h00000160;  wr_data_rom[   88]='h000001c8;
    rd_cycle[   89] = 1'b0;  wr_cycle[   89] = 1'b1;  addr_rom[   89]='h00000164;  wr_data_rom[   89]='h000002c1;
    rd_cycle[   90] = 1'b0;  wr_cycle[   90] = 1'b1;  addr_rom[   90]='h00000168;  wr_data_rom[   90]='h000003a2;
    rd_cycle[   91] = 1'b0;  wr_cycle[   91] = 1'b1;  addr_rom[   91]='h0000016c;  wr_data_rom[   91]='h0000047d;
    rd_cycle[   92] = 1'b0;  wr_cycle[   92] = 1'b1;  addr_rom[   92]='h00000170;  wr_data_rom[   92]='h000004a3;
    rd_cycle[   93] = 1'b0;  wr_cycle[   93] = 1'b1;  addr_rom[   93]='h00000174;  wr_data_rom[   93]='h00000814;
    rd_cycle[   94] = 1'b0;  wr_cycle[   94] = 1'b1;  addr_rom[   94]='h00000178;  wr_data_rom[   94]='h0000004f;
    rd_cycle[   95] = 1'b0;  wr_cycle[   95] = 1'b1;  addr_rom[   95]='h0000017c;  wr_data_rom[   95]='h00000b42;
    rd_cycle[   96] = 1'b0;  wr_cycle[   96] = 1'b1;  addr_rom[   96]='h00000180;  wr_data_rom[   96]='h000002cd;
    rd_cycle[   97] = 1'b0;  wr_cycle[   97] = 1'b1;  addr_rom[   97]='h00000184;  wr_data_rom[   97]='h0000091f;
    rd_cycle[   98] = 1'b0;  wr_cycle[   98] = 1'b1;  addr_rom[   98]='h00000188;  wr_data_rom[   98]='h00000496;
    rd_cycle[   99] = 1'b0;  wr_cycle[   99] = 1'b1;  addr_rom[   99]='h0000018c;  wr_data_rom[   99]='h0000007f;
    rd_cycle[  100] = 1'b0;  wr_cycle[  100] = 1'b1;  addr_rom[  100]='h00000190;  wr_data_rom[  100]='h000007b1;
    rd_cycle[  101] = 1'b0;  wr_cycle[  101] = 1'b1;  addr_rom[  101]='h00000194;  wr_data_rom[  101]='h00000c26;
    rd_cycle[  102] = 1'b0;  wr_cycle[  102] = 1'b1;  addr_rom[  102]='h00000198;  wr_data_rom[  102]='h000009b1;
    rd_cycle[  103] = 1'b0;  wr_cycle[  103] = 1'b1;  addr_rom[  103]='h0000019c;  wr_data_rom[  103]='h00000608;
    rd_cycle[  104] = 1'b0;  wr_cycle[  104] = 1'b1;  addr_rom[  104]='h000001a0;  wr_data_rom[  104]='h000003cd;
    rd_cycle[  105] = 1'b0;  wr_cycle[  105] = 1'b1;  addr_rom[  105]='h000001a4;  wr_data_rom[  105]='h00000d3e;
    rd_cycle[  106] = 1'b0;  wr_cycle[  106] = 1'b1;  addr_rom[  106]='h000001a8;  wr_data_rom[  106]='h000000e9;
    rd_cycle[  107] = 1'b0;  wr_cycle[  107] = 1'b1;  addr_rom[  107]='h000001ac;  wr_data_rom[  107]='h000006d0;
    rd_cycle[  108] = 1'b0;  wr_cycle[  108] = 1'b1;  addr_rom[  108]='h000001b0;  wr_data_rom[  108]='h00000aa2;
    rd_cycle[  109] = 1'b0;  wr_cycle[  109] = 1'b1;  addr_rom[  109]='h000001b4;  wr_data_rom[  109]='h00000a88;
    rd_cycle[  110] = 1'b0;  wr_cycle[  110] = 1'b1;  addr_rom[  110]='h000001b8;  wr_data_rom[  110]='h00000763;
    rd_cycle[  111] = 1'b0;  wr_cycle[  111] = 1'b1;  addr_rom[  111]='h000001bc;  wr_data_rom[  111]='h000001a8;
    rd_cycle[  112] = 1'b0;  wr_cycle[  112] = 1'b1;  addr_rom[  112]='h000001c0;  wr_data_rom[  112]='h000009ad;
    rd_cycle[  113] = 1'b0;  wr_cycle[  113] = 1'b1;  addr_rom[  113]='h000001c4;  wr_data_rom[  113]='h00000611;
    rd_cycle[  114] = 1'b0;  wr_cycle[  114] = 1'b1;  addr_rom[  114]='h000001c8;  wr_data_rom[  114]='h00000d5f;
    rd_cycle[  115] = 1'b0;  wr_cycle[  115] = 1'b1;  addr_rom[  115]='h000001cc;  wr_data_rom[  115]='h00000730;
    rd_cycle[  116] = 1'b0;  wr_cycle[  116] = 1'b1;  addr_rom[  116]='h000001d0;  wr_data_rom[  116]='h000007e2;
    rd_cycle[  117] = 1'b0;  wr_cycle[  117] = 1'b1;  addr_rom[  117]='h000001d4;  wr_data_rom[  117]='h000008bb;
    rd_cycle[  118] = 1'b0;  wr_cycle[  118] = 1'b1;  addr_rom[  118]='h000001d8;  wr_data_rom[  118]='h0000034e;
    rd_cycle[  119] = 1'b0;  wr_cycle[  119] = 1'b1;  addr_rom[  119]='h000001dc;  wr_data_rom[  119]='h000001c3;
    rd_cycle[  120] = 1'b0;  wr_cycle[  120] = 1'b1;  addr_rom[  120]='h000001e0;  wr_data_rom[  120]='h0000067c;
    rd_cycle[  121] = 1'b0;  wr_cycle[  121] = 1'b1;  addr_rom[  121]='h000001e4;  wr_data_rom[  121]='h000008f2;
    rd_cycle[  122] = 1'b0;  wr_cycle[  122] = 1'b1;  addr_rom[  122]='h000001e8;  wr_data_rom[  122]='h0000001c;
    rd_cycle[  123] = 1'b0;  wr_cycle[  123] = 1'b1;  addr_rom[  123]='h000001ec;  wr_data_rom[  123]='h0000059e;
    rd_cycle[  124] = 1'b0;  wr_cycle[  124] = 1'b1;  addr_rom[  124]='h000001f0;  wr_data_rom[  124]='h00000a85;
    rd_cycle[  125] = 1'b0;  wr_cycle[  125] = 1'b1;  addr_rom[  125]='h000001f4;  wr_data_rom[  125]='h00000572;
    rd_cycle[  126] = 1'b0;  wr_cycle[  126] = 1'b1;  addr_rom[  126]='h000001f8;  wr_data_rom[  126]='h00000ea5;
    rd_cycle[  127] = 1'b0;  wr_cycle[  127] = 1'b1;  addr_rom[  127]='h000001fc;  wr_data_rom[  127]='h000003ec;
    rd_cycle[  128] = 1'b0;  wr_cycle[  128] = 1'b1;  addr_rom[  128]='h00000200;  wr_data_rom[  128]='h00000a51;
    rd_cycle[  129] = 1'b0;  wr_cycle[  129] = 1'b1;  addr_rom[  129]='h00000204;  wr_data_rom[  129]='h0000082a;
    rd_cycle[  130] = 1'b0;  wr_cycle[  130] = 1'b1;  addr_rom[  130]='h00000208;  wr_data_rom[  130]='h00000e30;
    rd_cycle[  131] = 1'b0;  wr_cycle[  131] = 1'b1;  addr_rom[  131]='h0000020c;  wr_data_rom[  131]='h00000d19;
    rd_cycle[  132] = 1'b0;  wr_cycle[  132] = 1'b1;  addr_rom[  132]='h00000210;  wr_data_rom[  132]='h0000001b;
    rd_cycle[  133] = 1'b0;  wr_cycle[  133] = 1'b1;  addr_rom[  133]='h00000214;  wr_data_rom[  133]='h000003d0;
    rd_cycle[  134] = 1'b0;  wr_cycle[  134] = 1'b1;  addr_rom[  134]='h00000218;  wr_data_rom[  134]='h000003b5;
    rd_cycle[  135] = 1'b0;  wr_cycle[  135] = 1'b1;  addr_rom[  135]='h0000021c;  wr_data_rom[  135]='h00000da9;
    rd_cycle[  136] = 1'b0;  wr_cycle[  136] = 1'b1;  addr_rom[  136]='h00000220;  wr_data_rom[  136]='h00000c60;
    rd_cycle[  137] = 1'b0;  wr_cycle[  137] = 1'b1;  addr_rom[  137]='h00000224;  wr_data_rom[  137]='h000007e9;
    rd_cycle[  138] = 1'b0;  wr_cycle[  138] = 1'b1;  addr_rom[  138]='h00000228;  wr_data_rom[  138]='h00000749;
    rd_cycle[  139] = 1'b0;  wr_cycle[  139] = 1'b1;  addr_rom[  139]='h0000022c;  wr_data_rom[  139]='h0000099b;
    rd_cycle[  140] = 1'b0;  wr_cycle[  140] = 1'b1;  addr_rom[  140]='h00000230;  wr_data_rom[  140]='h00000c25;
    rd_cycle[  141] = 1'b0;  wr_cycle[  141] = 1'b1;  addr_rom[  141]='h00000234;  wr_data_rom[  141]='h00000158;
    rd_cycle[  142] = 1'b0;  wr_cycle[  142] = 1'b1;  addr_rom[  142]='h00000238;  wr_data_rom[  142]='h0000044e;
    rd_cycle[  143] = 1'b0;  wr_cycle[  143] = 1'b1;  addr_rom[  143]='h0000023c;  wr_data_rom[  143]='h000007e8;
    rd_cycle[  144] = 1'b0;  wr_cycle[  144] = 1'b1;  addr_rom[  144]='h00000240;  wr_data_rom[  144]='h00000967;
    rd_cycle[  145] = 1'b0;  wr_cycle[  145] = 1'b1;  addr_rom[  145]='h00000244;  wr_data_rom[  145]='h000006b9;
    rd_cycle[  146] = 1'b0;  wr_cycle[  146] = 1'b1;  addr_rom[  146]='h00000248;  wr_data_rom[  146]='h00000c99;
    rd_cycle[  147] = 1'b0;  wr_cycle[  147] = 1'b1;  addr_rom[  147]='h0000024c;  wr_data_rom[  147]='h00000cc4;
    rd_cycle[  148] = 1'b0;  wr_cycle[  148] = 1'b1;  addr_rom[  148]='h00000250;  wr_data_rom[  148]='h00000a6f;
    rd_cycle[  149] = 1'b0;  wr_cycle[  149] = 1'b1;  addr_rom[  149]='h00000254;  wr_data_rom[  149]='h000003a0;
    rd_cycle[  150] = 1'b0;  wr_cycle[  150] = 1'b1;  addr_rom[  150]='h00000258;  wr_data_rom[  150]='h0000014e;
    rd_cycle[  151] = 1'b0;  wr_cycle[  151] = 1'b1;  addr_rom[  151]='h0000025c;  wr_data_rom[  151]='h00000f2f;
    rd_cycle[  152] = 1'b0;  wr_cycle[  152] = 1'b1;  addr_rom[  152]='h00000260;  wr_data_rom[  152]='h00000588;
    rd_cycle[  153] = 1'b0;  wr_cycle[  153] = 1'b1;  addr_rom[  153]='h00000264;  wr_data_rom[  153]='h000007a6;
    rd_cycle[  154] = 1'b0;  wr_cycle[  154] = 1'b1;  addr_rom[  154]='h00000268;  wr_data_rom[  154]='h000006df;
    rd_cycle[  155] = 1'b0;  wr_cycle[  155] = 1'b1;  addr_rom[  155]='h0000026c;  wr_data_rom[  155]='h00000ad4;
    rd_cycle[  156] = 1'b0;  wr_cycle[  156] = 1'b1;  addr_rom[  156]='h00000270;  wr_data_rom[  156]='h00000604;
    rd_cycle[  157] = 1'b0;  wr_cycle[  157] = 1'b1;  addr_rom[  157]='h00000274;  wr_data_rom[  157]='h00000717;
    rd_cycle[  158] = 1'b0;  wr_cycle[  158] = 1'b1;  addr_rom[  158]='h00000278;  wr_data_rom[  158]='h00000243;
    rd_cycle[  159] = 1'b0;  wr_cycle[  159] = 1'b1;  addr_rom[  159]='h0000027c;  wr_data_rom[  159]='h000001bf;
    rd_cycle[  160] = 1'b0;  wr_cycle[  160] = 1'b1;  addr_rom[  160]='h00000280;  wr_data_rom[  160]='h000004dc;
    rd_cycle[  161] = 1'b0;  wr_cycle[  161] = 1'b1;  addr_rom[  161]='h00000284;  wr_data_rom[  161]='h00000102;
    rd_cycle[  162] = 1'b0;  wr_cycle[  162] = 1'b1;  addr_rom[  162]='h00000288;  wr_data_rom[  162]='h0000020b;
    rd_cycle[  163] = 1'b0;  wr_cycle[  163] = 1'b1;  addr_rom[  163]='h0000028c;  wr_data_rom[  163]='h00000165;
    rd_cycle[  164] = 1'b0;  wr_cycle[  164] = 1'b1;  addr_rom[  164]='h00000290;  wr_data_rom[  164]='h000009fd;
    rd_cycle[  165] = 1'b0;  wr_cycle[  165] = 1'b1;  addr_rom[  165]='h00000294;  wr_data_rom[  165]='h00000117;
    rd_cycle[  166] = 1'b0;  wr_cycle[  166] = 1'b1;  addr_rom[  166]='h00000298;  wr_data_rom[  166]='h00000495;
    rd_cycle[  167] = 1'b0;  wr_cycle[  167] = 1'b1;  addr_rom[  167]='h0000029c;  wr_data_rom[  167]='h00000af4;
    rd_cycle[  168] = 1'b0;  wr_cycle[  168] = 1'b1;  addr_rom[  168]='h000002a0;  wr_data_rom[  168]='h000002c0;
    rd_cycle[  169] = 1'b0;  wr_cycle[  169] = 1'b1;  addr_rom[  169]='h000002a4;  wr_data_rom[  169]='h000007e5;
    rd_cycle[  170] = 1'b0;  wr_cycle[  170] = 1'b1;  addr_rom[  170]='h000002a8;  wr_data_rom[  170]='h00000b7b;
    rd_cycle[  171] = 1'b0;  wr_cycle[  171] = 1'b1;  addr_rom[  171]='h000002ac;  wr_data_rom[  171]='h00000c11;
    rd_cycle[  172] = 1'b0;  wr_cycle[  172] = 1'b1;  addr_rom[  172]='h000002b0;  wr_data_rom[  172]='h00000d81;
    rd_cycle[  173] = 1'b0;  wr_cycle[  173] = 1'b1;  addr_rom[  173]='h000002b4;  wr_data_rom[  173]='h00000d4c;
    rd_cycle[  174] = 1'b0;  wr_cycle[  174] = 1'b1;  addr_rom[  174]='h000002b8;  wr_data_rom[  174]='h000008d9;
    rd_cycle[  175] = 1'b0;  wr_cycle[  175] = 1'b1;  addr_rom[  175]='h000002bc;  wr_data_rom[  175]='h00000e6d;
    rd_cycle[  176] = 1'b0;  wr_cycle[  176] = 1'b1;  addr_rom[  176]='h000002c0;  wr_data_rom[  176]='h00000f4a;
    rd_cycle[  177] = 1'b0;  wr_cycle[  177] = 1'b1;  addr_rom[  177]='h000002c4;  wr_data_rom[  177]='h00000713;
    rd_cycle[  178] = 1'b0;  wr_cycle[  178] = 1'b1;  addr_rom[  178]='h000002c8;  wr_data_rom[  178]='h00000698;
    rd_cycle[  179] = 1'b0;  wr_cycle[  179] = 1'b1;  addr_rom[  179]='h000002cc;  wr_data_rom[  179]='h00000e2e;
    rd_cycle[  180] = 1'b0;  wr_cycle[  180] = 1'b1;  addr_rom[  180]='h000002d0;  wr_data_rom[  180]='h00000056;
    rd_cycle[  181] = 1'b0;  wr_cycle[  181] = 1'b1;  addr_rom[  181]='h000002d4;  wr_data_rom[  181]='h0000090e;
    rd_cycle[  182] = 1'b0;  wr_cycle[  182] = 1'b1;  addr_rom[  182]='h000002d8;  wr_data_rom[  182]='h0000037b;
    rd_cycle[  183] = 1'b0;  wr_cycle[  183] = 1'b1;  addr_rom[  183]='h000002dc;  wr_data_rom[  183]='h00000979;
    rd_cycle[  184] = 1'b0;  wr_cycle[  184] = 1'b1;  addr_rom[  184]='h000002e0;  wr_data_rom[  184]='h00000a02;
    rd_cycle[  185] = 1'b0;  wr_cycle[  185] = 1'b1;  addr_rom[  185]='h000002e4;  wr_data_rom[  185]='h00000c53;
    rd_cycle[  186] = 1'b0;  wr_cycle[  186] = 1'b1;  addr_rom[  186]='h000002e8;  wr_data_rom[  186]='h00000c71;
    rd_cycle[  187] = 1'b0;  wr_cycle[  187] = 1'b1;  addr_rom[  187]='h000002ec;  wr_data_rom[  187]='h00000750;
    rd_cycle[  188] = 1'b0;  wr_cycle[  188] = 1'b1;  addr_rom[  188]='h000002f0;  wr_data_rom[  188]='h0000093b;
    rd_cycle[  189] = 1'b0;  wr_cycle[  189] = 1'b1;  addr_rom[  189]='h000002f4;  wr_data_rom[  189]='h00000ce9;
    rd_cycle[  190] = 1'b0;  wr_cycle[  190] = 1'b1;  addr_rom[  190]='h000002f8;  wr_data_rom[  190]='h00000609;
    rd_cycle[  191] = 1'b0;  wr_cycle[  191] = 1'b1;  addr_rom[  191]='h000002fc;  wr_data_rom[  191]='h00000b83;
    rd_cycle[  192] = 1'b0;  wr_cycle[  192] = 1'b1;  addr_rom[  192]='h00000300;  wr_data_rom[  192]='h00000115;
    rd_cycle[  193] = 1'b0;  wr_cycle[  193] = 1'b1;  addr_rom[  193]='h00000304;  wr_data_rom[  193]='h00000bb3;
    rd_cycle[  194] = 1'b0;  wr_cycle[  194] = 1'b1;  addr_rom[  194]='h00000308;  wr_data_rom[  194]='h0000086a;
    rd_cycle[  195] = 1'b0;  wr_cycle[  195] = 1'b1;  addr_rom[  195]='h0000030c;  wr_data_rom[  195]='h00000ee5;
    rd_cycle[  196] = 1'b0;  wr_cycle[  196] = 1'b1;  addr_rom[  196]='h00000310;  wr_data_rom[  196]='h000001fb;
    rd_cycle[  197] = 1'b0;  wr_cycle[  197] = 1'b1;  addr_rom[  197]='h00000314;  wr_data_rom[  197]='h0000065d;
    rd_cycle[  198] = 1'b0;  wr_cycle[  198] = 1'b1;  addr_rom[  198]='h00000318;  wr_data_rom[  198]='h00000b63;
    rd_cycle[  199] = 1'b0;  wr_cycle[  199] = 1'b1;  addr_rom[  199]='h0000031c;  wr_data_rom[  199]='h00000915;
    rd_cycle[  200] = 1'b0;  wr_cycle[  200] = 1'b1;  addr_rom[  200]='h00000320;  wr_data_rom[  200]='h0000095c;
    rd_cycle[  201] = 1'b0;  wr_cycle[  201] = 1'b1;  addr_rom[  201]='h00000324;  wr_data_rom[  201]='h0000064a;
    rd_cycle[  202] = 1'b0;  wr_cycle[  202] = 1'b1;  addr_rom[  202]='h00000328;  wr_data_rom[  202]='h00000c55;
    rd_cycle[  203] = 1'b0;  wr_cycle[  203] = 1'b1;  addr_rom[  203]='h0000032c;  wr_data_rom[  203]='h00000224;
    rd_cycle[  204] = 1'b0;  wr_cycle[  204] = 1'b1;  addr_rom[  204]='h00000330;  wr_data_rom[  204]='h00000462;
    rd_cycle[  205] = 1'b0;  wr_cycle[  205] = 1'b1;  addr_rom[  205]='h00000334;  wr_data_rom[  205]='h000006e9;
    rd_cycle[  206] = 1'b0;  wr_cycle[  206] = 1'b1;  addr_rom[  206]='h00000338;  wr_data_rom[  206]='h00000133;
    rd_cycle[  207] = 1'b0;  wr_cycle[  207] = 1'b1;  addr_rom[  207]='h0000033c;  wr_data_rom[  207]='h000009c4;
    rd_cycle[  208] = 1'b0;  wr_cycle[  208] = 1'b1;  addr_rom[  208]='h00000340;  wr_data_rom[  208]='h00000877;
    rd_cycle[  209] = 1'b0;  wr_cycle[  209] = 1'b1;  addr_rom[  209]='h00000344;  wr_data_rom[  209]='h0000091a;
    rd_cycle[  210] = 1'b0;  wr_cycle[  210] = 1'b1;  addr_rom[  210]='h00000348;  wr_data_rom[  210]='h00000c67;
    rd_cycle[  211] = 1'b0;  wr_cycle[  211] = 1'b1;  addr_rom[  211]='h0000034c;  wr_data_rom[  211]='h00000692;
    rd_cycle[  212] = 1'b0;  wr_cycle[  212] = 1'b1;  addr_rom[  212]='h00000350;  wr_data_rom[  212]='h00000383;
    rd_cycle[  213] = 1'b0;  wr_cycle[  213] = 1'b1;  addr_rom[  213]='h00000354;  wr_data_rom[  213]='h000003e8;
    rd_cycle[  214] = 1'b0;  wr_cycle[  214] = 1'b1;  addr_rom[  214]='h00000358;  wr_data_rom[  214]='h00000d38;
    rd_cycle[  215] = 1'b0;  wr_cycle[  215] = 1'b1;  addr_rom[  215]='h0000035c;  wr_data_rom[  215]='h00000118;
    rd_cycle[  216] = 1'b0;  wr_cycle[  216] = 1'b1;  addr_rom[  216]='h00000360;  wr_data_rom[  216]='h0000088f;
    rd_cycle[  217] = 1'b0;  wr_cycle[  217] = 1'b1;  addr_rom[  217]='h00000364;  wr_data_rom[  217]='h0000012c;
    rd_cycle[  218] = 1'b0;  wr_cycle[  218] = 1'b1;  addr_rom[  218]='h00000368;  wr_data_rom[  218]='h00000117;
    rd_cycle[  219] = 1'b0;  wr_cycle[  219] = 1'b1;  addr_rom[  219]='h0000036c;  wr_data_rom[  219]='h00000a71;
    rd_cycle[  220] = 1'b0;  wr_cycle[  220] = 1'b1;  addr_rom[  220]='h00000370;  wr_data_rom[  220]='h00000d32;
    rd_cycle[  221] = 1'b0;  wr_cycle[  221] = 1'b1;  addr_rom[  221]='h00000374;  wr_data_rom[  221]='h00000f07;
    rd_cycle[  222] = 1'b0;  wr_cycle[  222] = 1'b1;  addr_rom[  222]='h00000378;  wr_data_rom[  222]='h000006de;
    rd_cycle[  223] = 1'b0;  wr_cycle[  223] = 1'b1;  addr_rom[  223]='h0000037c;  wr_data_rom[  223]='h00000932;
    rd_cycle[  224] = 1'b0;  wr_cycle[  224] = 1'b1;  addr_rom[  224]='h00000380;  wr_data_rom[  224]='h00000233;
    rd_cycle[  225] = 1'b0;  wr_cycle[  225] = 1'b1;  addr_rom[  225]='h00000384;  wr_data_rom[  225]='h000006e1;
    rd_cycle[  226] = 1'b0;  wr_cycle[  226] = 1'b1;  addr_rom[  226]='h00000388;  wr_data_rom[  226]='h00000d5f;
    rd_cycle[  227] = 1'b0;  wr_cycle[  227] = 1'b1;  addr_rom[  227]='h0000038c;  wr_data_rom[  227]='h0000028a;
    rd_cycle[  228] = 1'b0;  wr_cycle[  228] = 1'b1;  addr_rom[  228]='h00000390;  wr_data_rom[  228]='h000009f1;
    rd_cycle[  229] = 1'b0;  wr_cycle[  229] = 1'b1;  addr_rom[  229]='h00000394;  wr_data_rom[  229]='h000007b4;
    rd_cycle[  230] = 1'b0;  wr_cycle[  230] = 1'b1;  addr_rom[  230]='h00000398;  wr_data_rom[  230]='h00000c7c;
    rd_cycle[  231] = 1'b0;  wr_cycle[  231] = 1'b1;  addr_rom[  231]='h0000039c;  wr_data_rom[  231]='h0000055f;
    rd_cycle[  232] = 1'b0;  wr_cycle[  232] = 1'b1;  addr_rom[  232]='h000003a0;  wr_data_rom[  232]='h00000082;
    rd_cycle[  233] = 1'b0;  wr_cycle[  233] = 1'b1;  addr_rom[  233]='h000003a4;  wr_data_rom[  233]='h00000679;
    rd_cycle[  234] = 1'b0;  wr_cycle[  234] = 1'b1;  addr_rom[  234]='h000003a8;  wr_data_rom[  234]='h0000028f;
    rd_cycle[  235] = 1'b0;  wr_cycle[  235] = 1'b1;  addr_rom[  235]='h000003ac;  wr_data_rom[  235]='h000009a0;
    rd_cycle[  236] = 1'b0;  wr_cycle[  236] = 1'b1;  addr_rom[  236]='h000003b0;  wr_data_rom[  236]='h00000f25;
    rd_cycle[  237] = 1'b0;  wr_cycle[  237] = 1'b1;  addr_rom[  237]='h000003b4;  wr_data_rom[  237]='h00000085;
    rd_cycle[  238] = 1'b0;  wr_cycle[  238] = 1'b1;  addr_rom[  238]='h000003b8;  wr_data_rom[  238]='h000006a7;
    rd_cycle[  239] = 1'b0;  wr_cycle[  239] = 1'b1;  addr_rom[  239]='h000003bc;  wr_data_rom[  239]='h00000519;
    rd_cycle[  240] = 1'b0;  wr_cycle[  240] = 1'b1;  addr_rom[  240]='h000003c0;  wr_data_rom[  240]='h00000f33;
    rd_cycle[  241] = 1'b0;  wr_cycle[  241] = 1'b1;  addr_rom[  241]='h000003c4;  wr_data_rom[  241]='h000007a4;
    rd_cycle[  242] = 1'b0;  wr_cycle[  242] = 1'b1;  addr_rom[  242]='h000003c8;  wr_data_rom[  242]='h00000508;
    rd_cycle[  243] = 1'b0;  wr_cycle[  243] = 1'b1;  addr_rom[  243]='h000003cc;  wr_data_rom[  243]='h00000185;
    rd_cycle[  244] = 1'b0;  wr_cycle[  244] = 1'b1;  addr_rom[  244]='h000003d0;  wr_data_rom[  244]='h00000948;
    rd_cycle[  245] = 1'b0;  wr_cycle[  245] = 1'b1;  addr_rom[  245]='h000003d4;  wr_data_rom[  245]='h000000e1;
    rd_cycle[  246] = 1'b0;  wr_cycle[  246] = 1'b1;  addr_rom[  246]='h000003d8;  wr_data_rom[  246]='h000008d3;
    rd_cycle[  247] = 1'b0;  wr_cycle[  247] = 1'b1;  addr_rom[  247]='h000003dc;  wr_data_rom[  247]='h000008bb;
    rd_cycle[  248] = 1'b0;  wr_cycle[  248] = 1'b1;  addr_rom[  248]='h000003e0;  wr_data_rom[  248]='h00000cc8;
    rd_cycle[  249] = 1'b0;  wr_cycle[  249] = 1'b1;  addr_rom[  249]='h000003e4;  wr_data_rom[  249]='h00000d1c;
    rd_cycle[  250] = 1'b0;  wr_cycle[  250] = 1'b1;  addr_rom[  250]='h000003e8;  wr_data_rom[  250]='h00000908;
    rd_cycle[  251] = 1'b0;  wr_cycle[  251] = 1'b1;  addr_rom[  251]='h000003ec;  wr_data_rom[  251]='h000006ac;
    rd_cycle[  252] = 1'b0;  wr_cycle[  252] = 1'b1;  addr_rom[  252]='h000003f0;  wr_data_rom[  252]='h00000f88;
    rd_cycle[  253] = 1'b0;  wr_cycle[  253] = 1'b1;  addr_rom[  253]='h000003f4;  wr_data_rom[  253]='h000003bb;
    rd_cycle[  254] = 1'b0;  wr_cycle[  254] = 1'b1;  addr_rom[  254]='h000003f8;  wr_data_rom[  254]='h00000489;
    rd_cycle[  255] = 1'b0;  wr_cycle[  255] = 1'b1;  addr_rom[  255]='h000003fc;  wr_data_rom[  255]='h00000b11;
    rd_cycle[  256] = 1'b0;  wr_cycle[  256] = 1'b1;  addr_rom[  256]='h00000400;  wr_data_rom[  256]='h00000e34;
    rd_cycle[  257] = 1'b0;  wr_cycle[  257] = 1'b1;  addr_rom[  257]='h00000404;  wr_data_rom[  257]='h00000786;
    rd_cycle[  258] = 1'b0;  wr_cycle[  258] = 1'b1;  addr_rom[  258]='h00000408;  wr_data_rom[  258]='h0000050d;
    rd_cycle[  259] = 1'b0;  wr_cycle[  259] = 1'b1;  addr_rom[  259]='h0000040c;  wr_data_rom[  259]='h000009b7;
    rd_cycle[  260] = 1'b0;  wr_cycle[  260] = 1'b1;  addr_rom[  260]='h00000410;  wr_data_rom[  260]='h00000560;
    rd_cycle[  261] = 1'b0;  wr_cycle[  261] = 1'b1;  addr_rom[  261]='h00000414;  wr_data_rom[  261]='h000005c3;
    rd_cycle[  262] = 1'b0;  wr_cycle[  262] = 1'b1;  addr_rom[  262]='h00000418;  wr_data_rom[  262]='h000008cd;
    rd_cycle[  263] = 1'b0;  wr_cycle[  263] = 1'b1;  addr_rom[  263]='h0000041c;  wr_data_rom[  263]='h00000973;
    rd_cycle[  264] = 1'b0;  wr_cycle[  264] = 1'b1;  addr_rom[  264]='h00000420;  wr_data_rom[  264]='h00000715;
    rd_cycle[  265] = 1'b0;  wr_cycle[  265] = 1'b1;  addr_rom[  265]='h00000424;  wr_data_rom[  265]='h00000933;
    rd_cycle[  266] = 1'b0;  wr_cycle[  266] = 1'b1;  addr_rom[  266]='h00000428;  wr_data_rom[  266]='h00000900;
    rd_cycle[  267] = 1'b0;  wr_cycle[  267] = 1'b1;  addr_rom[  267]='h0000042c;  wr_data_rom[  267]='h000009b2;
    rd_cycle[  268] = 1'b0;  wr_cycle[  268] = 1'b1;  addr_rom[  268]='h00000430;  wr_data_rom[  268]='h00000d6c;
    rd_cycle[  269] = 1'b0;  wr_cycle[  269] = 1'b1;  addr_rom[  269]='h00000434;  wr_data_rom[  269]='h00000381;
    rd_cycle[  270] = 1'b0;  wr_cycle[  270] = 1'b1;  addr_rom[  270]='h00000438;  wr_data_rom[  270]='h00000c9a;
    rd_cycle[  271] = 1'b0;  wr_cycle[  271] = 1'b1;  addr_rom[  271]='h0000043c;  wr_data_rom[  271]='h00000268;
    rd_cycle[  272] = 1'b0;  wr_cycle[  272] = 1'b1;  addr_rom[  272]='h00000440;  wr_data_rom[  272]='h0000060a;
    rd_cycle[  273] = 1'b0;  wr_cycle[  273] = 1'b1;  addr_rom[  273]='h00000444;  wr_data_rom[  273]='h00000aa1;
    rd_cycle[  274] = 1'b0;  wr_cycle[  274] = 1'b1;  addr_rom[  274]='h00000448;  wr_data_rom[  274]='h00000b26;
    rd_cycle[  275] = 1'b0;  wr_cycle[  275] = 1'b1;  addr_rom[  275]='h0000044c;  wr_data_rom[  275]='h00000f00;
    rd_cycle[  276] = 1'b0;  wr_cycle[  276] = 1'b1;  addr_rom[  276]='h00000450;  wr_data_rom[  276]='h00000efd;
    rd_cycle[  277] = 1'b0;  wr_cycle[  277] = 1'b1;  addr_rom[  277]='h00000454;  wr_data_rom[  277]='h0000039c;
    rd_cycle[  278] = 1'b0;  wr_cycle[  278] = 1'b1;  addr_rom[  278]='h00000458;  wr_data_rom[  278]='h00000100;
    rd_cycle[  279] = 1'b0;  wr_cycle[  279] = 1'b1;  addr_rom[  279]='h0000045c;  wr_data_rom[  279]='h00000919;
    rd_cycle[  280] = 1'b0;  wr_cycle[  280] = 1'b1;  addr_rom[  280]='h00000460;  wr_data_rom[  280]='h00000333;
    rd_cycle[  281] = 1'b0;  wr_cycle[  281] = 1'b1;  addr_rom[  281]='h00000464;  wr_data_rom[  281]='h00000a93;
    rd_cycle[  282] = 1'b0;  wr_cycle[  282] = 1'b1;  addr_rom[  282]='h00000468;  wr_data_rom[  282]='h00000b0d;
    rd_cycle[  283] = 1'b0;  wr_cycle[  283] = 1'b1;  addr_rom[  283]='h0000046c;  wr_data_rom[  283]='h0000097c;
    rd_cycle[  284] = 1'b0;  wr_cycle[  284] = 1'b1;  addr_rom[  284]='h00000470;  wr_data_rom[  284]='h000000d6;
    rd_cycle[  285] = 1'b0;  wr_cycle[  285] = 1'b1;  addr_rom[  285]='h00000474;  wr_data_rom[  285]='h000009d6;
    rd_cycle[  286] = 1'b0;  wr_cycle[  286] = 1'b1;  addr_rom[  286]='h00000478;  wr_data_rom[  286]='h00000de4;
    rd_cycle[  287] = 1'b0;  wr_cycle[  287] = 1'b1;  addr_rom[  287]='h0000047c;  wr_data_rom[  287]='h0000085e;
    rd_cycle[  288] = 1'b0;  wr_cycle[  288] = 1'b1;  addr_rom[  288]='h00000480;  wr_data_rom[  288]='h000004da;
    rd_cycle[  289] = 1'b0;  wr_cycle[  289] = 1'b1;  addr_rom[  289]='h00000484;  wr_data_rom[  289]='h00000dc9;
    rd_cycle[  290] = 1'b0;  wr_cycle[  290] = 1'b1;  addr_rom[  290]='h00000488;  wr_data_rom[  290]='h00000b36;
    rd_cycle[  291] = 1'b0;  wr_cycle[  291] = 1'b1;  addr_rom[  291]='h0000048c;  wr_data_rom[  291]='h000008cf;
    rd_cycle[  292] = 1'b0;  wr_cycle[  292] = 1'b1;  addr_rom[  292]='h00000490;  wr_data_rom[  292]='h000007ea;
    rd_cycle[  293] = 1'b0;  wr_cycle[  293] = 1'b1;  addr_rom[  293]='h00000494;  wr_data_rom[  293]='h00000653;
    rd_cycle[  294] = 1'b0;  wr_cycle[  294] = 1'b1;  addr_rom[  294]='h00000498;  wr_data_rom[  294]='h000005a7;
    rd_cycle[  295] = 1'b0;  wr_cycle[  295] = 1'b1;  addr_rom[  295]='h0000049c;  wr_data_rom[  295]='h00000681;
    rd_cycle[  296] = 1'b0;  wr_cycle[  296] = 1'b1;  addr_rom[  296]='h000004a0;  wr_data_rom[  296]='h0000005f;
    rd_cycle[  297] = 1'b0;  wr_cycle[  297] = 1'b1;  addr_rom[  297]='h000004a4;  wr_data_rom[  297]='h00000315;
    rd_cycle[  298] = 1'b0;  wr_cycle[  298] = 1'b1;  addr_rom[  298]='h000004a8;  wr_data_rom[  298]='h000003aa;
    rd_cycle[  299] = 1'b0;  wr_cycle[  299] = 1'b1;  addr_rom[  299]='h000004ac;  wr_data_rom[  299]='h00000564;
    rd_cycle[  300] = 1'b0;  wr_cycle[  300] = 1'b1;  addr_rom[  300]='h000004b0;  wr_data_rom[  300]='h00000b43;
    rd_cycle[  301] = 1'b0;  wr_cycle[  301] = 1'b1;  addr_rom[  301]='h000004b4;  wr_data_rom[  301]='h00000040;
    rd_cycle[  302] = 1'b0;  wr_cycle[  302] = 1'b1;  addr_rom[  302]='h000004b8;  wr_data_rom[  302]='h00000d76;
    rd_cycle[  303] = 1'b0;  wr_cycle[  303] = 1'b1;  addr_rom[  303]='h000004bc;  wr_data_rom[  303]='h00000ae6;
    rd_cycle[  304] = 1'b0;  wr_cycle[  304] = 1'b1;  addr_rom[  304]='h000004c0;  wr_data_rom[  304]='h00000a3d;
    rd_cycle[  305] = 1'b0;  wr_cycle[  305] = 1'b1;  addr_rom[  305]='h000004c4;  wr_data_rom[  305]='h00000a1d;
    rd_cycle[  306] = 1'b0;  wr_cycle[  306] = 1'b1;  addr_rom[  306]='h000004c8;  wr_data_rom[  306]='h00000a75;
    rd_cycle[  307] = 1'b0;  wr_cycle[  307] = 1'b1;  addr_rom[  307]='h000004cc;  wr_data_rom[  307]='h000003d2;
    rd_cycle[  308] = 1'b0;  wr_cycle[  308] = 1'b1;  addr_rom[  308]='h000004d0;  wr_data_rom[  308]='h00000d55;
    rd_cycle[  309] = 1'b0;  wr_cycle[  309] = 1'b1;  addr_rom[  309]='h000004d4;  wr_data_rom[  309]='h00000563;
    rd_cycle[  310] = 1'b0;  wr_cycle[  310] = 1'b1;  addr_rom[  310]='h000004d8;  wr_data_rom[  310]='h00000ac5;
    rd_cycle[  311] = 1'b0;  wr_cycle[  311] = 1'b1;  addr_rom[  311]='h000004dc;  wr_data_rom[  311]='h00000404;
    rd_cycle[  312] = 1'b0;  wr_cycle[  312] = 1'b1;  addr_rom[  312]='h000004e0;  wr_data_rom[  312]='h00000d33;
    rd_cycle[  313] = 1'b0;  wr_cycle[  313] = 1'b1;  addr_rom[  313]='h000004e4;  wr_data_rom[  313]='h000006c6;
    rd_cycle[  314] = 1'b0;  wr_cycle[  314] = 1'b1;  addr_rom[  314]='h000004e8;  wr_data_rom[  314]='h00000b60;
    rd_cycle[  315] = 1'b0;  wr_cycle[  315] = 1'b1;  addr_rom[  315]='h000004ec;  wr_data_rom[  315]='h000008d3;
    rd_cycle[  316] = 1'b0;  wr_cycle[  316] = 1'b1;  addr_rom[  316]='h000004f0;  wr_data_rom[  316]='h000000ac;
    rd_cycle[  317] = 1'b0;  wr_cycle[  317] = 1'b1;  addr_rom[  317]='h000004f4;  wr_data_rom[  317]='h000003a0;
    rd_cycle[  318] = 1'b0;  wr_cycle[  318] = 1'b1;  addr_rom[  318]='h000004f8;  wr_data_rom[  318]='h00000737;
    rd_cycle[  319] = 1'b0;  wr_cycle[  319] = 1'b1;  addr_rom[  319]='h000004fc;  wr_data_rom[  319]='h00000631;
    rd_cycle[  320] = 1'b0;  wr_cycle[  320] = 1'b1;  addr_rom[  320]='h00000500;  wr_data_rom[  320]='h0000099b;
    rd_cycle[  321] = 1'b0;  wr_cycle[  321] = 1'b1;  addr_rom[  321]='h00000504;  wr_data_rom[  321]='h00000539;
    rd_cycle[  322] = 1'b0;  wr_cycle[  322] = 1'b1;  addr_rom[  322]='h00000508;  wr_data_rom[  322]='h000000ab;
    rd_cycle[  323] = 1'b0;  wr_cycle[  323] = 1'b1;  addr_rom[  323]='h0000050c;  wr_data_rom[  323]='h00000e7b;
    rd_cycle[  324] = 1'b0;  wr_cycle[  324] = 1'b1;  addr_rom[  324]='h00000510;  wr_data_rom[  324]='h00000d9d;
    rd_cycle[  325] = 1'b0;  wr_cycle[  325] = 1'b1;  addr_rom[  325]='h00000514;  wr_data_rom[  325]='h00000278;
    rd_cycle[  326] = 1'b0;  wr_cycle[  326] = 1'b1;  addr_rom[  326]='h00000518;  wr_data_rom[  326]='h00000ede;
    rd_cycle[  327] = 1'b0;  wr_cycle[  327] = 1'b1;  addr_rom[  327]='h0000051c;  wr_data_rom[  327]='h00000ef5;
    rd_cycle[  328] = 1'b0;  wr_cycle[  328] = 1'b1;  addr_rom[  328]='h00000520;  wr_data_rom[  328]='h00000004;
    rd_cycle[  329] = 1'b0;  wr_cycle[  329] = 1'b1;  addr_rom[  329]='h00000524;  wr_data_rom[  329]='h00000238;
    rd_cycle[  330] = 1'b0;  wr_cycle[  330] = 1'b1;  addr_rom[  330]='h00000528;  wr_data_rom[  330]='h000009af;
    rd_cycle[  331] = 1'b0;  wr_cycle[  331] = 1'b1;  addr_rom[  331]='h0000052c;  wr_data_rom[  331]='h0000071b;
    rd_cycle[  332] = 1'b0;  wr_cycle[  332] = 1'b1;  addr_rom[  332]='h00000530;  wr_data_rom[  332]='h00000c62;
    rd_cycle[  333] = 1'b0;  wr_cycle[  333] = 1'b1;  addr_rom[  333]='h00000534;  wr_data_rom[  333]='h00000d6d;
    rd_cycle[  334] = 1'b0;  wr_cycle[  334] = 1'b1;  addr_rom[  334]='h00000538;  wr_data_rom[  334]='h00000cf7;
    rd_cycle[  335] = 1'b0;  wr_cycle[  335] = 1'b1;  addr_rom[  335]='h0000053c;  wr_data_rom[  335]='h00000828;
    rd_cycle[  336] = 1'b0;  wr_cycle[  336] = 1'b1;  addr_rom[  336]='h00000540;  wr_data_rom[  336]='h0000061c;
    rd_cycle[  337] = 1'b0;  wr_cycle[  337] = 1'b1;  addr_rom[  337]='h00000544;  wr_data_rom[  337]='h00000f79;
    rd_cycle[  338] = 1'b0;  wr_cycle[  338] = 1'b1;  addr_rom[  338]='h00000548;  wr_data_rom[  338]='h00000f78;
    rd_cycle[  339] = 1'b0;  wr_cycle[  339] = 1'b1;  addr_rom[  339]='h0000054c;  wr_data_rom[  339]='h000001cf;
    rd_cycle[  340] = 1'b0;  wr_cycle[  340] = 1'b1;  addr_rom[  340]='h00000550;  wr_data_rom[  340]='h00000944;
    rd_cycle[  341] = 1'b0;  wr_cycle[  341] = 1'b1;  addr_rom[  341]='h00000554;  wr_data_rom[  341]='h000008ba;
    rd_cycle[  342] = 1'b0;  wr_cycle[  342] = 1'b1;  addr_rom[  342]='h00000558;  wr_data_rom[  342]='h000001dc;
    rd_cycle[  343] = 1'b0;  wr_cycle[  343] = 1'b1;  addr_rom[  343]='h0000055c;  wr_data_rom[  343]='h000004ca;
    rd_cycle[  344] = 1'b0;  wr_cycle[  344] = 1'b1;  addr_rom[  344]='h00000560;  wr_data_rom[  344]='h00000228;
    rd_cycle[  345] = 1'b0;  wr_cycle[  345] = 1'b1;  addr_rom[  345]='h00000564;  wr_data_rom[  345]='h000007a7;
    rd_cycle[  346] = 1'b0;  wr_cycle[  346] = 1'b1;  addr_rom[  346]='h00000568;  wr_data_rom[  346]='h0000023f;
    rd_cycle[  347] = 1'b0;  wr_cycle[  347] = 1'b1;  addr_rom[  347]='h0000056c;  wr_data_rom[  347]='h0000078b;
    rd_cycle[  348] = 1'b0;  wr_cycle[  348] = 1'b1;  addr_rom[  348]='h00000570;  wr_data_rom[  348]='h00000323;
    rd_cycle[  349] = 1'b0;  wr_cycle[  349] = 1'b1;  addr_rom[  349]='h00000574;  wr_data_rom[  349]='h00000444;
    rd_cycle[  350] = 1'b0;  wr_cycle[  350] = 1'b1;  addr_rom[  350]='h00000578;  wr_data_rom[  350]='h00000c69;
    rd_cycle[  351] = 1'b0;  wr_cycle[  351] = 1'b1;  addr_rom[  351]='h0000057c;  wr_data_rom[  351]='h000001dd;
    rd_cycle[  352] = 1'b0;  wr_cycle[  352] = 1'b1;  addr_rom[  352]='h00000580;  wr_data_rom[  352]='h00000cf4;
    rd_cycle[  353] = 1'b0;  wr_cycle[  353] = 1'b1;  addr_rom[  353]='h00000584;  wr_data_rom[  353]='h00000b2d;
    rd_cycle[  354] = 1'b0;  wr_cycle[  354] = 1'b1;  addr_rom[  354]='h00000588;  wr_data_rom[  354]='h0000094c;
    rd_cycle[  355] = 1'b0;  wr_cycle[  355] = 1'b1;  addr_rom[  355]='h0000058c;  wr_data_rom[  355]='h00000e81;
    rd_cycle[  356] = 1'b0;  wr_cycle[  356] = 1'b1;  addr_rom[  356]='h00000590;  wr_data_rom[  356]='h00000db5;
    rd_cycle[  357] = 1'b0;  wr_cycle[  357] = 1'b1;  addr_rom[  357]='h00000594;  wr_data_rom[  357]='h00000f8d;
    rd_cycle[  358] = 1'b0;  wr_cycle[  358] = 1'b1;  addr_rom[  358]='h00000598;  wr_data_rom[  358]='h000008fa;
    rd_cycle[  359] = 1'b0;  wr_cycle[  359] = 1'b1;  addr_rom[  359]='h0000059c;  wr_data_rom[  359]='h000000f9;
    rd_cycle[  360] = 1'b0;  wr_cycle[  360] = 1'b1;  addr_rom[  360]='h000005a0;  wr_data_rom[  360]='h00000e8c;
    rd_cycle[  361] = 1'b0;  wr_cycle[  361] = 1'b1;  addr_rom[  361]='h000005a4;  wr_data_rom[  361]='h000004a8;
    rd_cycle[  362] = 1'b0;  wr_cycle[  362] = 1'b1;  addr_rom[  362]='h000005a8;  wr_data_rom[  362]='h000002b7;
    rd_cycle[  363] = 1'b0;  wr_cycle[  363] = 1'b1;  addr_rom[  363]='h000005ac;  wr_data_rom[  363]='h000003ce;
    rd_cycle[  364] = 1'b0;  wr_cycle[  364] = 1'b1;  addr_rom[  364]='h000005b0;  wr_data_rom[  364]='h000003ca;
    rd_cycle[  365] = 1'b0;  wr_cycle[  365] = 1'b1;  addr_rom[  365]='h000005b4;  wr_data_rom[  365]='h00000a04;
    rd_cycle[  366] = 1'b0;  wr_cycle[  366] = 1'b1;  addr_rom[  366]='h000005b8;  wr_data_rom[  366]='h0000024e;
    rd_cycle[  367] = 1'b0;  wr_cycle[  367] = 1'b1;  addr_rom[  367]='h000005bc;  wr_data_rom[  367]='h000002f1;
    rd_cycle[  368] = 1'b0;  wr_cycle[  368] = 1'b1;  addr_rom[  368]='h000005c0;  wr_data_rom[  368]='h00000a0b;
    rd_cycle[  369] = 1'b0;  wr_cycle[  369] = 1'b1;  addr_rom[  369]='h000005c4;  wr_data_rom[  369]='h0000089c;
    rd_cycle[  370] = 1'b0;  wr_cycle[  370] = 1'b1;  addr_rom[  370]='h000005c8;  wr_data_rom[  370]='h00000e5c;
    rd_cycle[  371] = 1'b0;  wr_cycle[  371] = 1'b1;  addr_rom[  371]='h000005cc;  wr_data_rom[  371]='h0000041d;
    rd_cycle[  372] = 1'b0;  wr_cycle[  372] = 1'b1;  addr_rom[  372]='h000005d0;  wr_data_rom[  372]='h000002bd;
    rd_cycle[  373] = 1'b0;  wr_cycle[  373] = 1'b1;  addr_rom[  373]='h000005d4;  wr_data_rom[  373]='h0000020c;
    rd_cycle[  374] = 1'b0;  wr_cycle[  374] = 1'b1;  addr_rom[  374]='h000005d8;  wr_data_rom[  374]='h000007ea;
    rd_cycle[  375] = 1'b0;  wr_cycle[  375] = 1'b1;  addr_rom[  375]='h000005dc;  wr_data_rom[  375]='h0000038d;
    rd_cycle[  376] = 1'b0;  wr_cycle[  376] = 1'b1;  addr_rom[  376]='h000005e0;  wr_data_rom[  376]='h00000e2c;
    rd_cycle[  377] = 1'b0;  wr_cycle[  377] = 1'b1;  addr_rom[  377]='h000005e4;  wr_data_rom[  377]='h000002cd;
    rd_cycle[  378] = 1'b0;  wr_cycle[  378] = 1'b1;  addr_rom[  378]='h000005e8;  wr_data_rom[  378]='h000008a0;
    rd_cycle[  379] = 1'b0;  wr_cycle[  379] = 1'b1;  addr_rom[  379]='h000005ec;  wr_data_rom[  379]='h00000f61;
    rd_cycle[  380] = 1'b0;  wr_cycle[  380] = 1'b1;  addr_rom[  380]='h000005f0;  wr_data_rom[  380]='h0000049b;
    rd_cycle[  381] = 1'b0;  wr_cycle[  381] = 1'b1;  addr_rom[  381]='h000005f4;  wr_data_rom[  381]='h00000def;
    rd_cycle[  382] = 1'b0;  wr_cycle[  382] = 1'b1;  addr_rom[  382]='h000005f8;  wr_data_rom[  382]='h0000000d;
    rd_cycle[  383] = 1'b0;  wr_cycle[  383] = 1'b1;  addr_rom[  383]='h000005fc;  wr_data_rom[  383]='h00000d35;
    rd_cycle[  384] = 1'b0;  wr_cycle[  384] = 1'b1;  addr_rom[  384]='h00000600;  wr_data_rom[  384]='h00000b4a;
    rd_cycle[  385] = 1'b0;  wr_cycle[  385] = 1'b1;  addr_rom[  385]='h00000604;  wr_data_rom[  385]='h000003d4;
    rd_cycle[  386] = 1'b0;  wr_cycle[  386] = 1'b1;  addr_rom[  386]='h00000608;  wr_data_rom[  386]='h00000298;
    rd_cycle[  387] = 1'b0;  wr_cycle[  387] = 1'b1;  addr_rom[  387]='h0000060c;  wr_data_rom[  387]='h0000059c;
    rd_cycle[  388] = 1'b0;  wr_cycle[  388] = 1'b1;  addr_rom[  388]='h00000610;  wr_data_rom[  388]='h000002f3;
    rd_cycle[  389] = 1'b0;  wr_cycle[  389] = 1'b1;  addr_rom[  389]='h00000614;  wr_data_rom[  389]='h0000078a;
    rd_cycle[  390] = 1'b0;  wr_cycle[  390] = 1'b1;  addr_rom[  390]='h00000618;  wr_data_rom[  390]='h000009c1;
    rd_cycle[  391] = 1'b0;  wr_cycle[  391] = 1'b1;  addr_rom[  391]='h0000061c;  wr_data_rom[  391]='h0000025b;
    rd_cycle[  392] = 1'b0;  wr_cycle[  392] = 1'b1;  addr_rom[  392]='h00000620;  wr_data_rom[  392]='h0000091b;
    rd_cycle[  393] = 1'b0;  wr_cycle[  393] = 1'b1;  addr_rom[  393]='h00000624;  wr_data_rom[  393]='h00000f3d;
    rd_cycle[  394] = 1'b0;  wr_cycle[  394] = 1'b1;  addr_rom[  394]='h00000628;  wr_data_rom[  394]='h000005c1;
    rd_cycle[  395] = 1'b0;  wr_cycle[  395] = 1'b1;  addr_rom[  395]='h0000062c;  wr_data_rom[  395]='h0000061d;
    rd_cycle[  396] = 1'b0;  wr_cycle[  396] = 1'b1;  addr_rom[  396]='h00000630;  wr_data_rom[  396]='h00000ebc;
    rd_cycle[  397] = 1'b0;  wr_cycle[  397] = 1'b1;  addr_rom[  397]='h00000634;  wr_data_rom[  397]='h00000513;
    rd_cycle[  398] = 1'b0;  wr_cycle[  398] = 1'b1;  addr_rom[  398]='h00000638;  wr_data_rom[  398]='h00000958;
    rd_cycle[  399] = 1'b0;  wr_cycle[  399] = 1'b1;  addr_rom[  399]='h0000063c;  wr_data_rom[  399]='h0000032c;
    rd_cycle[  400] = 1'b0;  wr_cycle[  400] = 1'b1;  addr_rom[  400]='h00000640;  wr_data_rom[  400]='h00000d85;
    rd_cycle[  401] = 1'b0;  wr_cycle[  401] = 1'b1;  addr_rom[  401]='h00000644;  wr_data_rom[  401]='h00000c12;
    rd_cycle[  402] = 1'b0;  wr_cycle[  402] = 1'b1;  addr_rom[  402]='h00000648;  wr_data_rom[  402]='h00000c65;
    rd_cycle[  403] = 1'b0;  wr_cycle[  403] = 1'b1;  addr_rom[  403]='h0000064c;  wr_data_rom[  403]='h000004c9;
    rd_cycle[  404] = 1'b0;  wr_cycle[  404] = 1'b1;  addr_rom[  404]='h00000650;  wr_data_rom[  404]='h00000487;
    rd_cycle[  405] = 1'b0;  wr_cycle[  405] = 1'b1;  addr_rom[  405]='h00000654;  wr_data_rom[  405]='h00000aa0;
    rd_cycle[  406] = 1'b0;  wr_cycle[  406] = 1'b1;  addr_rom[  406]='h00000658;  wr_data_rom[  406]='h00000b43;
    rd_cycle[  407] = 1'b0;  wr_cycle[  407] = 1'b1;  addr_rom[  407]='h0000065c;  wr_data_rom[  407]='h00000af6;
    rd_cycle[  408] = 1'b0;  wr_cycle[  408] = 1'b1;  addr_rom[  408]='h00000660;  wr_data_rom[  408]='h000008b0;
    rd_cycle[  409] = 1'b0;  wr_cycle[  409] = 1'b1;  addr_rom[  409]='h00000664;  wr_data_rom[  409]='h000006e7;
    rd_cycle[  410] = 1'b0;  wr_cycle[  410] = 1'b1;  addr_rom[  410]='h00000668;  wr_data_rom[  410]='h0000011e;
    rd_cycle[  411] = 1'b0;  wr_cycle[  411] = 1'b1;  addr_rom[  411]='h0000066c;  wr_data_rom[  411]='h00000f86;
    rd_cycle[  412] = 1'b0;  wr_cycle[  412] = 1'b1;  addr_rom[  412]='h00000670;  wr_data_rom[  412]='h00000ca2;
    rd_cycle[  413] = 1'b0;  wr_cycle[  413] = 1'b1;  addr_rom[  413]='h00000674;  wr_data_rom[  413]='h00000ae0;
    rd_cycle[  414] = 1'b0;  wr_cycle[  414] = 1'b1;  addr_rom[  414]='h00000678;  wr_data_rom[  414]='h00000843;
    rd_cycle[  415] = 1'b0;  wr_cycle[  415] = 1'b1;  addr_rom[  415]='h0000067c;  wr_data_rom[  415]='h00000634;
    rd_cycle[  416] = 1'b0;  wr_cycle[  416] = 1'b1;  addr_rom[  416]='h00000680;  wr_data_rom[  416]='h00000684;
    rd_cycle[  417] = 1'b0;  wr_cycle[  417] = 1'b1;  addr_rom[  417]='h00000684;  wr_data_rom[  417]='h00000619;
    rd_cycle[  418] = 1'b0;  wr_cycle[  418] = 1'b1;  addr_rom[  418]='h00000688;  wr_data_rom[  418]='h0000024d;
    rd_cycle[  419] = 1'b0;  wr_cycle[  419] = 1'b1;  addr_rom[  419]='h0000068c;  wr_data_rom[  419]='h00000f94;
    rd_cycle[  420] = 1'b0;  wr_cycle[  420] = 1'b1;  addr_rom[  420]='h00000690;  wr_data_rom[  420]='h00000506;
    rd_cycle[  421] = 1'b0;  wr_cycle[  421] = 1'b1;  addr_rom[  421]='h00000694;  wr_data_rom[  421]='h00000a7b;
    rd_cycle[  422] = 1'b0;  wr_cycle[  422] = 1'b1;  addr_rom[  422]='h00000698;  wr_data_rom[  422]='h00000eeb;
    rd_cycle[  423] = 1'b0;  wr_cycle[  423] = 1'b1;  addr_rom[  423]='h0000069c;  wr_data_rom[  423]='h000004c7;
    rd_cycle[  424] = 1'b0;  wr_cycle[  424] = 1'b1;  addr_rom[  424]='h000006a0;  wr_data_rom[  424]='h000001e4;
    rd_cycle[  425] = 1'b0;  wr_cycle[  425] = 1'b1;  addr_rom[  425]='h000006a4;  wr_data_rom[  425]='h00000a81;
    rd_cycle[  426] = 1'b0;  wr_cycle[  426] = 1'b1;  addr_rom[  426]='h000006a8;  wr_data_rom[  426]='h00000502;
    rd_cycle[  427] = 1'b0;  wr_cycle[  427] = 1'b1;  addr_rom[  427]='h000006ac;  wr_data_rom[  427]='h0000029f;
    rd_cycle[  428] = 1'b0;  wr_cycle[  428] = 1'b1;  addr_rom[  428]='h000006b0;  wr_data_rom[  428]='h00000071;
    rd_cycle[  429] = 1'b0;  wr_cycle[  429] = 1'b1;  addr_rom[  429]='h000006b4;  wr_data_rom[  429]='h000004d1;
    rd_cycle[  430] = 1'b0;  wr_cycle[  430] = 1'b1;  addr_rom[  430]='h000006b8;  wr_data_rom[  430]='h00000f63;
    rd_cycle[  431] = 1'b0;  wr_cycle[  431] = 1'b1;  addr_rom[  431]='h000006bc;  wr_data_rom[  431]='h00000bdb;
    rd_cycle[  432] = 1'b0;  wr_cycle[  432] = 1'b1;  addr_rom[  432]='h000006c0;  wr_data_rom[  432]='h00000c8d;
    rd_cycle[  433] = 1'b0;  wr_cycle[  433] = 1'b1;  addr_rom[  433]='h000006c4;  wr_data_rom[  433]='h000006a6;
    rd_cycle[  434] = 1'b0;  wr_cycle[  434] = 1'b1;  addr_rom[  434]='h000006c8;  wr_data_rom[  434]='h00000318;
    rd_cycle[  435] = 1'b0;  wr_cycle[  435] = 1'b1;  addr_rom[  435]='h000006cc;  wr_data_rom[  435]='h0000006b;
    rd_cycle[  436] = 1'b0;  wr_cycle[  436] = 1'b1;  addr_rom[  436]='h000006d0;  wr_data_rom[  436]='h00000378;
    rd_cycle[  437] = 1'b0;  wr_cycle[  437] = 1'b1;  addr_rom[  437]='h000006d4;  wr_data_rom[  437]='h0000000a;
    rd_cycle[  438] = 1'b0;  wr_cycle[  438] = 1'b1;  addr_rom[  438]='h000006d8;  wr_data_rom[  438]='h0000093b;
    rd_cycle[  439] = 1'b0;  wr_cycle[  439] = 1'b1;  addr_rom[  439]='h000006dc;  wr_data_rom[  439]='h00000115;
    rd_cycle[  440] = 1'b0;  wr_cycle[  440] = 1'b1;  addr_rom[  440]='h000006e0;  wr_data_rom[  440]='h00000f75;
    rd_cycle[  441] = 1'b0;  wr_cycle[  441] = 1'b1;  addr_rom[  441]='h000006e4;  wr_data_rom[  441]='h00000166;
    rd_cycle[  442] = 1'b0;  wr_cycle[  442] = 1'b1;  addr_rom[  442]='h000006e8;  wr_data_rom[  442]='h000008a9;
    rd_cycle[  443] = 1'b0;  wr_cycle[  443] = 1'b1;  addr_rom[  443]='h000006ec;  wr_data_rom[  443]='h00000347;
    rd_cycle[  444] = 1'b0;  wr_cycle[  444] = 1'b1;  addr_rom[  444]='h000006f0;  wr_data_rom[  444]='h00000d28;
    rd_cycle[  445] = 1'b0;  wr_cycle[  445] = 1'b1;  addr_rom[  445]='h000006f4;  wr_data_rom[  445]='h00000752;
    rd_cycle[  446] = 1'b0;  wr_cycle[  446] = 1'b1;  addr_rom[  446]='h000006f8;  wr_data_rom[  446]='h00000046;
    rd_cycle[  447] = 1'b0;  wr_cycle[  447] = 1'b1;  addr_rom[  447]='h000006fc;  wr_data_rom[  447]='h00000d4d;
    rd_cycle[  448] = 1'b0;  wr_cycle[  448] = 1'b1;  addr_rom[  448]='h00000700;  wr_data_rom[  448]='h00000591;
    rd_cycle[  449] = 1'b0;  wr_cycle[  449] = 1'b1;  addr_rom[  449]='h00000704;  wr_data_rom[  449]='h000009c4;
    rd_cycle[  450] = 1'b0;  wr_cycle[  450] = 1'b1;  addr_rom[  450]='h00000708;  wr_data_rom[  450]='h000000e9;
    rd_cycle[  451] = 1'b0;  wr_cycle[  451] = 1'b1;  addr_rom[  451]='h0000070c;  wr_data_rom[  451]='h00000892;
    rd_cycle[  452] = 1'b0;  wr_cycle[  452] = 1'b1;  addr_rom[  452]='h00000710;  wr_data_rom[  452]='h00000aee;
    rd_cycle[  453] = 1'b0;  wr_cycle[  453] = 1'b1;  addr_rom[  453]='h00000714;  wr_data_rom[  453]='h000004e5;
    rd_cycle[  454] = 1'b0;  wr_cycle[  454] = 1'b1;  addr_rom[  454]='h00000718;  wr_data_rom[  454]='h00000df5;
    rd_cycle[  455] = 1'b0;  wr_cycle[  455] = 1'b1;  addr_rom[  455]='h0000071c;  wr_data_rom[  455]='h0000073e;
    rd_cycle[  456] = 1'b0;  wr_cycle[  456] = 1'b1;  addr_rom[  456]='h00000720;  wr_data_rom[  456]='h000004ea;
    rd_cycle[  457] = 1'b0;  wr_cycle[  457] = 1'b1;  addr_rom[  457]='h00000724;  wr_data_rom[  457]='h0000027e;
    rd_cycle[  458] = 1'b0;  wr_cycle[  458] = 1'b1;  addr_rom[  458]='h00000728;  wr_data_rom[  458]='h0000084f;
    rd_cycle[  459] = 1'b0;  wr_cycle[  459] = 1'b1;  addr_rom[  459]='h0000072c;  wr_data_rom[  459]='h00000ee2;
    rd_cycle[  460] = 1'b0;  wr_cycle[  460] = 1'b1;  addr_rom[  460]='h00000730;  wr_data_rom[  460]='h00000dc8;
    rd_cycle[  461] = 1'b0;  wr_cycle[  461] = 1'b1;  addr_rom[  461]='h00000734;  wr_data_rom[  461]='h00000059;
    rd_cycle[  462] = 1'b0;  wr_cycle[  462] = 1'b1;  addr_rom[  462]='h00000738;  wr_data_rom[  462]='h00000c08;
    rd_cycle[  463] = 1'b0;  wr_cycle[  463] = 1'b1;  addr_rom[  463]='h0000073c;  wr_data_rom[  463]='h00000f56;
    rd_cycle[  464] = 1'b0;  wr_cycle[  464] = 1'b1;  addr_rom[  464]='h00000740;  wr_data_rom[  464]='h00000d5b;
    rd_cycle[  465] = 1'b0;  wr_cycle[  465] = 1'b1;  addr_rom[  465]='h00000744;  wr_data_rom[  465]='h00000bd2;
    rd_cycle[  466] = 1'b0;  wr_cycle[  466] = 1'b1;  addr_rom[  466]='h00000748;  wr_data_rom[  466]='h00000791;
    rd_cycle[  467] = 1'b0;  wr_cycle[  467] = 1'b1;  addr_rom[  467]='h0000074c;  wr_data_rom[  467]='h00000b36;
    rd_cycle[  468] = 1'b0;  wr_cycle[  468] = 1'b1;  addr_rom[  468]='h00000750;  wr_data_rom[  468]='h00000bb0;
    rd_cycle[  469] = 1'b0;  wr_cycle[  469] = 1'b1;  addr_rom[  469]='h00000754;  wr_data_rom[  469]='h00000330;
    rd_cycle[  470] = 1'b0;  wr_cycle[  470] = 1'b1;  addr_rom[  470]='h00000758;  wr_data_rom[  470]='h0000050f;
    rd_cycle[  471] = 1'b0;  wr_cycle[  471] = 1'b1;  addr_rom[  471]='h0000075c;  wr_data_rom[  471]='h00000420;
    rd_cycle[  472] = 1'b0;  wr_cycle[  472] = 1'b1;  addr_rom[  472]='h00000760;  wr_data_rom[  472]='h000008fc;
    rd_cycle[  473] = 1'b0;  wr_cycle[  473] = 1'b1;  addr_rom[  473]='h00000764;  wr_data_rom[  473]='h00000f92;
    rd_cycle[  474] = 1'b0;  wr_cycle[  474] = 1'b1;  addr_rom[  474]='h00000768;  wr_data_rom[  474]='h00000945;
    rd_cycle[  475] = 1'b0;  wr_cycle[  475] = 1'b1;  addr_rom[  475]='h0000076c;  wr_data_rom[  475]='h000000c1;
    rd_cycle[  476] = 1'b0;  wr_cycle[  476] = 1'b1;  addr_rom[  476]='h00000770;  wr_data_rom[  476]='h00000b04;
    rd_cycle[  477] = 1'b0;  wr_cycle[  477] = 1'b1;  addr_rom[  477]='h00000774;  wr_data_rom[  477]='h00000e3e;
    rd_cycle[  478] = 1'b0;  wr_cycle[  478] = 1'b1;  addr_rom[  478]='h00000778;  wr_data_rom[  478]='h000004fc;
    rd_cycle[  479] = 1'b0;  wr_cycle[  479] = 1'b1;  addr_rom[  479]='h0000077c;  wr_data_rom[  479]='h00000352;
    rd_cycle[  480] = 1'b0;  wr_cycle[  480] = 1'b1;  addr_rom[  480]='h00000780;  wr_data_rom[  480]='h0000058e;
    rd_cycle[  481] = 1'b0;  wr_cycle[  481] = 1'b1;  addr_rom[  481]='h00000784;  wr_data_rom[  481]='h000001d7;
    rd_cycle[  482] = 1'b0;  wr_cycle[  482] = 1'b1;  addr_rom[  482]='h00000788;  wr_data_rom[  482]='h00000b02;
    rd_cycle[  483] = 1'b0;  wr_cycle[  483] = 1'b1;  addr_rom[  483]='h0000078c;  wr_data_rom[  483]='h00000d60;
    rd_cycle[  484] = 1'b0;  wr_cycle[  484] = 1'b1;  addr_rom[  484]='h00000790;  wr_data_rom[  484]='h000004c3;
    rd_cycle[  485] = 1'b0;  wr_cycle[  485] = 1'b1;  addr_rom[  485]='h00000794;  wr_data_rom[  485]='h0000096c;
    rd_cycle[  486] = 1'b0;  wr_cycle[  486] = 1'b1;  addr_rom[  486]='h00000798;  wr_data_rom[  486]='h000006b1;
    rd_cycle[  487] = 1'b0;  wr_cycle[  487] = 1'b1;  addr_rom[  487]='h0000079c;  wr_data_rom[  487]='h00000200;
    rd_cycle[  488] = 1'b0;  wr_cycle[  488] = 1'b1;  addr_rom[  488]='h000007a0;  wr_data_rom[  488]='h0000002e;
    rd_cycle[  489] = 1'b0;  wr_cycle[  489] = 1'b1;  addr_rom[  489]='h000007a4;  wr_data_rom[  489]='h00000738;
    rd_cycle[  490] = 1'b0;  wr_cycle[  490] = 1'b1;  addr_rom[  490]='h000007a8;  wr_data_rom[  490]='h00000ad7;
    rd_cycle[  491] = 1'b0;  wr_cycle[  491] = 1'b1;  addr_rom[  491]='h000007ac;  wr_data_rom[  491]='h000002b5;
    rd_cycle[  492] = 1'b0;  wr_cycle[  492] = 1'b1;  addr_rom[  492]='h000007b0;  wr_data_rom[  492]='h00000a78;
    rd_cycle[  493] = 1'b0;  wr_cycle[  493] = 1'b1;  addr_rom[  493]='h000007b4;  wr_data_rom[  493]='h000004d8;
    rd_cycle[  494] = 1'b0;  wr_cycle[  494] = 1'b1;  addr_rom[  494]='h000007b8;  wr_data_rom[  494]='h00000834;
    rd_cycle[  495] = 1'b0;  wr_cycle[  495] = 1'b1;  addr_rom[  495]='h000007bc;  wr_data_rom[  495]='h0000088f;
    rd_cycle[  496] = 1'b0;  wr_cycle[  496] = 1'b1;  addr_rom[  496]='h000007c0;  wr_data_rom[  496]='h0000014d;
    rd_cycle[  497] = 1'b0;  wr_cycle[  497] = 1'b1;  addr_rom[  497]='h000007c4;  wr_data_rom[  497]='h00000ceb;
    rd_cycle[  498] = 1'b0;  wr_cycle[  498] = 1'b1;  addr_rom[  498]='h000007c8;  wr_data_rom[  498]='h0000082c;
    rd_cycle[  499] = 1'b0;  wr_cycle[  499] = 1'b1;  addr_rom[  499]='h000007cc;  wr_data_rom[  499]='h000008f8;
    rd_cycle[  500] = 1'b0;  wr_cycle[  500] = 1'b1;  addr_rom[  500]='h000007d0;  wr_data_rom[  500]='h00000292;
    rd_cycle[  501] = 1'b0;  wr_cycle[  501] = 1'b1;  addr_rom[  501]='h000007d4;  wr_data_rom[  501]='h0000022c;
    rd_cycle[  502] = 1'b0;  wr_cycle[  502] = 1'b1;  addr_rom[  502]='h000007d8;  wr_data_rom[  502]='h00000334;
    rd_cycle[  503] = 1'b0;  wr_cycle[  503] = 1'b1;  addr_rom[  503]='h000007dc;  wr_data_rom[  503]='h00000209;
    rd_cycle[  504] = 1'b0;  wr_cycle[  504] = 1'b1;  addr_rom[  504]='h000007e0;  wr_data_rom[  504]='h00000c56;
    rd_cycle[  505] = 1'b0;  wr_cycle[  505] = 1'b1;  addr_rom[  505]='h000007e4;  wr_data_rom[  505]='h00000c9d;
    rd_cycle[  506] = 1'b0;  wr_cycle[  506] = 1'b1;  addr_rom[  506]='h000007e8;  wr_data_rom[  506]='h00000757;
    rd_cycle[  507] = 1'b0;  wr_cycle[  507] = 1'b1;  addr_rom[  507]='h000007ec;  wr_data_rom[  507]='h00000077;
    rd_cycle[  508] = 1'b0;  wr_cycle[  508] = 1'b1;  addr_rom[  508]='h000007f0;  wr_data_rom[  508]='h00000977;
    rd_cycle[  509] = 1'b0;  wr_cycle[  509] = 1'b1;  addr_rom[  509]='h000007f4;  wr_data_rom[  509]='h00000445;
    rd_cycle[  510] = 1'b0;  wr_cycle[  510] = 1'b1;  addr_rom[  510]='h000007f8;  wr_data_rom[  510]='h00000c26;
    rd_cycle[  511] = 1'b0;  wr_cycle[  511] = 1'b1;  addr_rom[  511]='h000007fc;  wr_data_rom[  511]='h00000331;
    rd_cycle[  512] = 1'b0;  wr_cycle[  512] = 1'b1;  addr_rom[  512]='h00000800;  wr_data_rom[  512]='h00000dde;
    rd_cycle[  513] = 1'b0;  wr_cycle[  513] = 1'b1;  addr_rom[  513]='h00000804;  wr_data_rom[  513]='h000009fb;
    rd_cycle[  514] = 1'b0;  wr_cycle[  514] = 1'b1;  addr_rom[  514]='h00000808;  wr_data_rom[  514]='h00000595;
    rd_cycle[  515] = 1'b0;  wr_cycle[  515] = 1'b1;  addr_rom[  515]='h0000080c;  wr_data_rom[  515]='h00000772;
    rd_cycle[  516] = 1'b0;  wr_cycle[  516] = 1'b1;  addr_rom[  516]='h00000810;  wr_data_rom[  516]='h00000bd9;
    rd_cycle[  517] = 1'b0;  wr_cycle[  517] = 1'b1;  addr_rom[  517]='h00000814;  wr_data_rom[  517]='h000006a0;
    rd_cycle[  518] = 1'b0;  wr_cycle[  518] = 1'b1;  addr_rom[  518]='h00000818;  wr_data_rom[  518]='h00000162;
    rd_cycle[  519] = 1'b0;  wr_cycle[  519] = 1'b1;  addr_rom[  519]='h0000081c;  wr_data_rom[  519]='h00000e70;
    rd_cycle[  520] = 1'b0;  wr_cycle[  520] = 1'b1;  addr_rom[  520]='h00000820;  wr_data_rom[  520]='h000002b9;
    rd_cycle[  521] = 1'b0;  wr_cycle[  521] = 1'b1;  addr_rom[  521]='h00000824;  wr_data_rom[  521]='h00000a46;
    rd_cycle[  522] = 1'b0;  wr_cycle[  522] = 1'b1;  addr_rom[  522]='h00000828;  wr_data_rom[  522]='h0000035a;
    rd_cycle[  523] = 1'b0;  wr_cycle[  523] = 1'b1;  addr_rom[  523]='h0000082c;  wr_data_rom[  523]='h00000bf2;
    rd_cycle[  524] = 1'b0;  wr_cycle[  524] = 1'b1;  addr_rom[  524]='h00000830;  wr_data_rom[  524]='h0000028c;
    rd_cycle[  525] = 1'b0;  wr_cycle[  525] = 1'b1;  addr_rom[  525]='h00000834;  wr_data_rom[  525]='h00000779;
    rd_cycle[  526] = 1'b0;  wr_cycle[  526] = 1'b1;  addr_rom[  526]='h00000838;  wr_data_rom[  526]='h00000614;
    rd_cycle[  527] = 1'b0;  wr_cycle[  527] = 1'b1;  addr_rom[  527]='h0000083c;  wr_data_rom[  527]='h00000371;
    rd_cycle[  528] = 1'b0;  wr_cycle[  528] = 1'b1;  addr_rom[  528]='h00000840;  wr_data_rom[  528]='h000004ec;
    rd_cycle[  529] = 1'b0;  wr_cycle[  529] = 1'b1;  addr_rom[  529]='h00000844;  wr_data_rom[  529]='h00000ad6;
    rd_cycle[  530] = 1'b0;  wr_cycle[  530] = 1'b1;  addr_rom[  530]='h00000848;  wr_data_rom[  530]='h00000e05;
    rd_cycle[  531] = 1'b0;  wr_cycle[  531] = 1'b1;  addr_rom[  531]='h0000084c;  wr_data_rom[  531]='h00000ba7;
    rd_cycle[  532] = 1'b0;  wr_cycle[  532] = 1'b1;  addr_rom[  532]='h00000850;  wr_data_rom[  532]='h00000a0d;
    rd_cycle[  533] = 1'b0;  wr_cycle[  533] = 1'b1;  addr_rom[  533]='h00000854;  wr_data_rom[  533]='h00000027;
    rd_cycle[  534] = 1'b0;  wr_cycle[  534] = 1'b1;  addr_rom[  534]='h00000858;  wr_data_rom[  534]='h00000031;
    rd_cycle[  535] = 1'b0;  wr_cycle[  535] = 1'b1;  addr_rom[  535]='h0000085c;  wr_data_rom[  535]='h00000077;
    rd_cycle[  536] = 1'b0;  wr_cycle[  536] = 1'b1;  addr_rom[  536]='h00000860;  wr_data_rom[  536]='h000007c6;
    rd_cycle[  537] = 1'b0;  wr_cycle[  537] = 1'b1;  addr_rom[  537]='h00000864;  wr_data_rom[  537]='h000003a6;
    rd_cycle[  538] = 1'b0;  wr_cycle[  538] = 1'b1;  addr_rom[  538]='h00000868;  wr_data_rom[  538]='h000002a1;
    rd_cycle[  539] = 1'b0;  wr_cycle[  539] = 1'b1;  addr_rom[  539]='h0000086c;  wr_data_rom[  539]='h00000180;
    rd_cycle[  540] = 1'b0;  wr_cycle[  540] = 1'b1;  addr_rom[  540]='h00000870;  wr_data_rom[  540]='h000007d4;
    rd_cycle[  541] = 1'b0;  wr_cycle[  541] = 1'b1;  addr_rom[  541]='h00000874;  wr_data_rom[  541]='h000000fd;
    rd_cycle[  542] = 1'b0;  wr_cycle[  542] = 1'b1;  addr_rom[  542]='h00000878;  wr_data_rom[  542]='h00000357;
    rd_cycle[  543] = 1'b0;  wr_cycle[  543] = 1'b1;  addr_rom[  543]='h0000087c;  wr_data_rom[  543]='h00000614;
    rd_cycle[  544] = 1'b0;  wr_cycle[  544] = 1'b1;  addr_rom[  544]='h00000880;  wr_data_rom[  544]='h00000e96;
    rd_cycle[  545] = 1'b0;  wr_cycle[  545] = 1'b1;  addr_rom[  545]='h00000884;  wr_data_rom[  545]='h00000c3f;
    rd_cycle[  546] = 1'b0;  wr_cycle[  546] = 1'b1;  addr_rom[  546]='h00000888;  wr_data_rom[  546]='h000008b0;
    rd_cycle[  547] = 1'b0;  wr_cycle[  547] = 1'b1;  addr_rom[  547]='h0000088c;  wr_data_rom[  547]='h0000096e;
    rd_cycle[  548] = 1'b0;  wr_cycle[  548] = 1'b1;  addr_rom[  548]='h00000890;  wr_data_rom[  548]='h0000063f;
    rd_cycle[  549] = 1'b0;  wr_cycle[  549] = 1'b1;  addr_rom[  549]='h00000894;  wr_data_rom[  549]='h00000bad;
    rd_cycle[  550] = 1'b0;  wr_cycle[  550] = 1'b1;  addr_rom[  550]='h00000898;  wr_data_rom[  550]='h00000abd;
    rd_cycle[  551] = 1'b0;  wr_cycle[  551] = 1'b1;  addr_rom[  551]='h0000089c;  wr_data_rom[  551]='h00000256;
    rd_cycle[  552] = 1'b0;  wr_cycle[  552] = 1'b1;  addr_rom[  552]='h000008a0;  wr_data_rom[  552]='h00000c28;
    rd_cycle[  553] = 1'b0;  wr_cycle[  553] = 1'b1;  addr_rom[  553]='h000008a4;  wr_data_rom[  553]='h000004f4;
    rd_cycle[  554] = 1'b0;  wr_cycle[  554] = 1'b1;  addr_rom[  554]='h000008a8;  wr_data_rom[  554]='h00000195;
    rd_cycle[  555] = 1'b0;  wr_cycle[  555] = 1'b1;  addr_rom[  555]='h000008ac;  wr_data_rom[  555]='h000004c9;
    rd_cycle[  556] = 1'b0;  wr_cycle[  556] = 1'b1;  addr_rom[  556]='h000008b0;  wr_data_rom[  556]='h00000a3c;
    rd_cycle[  557] = 1'b0;  wr_cycle[  557] = 1'b1;  addr_rom[  557]='h000008b4;  wr_data_rom[  557]='h00000892;
    rd_cycle[  558] = 1'b0;  wr_cycle[  558] = 1'b1;  addr_rom[  558]='h000008b8;  wr_data_rom[  558]='h00000af1;
    rd_cycle[  559] = 1'b0;  wr_cycle[  559] = 1'b1;  addr_rom[  559]='h000008bc;  wr_data_rom[  559]='h00000186;
    rd_cycle[  560] = 1'b0;  wr_cycle[  560] = 1'b1;  addr_rom[  560]='h000008c0;  wr_data_rom[  560]='h00000b0a;
    rd_cycle[  561] = 1'b0;  wr_cycle[  561] = 1'b1;  addr_rom[  561]='h000008c4;  wr_data_rom[  561]='h000008f3;
    rd_cycle[  562] = 1'b0;  wr_cycle[  562] = 1'b1;  addr_rom[  562]='h000008c8;  wr_data_rom[  562]='h00000875;
    rd_cycle[  563] = 1'b0;  wr_cycle[  563] = 1'b1;  addr_rom[  563]='h000008cc;  wr_data_rom[  563]='h000008a7;
    rd_cycle[  564] = 1'b0;  wr_cycle[  564] = 1'b1;  addr_rom[  564]='h000008d0;  wr_data_rom[  564]='h00000280;
    rd_cycle[  565] = 1'b0;  wr_cycle[  565] = 1'b1;  addr_rom[  565]='h000008d4;  wr_data_rom[  565]='h000002f8;
    rd_cycle[  566] = 1'b0;  wr_cycle[  566] = 1'b1;  addr_rom[  566]='h000008d8;  wr_data_rom[  566]='h00000c42;
    rd_cycle[  567] = 1'b0;  wr_cycle[  567] = 1'b1;  addr_rom[  567]='h000008dc;  wr_data_rom[  567]='h0000048a;
    rd_cycle[  568] = 1'b0;  wr_cycle[  568] = 1'b1;  addr_rom[  568]='h000008e0;  wr_data_rom[  568]='h00000438;
    rd_cycle[  569] = 1'b0;  wr_cycle[  569] = 1'b1;  addr_rom[  569]='h000008e4;  wr_data_rom[  569]='h0000048d;
    rd_cycle[  570] = 1'b0;  wr_cycle[  570] = 1'b1;  addr_rom[  570]='h000008e8;  wr_data_rom[  570]='h00000e5f;
    rd_cycle[  571] = 1'b0;  wr_cycle[  571] = 1'b1;  addr_rom[  571]='h000008ec;  wr_data_rom[  571]='h00000609;
    rd_cycle[  572] = 1'b0;  wr_cycle[  572] = 1'b1;  addr_rom[  572]='h000008f0;  wr_data_rom[  572]='h00000c7f;
    rd_cycle[  573] = 1'b0;  wr_cycle[  573] = 1'b1;  addr_rom[  573]='h000008f4;  wr_data_rom[  573]='h000006be;
    rd_cycle[  574] = 1'b0;  wr_cycle[  574] = 1'b1;  addr_rom[  574]='h000008f8;  wr_data_rom[  574]='h000008c5;
    rd_cycle[  575] = 1'b0;  wr_cycle[  575] = 1'b1;  addr_rom[  575]='h000008fc;  wr_data_rom[  575]='h000006f1;
    rd_cycle[  576] = 1'b0;  wr_cycle[  576] = 1'b1;  addr_rom[  576]='h00000900;  wr_data_rom[  576]='h00000636;
    rd_cycle[  577] = 1'b0;  wr_cycle[  577] = 1'b1;  addr_rom[  577]='h00000904;  wr_data_rom[  577]='h000000ff;
    rd_cycle[  578] = 1'b0;  wr_cycle[  578] = 1'b1;  addr_rom[  578]='h00000908;  wr_data_rom[  578]='h0000059d;
    rd_cycle[  579] = 1'b0;  wr_cycle[  579] = 1'b1;  addr_rom[  579]='h0000090c;  wr_data_rom[  579]='h000000ae;
    rd_cycle[  580] = 1'b0;  wr_cycle[  580] = 1'b1;  addr_rom[  580]='h00000910;  wr_data_rom[  580]='h00000244;
    rd_cycle[  581] = 1'b0;  wr_cycle[  581] = 1'b1;  addr_rom[  581]='h00000914;  wr_data_rom[  581]='h00000439;
    rd_cycle[  582] = 1'b0;  wr_cycle[  582] = 1'b1;  addr_rom[  582]='h00000918;  wr_data_rom[  582]='h00000e60;
    rd_cycle[  583] = 1'b0;  wr_cycle[  583] = 1'b1;  addr_rom[  583]='h0000091c;  wr_data_rom[  583]='h000004cb;
    rd_cycle[  584] = 1'b0;  wr_cycle[  584] = 1'b1;  addr_rom[  584]='h00000920;  wr_data_rom[  584]='h00000209;
    rd_cycle[  585] = 1'b0;  wr_cycle[  585] = 1'b1;  addr_rom[  585]='h00000924;  wr_data_rom[  585]='h00000a41;
    rd_cycle[  586] = 1'b0;  wr_cycle[  586] = 1'b1;  addr_rom[  586]='h00000928;  wr_data_rom[  586]='h00000685;
    rd_cycle[  587] = 1'b0;  wr_cycle[  587] = 1'b1;  addr_rom[  587]='h0000092c;  wr_data_rom[  587]='h00000f91;
    rd_cycle[  588] = 1'b0;  wr_cycle[  588] = 1'b1;  addr_rom[  588]='h00000930;  wr_data_rom[  588]='h00000ba8;
    rd_cycle[  589] = 1'b0;  wr_cycle[  589] = 1'b1;  addr_rom[  589]='h00000934;  wr_data_rom[  589]='h00000309;
    rd_cycle[  590] = 1'b0;  wr_cycle[  590] = 1'b1;  addr_rom[  590]='h00000938;  wr_data_rom[  590]='h000005a8;
    rd_cycle[  591] = 1'b0;  wr_cycle[  591] = 1'b1;  addr_rom[  591]='h0000093c;  wr_data_rom[  591]='h00000a42;
    rd_cycle[  592] = 1'b0;  wr_cycle[  592] = 1'b1;  addr_rom[  592]='h00000940;  wr_data_rom[  592]='h00000a9b;
    rd_cycle[  593] = 1'b0;  wr_cycle[  593] = 1'b1;  addr_rom[  593]='h00000944;  wr_data_rom[  593]='h0000010d;
    rd_cycle[  594] = 1'b0;  wr_cycle[  594] = 1'b1;  addr_rom[  594]='h00000948;  wr_data_rom[  594]='h00000bf9;
    rd_cycle[  595] = 1'b0;  wr_cycle[  595] = 1'b1;  addr_rom[  595]='h0000094c;  wr_data_rom[  595]='h00000176;
    rd_cycle[  596] = 1'b0;  wr_cycle[  596] = 1'b1;  addr_rom[  596]='h00000950;  wr_data_rom[  596]='h00000b6e;
    rd_cycle[  597] = 1'b0;  wr_cycle[  597] = 1'b1;  addr_rom[  597]='h00000954;  wr_data_rom[  597]='h000007da;
    rd_cycle[  598] = 1'b0;  wr_cycle[  598] = 1'b1;  addr_rom[  598]='h00000958;  wr_data_rom[  598]='h00000113;
    rd_cycle[  599] = 1'b0;  wr_cycle[  599] = 1'b1;  addr_rom[  599]='h0000095c;  wr_data_rom[  599]='h000001b5;
    rd_cycle[  600] = 1'b0;  wr_cycle[  600] = 1'b1;  addr_rom[  600]='h00000960;  wr_data_rom[  600]='h00000d24;
    rd_cycle[  601] = 1'b0;  wr_cycle[  601] = 1'b1;  addr_rom[  601]='h00000964;  wr_data_rom[  601]='h000001a4;
    rd_cycle[  602] = 1'b0;  wr_cycle[  602] = 1'b1;  addr_rom[  602]='h00000968;  wr_data_rom[  602]='h000002c1;
    rd_cycle[  603] = 1'b0;  wr_cycle[  603] = 1'b1;  addr_rom[  603]='h0000096c;  wr_data_rom[  603]='h0000072d;
    rd_cycle[  604] = 1'b0;  wr_cycle[  604] = 1'b1;  addr_rom[  604]='h00000970;  wr_data_rom[  604]='h000007d4;
    rd_cycle[  605] = 1'b0;  wr_cycle[  605] = 1'b1;  addr_rom[  605]='h00000974;  wr_data_rom[  605]='h00000567;
    rd_cycle[  606] = 1'b0;  wr_cycle[  606] = 1'b1;  addr_rom[  606]='h00000978;  wr_data_rom[  606]='h0000060e;
    rd_cycle[  607] = 1'b0;  wr_cycle[  607] = 1'b1;  addr_rom[  607]='h0000097c;  wr_data_rom[  607]='h00000c03;
    rd_cycle[  608] = 1'b0;  wr_cycle[  608] = 1'b1;  addr_rom[  608]='h00000980;  wr_data_rom[  608]='h00000ab8;
    rd_cycle[  609] = 1'b0;  wr_cycle[  609] = 1'b1;  addr_rom[  609]='h00000984;  wr_data_rom[  609]='h000001f6;
    rd_cycle[  610] = 1'b0;  wr_cycle[  610] = 1'b1;  addr_rom[  610]='h00000988;  wr_data_rom[  610]='h0000095e;
    rd_cycle[  611] = 1'b0;  wr_cycle[  611] = 1'b1;  addr_rom[  611]='h0000098c;  wr_data_rom[  611]='h0000077b;
    rd_cycle[  612] = 1'b0;  wr_cycle[  612] = 1'b1;  addr_rom[  612]='h00000990;  wr_data_rom[  612]='h00000017;
    rd_cycle[  613] = 1'b0;  wr_cycle[  613] = 1'b1;  addr_rom[  613]='h00000994;  wr_data_rom[  613]='h000003ba;
    rd_cycle[  614] = 1'b0;  wr_cycle[  614] = 1'b1;  addr_rom[  614]='h00000998;  wr_data_rom[  614]='h0000034f;
    rd_cycle[  615] = 1'b0;  wr_cycle[  615] = 1'b1;  addr_rom[  615]='h0000099c;  wr_data_rom[  615]='h00000972;
    rd_cycle[  616] = 1'b0;  wr_cycle[  616] = 1'b1;  addr_rom[  616]='h000009a0;  wr_data_rom[  616]='h00000dc0;
    rd_cycle[  617] = 1'b0;  wr_cycle[  617] = 1'b1;  addr_rom[  617]='h000009a4;  wr_data_rom[  617]='h00000709;
    rd_cycle[  618] = 1'b0;  wr_cycle[  618] = 1'b1;  addr_rom[  618]='h000009a8;  wr_data_rom[  618]='h00000c71;
    rd_cycle[  619] = 1'b0;  wr_cycle[  619] = 1'b1;  addr_rom[  619]='h000009ac;  wr_data_rom[  619]='h00000f9b;
    rd_cycle[  620] = 1'b0;  wr_cycle[  620] = 1'b1;  addr_rom[  620]='h000009b0;  wr_data_rom[  620]='h000009b5;
    rd_cycle[  621] = 1'b0;  wr_cycle[  621] = 1'b1;  addr_rom[  621]='h000009b4;  wr_data_rom[  621]='h00000990;
    rd_cycle[  622] = 1'b0;  wr_cycle[  622] = 1'b1;  addr_rom[  622]='h000009b8;  wr_data_rom[  622]='h000008f1;
    rd_cycle[  623] = 1'b0;  wr_cycle[  623] = 1'b1;  addr_rom[  623]='h000009bc;  wr_data_rom[  623]='h00000037;
    rd_cycle[  624] = 1'b0;  wr_cycle[  624] = 1'b1;  addr_rom[  624]='h000009c0;  wr_data_rom[  624]='h000003c8;
    rd_cycle[  625] = 1'b0;  wr_cycle[  625] = 1'b1;  addr_rom[  625]='h000009c4;  wr_data_rom[  625]='h00000524;
    rd_cycle[  626] = 1'b0;  wr_cycle[  626] = 1'b1;  addr_rom[  626]='h000009c8;  wr_data_rom[  626]='h00000543;
    rd_cycle[  627] = 1'b0;  wr_cycle[  627] = 1'b1;  addr_rom[  627]='h000009cc;  wr_data_rom[  627]='h0000000b;
    rd_cycle[  628] = 1'b0;  wr_cycle[  628] = 1'b1;  addr_rom[  628]='h000009d0;  wr_data_rom[  628]='h000008fc;
    rd_cycle[  629] = 1'b0;  wr_cycle[  629] = 1'b1;  addr_rom[  629]='h000009d4;  wr_data_rom[  629]='h00000e0a;
    rd_cycle[  630] = 1'b0;  wr_cycle[  630] = 1'b1;  addr_rom[  630]='h000009d8;  wr_data_rom[  630]='h00000d75;
    rd_cycle[  631] = 1'b0;  wr_cycle[  631] = 1'b1;  addr_rom[  631]='h000009dc;  wr_data_rom[  631]='h000008f2;
    rd_cycle[  632] = 1'b0;  wr_cycle[  632] = 1'b1;  addr_rom[  632]='h000009e0;  wr_data_rom[  632]='h000007fc;
    rd_cycle[  633] = 1'b0;  wr_cycle[  633] = 1'b1;  addr_rom[  633]='h000009e4;  wr_data_rom[  633]='h00000590;
    rd_cycle[  634] = 1'b0;  wr_cycle[  634] = 1'b1;  addr_rom[  634]='h000009e8;  wr_data_rom[  634]='h00000473;
    rd_cycle[  635] = 1'b0;  wr_cycle[  635] = 1'b1;  addr_rom[  635]='h000009ec;  wr_data_rom[  635]='h000004ea;
    rd_cycle[  636] = 1'b0;  wr_cycle[  636] = 1'b1;  addr_rom[  636]='h000009f0;  wr_data_rom[  636]='h00000a8e;
    rd_cycle[  637] = 1'b0;  wr_cycle[  637] = 1'b1;  addr_rom[  637]='h000009f4;  wr_data_rom[  637]='h000009de;
    rd_cycle[  638] = 1'b0;  wr_cycle[  638] = 1'b1;  addr_rom[  638]='h000009f8;  wr_data_rom[  638]='h00000774;
    rd_cycle[  639] = 1'b0;  wr_cycle[  639] = 1'b1;  addr_rom[  639]='h000009fc;  wr_data_rom[  639]='h000006fd;
    rd_cycle[  640] = 1'b0;  wr_cycle[  640] = 1'b1;  addr_rom[  640]='h00000a00;  wr_data_rom[  640]='h00000a09;
    rd_cycle[  641] = 1'b0;  wr_cycle[  641] = 1'b1;  addr_rom[  641]='h00000a04;  wr_data_rom[  641]='h00000d17;
    rd_cycle[  642] = 1'b0;  wr_cycle[  642] = 1'b1;  addr_rom[  642]='h00000a08;  wr_data_rom[  642]='h00000a98;
    rd_cycle[  643] = 1'b0;  wr_cycle[  643] = 1'b1;  addr_rom[  643]='h00000a0c;  wr_data_rom[  643]='h000004e3;
    rd_cycle[  644] = 1'b0;  wr_cycle[  644] = 1'b1;  addr_rom[  644]='h00000a10;  wr_data_rom[  644]='h0000078f;
    rd_cycle[  645] = 1'b0;  wr_cycle[  645] = 1'b1;  addr_rom[  645]='h00000a14;  wr_data_rom[  645]='h0000088d;
    rd_cycle[  646] = 1'b0;  wr_cycle[  646] = 1'b1;  addr_rom[  646]='h00000a18;  wr_data_rom[  646]='h00000dcb;
    rd_cycle[  647] = 1'b0;  wr_cycle[  647] = 1'b1;  addr_rom[  647]='h00000a1c;  wr_data_rom[  647]='h000006cb;
    rd_cycle[  648] = 1'b0;  wr_cycle[  648] = 1'b1;  addr_rom[  648]='h00000a20;  wr_data_rom[  648]='h00000395;
    rd_cycle[  649] = 1'b0;  wr_cycle[  649] = 1'b1;  addr_rom[  649]='h00000a24;  wr_data_rom[  649]='h00000d5c;
    rd_cycle[  650] = 1'b0;  wr_cycle[  650] = 1'b1;  addr_rom[  650]='h00000a28;  wr_data_rom[  650]='h000007ec;
    rd_cycle[  651] = 1'b0;  wr_cycle[  651] = 1'b1;  addr_rom[  651]='h00000a2c;  wr_data_rom[  651]='h00000981;
    rd_cycle[  652] = 1'b0;  wr_cycle[  652] = 1'b1;  addr_rom[  652]='h00000a30;  wr_data_rom[  652]='h00000453;
    rd_cycle[  653] = 1'b0;  wr_cycle[  653] = 1'b1;  addr_rom[  653]='h00000a34;  wr_data_rom[  653]='h000009ad;
    rd_cycle[  654] = 1'b0;  wr_cycle[  654] = 1'b1;  addr_rom[  654]='h00000a38;  wr_data_rom[  654]='h000006ea;
    rd_cycle[  655] = 1'b0;  wr_cycle[  655] = 1'b1;  addr_rom[  655]='h00000a3c;  wr_data_rom[  655]='h0000086c;
    rd_cycle[  656] = 1'b0;  wr_cycle[  656] = 1'b1;  addr_rom[  656]='h00000a40;  wr_data_rom[  656]='h000009a6;
    rd_cycle[  657] = 1'b0;  wr_cycle[  657] = 1'b1;  addr_rom[  657]='h00000a44;  wr_data_rom[  657]='h00000f0d;
    rd_cycle[  658] = 1'b0;  wr_cycle[  658] = 1'b1;  addr_rom[  658]='h00000a48;  wr_data_rom[  658]='h00000686;
    rd_cycle[  659] = 1'b0;  wr_cycle[  659] = 1'b1;  addr_rom[  659]='h00000a4c;  wr_data_rom[  659]='h00000f8e;
    rd_cycle[  660] = 1'b0;  wr_cycle[  660] = 1'b1;  addr_rom[  660]='h00000a50;  wr_data_rom[  660]='h00000041;
    rd_cycle[  661] = 1'b0;  wr_cycle[  661] = 1'b1;  addr_rom[  661]='h00000a54;  wr_data_rom[  661]='h00000d57;
    rd_cycle[  662] = 1'b0;  wr_cycle[  662] = 1'b1;  addr_rom[  662]='h00000a58;  wr_data_rom[  662]='h00000d7a;
    rd_cycle[  663] = 1'b0;  wr_cycle[  663] = 1'b1;  addr_rom[  663]='h00000a5c;  wr_data_rom[  663]='h00000d8b;
    rd_cycle[  664] = 1'b0;  wr_cycle[  664] = 1'b1;  addr_rom[  664]='h00000a60;  wr_data_rom[  664]='h000004cd;
    rd_cycle[  665] = 1'b0;  wr_cycle[  665] = 1'b1;  addr_rom[  665]='h00000a64;  wr_data_rom[  665]='h00000c9b;
    rd_cycle[  666] = 1'b0;  wr_cycle[  666] = 1'b1;  addr_rom[  666]='h00000a68;  wr_data_rom[  666]='h00000810;
    rd_cycle[  667] = 1'b0;  wr_cycle[  667] = 1'b1;  addr_rom[  667]='h00000a6c;  wr_data_rom[  667]='h00000d5b;
    rd_cycle[  668] = 1'b0;  wr_cycle[  668] = 1'b1;  addr_rom[  668]='h00000a70;  wr_data_rom[  668]='h00000939;
    rd_cycle[  669] = 1'b0;  wr_cycle[  669] = 1'b1;  addr_rom[  669]='h00000a74;  wr_data_rom[  669]='h00000e20;
    rd_cycle[  670] = 1'b0;  wr_cycle[  670] = 1'b1;  addr_rom[  670]='h00000a78;  wr_data_rom[  670]='h0000089b;
    rd_cycle[  671] = 1'b0;  wr_cycle[  671] = 1'b1;  addr_rom[  671]='h00000a7c;  wr_data_rom[  671]='h00000b06;
    rd_cycle[  672] = 1'b0;  wr_cycle[  672] = 1'b1;  addr_rom[  672]='h00000a80;  wr_data_rom[  672]='h00000736;
    rd_cycle[  673] = 1'b0;  wr_cycle[  673] = 1'b1;  addr_rom[  673]='h00000a84;  wr_data_rom[  673]='h00000b87;
    rd_cycle[  674] = 1'b0;  wr_cycle[  674] = 1'b1;  addr_rom[  674]='h00000a88;  wr_data_rom[  674]='h00000401;
    rd_cycle[  675] = 1'b0;  wr_cycle[  675] = 1'b1;  addr_rom[  675]='h00000a8c;  wr_data_rom[  675]='h000009ad;
    rd_cycle[  676] = 1'b0;  wr_cycle[  676] = 1'b1;  addr_rom[  676]='h00000a90;  wr_data_rom[  676]='h00000d19;
    rd_cycle[  677] = 1'b0;  wr_cycle[  677] = 1'b1;  addr_rom[  677]='h00000a94;  wr_data_rom[  677]='h00000265;
    rd_cycle[  678] = 1'b0;  wr_cycle[  678] = 1'b1;  addr_rom[  678]='h00000a98;  wr_data_rom[  678]='h00000927;
    rd_cycle[  679] = 1'b0;  wr_cycle[  679] = 1'b1;  addr_rom[  679]='h00000a9c;  wr_data_rom[  679]='h000006f4;
    rd_cycle[  680] = 1'b0;  wr_cycle[  680] = 1'b1;  addr_rom[  680]='h00000aa0;  wr_data_rom[  680]='h00000c9d;
    rd_cycle[  681] = 1'b0;  wr_cycle[  681] = 1'b1;  addr_rom[  681]='h00000aa4;  wr_data_rom[  681]='h00000093;
    rd_cycle[  682] = 1'b0;  wr_cycle[  682] = 1'b1;  addr_rom[  682]='h00000aa8;  wr_data_rom[  682]='h00000879;
    rd_cycle[  683] = 1'b0;  wr_cycle[  683] = 1'b1;  addr_rom[  683]='h00000aac;  wr_data_rom[  683]='h0000084c;
    rd_cycle[  684] = 1'b0;  wr_cycle[  684] = 1'b1;  addr_rom[  684]='h00000ab0;  wr_data_rom[  684]='h00000570;
    rd_cycle[  685] = 1'b0;  wr_cycle[  685] = 1'b1;  addr_rom[  685]='h00000ab4;  wr_data_rom[  685]='h00000438;
    rd_cycle[  686] = 1'b0;  wr_cycle[  686] = 1'b1;  addr_rom[  686]='h00000ab8;  wr_data_rom[  686]='h000003cd;
    rd_cycle[  687] = 1'b0;  wr_cycle[  687] = 1'b1;  addr_rom[  687]='h00000abc;  wr_data_rom[  687]='h000006bc;
    rd_cycle[  688] = 1'b0;  wr_cycle[  688] = 1'b1;  addr_rom[  688]='h00000ac0;  wr_data_rom[  688]='h00000ae3;
    rd_cycle[  689] = 1'b0;  wr_cycle[  689] = 1'b1;  addr_rom[  689]='h00000ac4;  wr_data_rom[  689]='h0000025a;
    rd_cycle[  690] = 1'b0;  wr_cycle[  690] = 1'b1;  addr_rom[  690]='h00000ac8;  wr_data_rom[  690]='h00000160;
    rd_cycle[  691] = 1'b0;  wr_cycle[  691] = 1'b1;  addr_rom[  691]='h00000acc;  wr_data_rom[  691]='h00000b6e;
    rd_cycle[  692] = 1'b0;  wr_cycle[  692] = 1'b1;  addr_rom[  692]='h00000ad0;  wr_data_rom[  692]='h00000c51;
    rd_cycle[  693] = 1'b0;  wr_cycle[  693] = 1'b1;  addr_rom[  693]='h00000ad4;  wr_data_rom[  693]='h00000c44;
    rd_cycle[  694] = 1'b0;  wr_cycle[  694] = 1'b1;  addr_rom[  694]='h00000ad8;  wr_data_rom[  694]='h00000a4d;
    rd_cycle[  695] = 1'b0;  wr_cycle[  695] = 1'b1;  addr_rom[  695]='h00000adc;  wr_data_rom[  695]='h0000082f;
    rd_cycle[  696] = 1'b0;  wr_cycle[  696] = 1'b1;  addr_rom[  696]='h00000ae0;  wr_data_rom[  696]='h00000c2d;
    rd_cycle[  697] = 1'b0;  wr_cycle[  697] = 1'b1;  addr_rom[  697]='h00000ae4;  wr_data_rom[  697]='h00000bae;
    rd_cycle[  698] = 1'b0;  wr_cycle[  698] = 1'b1;  addr_rom[  698]='h00000ae8;  wr_data_rom[  698]='h00000cba;
    rd_cycle[  699] = 1'b0;  wr_cycle[  699] = 1'b1;  addr_rom[  699]='h00000aec;  wr_data_rom[  699]='h000001b8;
    rd_cycle[  700] = 1'b0;  wr_cycle[  700] = 1'b1;  addr_rom[  700]='h00000af0;  wr_data_rom[  700]='h00000065;
    rd_cycle[  701] = 1'b0;  wr_cycle[  701] = 1'b1;  addr_rom[  701]='h00000af4;  wr_data_rom[  701]='h00000a2d;
    rd_cycle[  702] = 1'b0;  wr_cycle[  702] = 1'b1;  addr_rom[  702]='h00000af8;  wr_data_rom[  702]='h00000e9b;
    rd_cycle[  703] = 1'b0;  wr_cycle[  703] = 1'b1;  addr_rom[  703]='h00000afc;  wr_data_rom[  703]='h000001cd;
    rd_cycle[  704] = 1'b0;  wr_cycle[  704] = 1'b1;  addr_rom[  704]='h00000b00;  wr_data_rom[  704]='h00000e4f;
    rd_cycle[  705] = 1'b0;  wr_cycle[  705] = 1'b1;  addr_rom[  705]='h00000b04;  wr_data_rom[  705]='h000000fb;
    rd_cycle[  706] = 1'b0;  wr_cycle[  706] = 1'b1;  addr_rom[  706]='h00000b08;  wr_data_rom[  706]='h00000ac7;
    rd_cycle[  707] = 1'b0;  wr_cycle[  707] = 1'b1;  addr_rom[  707]='h00000b0c;  wr_data_rom[  707]='h00000865;
    rd_cycle[  708] = 1'b0;  wr_cycle[  708] = 1'b1;  addr_rom[  708]='h00000b10;  wr_data_rom[  708]='h00000839;
    rd_cycle[  709] = 1'b0;  wr_cycle[  709] = 1'b1;  addr_rom[  709]='h00000b14;  wr_data_rom[  709]='h0000094c;
    rd_cycle[  710] = 1'b0;  wr_cycle[  710] = 1'b1;  addr_rom[  710]='h00000b18;  wr_data_rom[  710]='h000002ce;
    rd_cycle[  711] = 1'b0;  wr_cycle[  711] = 1'b1;  addr_rom[  711]='h00000b1c;  wr_data_rom[  711]='h00000f7a;
    rd_cycle[  712] = 1'b0;  wr_cycle[  712] = 1'b1;  addr_rom[  712]='h00000b20;  wr_data_rom[  712]='h0000017a;
    rd_cycle[  713] = 1'b0;  wr_cycle[  713] = 1'b1;  addr_rom[  713]='h00000b24;  wr_data_rom[  713]='h00000427;
    rd_cycle[  714] = 1'b0;  wr_cycle[  714] = 1'b1;  addr_rom[  714]='h00000b28;  wr_data_rom[  714]='h00000468;
    rd_cycle[  715] = 1'b0;  wr_cycle[  715] = 1'b1;  addr_rom[  715]='h00000b2c;  wr_data_rom[  715]='h00000bc7;
    rd_cycle[  716] = 1'b0;  wr_cycle[  716] = 1'b1;  addr_rom[  716]='h00000b30;  wr_data_rom[  716]='h0000004c;
    rd_cycle[  717] = 1'b0;  wr_cycle[  717] = 1'b1;  addr_rom[  717]='h00000b34;  wr_data_rom[  717]='h00000f9f;
    rd_cycle[  718] = 1'b0;  wr_cycle[  718] = 1'b1;  addr_rom[  718]='h00000b38;  wr_data_rom[  718]='h000006e2;
    rd_cycle[  719] = 1'b0;  wr_cycle[  719] = 1'b1;  addr_rom[  719]='h00000b3c;  wr_data_rom[  719]='h0000000a;
    rd_cycle[  720] = 1'b0;  wr_cycle[  720] = 1'b1;  addr_rom[  720]='h00000b40;  wr_data_rom[  720]='h00000a44;
    rd_cycle[  721] = 1'b0;  wr_cycle[  721] = 1'b1;  addr_rom[  721]='h00000b44;  wr_data_rom[  721]='h0000091c;
    rd_cycle[  722] = 1'b0;  wr_cycle[  722] = 1'b1;  addr_rom[  722]='h00000b48;  wr_data_rom[  722]='h000008ad;
    rd_cycle[  723] = 1'b0;  wr_cycle[  723] = 1'b1;  addr_rom[  723]='h00000b4c;  wr_data_rom[  723]='h00000f63;
    rd_cycle[  724] = 1'b0;  wr_cycle[  724] = 1'b1;  addr_rom[  724]='h00000b50;  wr_data_rom[  724]='h00000d49;
    rd_cycle[  725] = 1'b0;  wr_cycle[  725] = 1'b1;  addr_rom[  725]='h00000b54;  wr_data_rom[  725]='h00000dc6;
    rd_cycle[  726] = 1'b0;  wr_cycle[  726] = 1'b1;  addr_rom[  726]='h00000b58;  wr_data_rom[  726]='h000008c0;
    rd_cycle[  727] = 1'b0;  wr_cycle[  727] = 1'b1;  addr_rom[  727]='h00000b5c;  wr_data_rom[  727]='h00000ae7;
    rd_cycle[  728] = 1'b0;  wr_cycle[  728] = 1'b1;  addr_rom[  728]='h00000b60;  wr_data_rom[  728]='h00000431;
    rd_cycle[  729] = 1'b0;  wr_cycle[  729] = 1'b1;  addr_rom[  729]='h00000b64;  wr_data_rom[  729]='h00000683;
    rd_cycle[  730] = 1'b0;  wr_cycle[  730] = 1'b1;  addr_rom[  730]='h00000b68;  wr_data_rom[  730]='h000008d1;
    rd_cycle[  731] = 1'b0;  wr_cycle[  731] = 1'b1;  addr_rom[  731]='h00000b6c;  wr_data_rom[  731]='h00000190;
    rd_cycle[  732] = 1'b0;  wr_cycle[  732] = 1'b1;  addr_rom[  732]='h00000b70;  wr_data_rom[  732]='h00000478;
    rd_cycle[  733] = 1'b0;  wr_cycle[  733] = 1'b1;  addr_rom[  733]='h00000b74;  wr_data_rom[  733]='h000009ac;
    rd_cycle[  734] = 1'b0;  wr_cycle[  734] = 1'b1;  addr_rom[  734]='h00000b78;  wr_data_rom[  734]='h000004a2;
    rd_cycle[  735] = 1'b0;  wr_cycle[  735] = 1'b1;  addr_rom[  735]='h00000b7c;  wr_data_rom[  735]='h00000a1d;
    rd_cycle[  736] = 1'b0;  wr_cycle[  736] = 1'b1;  addr_rom[  736]='h00000b80;  wr_data_rom[  736]='h00000f9c;
    rd_cycle[  737] = 1'b0;  wr_cycle[  737] = 1'b1;  addr_rom[  737]='h00000b84;  wr_data_rom[  737]='h00000c61;
    rd_cycle[  738] = 1'b0;  wr_cycle[  738] = 1'b1;  addr_rom[  738]='h00000b88;  wr_data_rom[  738]='h00000a0d;
    rd_cycle[  739] = 1'b0;  wr_cycle[  739] = 1'b1;  addr_rom[  739]='h00000b8c;  wr_data_rom[  739]='h00000e95;
    rd_cycle[  740] = 1'b0;  wr_cycle[  740] = 1'b1;  addr_rom[  740]='h00000b90;  wr_data_rom[  740]='h00000f3c;
    rd_cycle[  741] = 1'b0;  wr_cycle[  741] = 1'b1;  addr_rom[  741]='h00000b94;  wr_data_rom[  741]='h00000549;
    rd_cycle[  742] = 1'b0;  wr_cycle[  742] = 1'b1;  addr_rom[  742]='h00000b98;  wr_data_rom[  742]='h00000be0;
    rd_cycle[  743] = 1'b0;  wr_cycle[  743] = 1'b1;  addr_rom[  743]='h00000b9c;  wr_data_rom[  743]='h00000851;
    rd_cycle[  744] = 1'b0;  wr_cycle[  744] = 1'b1;  addr_rom[  744]='h00000ba0;  wr_data_rom[  744]='h00000f8b;
    rd_cycle[  745] = 1'b0;  wr_cycle[  745] = 1'b1;  addr_rom[  745]='h00000ba4;  wr_data_rom[  745]='h00000bad;
    rd_cycle[  746] = 1'b0;  wr_cycle[  746] = 1'b1;  addr_rom[  746]='h00000ba8;  wr_data_rom[  746]='h00000867;
    rd_cycle[  747] = 1'b0;  wr_cycle[  747] = 1'b1;  addr_rom[  747]='h00000bac;  wr_data_rom[  747]='h00000ba2;
    rd_cycle[  748] = 1'b0;  wr_cycle[  748] = 1'b1;  addr_rom[  748]='h00000bb0;  wr_data_rom[  748]='h00000d1c;
    rd_cycle[  749] = 1'b0;  wr_cycle[  749] = 1'b1;  addr_rom[  749]='h00000bb4;  wr_data_rom[  749]='h000002fd;
    rd_cycle[  750] = 1'b0;  wr_cycle[  750] = 1'b1;  addr_rom[  750]='h00000bb8;  wr_data_rom[  750]='h00000a70;
    rd_cycle[  751] = 1'b0;  wr_cycle[  751] = 1'b1;  addr_rom[  751]='h00000bbc;  wr_data_rom[  751]='h00000b85;
    rd_cycle[  752] = 1'b0;  wr_cycle[  752] = 1'b1;  addr_rom[  752]='h00000bc0;  wr_data_rom[  752]='h00000978;
    rd_cycle[  753] = 1'b0;  wr_cycle[  753] = 1'b1;  addr_rom[  753]='h00000bc4;  wr_data_rom[  753]='h000007cb;
    rd_cycle[  754] = 1'b0;  wr_cycle[  754] = 1'b1;  addr_rom[  754]='h00000bc8;  wr_data_rom[  754]='h000009c2;
    rd_cycle[  755] = 1'b0;  wr_cycle[  755] = 1'b1;  addr_rom[  755]='h00000bcc;  wr_data_rom[  755]='h000001b4;
    rd_cycle[  756] = 1'b0;  wr_cycle[  756] = 1'b1;  addr_rom[  756]='h00000bd0;  wr_data_rom[  756]='h000005ca;
    rd_cycle[  757] = 1'b0;  wr_cycle[  757] = 1'b1;  addr_rom[  757]='h00000bd4;  wr_data_rom[  757]='h00000ce6;
    rd_cycle[  758] = 1'b0;  wr_cycle[  758] = 1'b1;  addr_rom[  758]='h00000bd8;  wr_data_rom[  758]='h000005dc;
    rd_cycle[  759] = 1'b0;  wr_cycle[  759] = 1'b1;  addr_rom[  759]='h00000bdc;  wr_data_rom[  759]='h0000024a;
    rd_cycle[  760] = 1'b0;  wr_cycle[  760] = 1'b1;  addr_rom[  760]='h00000be0;  wr_data_rom[  760]='h000001ee;
    rd_cycle[  761] = 1'b0;  wr_cycle[  761] = 1'b1;  addr_rom[  761]='h00000be4;  wr_data_rom[  761]='h00000476;
    rd_cycle[  762] = 1'b0;  wr_cycle[  762] = 1'b1;  addr_rom[  762]='h00000be8;  wr_data_rom[  762]='h0000055c;
    rd_cycle[  763] = 1'b0;  wr_cycle[  763] = 1'b1;  addr_rom[  763]='h00000bec;  wr_data_rom[  763]='h000000fb;
    rd_cycle[  764] = 1'b0;  wr_cycle[  764] = 1'b1;  addr_rom[  764]='h00000bf0;  wr_data_rom[  764]='h00000238;
    rd_cycle[  765] = 1'b0;  wr_cycle[  765] = 1'b1;  addr_rom[  765]='h00000bf4;  wr_data_rom[  765]='h0000029c;
    rd_cycle[  766] = 1'b0;  wr_cycle[  766] = 1'b1;  addr_rom[  766]='h00000bf8;  wr_data_rom[  766]='h00000a30;
    rd_cycle[  767] = 1'b0;  wr_cycle[  767] = 1'b1;  addr_rom[  767]='h00000bfc;  wr_data_rom[  767]='h00000cc6;
    rd_cycle[  768] = 1'b0;  wr_cycle[  768] = 1'b1;  addr_rom[  768]='h00000c00;  wr_data_rom[  768]='h00000684;
    rd_cycle[  769] = 1'b0;  wr_cycle[  769] = 1'b1;  addr_rom[  769]='h00000c04;  wr_data_rom[  769]='h00000a89;
    rd_cycle[  770] = 1'b0;  wr_cycle[  770] = 1'b1;  addr_rom[  770]='h00000c08;  wr_data_rom[  770]='h00000044;
    rd_cycle[  771] = 1'b0;  wr_cycle[  771] = 1'b1;  addr_rom[  771]='h00000c0c;  wr_data_rom[  771]='h00000db5;
    rd_cycle[  772] = 1'b0;  wr_cycle[  772] = 1'b1;  addr_rom[  772]='h00000c10;  wr_data_rom[  772]='h000004f1;
    rd_cycle[  773] = 1'b0;  wr_cycle[  773] = 1'b1;  addr_rom[  773]='h00000c14;  wr_data_rom[  773]='h000001ff;
    rd_cycle[  774] = 1'b0;  wr_cycle[  774] = 1'b1;  addr_rom[  774]='h00000c18;  wr_data_rom[  774]='h00000d8f;
    rd_cycle[  775] = 1'b0;  wr_cycle[  775] = 1'b1;  addr_rom[  775]='h00000c1c;  wr_data_rom[  775]='h00000f41;
    rd_cycle[  776] = 1'b0;  wr_cycle[  776] = 1'b1;  addr_rom[  776]='h00000c20;  wr_data_rom[  776]='h000005d3;
    rd_cycle[  777] = 1'b0;  wr_cycle[  777] = 1'b1;  addr_rom[  777]='h00000c24;  wr_data_rom[  777]='h00000bce;
    rd_cycle[  778] = 1'b0;  wr_cycle[  778] = 1'b1;  addr_rom[  778]='h00000c28;  wr_data_rom[  778]='h000006be;
    rd_cycle[  779] = 1'b0;  wr_cycle[  779] = 1'b1;  addr_rom[  779]='h00000c2c;  wr_data_rom[  779]='h00000531;
    rd_cycle[  780] = 1'b0;  wr_cycle[  780] = 1'b1;  addr_rom[  780]='h00000c30;  wr_data_rom[  780]='h000008ea;
    rd_cycle[  781] = 1'b0;  wr_cycle[  781] = 1'b1;  addr_rom[  781]='h00000c34;  wr_data_rom[  781]='h00000418;
    rd_cycle[  782] = 1'b0;  wr_cycle[  782] = 1'b1;  addr_rom[  782]='h00000c38;  wr_data_rom[  782]='h0000071e;
    rd_cycle[  783] = 1'b0;  wr_cycle[  783] = 1'b1;  addr_rom[  783]='h00000c3c;  wr_data_rom[  783]='h00000269;
    rd_cycle[  784] = 1'b0;  wr_cycle[  784] = 1'b1;  addr_rom[  784]='h00000c40;  wr_data_rom[  784]='h000008a9;
    rd_cycle[  785] = 1'b0;  wr_cycle[  785] = 1'b1;  addr_rom[  785]='h00000c44;  wr_data_rom[  785]='h00000a80;
    rd_cycle[  786] = 1'b0;  wr_cycle[  786] = 1'b1;  addr_rom[  786]='h00000c48;  wr_data_rom[  786]='h00000901;
    rd_cycle[  787] = 1'b0;  wr_cycle[  787] = 1'b1;  addr_rom[  787]='h00000c4c;  wr_data_rom[  787]='h00000f52;
    rd_cycle[  788] = 1'b0;  wr_cycle[  788] = 1'b1;  addr_rom[  788]='h00000c50;  wr_data_rom[  788]='h00000bc7;
    rd_cycle[  789] = 1'b0;  wr_cycle[  789] = 1'b1;  addr_rom[  789]='h00000c54;  wr_data_rom[  789]='h0000040a;
    rd_cycle[  790] = 1'b0;  wr_cycle[  790] = 1'b1;  addr_rom[  790]='h00000c58;  wr_data_rom[  790]='h0000019c;
    rd_cycle[  791] = 1'b0;  wr_cycle[  791] = 1'b1;  addr_rom[  791]='h00000c5c;  wr_data_rom[  791]='h00000b5d;
    rd_cycle[  792] = 1'b0;  wr_cycle[  792] = 1'b1;  addr_rom[  792]='h00000c60;  wr_data_rom[  792]='h0000085f;
    rd_cycle[  793] = 1'b0;  wr_cycle[  793] = 1'b1;  addr_rom[  793]='h00000c64;  wr_data_rom[  793]='h0000098e;
    rd_cycle[  794] = 1'b0;  wr_cycle[  794] = 1'b1;  addr_rom[  794]='h00000c68;  wr_data_rom[  794]='h00000501;
    rd_cycle[  795] = 1'b0;  wr_cycle[  795] = 1'b1;  addr_rom[  795]='h00000c6c;  wr_data_rom[  795]='h0000095a;
    rd_cycle[  796] = 1'b0;  wr_cycle[  796] = 1'b1;  addr_rom[  796]='h00000c70;  wr_data_rom[  796]='h0000049f;
    rd_cycle[  797] = 1'b0;  wr_cycle[  797] = 1'b1;  addr_rom[  797]='h00000c74;  wr_data_rom[  797]='h00000e8a;
    rd_cycle[  798] = 1'b0;  wr_cycle[  798] = 1'b1;  addr_rom[  798]='h00000c78;  wr_data_rom[  798]='h00000f24;
    rd_cycle[  799] = 1'b0;  wr_cycle[  799] = 1'b1;  addr_rom[  799]='h00000c7c;  wr_data_rom[  799]='h00000054;
    rd_cycle[  800] = 1'b0;  wr_cycle[  800] = 1'b1;  addr_rom[  800]='h00000c80;  wr_data_rom[  800]='h0000061d;
    rd_cycle[  801] = 1'b0;  wr_cycle[  801] = 1'b1;  addr_rom[  801]='h00000c84;  wr_data_rom[  801]='h00000894;
    rd_cycle[  802] = 1'b0;  wr_cycle[  802] = 1'b1;  addr_rom[  802]='h00000c88;  wr_data_rom[  802]='h00000401;
    rd_cycle[  803] = 1'b0;  wr_cycle[  803] = 1'b1;  addr_rom[  803]='h00000c8c;  wr_data_rom[  803]='h0000084e;
    rd_cycle[  804] = 1'b0;  wr_cycle[  804] = 1'b1;  addr_rom[  804]='h00000c90;  wr_data_rom[  804]='h00000762;
    rd_cycle[  805] = 1'b0;  wr_cycle[  805] = 1'b1;  addr_rom[  805]='h00000c94;  wr_data_rom[  805]='h0000013b;
    rd_cycle[  806] = 1'b0;  wr_cycle[  806] = 1'b1;  addr_rom[  806]='h00000c98;  wr_data_rom[  806]='h00000ee1;
    rd_cycle[  807] = 1'b0;  wr_cycle[  807] = 1'b1;  addr_rom[  807]='h00000c9c;  wr_data_rom[  807]='h00000d43;
    rd_cycle[  808] = 1'b0;  wr_cycle[  808] = 1'b1;  addr_rom[  808]='h00000ca0;  wr_data_rom[  808]='h000006e5;
    rd_cycle[  809] = 1'b0;  wr_cycle[  809] = 1'b1;  addr_rom[  809]='h00000ca4;  wr_data_rom[  809]='h0000039b;
    rd_cycle[  810] = 1'b0;  wr_cycle[  810] = 1'b1;  addr_rom[  810]='h00000ca8;  wr_data_rom[  810]='h0000050f;
    rd_cycle[  811] = 1'b0;  wr_cycle[  811] = 1'b1;  addr_rom[  811]='h00000cac;  wr_data_rom[  811]='h000003cd;
    rd_cycle[  812] = 1'b0;  wr_cycle[  812] = 1'b1;  addr_rom[  812]='h00000cb0;  wr_data_rom[  812]='h0000077d;
    rd_cycle[  813] = 1'b0;  wr_cycle[  813] = 1'b1;  addr_rom[  813]='h00000cb4;  wr_data_rom[  813]='h000000f3;
    rd_cycle[  814] = 1'b0;  wr_cycle[  814] = 1'b1;  addr_rom[  814]='h00000cb8;  wr_data_rom[  814]='h00000393;
    rd_cycle[  815] = 1'b0;  wr_cycle[  815] = 1'b1;  addr_rom[  815]='h00000cbc;  wr_data_rom[  815]='h00000d76;
    rd_cycle[  816] = 1'b0;  wr_cycle[  816] = 1'b1;  addr_rom[  816]='h00000cc0;  wr_data_rom[  816]='h00000b38;
    rd_cycle[  817] = 1'b0;  wr_cycle[  817] = 1'b1;  addr_rom[  817]='h00000cc4;  wr_data_rom[  817]='h00000834;
    rd_cycle[  818] = 1'b0;  wr_cycle[  818] = 1'b1;  addr_rom[  818]='h00000cc8;  wr_data_rom[  818]='h00000296;
    rd_cycle[  819] = 1'b0;  wr_cycle[  819] = 1'b1;  addr_rom[  819]='h00000ccc;  wr_data_rom[  819]='h00000d36;
    rd_cycle[  820] = 1'b0;  wr_cycle[  820] = 1'b1;  addr_rom[  820]='h00000cd0;  wr_data_rom[  820]='h00000f22;
    rd_cycle[  821] = 1'b0;  wr_cycle[  821] = 1'b1;  addr_rom[  821]='h00000cd4;  wr_data_rom[  821]='h000008c2;
    rd_cycle[  822] = 1'b0;  wr_cycle[  822] = 1'b1;  addr_rom[  822]='h00000cd8;  wr_data_rom[  822]='h00000d95;
    rd_cycle[  823] = 1'b0;  wr_cycle[  823] = 1'b1;  addr_rom[  823]='h00000cdc;  wr_data_rom[  823]='h00000edd;
    rd_cycle[  824] = 1'b0;  wr_cycle[  824] = 1'b1;  addr_rom[  824]='h00000ce0;  wr_data_rom[  824]='h00000209;
    rd_cycle[  825] = 1'b0;  wr_cycle[  825] = 1'b1;  addr_rom[  825]='h00000ce4;  wr_data_rom[  825]='h00000436;
    rd_cycle[  826] = 1'b0;  wr_cycle[  826] = 1'b1;  addr_rom[  826]='h00000ce8;  wr_data_rom[  826]='h0000016b;
    rd_cycle[  827] = 1'b0;  wr_cycle[  827] = 1'b1;  addr_rom[  827]='h00000cec;  wr_data_rom[  827]='h00000084;
    rd_cycle[  828] = 1'b0;  wr_cycle[  828] = 1'b1;  addr_rom[  828]='h00000cf0;  wr_data_rom[  828]='h00000752;
    rd_cycle[  829] = 1'b0;  wr_cycle[  829] = 1'b1;  addr_rom[  829]='h00000cf4;  wr_data_rom[  829]='h000006bb;
    rd_cycle[  830] = 1'b0;  wr_cycle[  830] = 1'b1;  addr_rom[  830]='h00000cf8;  wr_data_rom[  830]='h00000b62;
    rd_cycle[  831] = 1'b0;  wr_cycle[  831] = 1'b1;  addr_rom[  831]='h00000cfc;  wr_data_rom[  831]='h00000e4e;
    rd_cycle[  832] = 1'b0;  wr_cycle[  832] = 1'b1;  addr_rom[  832]='h00000d00;  wr_data_rom[  832]='h000002f8;
    rd_cycle[  833] = 1'b0;  wr_cycle[  833] = 1'b1;  addr_rom[  833]='h00000d04;  wr_data_rom[  833]='h0000011e;
    rd_cycle[  834] = 1'b0;  wr_cycle[  834] = 1'b1;  addr_rom[  834]='h00000d08;  wr_data_rom[  834]='h00000f74;
    rd_cycle[  835] = 1'b0;  wr_cycle[  835] = 1'b1;  addr_rom[  835]='h00000d0c;  wr_data_rom[  835]='h00000cee;
    rd_cycle[  836] = 1'b0;  wr_cycle[  836] = 1'b1;  addr_rom[  836]='h00000d10;  wr_data_rom[  836]='h0000004a;
    rd_cycle[  837] = 1'b0;  wr_cycle[  837] = 1'b1;  addr_rom[  837]='h00000d14;  wr_data_rom[  837]='h00000500;
    rd_cycle[  838] = 1'b0;  wr_cycle[  838] = 1'b1;  addr_rom[  838]='h00000d18;  wr_data_rom[  838]='h00000771;
    rd_cycle[  839] = 1'b0;  wr_cycle[  839] = 1'b1;  addr_rom[  839]='h00000d1c;  wr_data_rom[  839]='h000007f4;
    rd_cycle[  840] = 1'b0;  wr_cycle[  840] = 1'b1;  addr_rom[  840]='h00000d20;  wr_data_rom[  840]='h00000789;
    rd_cycle[  841] = 1'b0;  wr_cycle[  841] = 1'b1;  addr_rom[  841]='h00000d24;  wr_data_rom[  841]='h00000120;
    rd_cycle[  842] = 1'b0;  wr_cycle[  842] = 1'b1;  addr_rom[  842]='h00000d28;  wr_data_rom[  842]='h00000604;
    rd_cycle[  843] = 1'b0;  wr_cycle[  843] = 1'b1;  addr_rom[  843]='h00000d2c;  wr_data_rom[  843]='h00000276;
    rd_cycle[  844] = 1'b0;  wr_cycle[  844] = 1'b1;  addr_rom[  844]='h00000d30;  wr_data_rom[  844]='h00000f26;
    rd_cycle[  845] = 1'b0;  wr_cycle[  845] = 1'b1;  addr_rom[  845]='h00000d34;  wr_data_rom[  845]='h00000113;
    rd_cycle[  846] = 1'b0;  wr_cycle[  846] = 1'b1;  addr_rom[  846]='h00000d38;  wr_data_rom[  846]='h00000dd4;
    rd_cycle[  847] = 1'b0;  wr_cycle[  847] = 1'b1;  addr_rom[  847]='h00000d3c;  wr_data_rom[  847]='h00000dbe;
    rd_cycle[  848] = 1'b0;  wr_cycle[  848] = 1'b1;  addr_rom[  848]='h00000d40;  wr_data_rom[  848]='h000001b9;
    rd_cycle[  849] = 1'b0;  wr_cycle[  849] = 1'b1;  addr_rom[  849]='h00000d44;  wr_data_rom[  849]='h00000c13;
    rd_cycle[  850] = 1'b0;  wr_cycle[  850] = 1'b1;  addr_rom[  850]='h00000d48;  wr_data_rom[  850]='h00000c00;
    rd_cycle[  851] = 1'b0;  wr_cycle[  851] = 1'b1;  addr_rom[  851]='h00000d4c;  wr_data_rom[  851]='h0000016e;
    rd_cycle[  852] = 1'b0;  wr_cycle[  852] = 1'b1;  addr_rom[  852]='h00000d50;  wr_data_rom[  852]='h00000e14;
    rd_cycle[  853] = 1'b0;  wr_cycle[  853] = 1'b1;  addr_rom[  853]='h00000d54;  wr_data_rom[  853]='h00000dc3;
    rd_cycle[  854] = 1'b0;  wr_cycle[  854] = 1'b1;  addr_rom[  854]='h00000d58;  wr_data_rom[  854]='h0000081a;
    rd_cycle[  855] = 1'b0;  wr_cycle[  855] = 1'b1;  addr_rom[  855]='h00000d5c;  wr_data_rom[  855]='h000009b5;
    rd_cycle[  856] = 1'b0;  wr_cycle[  856] = 1'b1;  addr_rom[  856]='h00000d60;  wr_data_rom[  856]='h00000cb6;
    rd_cycle[  857] = 1'b0;  wr_cycle[  857] = 1'b1;  addr_rom[  857]='h00000d64;  wr_data_rom[  857]='h00000e41;
    rd_cycle[  858] = 1'b0;  wr_cycle[  858] = 1'b1;  addr_rom[  858]='h00000d68;  wr_data_rom[  858]='h00000f73;
    rd_cycle[  859] = 1'b0;  wr_cycle[  859] = 1'b1;  addr_rom[  859]='h00000d6c;  wr_data_rom[  859]='h00000713;
    rd_cycle[  860] = 1'b0;  wr_cycle[  860] = 1'b1;  addr_rom[  860]='h00000d70;  wr_data_rom[  860]='h00000e4c;
    rd_cycle[  861] = 1'b0;  wr_cycle[  861] = 1'b1;  addr_rom[  861]='h00000d74;  wr_data_rom[  861]='h0000021a;
    rd_cycle[  862] = 1'b0;  wr_cycle[  862] = 1'b1;  addr_rom[  862]='h00000d78;  wr_data_rom[  862]='h000006ee;
    rd_cycle[  863] = 1'b0;  wr_cycle[  863] = 1'b1;  addr_rom[  863]='h00000d7c;  wr_data_rom[  863]='h00000b90;
    rd_cycle[  864] = 1'b0;  wr_cycle[  864] = 1'b1;  addr_rom[  864]='h00000d80;  wr_data_rom[  864]='h00000c43;
    rd_cycle[  865] = 1'b0;  wr_cycle[  865] = 1'b1;  addr_rom[  865]='h00000d84;  wr_data_rom[  865]='h00000b6a;
    rd_cycle[  866] = 1'b0;  wr_cycle[  866] = 1'b1;  addr_rom[  866]='h00000d88;  wr_data_rom[  866]='h00000212;
    rd_cycle[  867] = 1'b0;  wr_cycle[  867] = 1'b1;  addr_rom[  867]='h00000d8c;  wr_data_rom[  867]='h00000655;
    rd_cycle[  868] = 1'b0;  wr_cycle[  868] = 1'b1;  addr_rom[  868]='h00000d90;  wr_data_rom[  868]='h00000a7c;
    rd_cycle[  869] = 1'b0;  wr_cycle[  869] = 1'b1;  addr_rom[  869]='h00000d94;  wr_data_rom[  869]='h00000594;
    rd_cycle[  870] = 1'b0;  wr_cycle[  870] = 1'b1;  addr_rom[  870]='h00000d98;  wr_data_rom[  870]='h00000f8c;
    rd_cycle[  871] = 1'b0;  wr_cycle[  871] = 1'b1;  addr_rom[  871]='h00000d9c;  wr_data_rom[  871]='h00000937;
    rd_cycle[  872] = 1'b0;  wr_cycle[  872] = 1'b1;  addr_rom[  872]='h00000da0;  wr_data_rom[  872]='h00000a10;
    rd_cycle[  873] = 1'b0;  wr_cycle[  873] = 1'b1;  addr_rom[  873]='h00000da4;  wr_data_rom[  873]='h00000b61;
    rd_cycle[  874] = 1'b0;  wr_cycle[  874] = 1'b1;  addr_rom[  874]='h00000da8;  wr_data_rom[  874]='h00000078;
    rd_cycle[  875] = 1'b0;  wr_cycle[  875] = 1'b1;  addr_rom[  875]='h00000dac;  wr_data_rom[  875]='h00000af4;
    rd_cycle[  876] = 1'b0;  wr_cycle[  876] = 1'b1;  addr_rom[  876]='h00000db0;  wr_data_rom[  876]='h00000313;
    rd_cycle[  877] = 1'b0;  wr_cycle[  877] = 1'b1;  addr_rom[  877]='h00000db4;  wr_data_rom[  877]='h00000a85;
    rd_cycle[  878] = 1'b0;  wr_cycle[  878] = 1'b1;  addr_rom[  878]='h00000db8;  wr_data_rom[  878]='h0000085b;
    rd_cycle[  879] = 1'b0;  wr_cycle[  879] = 1'b1;  addr_rom[  879]='h00000dbc;  wr_data_rom[  879]='h00000dd1;
    rd_cycle[  880] = 1'b0;  wr_cycle[  880] = 1'b1;  addr_rom[  880]='h00000dc0;  wr_data_rom[  880]='h00000a3b;
    rd_cycle[  881] = 1'b0;  wr_cycle[  881] = 1'b1;  addr_rom[  881]='h00000dc4;  wr_data_rom[  881]='h00000ad2;
    rd_cycle[  882] = 1'b0;  wr_cycle[  882] = 1'b1;  addr_rom[  882]='h00000dc8;  wr_data_rom[  882]='h00000ab6;
    rd_cycle[  883] = 1'b0;  wr_cycle[  883] = 1'b1;  addr_rom[  883]='h00000dcc;  wr_data_rom[  883]='h0000080d;
    rd_cycle[  884] = 1'b0;  wr_cycle[  884] = 1'b1;  addr_rom[  884]='h00000dd0;  wr_data_rom[  884]='h000000f1;
    rd_cycle[  885] = 1'b0;  wr_cycle[  885] = 1'b1;  addr_rom[  885]='h00000dd4;  wr_data_rom[  885]='h0000064f;
    rd_cycle[  886] = 1'b0;  wr_cycle[  886] = 1'b1;  addr_rom[  886]='h00000dd8;  wr_data_rom[  886]='h0000097e;
    rd_cycle[  887] = 1'b0;  wr_cycle[  887] = 1'b1;  addr_rom[  887]='h00000ddc;  wr_data_rom[  887]='h00000e27;
    rd_cycle[  888] = 1'b0;  wr_cycle[  888] = 1'b1;  addr_rom[  888]='h00000de0;  wr_data_rom[  888]='h00000bea;
    rd_cycle[  889] = 1'b0;  wr_cycle[  889] = 1'b1;  addr_rom[  889]='h00000de4;  wr_data_rom[  889]='h00000648;
    rd_cycle[  890] = 1'b0;  wr_cycle[  890] = 1'b1;  addr_rom[  890]='h00000de8;  wr_data_rom[  890]='h000007f3;
    rd_cycle[  891] = 1'b0;  wr_cycle[  891] = 1'b1;  addr_rom[  891]='h00000dec;  wr_data_rom[  891]='h00000e44;
    rd_cycle[  892] = 1'b0;  wr_cycle[  892] = 1'b1;  addr_rom[  892]='h00000df0;  wr_data_rom[  892]='h00000f3e;
    rd_cycle[  893] = 1'b0;  wr_cycle[  893] = 1'b1;  addr_rom[  893]='h00000df4;  wr_data_rom[  893]='h0000044a;
    rd_cycle[  894] = 1'b0;  wr_cycle[  894] = 1'b1;  addr_rom[  894]='h00000df8;  wr_data_rom[  894]='h00000e65;
    rd_cycle[  895] = 1'b0;  wr_cycle[  895] = 1'b1;  addr_rom[  895]='h00000dfc;  wr_data_rom[  895]='h00000629;
    rd_cycle[  896] = 1'b0;  wr_cycle[  896] = 1'b1;  addr_rom[  896]='h00000e00;  wr_data_rom[  896]='h000002f8;
    rd_cycle[  897] = 1'b0;  wr_cycle[  897] = 1'b1;  addr_rom[  897]='h00000e04;  wr_data_rom[  897]='h00000492;
    rd_cycle[  898] = 1'b0;  wr_cycle[  898] = 1'b1;  addr_rom[  898]='h00000e08;  wr_data_rom[  898]='h00000d3d;
    rd_cycle[  899] = 1'b0;  wr_cycle[  899] = 1'b1;  addr_rom[  899]='h00000e0c;  wr_data_rom[  899]='h00000a75;
    rd_cycle[  900] = 1'b0;  wr_cycle[  900] = 1'b1;  addr_rom[  900]='h00000e10;  wr_data_rom[  900]='h00000312;
    rd_cycle[  901] = 1'b0;  wr_cycle[  901] = 1'b1;  addr_rom[  901]='h00000e14;  wr_data_rom[  901]='h00000010;
    rd_cycle[  902] = 1'b0;  wr_cycle[  902] = 1'b1;  addr_rom[  902]='h00000e18;  wr_data_rom[  902]='h00000201;
    rd_cycle[  903] = 1'b0;  wr_cycle[  903] = 1'b1;  addr_rom[  903]='h00000e1c;  wr_data_rom[  903]='h00000a07;
    rd_cycle[  904] = 1'b0;  wr_cycle[  904] = 1'b1;  addr_rom[  904]='h00000e20;  wr_data_rom[  904]='h00000654;
    rd_cycle[  905] = 1'b0;  wr_cycle[  905] = 1'b1;  addr_rom[  905]='h00000e24;  wr_data_rom[  905]='h0000083a;
    rd_cycle[  906] = 1'b0;  wr_cycle[  906] = 1'b1;  addr_rom[  906]='h00000e28;  wr_data_rom[  906]='h000007b2;
    rd_cycle[  907] = 1'b0;  wr_cycle[  907] = 1'b1;  addr_rom[  907]='h00000e2c;  wr_data_rom[  907]='h00000546;
    rd_cycle[  908] = 1'b0;  wr_cycle[  908] = 1'b1;  addr_rom[  908]='h00000e30;  wr_data_rom[  908]='h00000a8a;
    rd_cycle[  909] = 1'b0;  wr_cycle[  909] = 1'b1;  addr_rom[  909]='h00000e34;  wr_data_rom[  909]='h00000869;
    rd_cycle[  910] = 1'b0;  wr_cycle[  910] = 1'b1;  addr_rom[  910]='h00000e38;  wr_data_rom[  910]='h000009fa;
    rd_cycle[  911] = 1'b0;  wr_cycle[  911] = 1'b1;  addr_rom[  911]='h00000e3c;  wr_data_rom[  911]='h00000525;
    rd_cycle[  912] = 1'b0;  wr_cycle[  912] = 1'b1;  addr_rom[  912]='h00000e40;  wr_data_rom[  912]='h00000266;
    rd_cycle[  913] = 1'b0;  wr_cycle[  913] = 1'b1;  addr_rom[  913]='h00000e44;  wr_data_rom[  913]='h00000b40;
    rd_cycle[  914] = 1'b0;  wr_cycle[  914] = 1'b1;  addr_rom[  914]='h00000e48;  wr_data_rom[  914]='h000005b0;
    rd_cycle[  915] = 1'b0;  wr_cycle[  915] = 1'b1;  addr_rom[  915]='h00000e4c;  wr_data_rom[  915]='h00000f76;
    rd_cycle[  916] = 1'b0;  wr_cycle[  916] = 1'b1;  addr_rom[  916]='h00000e50;  wr_data_rom[  916]='h00000460;
    rd_cycle[  917] = 1'b0;  wr_cycle[  917] = 1'b1;  addr_rom[  917]='h00000e54;  wr_data_rom[  917]='h00000153;
    rd_cycle[  918] = 1'b0;  wr_cycle[  918] = 1'b1;  addr_rom[  918]='h00000e58;  wr_data_rom[  918]='h0000049f;
    rd_cycle[  919] = 1'b0;  wr_cycle[  919] = 1'b1;  addr_rom[  919]='h00000e5c;  wr_data_rom[  919]='h00000a96;
    rd_cycle[  920] = 1'b0;  wr_cycle[  920] = 1'b1;  addr_rom[  920]='h00000e60;  wr_data_rom[  920]='h000009f5;
    rd_cycle[  921] = 1'b0;  wr_cycle[  921] = 1'b1;  addr_rom[  921]='h00000e64;  wr_data_rom[  921]='h0000008c;
    rd_cycle[  922] = 1'b0;  wr_cycle[  922] = 1'b1;  addr_rom[  922]='h00000e68;  wr_data_rom[  922]='h00000644;
    rd_cycle[  923] = 1'b0;  wr_cycle[  923] = 1'b1;  addr_rom[  923]='h00000e6c;  wr_data_rom[  923]='h000008b9;
    rd_cycle[  924] = 1'b0;  wr_cycle[  924] = 1'b1;  addr_rom[  924]='h00000e70;  wr_data_rom[  924]='h00000f45;
    rd_cycle[  925] = 1'b0;  wr_cycle[  925] = 1'b1;  addr_rom[  925]='h00000e74;  wr_data_rom[  925]='h0000061a;
    rd_cycle[  926] = 1'b0;  wr_cycle[  926] = 1'b1;  addr_rom[  926]='h00000e78;  wr_data_rom[  926]='h00000693;
    rd_cycle[  927] = 1'b0;  wr_cycle[  927] = 1'b1;  addr_rom[  927]='h00000e7c;  wr_data_rom[  927]='h000008c9;
    rd_cycle[  928] = 1'b0;  wr_cycle[  928] = 1'b1;  addr_rom[  928]='h00000e80;  wr_data_rom[  928]='h000006b0;
    rd_cycle[  929] = 1'b0;  wr_cycle[  929] = 1'b1;  addr_rom[  929]='h00000e84;  wr_data_rom[  929]='h00000bd7;
    rd_cycle[  930] = 1'b0;  wr_cycle[  930] = 1'b1;  addr_rom[  930]='h00000e88;  wr_data_rom[  930]='h0000003b;
    rd_cycle[  931] = 1'b0;  wr_cycle[  931] = 1'b1;  addr_rom[  931]='h00000e8c;  wr_data_rom[  931]='h00000f7f;
    rd_cycle[  932] = 1'b0;  wr_cycle[  932] = 1'b1;  addr_rom[  932]='h00000e90;  wr_data_rom[  932]='h00000294;
    rd_cycle[  933] = 1'b0;  wr_cycle[  933] = 1'b1;  addr_rom[  933]='h00000e94;  wr_data_rom[  933]='h000007e7;
    rd_cycle[  934] = 1'b0;  wr_cycle[  934] = 1'b1;  addr_rom[  934]='h00000e98;  wr_data_rom[  934]='h00000f23;
    rd_cycle[  935] = 1'b0;  wr_cycle[  935] = 1'b1;  addr_rom[  935]='h00000e9c;  wr_data_rom[  935]='h000007fc;
    rd_cycle[  936] = 1'b0;  wr_cycle[  936] = 1'b1;  addr_rom[  936]='h00000ea0;  wr_data_rom[  936]='h00000352;
    rd_cycle[  937] = 1'b0;  wr_cycle[  937] = 1'b1;  addr_rom[  937]='h00000ea4;  wr_data_rom[  937]='h00000626;
    rd_cycle[  938] = 1'b0;  wr_cycle[  938] = 1'b1;  addr_rom[  938]='h00000ea8;  wr_data_rom[  938]='h000001b2;
    rd_cycle[  939] = 1'b0;  wr_cycle[  939] = 1'b1;  addr_rom[  939]='h00000eac;  wr_data_rom[  939]='h000008e9;
    rd_cycle[  940] = 1'b0;  wr_cycle[  940] = 1'b1;  addr_rom[  940]='h00000eb0;  wr_data_rom[  940]='h00000a1d;
    rd_cycle[  941] = 1'b0;  wr_cycle[  941] = 1'b1;  addr_rom[  941]='h00000eb4;  wr_data_rom[  941]='h0000037f;
    rd_cycle[  942] = 1'b0;  wr_cycle[  942] = 1'b1;  addr_rom[  942]='h00000eb8;  wr_data_rom[  942]='h000006a6;
    rd_cycle[  943] = 1'b0;  wr_cycle[  943] = 1'b1;  addr_rom[  943]='h00000ebc;  wr_data_rom[  943]='h0000021d;
    rd_cycle[  944] = 1'b0;  wr_cycle[  944] = 1'b1;  addr_rom[  944]='h00000ec0;  wr_data_rom[  944]='h00000835;
    rd_cycle[  945] = 1'b0;  wr_cycle[  945] = 1'b1;  addr_rom[  945]='h00000ec4;  wr_data_rom[  945]='h00000f73;
    rd_cycle[  946] = 1'b0;  wr_cycle[  946] = 1'b1;  addr_rom[  946]='h00000ec8;  wr_data_rom[  946]='h00000442;
    rd_cycle[  947] = 1'b0;  wr_cycle[  947] = 1'b1;  addr_rom[  947]='h00000ecc;  wr_data_rom[  947]='h00000b2c;
    rd_cycle[  948] = 1'b0;  wr_cycle[  948] = 1'b1;  addr_rom[  948]='h00000ed0;  wr_data_rom[  948]='h000005e8;
    rd_cycle[  949] = 1'b0;  wr_cycle[  949] = 1'b1;  addr_rom[  949]='h00000ed4;  wr_data_rom[  949]='h00000a4c;
    rd_cycle[  950] = 1'b0;  wr_cycle[  950] = 1'b1;  addr_rom[  950]='h00000ed8;  wr_data_rom[  950]='h00000d6a;
    rd_cycle[  951] = 1'b0;  wr_cycle[  951] = 1'b1;  addr_rom[  951]='h00000edc;  wr_data_rom[  951]='h0000032f;
    rd_cycle[  952] = 1'b0;  wr_cycle[  952] = 1'b1;  addr_rom[  952]='h00000ee0;  wr_data_rom[  952]='h00000734;
    rd_cycle[  953] = 1'b0;  wr_cycle[  953] = 1'b1;  addr_rom[  953]='h00000ee4;  wr_data_rom[  953]='h00000d0f;
    rd_cycle[  954] = 1'b0;  wr_cycle[  954] = 1'b1;  addr_rom[  954]='h00000ee8;  wr_data_rom[  954]='h00000dfb;
    rd_cycle[  955] = 1'b0;  wr_cycle[  955] = 1'b1;  addr_rom[  955]='h00000eec;  wr_data_rom[  955]='h000006b5;
    rd_cycle[  956] = 1'b0;  wr_cycle[  956] = 1'b1;  addr_rom[  956]='h00000ef0;  wr_data_rom[  956]='h00000e93;
    rd_cycle[  957] = 1'b0;  wr_cycle[  957] = 1'b1;  addr_rom[  957]='h00000ef4;  wr_data_rom[  957]='h00000f35;
    rd_cycle[  958] = 1'b0;  wr_cycle[  958] = 1'b1;  addr_rom[  958]='h00000ef8;  wr_data_rom[  958]='h00000f7c;
    rd_cycle[  959] = 1'b0;  wr_cycle[  959] = 1'b1;  addr_rom[  959]='h00000efc;  wr_data_rom[  959]='h000002c8;
    rd_cycle[  960] = 1'b0;  wr_cycle[  960] = 1'b1;  addr_rom[  960]='h00000f00;  wr_data_rom[  960]='h0000051b;
    rd_cycle[  961] = 1'b0;  wr_cycle[  961] = 1'b1;  addr_rom[  961]='h00000f04;  wr_data_rom[  961]='h000006f3;
    rd_cycle[  962] = 1'b0;  wr_cycle[  962] = 1'b1;  addr_rom[  962]='h00000f08;  wr_data_rom[  962]='h000002d7;
    rd_cycle[  963] = 1'b0;  wr_cycle[  963] = 1'b1;  addr_rom[  963]='h00000f0c;  wr_data_rom[  963]='h00000c18;
    rd_cycle[  964] = 1'b0;  wr_cycle[  964] = 1'b1;  addr_rom[  964]='h00000f10;  wr_data_rom[  964]='h00000ed0;
    rd_cycle[  965] = 1'b0;  wr_cycle[  965] = 1'b1;  addr_rom[  965]='h00000f14;  wr_data_rom[  965]='h00000057;
    rd_cycle[  966] = 1'b0;  wr_cycle[  966] = 1'b1;  addr_rom[  966]='h00000f18;  wr_data_rom[  966]='h000000b9;
    rd_cycle[  967] = 1'b0;  wr_cycle[  967] = 1'b1;  addr_rom[  967]='h00000f1c;  wr_data_rom[  967]='h00000729;
    rd_cycle[  968] = 1'b0;  wr_cycle[  968] = 1'b1;  addr_rom[  968]='h00000f20;  wr_data_rom[  968]='h00000922;
    rd_cycle[  969] = 1'b0;  wr_cycle[  969] = 1'b1;  addr_rom[  969]='h00000f24;  wr_data_rom[  969]='h00000392;
    rd_cycle[  970] = 1'b0;  wr_cycle[  970] = 1'b1;  addr_rom[  970]='h00000f28;  wr_data_rom[  970]='h000001e6;
    rd_cycle[  971] = 1'b0;  wr_cycle[  971] = 1'b1;  addr_rom[  971]='h00000f2c;  wr_data_rom[  971]='h000006b6;
    rd_cycle[  972] = 1'b0;  wr_cycle[  972] = 1'b1;  addr_rom[  972]='h00000f30;  wr_data_rom[  972]='h00000ebb;
    rd_cycle[  973] = 1'b0;  wr_cycle[  973] = 1'b1;  addr_rom[  973]='h00000f34;  wr_data_rom[  973]='h0000002e;
    rd_cycle[  974] = 1'b0;  wr_cycle[  974] = 1'b1;  addr_rom[  974]='h00000f38;  wr_data_rom[  974]='h00000ced;
    rd_cycle[  975] = 1'b0;  wr_cycle[  975] = 1'b1;  addr_rom[  975]='h00000f3c;  wr_data_rom[  975]='h00000433;
    rd_cycle[  976] = 1'b0;  wr_cycle[  976] = 1'b1;  addr_rom[  976]='h00000f40;  wr_data_rom[  976]='h000004e5;
    rd_cycle[  977] = 1'b0;  wr_cycle[  977] = 1'b1;  addr_rom[  977]='h00000f44;  wr_data_rom[  977]='h00000354;
    rd_cycle[  978] = 1'b0;  wr_cycle[  978] = 1'b1;  addr_rom[  978]='h00000f48;  wr_data_rom[  978]='h00000c89;
    rd_cycle[  979] = 1'b0;  wr_cycle[  979] = 1'b1;  addr_rom[  979]='h00000f4c;  wr_data_rom[  979]='h000006db;
    rd_cycle[  980] = 1'b0;  wr_cycle[  980] = 1'b1;  addr_rom[  980]='h00000f50;  wr_data_rom[  980]='h00000f16;
    rd_cycle[  981] = 1'b0;  wr_cycle[  981] = 1'b1;  addr_rom[  981]='h00000f54;  wr_data_rom[  981]='h000008e6;
    rd_cycle[  982] = 1'b0;  wr_cycle[  982] = 1'b1;  addr_rom[  982]='h00000f58;  wr_data_rom[  982]='h00000537;
    rd_cycle[  983] = 1'b0;  wr_cycle[  983] = 1'b1;  addr_rom[  983]='h00000f5c;  wr_data_rom[  983]='h00000072;
    rd_cycle[  984] = 1'b0;  wr_cycle[  984] = 1'b1;  addr_rom[  984]='h00000f60;  wr_data_rom[  984]='h00000f6e;
    rd_cycle[  985] = 1'b0;  wr_cycle[  985] = 1'b1;  addr_rom[  985]='h00000f64;  wr_data_rom[  985]='h000003fc;
    rd_cycle[  986] = 1'b0;  wr_cycle[  986] = 1'b1;  addr_rom[  986]='h00000f68;  wr_data_rom[  986]='h00000bc1;
    rd_cycle[  987] = 1'b0;  wr_cycle[  987] = 1'b1;  addr_rom[  987]='h00000f6c;  wr_data_rom[  987]='h0000096f;
    rd_cycle[  988] = 1'b0;  wr_cycle[  988] = 1'b1;  addr_rom[  988]='h00000f70;  wr_data_rom[  988]='h00000d0c;
    rd_cycle[  989] = 1'b0;  wr_cycle[  989] = 1'b1;  addr_rom[  989]='h00000f74;  wr_data_rom[  989]='h00000298;
    rd_cycle[  990] = 1'b0;  wr_cycle[  990] = 1'b1;  addr_rom[  990]='h00000f78;  wr_data_rom[  990]='h00000f71;
    rd_cycle[  991] = 1'b0;  wr_cycle[  991] = 1'b1;  addr_rom[  991]='h00000f7c;  wr_data_rom[  991]='h00000e93;
    rd_cycle[  992] = 1'b0;  wr_cycle[  992] = 1'b1;  addr_rom[  992]='h00000f80;  wr_data_rom[  992]='h000005e8;
    rd_cycle[  993] = 1'b0;  wr_cycle[  993] = 1'b1;  addr_rom[  993]='h00000f84;  wr_data_rom[  993]='h00000f27;
    rd_cycle[  994] = 1'b0;  wr_cycle[  994] = 1'b1;  addr_rom[  994]='h00000f88;  wr_data_rom[  994]='h00000262;
    rd_cycle[  995] = 1'b0;  wr_cycle[  995] = 1'b1;  addr_rom[  995]='h00000f8c;  wr_data_rom[  995]='h00000d7d;
    rd_cycle[  996] = 1'b0;  wr_cycle[  996] = 1'b1;  addr_rom[  996]='h00000f90;  wr_data_rom[  996]='h000006b4;
    rd_cycle[  997] = 1'b0;  wr_cycle[  997] = 1'b1;  addr_rom[  997]='h00000f94;  wr_data_rom[  997]='h000004ac;
    rd_cycle[  998] = 1'b0;  wr_cycle[  998] = 1'b1;  addr_rom[  998]='h00000f98;  wr_data_rom[  998]='h0000066d;
    rd_cycle[  999] = 1'b0;  wr_cycle[  999] = 1'b1;  addr_rom[  999]='h00000f9c;  wr_data_rom[  999]='h00000acf;
    // 3000 random read and write cycles
    rd_cycle[ 1000] = 1'b1;  wr_cycle[ 1000] = 1'b0;  addr_rom[ 1000]='h0000073c;  wr_data_rom[ 1000]='h00000000;
    rd_cycle[ 1001] = 1'b0;  wr_cycle[ 1001] = 1'b1;  addr_rom[ 1001]='h00000638;  wr_data_rom[ 1001]='h000003f3;
    rd_cycle[ 1002] = 1'b0;  wr_cycle[ 1002] = 1'b1;  addr_rom[ 1002]='h000004c4;  wr_data_rom[ 1002]='h000005a1;
    rd_cycle[ 1003] = 1'b0;  wr_cycle[ 1003] = 1'b1;  addr_rom[ 1003]='h00000898;  wr_data_rom[ 1003]='h0000014b;
    rd_cycle[ 1004] = 1'b0;  wr_cycle[ 1004] = 1'b1;  addr_rom[ 1004]='h00000ea8;  wr_data_rom[ 1004]='h00000830;
    rd_cycle[ 1005] = 1'b1;  wr_cycle[ 1005] = 1'b0;  addr_rom[ 1005]='h00000df4;  wr_data_rom[ 1005]='h00000000;
    rd_cycle[ 1006] = 1'b0;  wr_cycle[ 1006] = 1'b1;  addr_rom[ 1006]='h000007a0;  wr_data_rom[ 1006]='h00000994;
    rd_cycle[ 1007] = 1'b0;  wr_cycle[ 1007] = 1'b1;  addr_rom[ 1007]='h00000390;  wr_data_rom[ 1007]='h00000f63;
    rd_cycle[ 1008] = 1'b1;  wr_cycle[ 1008] = 1'b0;  addr_rom[ 1008]='h00000100;  wr_data_rom[ 1008]='h00000000;
    rd_cycle[ 1009] = 1'b1;  wr_cycle[ 1009] = 1'b0;  addr_rom[ 1009]='h0000065c;  wr_data_rom[ 1009]='h00000000;
    rd_cycle[ 1010] = 1'b0;  wr_cycle[ 1010] = 1'b1;  addr_rom[ 1010]='h00000738;  wr_data_rom[ 1010]='h00000e4a;
    rd_cycle[ 1011] = 1'b0;  wr_cycle[ 1011] = 1'b1;  addr_rom[ 1011]='h0000099c;  wr_data_rom[ 1011]='h00000a1c;
    rd_cycle[ 1012] = 1'b1;  wr_cycle[ 1012] = 1'b0;  addr_rom[ 1012]='h00000d14;  wr_data_rom[ 1012]='h00000000;
    rd_cycle[ 1013] = 1'b1;  wr_cycle[ 1013] = 1'b0;  addr_rom[ 1013]='h00000968;  wr_data_rom[ 1013]='h00000000;
    rd_cycle[ 1014] = 1'b0;  wr_cycle[ 1014] = 1'b1;  addr_rom[ 1014]='h000008dc;  wr_data_rom[ 1014]='h00000a0a;
    rd_cycle[ 1015] = 1'b1;  wr_cycle[ 1015] = 1'b0;  addr_rom[ 1015]='h00000c3c;  wr_data_rom[ 1015]='h00000000;
    rd_cycle[ 1016] = 1'b0;  wr_cycle[ 1016] = 1'b1;  addr_rom[ 1016]='h00000714;  wr_data_rom[ 1016]='h00000932;
    rd_cycle[ 1017] = 1'b0;  wr_cycle[ 1017] = 1'b1;  addr_rom[ 1017]='h00000a70;  wr_data_rom[ 1017]='h00000e55;
    rd_cycle[ 1018] = 1'b0;  wr_cycle[ 1018] = 1'b1;  addr_rom[ 1018]='h00000a18;  wr_data_rom[ 1018]='h00000755;
    rd_cycle[ 1019] = 1'b0;  wr_cycle[ 1019] = 1'b1;  addr_rom[ 1019]='h00000914;  wr_data_rom[ 1019]='h00000b3c;
    rd_cycle[ 1020] = 1'b0;  wr_cycle[ 1020] = 1'b1;  addr_rom[ 1020]='h00000788;  wr_data_rom[ 1020]='h00000040;
    rd_cycle[ 1021] = 1'b1;  wr_cycle[ 1021] = 1'b0;  addr_rom[ 1021]='h00000ac0;  wr_data_rom[ 1021]='h00000000;
    rd_cycle[ 1022] = 1'b1;  wr_cycle[ 1022] = 1'b0;  addr_rom[ 1022]='h000002ac;  wr_data_rom[ 1022]='h00000000;
    rd_cycle[ 1023] = 1'b1;  wr_cycle[ 1023] = 1'b0;  addr_rom[ 1023]='h00000420;  wr_data_rom[ 1023]='h00000000;
    rd_cycle[ 1024] = 1'b0;  wr_cycle[ 1024] = 1'b1;  addr_rom[ 1024]='h00000074;  wr_data_rom[ 1024]='h000001c8;
    rd_cycle[ 1025] = 1'b0;  wr_cycle[ 1025] = 1'b1;  addr_rom[ 1025]='h0000015c;  wr_data_rom[ 1025]='h0000031d;
    rd_cycle[ 1026] = 1'b0;  wr_cycle[ 1026] = 1'b1;  addr_rom[ 1026]='h0000027c;  wr_data_rom[ 1026]='h000001f3;
    rd_cycle[ 1027] = 1'b0;  wr_cycle[ 1027] = 1'b1;  addr_rom[ 1027]='h00000cdc;  wr_data_rom[ 1027]='h00000c96;
    rd_cycle[ 1028] = 1'b0;  wr_cycle[ 1028] = 1'b1;  addr_rom[ 1028]='h0000078c;  wr_data_rom[ 1028]='h00000607;
    rd_cycle[ 1029] = 1'b0;  wr_cycle[ 1029] = 1'b1;  addr_rom[ 1029]='h000005c4;  wr_data_rom[ 1029]='h00000128;
    rd_cycle[ 1030] = 1'b0;  wr_cycle[ 1030] = 1'b1;  addr_rom[ 1030]='h00000558;  wr_data_rom[ 1030]='h00000404;
    rd_cycle[ 1031] = 1'b1;  wr_cycle[ 1031] = 1'b0;  addr_rom[ 1031]='h000009a8;  wr_data_rom[ 1031]='h00000000;
    rd_cycle[ 1032] = 1'b1;  wr_cycle[ 1032] = 1'b0;  addr_rom[ 1032]='h00000838;  wr_data_rom[ 1032]='h00000000;
    rd_cycle[ 1033] = 1'b1;  wr_cycle[ 1033] = 1'b0;  addr_rom[ 1033]='h00000c4c;  wr_data_rom[ 1033]='h00000000;
    rd_cycle[ 1034] = 1'b1;  wr_cycle[ 1034] = 1'b0;  addr_rom[ 1034]='h00000360;  wr_data_rom[ 1034]='h00000000;
    rd_cycle[ 1035] = 1'b1;  wr_cycle[ 1035] = 1'b0;  addr_rom[ 1035]='h000006c0;  wr_data_rom[ 1035]='h00000000;
    rd_cycle[ 1036] = 1'b0;  wr_cycle[ 1036] = 1'b1;  addr_rom[ 1036]='h00000364;  wr_data_rom[ 1036]='h00000e56;
    rd_cycle[ 1037] = 1'b0;  wr_cycle[ 1037] = 1'b1;  addr_rom[ 1037]='h00000934;  wr_data_rom[ 1037]='h00000d5b;
    rd_cycle[ 1038] = 1'b1;  wr_cycle[ 1038] = 1'b0;  addr_rom[ 1038]='h00000658;  wr_data_rom[ 1038]='h00000000;
    rd_cycle[ 1039] = 1'b1;  wr_cycle[ 1039] = 1'b0;  addr_rom[ 1039]='h000009f8;  wr_data_rom[ 1039]='h00000000;
    rd_cycle[ 1040] = 1'b1;  wr_cycle[ 1040] = 1'b0;  addr_rom[ 1040]='h00000b9c;  wr_data_rom[ 1040]='h00000000;
    rd_cycle[ 1041] = 1'b1;  wr_cycle[ 1041] = 1'b0;  addr_rom[ 1041]='h00000f54;  wr_data_rom[ 1041]='h00000000;
    rd_cycle[ 1042] = 1'b0;  wr_cycle[ 1042] = 1'b1;  addr_rom[ 1042]='h00000f90;  wr_data_rom[ 1042]='h0000076f;
    rd_cycle[ 1043] = 1'b1;  wr_cycle[ 1043] = 1'b0;  addr_rom[ 1043]='h0000082c;  wr_data_rom[ 1043]='h00000000;
    rd_cycle[ 1044] = 1'b1;  wr_cycle[ 1044] = 1'b0;  addr_rom[ 1044]='h00000244;  wr_data_rom[ 1044]='h00000000;
    rd_cycle[ 1045] = 1'b1;  wr_cycle[ 1045] = 1'b0;  addr_rom[ 1045]='h00000424;  wr_data_rom[ 1045]='h00000000;
    rd_cycle[ 1046] = 1'b0;  wr_cycle[ 1046] = 1'b1;  addr_rom[ 1046]='h00000afc;  wr_data_rom[ 1046]='h00000e67;
    rd_cycle[ 1047] = 1'b1;  wr_cycle[ 1047] = 1'b0;  addr_rom[ 1047]='h00000e54;  wr_data_rom[ 1047]='h00000000;
    rd_cycle[ 1048] = 1'b1;  wr_cycle[ 1048] = 1'b0;  addr_rom[ 1048]='h00000a58;  wr_data_rom[ 1048]='h00000000;
    rd_cycle[ 1049] = 1'b1;  wr_cycle[ 1049] = 1'b0;  addr_rom[ 1049]='h000008d8;  wr_data_rom[ 1049]='h00000000;
    rd_cycle[ 1050] = 1'b0;  wr_cycle[ 1050] = 1'b1;  addr_rom[ 1050]='h000003e0;  wr_data_rom[ 1050]='h00000467;
    rd_cycle[ 1051] = 1'b1;  wr_cycle[ 1051] = 1'b0;  addr_rom[ 1051]='h00000028;  wr_data_rom[ 1051]='h00000000;
    rd_cycle[ 1052] = 1'b1;  wr_cycle[ 1052] = 1'b0;  addr_rom[ 1052]='h00000980;  wr_data_rom[ 1052]='h00000000;
    rd_cycle[ 1053] = 1'b1;  wr_cycle[ 1053] = 1'b0;  addr_rom[ 1053]='h00000a38;  wr_data_rom[ 1053]='h00000000;
    rd_cycle[ 1054] = 1'b1;  wr_cycle[ 1054] = 1'b0;  addr_rom[ 1054]='h00000258;  wr_data_rom[ 1054]='h00000000;
    rd_cycle[ 1055] = 1'b1;  wr_cycle[ 1055] = 1'b0;  addr_rom[ 1055]='h00000b80;  wr_data_rom[ 1055]='h00000000;
    rd_cycle[ 1056] = 1'b1;  wr_cycle[ 1056] = 1'b0;  addr_rom[ 1056]='h00000688;  wr_data_rom[ 1056]='h00000000;
    rd_cycle[ 1057] = 1'b0;  wr_cycle[ 1057] = 1'b1;  addr_rom[ 1057]='h0000090c;  wr_data_rom[ 1057]='h000009a8;
    rd_cycle[ 1058] = 1'b0;  wr_cycle[ 1058] = 1'b1;  addr_rom[ 1058]='h00000104;  wr_data_rom[ 1058]='h00000818;
    rd_cycle[ 1059] = 1'b0;  wr_cycle[ 1059] = 1'b1;  addr_rom[ 1059]='h0000027c;  wr_data_rom[ 1059]='h00000d14;
    rd_cycle[ 1060] = 1'b0;  wr_cycle[ 1060] = 1'b1;  addr_rom[ 1060]='h000000a8;  wr_data_rom[ 1060]='h00000982;
    rd_cycle[ 1061] = 1'b1;  wr_cycle[ 1061] = 1'b0;  addr_rom[ 1061]='h00000f20;  wr_data_rom[ 1061]='h00000000;
    rd_cycle[ 1062] = 1'b0;  wr_cycle[ 1062] = 1'b1;  addr_rom[ 1062]='h00000f58;  wr_data_rom[ 1062]='h00000b07;
    rd_cycle[ 1063] = 1'b0;  wr_cycle[ 1063] = 1'b1;  addr_rom[ 1063]='h00000400;  wr_data_rom[ 1063]='h0000012e;
    rd_cycle[ 1064] = 1'b0;  wr_cycle[ 1064] = 1'b1;  addr_rom[ 1064]='h00000cb8;  wr_data_rom[ 1064]='h00000af5;
    rd_cycle[ 1065] = 1'b0;  wr_cycle[ 1065] = 1'b1;  addr_rom[ 1065]='h00000d48;  wr_data_rom[ 1065]='h0000062c;
    rd_cycle[ 1066] = 1'b1;  wr_cycle[ 1066] = 1'b0;  addr_rom[ 1066]='h000002cc;  wr_data_rom[ 1066]='h00000000;
    rd_cycle[ 1067] = 1'b0;  wr_cycle[ 1067] = 1'b1;  addr_rom[ 1067]='h00000800;  wr_data_rom[ 1067]='h000005a3;
    rd_cycle[ 1068] = 1'b0;  wr_cycle[ 1068] = 1'b1;  addr_rom[ 1068]='h000008d0;  wr_data_rom[ 1068]='h00000664;
    rd_cycle[ 1069] = 1'b1;  wr_cycle[ 1069] = 1'b0;  addr_rom[ 1069]='h0000006c;  wr_data_rom[ 1069]='h00000000;
    rd_cycle[ 1070] = 1'b1;  wr_cycle[ 1070] = 1'b0;  addr_rom[ 1070]='h00000390;  wr_data_rom[ 1070]='h00000000;
    rd_cycle[ 1071] = 1'b1;  wr_cycle[ 1071] = 1'b0;  addr_rom[ 1071]='h00000554;  wr_data_rom[ 1071]='h00000000;
    rd_cycle[ 1072] = 1'b1;  wr_cycle[ 1072] = 1'b0;  addr_rom[ 1072]='h000004c8;  wr_data_rom[ 1072]='h00000000;
    rd_cycle[ 1073] = 1'b1;  wr_cycle[ 1073] = 1'b0;  addr_rom[ 1073]='h000003c8;  wr_data_rom[ 1073]='h00000000;
    rd_cycle[ 1074] = 1'b0;  wr_cycle[ 1074] = 1'b1;  addr_rom[ 1074]='h00000edc;  wr_data_rom[ 1074]='h000005f3;
    rd_cycle[ 1075] = 1'b1;  wr_cycle[ 1075] = 1'b0;  addr_rom[ 1075]='h00000e74;  wr_data_rom[ 1075]='h00000000;
    rd_cycle[ 1076] = 1'b1;  wr_cycle[ 1076] = 1'b0;  addr_rom[ 1076]='h00000d28;  wr_data_rom[ 1076]='h00000000;
    rd_cycle[ 1077] = 1'b1;  wr_cycle[ 1077] = 1'b0;  addr_rom[ 1077]='h00000b4c;  wr_data_rom[ 1077]='h00000000;
    rd_cycle[ 1078] = 1'b1;  wr_cycle[ 1078] = 1'b0;  addr_rom[ 1078]='h00000738;  wr_data_rom[ 1078]='h00000000;
    rd_cycle[ 1079] = 1'b1;  wr_cycle[ 1079] = 1'b0;  addr_rom[ 1079]='h00000760;  wr_data_rom[ 1079]='h00000000;
    rd_cycle[ 1080] = 1'b0;  wr_cycle[ 1080] = 1'b1;  addr_rom[ 1080]='h00000a98;  wr_data_rom[ 1080]='h00000bcd;
    rd_cycle[ 1081] = 1'b1;  wr_cycle[ 1081] = 1'b0;  addr_rom[ 1081]='h00000f34;  wr_data_rom[ 1081]='h00000000;
    rd_cycle[ 1082] = 1'b1;  wr_cycle[ 1082] = 1'b0;  addr_rom[ 1082]='h00000f58;  wr_data_rom[ 1082]='h00000000;
    rd_cycle[ 1083] = 1'b0;  wr_cycle[ 1083] = 1'b1;  addr_rom[ 1083]='h00000dfc;  wr_data_rom[ 1083]='h00000623;
    rd_cycle[ 1084] = 1'b1;  wr_cycle[ 1084] = 1'b0;  addr_rom[ 1084]='h0000015c;  wr_data_rom[ 1084]='h00000000;
    rd_cycle[ 1085] = 1'b1;  wr_cycle[ 1085] = 1'b0;  addr_rom[ 1085]='h00000da0;  wr_data_rom[ 1085]='h00000000;
    rd_cycle[ 1086] = 1'b1;  wr_cycle[ 1086] = 1'b0;  addr_rom[ 1086]='h00000180;  wr_data_rom[ 1086]='h00000000;
    rd_cycle[ 1087] = 1'b0;  wr_cycle[ 1087] = 1'b1;  addr_rom[ 1087]='h00000d34;  wr_data_rom[ 1087]='h000001f5;
    rd_cycle[ 1088] = 1'b0;  wr_cycle[ 1088] = 1'b1;  addr_rom[ 1088]='h00000e38;  wr_data_rom[ 1088]='h00000512;
    rd_cycle[ 1089] = 1'b1;  wr_cycle[ 1089] = 1'b0;  addr_rom[ 1089]='h00000f28;  wr_data_rom[ 1089]='h00000000;
    rd_cycle[ 1090] = 1'b0;  wr_cycle[ 1090] = 1'b1;  addr_rom[ 1090]='h00000028;  wr_data_rom[ 1090]='h00000617;
    rd_cycle[ 1091] = 1'b0;  wr_cycle[ 1091] = 1'b1;  addr_rom[ 1091]='h0000065c;  wr_data_rom[ 1091]='h00000f13;
    rd_cycle[ 1092] = 1'b0;  wr_cycle[ 1092] = 1'b1;  addr_rom[ 1092]='h000006f8;  wr_data_rom[ 1092]='h0000043f;
    rd_cycle[ 1093] = 1'b1;  wr_cycle[ 1093] = 1'b0;  addr_rom[ 1093]='h000001b4;  wr_data_rom[ 1093]='h00000000;
    rd_cycle[ 1094] = 1'b0;  wr_cycle[ 1094] = 1'b1;  addr_rom[ 1094]='h00000be0;  wr_data_rom[ 1094]='h00000ae8;
    rd_cycle[ 1095] = 1'b0;  wr_cycle[ 1095] = 1'b1;  addr_rom[ 1095]='h00000ac4;  wr_data_rom[ 1095]='h000008a9;
    rd_cycle[ 1096] = 1'b0;  wr_cycle[ 1096] = 1'b1;  addr_rom[ 1096]='h00000758;  wr_data_rom[ 1096]='h000002cd;
    rd_cycle[ 1097] = 1'b0;  wr_cycle[ 1097] = 1'b1;  addr_rom[ 1097]='h00000970;  wr_data_rom[ 1097]='h0000052c;
    rd_cycle[ 1098] = 1'b0;  wr_cycle[ 1098] = 1'b1;  addr_rom[ 1098]='h000007ac;  wr_data_rom[ 1098]='h00000226;
    rd_cycle[ 1099] = 1'b0;  wr_cycle[ 1099] = 1'b1;  addr_rom[ 1099]='h00000274;  wr_data_rom[ 1099]='h000001cb;
    rd_cycle[ 1100] = 1'b1;  wr_cycle[ 1100] = 1'b0;  addr_rom[ 1100]='h00000160;  wr_data_rom[ 1100]='h00000000;
    rd_cycle[ 1101] = 1'b0;  wr_cycle[ 1101] = 1'b1;  addr_rom[ 1101]='h00000f9c;  wr_data_rom[ 1101]='h00000cf3;
    rd_cycle[ 1102] = 1'b0;  wr_cycle[ 1102] = 1'b1;  addr_rom[ 1102]='h000005a4;  wr_data_rom[ 1102]='h000001bc;
    rd_cycle[ 1103] = 1'b0;  wr_cycle[ 1103] = 1'b1;  addr_rom[ 1103]='h000004c8;  wr_data_rom[ 1103]='h0000009a;
    rd_cycle[ 1104] = 1'b0;  wr_cycle[ 1104] = 1'b1;  addr_rom[ 1104]='h00000e78;  wr_data_rom[ 1104]='h00000b36;
    rd_cycle[ 1105] = 1'b1;  wr_cycle[ 1105] = 1'b0;  addr_rom[ 1105]='h00000300;  wr_data_rom[ 1105]='h00000000;
    rd_cycle[ 1106] = 1'b0;  wr_cycle[ 1106] = 1'b1;  addr_rom[ 1106]='h00000eb4;  wr_data_rom[ 1106]='h000009be;
    rd_cycle[ 1107] = 1'b1;  wr_cycle[ 1107] = 1'b0;  addr_rom[ 1107]='h000000f0;  wr_data_rom[ 1107]='h00000000;
    rd_cycle[ 1108] = 1'b0;  wr_cycle[ 1108] = 1'b1;  addr_rom[ 1108]='h000003c8;  wr_data_rom[ 1108]='h0000045e;
    rd_cycle[ 1109] = 1'b0;  wr_cycle[ 1109] = 1'b1;  addr_rom[ 1109]='h0000096c;  wr_data_rom[ 1109]='h0000087d;
    rd_cycle[ 1110] = 1'b0;  wr_cycle[ 1110] = 1'b1;  addr_rom[ 1110]='h00000f40;  wr_data_rom[ 1110]='h00000cd7;
    rd_cycle[ 1111] = 1'b1;  wr_cycle[ 1111] = 1'b0;  addr_rom[ 1111]='h00000cd0;  wr_data_rom[ 1111]='h00000000;
    rd_cycle[ 1112] = 1'b0;  wr_cycle[ 1112] = 1'b1;  addr_rom[ 1112]='h00000960;  wr_data_rom[ 1112]='h00000ebf;
    rd_cycle[ 1113] = 1'b1;  wr_cycle[ 1113] = 1'b0;  addr_rom[ 1113]='h000007f4;  wr_data_rom[ 1113]='h00000000;
    rd_cycle[ 1114] = 1'b1;  wr_cycle[ 1114] = 1'b0;  addr_rom[ 1114]='h00000bd8;  wr_data_rom[ 1114]='h00000000;
    rd_cycle[ 1115] = 1'b1;  wr_cycle[ 1115] = 1'b0;  addr_rom[ 1115]='h00000c88;  wr_data_rom[ 1115]='h00000000;
    rd_cycle[ 1116] = 1'b1;  wr_cycle[ 1116] = 1'b0;  addr_rom[ 1116]='h000004a8;  wr_data_rom[ 1116]='h00000000;
    rd_cycle[ 1117] = 1'b1;  wr_cycle[ 1117] = 1'b0;  addr_rom[ 1117]='h00000884;  wr_data_rom[ 1117]='h00000000;
    rd_cycle[ 1118] = 1'b0;  wr_cycle[ 1118] = 1'b1;  addr_rom[ 1118]='h000004fc;  wr_data_rom[ 1118]='h000007e8;
    rd_cycle[ 1119] = 1'b1;  wr_cycle[ 1119] = 1'b0;  addr_rom[ 1119]='h00000d74;  wr_data_rom[ 1119]='h00000000;
    rd_cycle[ 1120] = 1'b1;  wr_cycle[ 1120] = 1'b0;  addr_rom[ 1120]='h00000c00;  wr_data_rom[ 1120]='h00000000;
    rd_cycle[ 1121] = 1'b0;  wr_cycle[ 1121] = 1'b1;  addr_rom[ 1121]='h00000cbc;  wr_data_rom[ 1121]='h00000878;
    rd_cycle[ 1122] = 1'b1;  wr_cycle[ 1122] = 1'b0;  addr_rom[ 1122]='h00000148;  wr_data_rom[ 1122]='h00000000;
    rd_cycle[ 1123] = 1'b1;  wr_cycle[ 1123] = 1'b0;  addr_rom[ 1123]='h0000063c;  wr_data_rom[ 1123]='h00000000;
    rd_cycle[ 1124] = 1'b0;  wr_cycle[ 1124] = 1'b1;  addr_rom[ 1124]='h000007d4;  wr_data_rom[ 1124]='h00000216;
    rd_cycle[ 1125] = 1'b0;  wr_cycle[ 1125] = 1'b1;  addr_rom[ 1125]='h00000b9c;  wr_data_rom[ 1125]='h00000d35;
    rd_cycle[ 1126] = 1'b1;  wr_cycle[ 1126] = 1'b0;  addr_rom[ 1126]='h00000e7c;  wr_data_rom[ 1126]='h00000000;
    rd_cycle[ 1127] = 1'b0;  wr_cycle[ 1127] = 1'b1;  addr_rom[ 1127]='h00000264;  wr_data_rom[ 1127]='h0000037c;
    rd_cycle[ 1128] = 1'b1;  wr_cycle[ 1128] = 1'b0;  addr_rom[ 1128]='h00000bf4;  wr_data_rom[ 1128]='h00000000;
    rd_cycle[ 1129] = 1'b1;  wr_cycle[ 1129] = 1'b0;  addr_rom[ 1129]='h00000994;  wr_data_rom[ 1129]='h00000000;
    rd_cycle[ 1130] = 1'b1;  wr_cycle[ 1130] = 1'b0;  addr_rom[ 1130]='h00000f84;  wr_data_rom[ 1130]='h00000000;
    rd_cycle[ 1131] = 1'b0;  wr_cycle[ 1131] = 1'b1;  addr_rom[ 1131]='h000003ac;  wr_data_rom[ 1131]='h000002ac;
    rd_cycle[ 1132] = 1'b1;  wr_cycle[ 1132] = 1'b0;  addr_rom[ 1132]='h000005f8;  wr_data_rom[ 1132]='h00000000;
    rd_cycle[ 1133] = 1'b0;  wr_cycle[ 1133] = 1'b1;  addr_rom[ 1133]='h00000668;  wr_data_rom[ 1133]='h0000053f;
    rd_cycle[ 1134] = 1'b0;  wr_cycle[ 1134] = 1'b1;  addr_rom[ 1134]='h00000ed8;  wr_data_rom[ 1134]='h000008bd;
    rd_cycle[ 1135] = 1'b0;  wr_cycle[ 1135] = 1'b1;  addr_rom[ 1135]='h000005d8;  wr_data_rom[ 1135]='h00000706;
    rd_cycle[ 1136] = 1'b0;  wr_cycle[ 1136] = 1'b1;  addr_rom[ 1136]='h00000100;  wr_data_rom[ 1136]='h00000be7;
    rd_cycle[ 1137] = 1'b0;  wr_cycle[ 1137] = 1'b1;  addr_rom[ 1137]='h00000648;  wr_data_rom[ 1137]='h0000002d;
    rd_cycle[ 1138] = 1'b1;  wr_cycle[ 1138] = 1'b0;  addr_rom[ 1138]='h00000a48;  wr_data_rom[ 1138]='h00000000;
    rd_cycle[ 1139] = 1'b0;  wr_cycle[ 1139] = 1'b1;  addr_rom[ 1139]='h000009a4;  wr_data_rom[ 1139]='h00000565;
    rd_cycle[ 1140] = 1'b0;  wr_cycle[ 1140] = 1'b1;  addr_rom[ 1140]='h000002bc;  wr_data_rom[ 1140]='h00000530;
    rd_cycle[ 1141] = 1'b1;  wr_cycle[ 1141] = 1'b0;  addr_rom[ 1141]='h000007e4;  wr_data_rom[ 1141]='h00000000;
    rd_cycle[ 1142] = 1'b0;  wr_cycle[ 1142] = 1'b1;  addr_rom[ 1142]='h00000488;  wr_data_rom[ 1142]='h000002f2;
    rd_cycle[ 1143] = 1'b1;  wr_cycle[ 1143] = 1'b0;  addr_rom[ 1143]='h00000598;  wr_data_rom[ 1143]='h00000000;
    rd_cycle[ 1144] = 1'b1;  wr_cycle[ 1144] = 1'b0;  addr_rom[ 1144]='h00000a98;  wr_data_rom[ 1144]='h00000000;
    rd_cycle[ 1145] = 1'b0;  wr_cycle[ 1145] = 1'b1;  addr_rom[ 1145]='h00000b68;  wr_data_rom[ 1145]='h000009e8;
    rd_cycle[ 1146] = 1'b0;  wr_cycle[ 1146] = 1'b1;  addr_rom[ 1146]='h00000498;  wr_data_rom[ 1146]='h00000627;
    rd_cycle[ 1147] = 1'b1;  wr_cycle[ 1147] = 1'b0;  addr_rom[ 1147]='h00000f90;  wr_data_rom[ 1147]='h00000000;
    rd_cycle[ 1148] = 1'b0;  wr_cycle[ 1148] = 1'b1;  addr_rom[ 1148]='h00000d48;  wr_data_rom[ 1148]='h00000ea0;
    rd_cycle[ 1149] = 1'b0;  wr_cycle[ 1149] = 1'b1;  addr_rom[ 1149]='h0000045c;  wr_data_rom[ 1149]='h00000135;
    rd_cycle[ 1150] = 1'b1;  wr_cycle[ 1150] = 1'b0;  addr_rom[ 1150]='h000009e4;  wr_data_rom[ 1150]='h00000000;
    rd_cycle[ 1151] = 1'b1;  wr_cycle[ 1151] = 1'b0;  addr_rom[ 1151]='h000001f4;  wr_data_rom[ 1151]='h00000000;
    rd_cycle[ 1152] = 1'b0;  wr_cycle[ 1152] = 1'b1;  addr_rom[ 1152]='h00000f98;  wr_data_rom[ 1152]='h00000ad7;
    rd_cycle[ 1153] = 1'b0;  wr_cycle[ 1153] = 1'b1;  addr_rom[ 1153]='h00000418;  wr_data_rom[ 1153]='h00000d25;
    rd_cycle[ 1154] = 1'b1;  wr_cycle[ 1154] = 1'b0;  addr_rom[ 1154]='h00000f54;  wr_data_rom[ 1154]='h00000000;
    rd_cycle[ 1155] = 1'b0;  wr_cycle[ 1155] = 1'b1;  addr_rom[ 1155]='h00000b6c;  wr_data_rom[ 1155]='h000008e2;
    rd_cycle[ 1156] = 1'b1;  wr_cycle[ 1156] = 1'b0;  addr_rom[ 1156]='h000003d8;  wr_data_rom[ 1156]='h00000000;
    rd_cycle[ 1157] = 1'b1;  wr_cycle[ 1157] = 1'b0;  addr_rom[ 1157]='h000001b8;  wr_data_rom[ 1157]='h00000000;
    rd_cycle[ 1158] = 1'b1;  wr_cycle[ 1158] = 1'b0;  addr_rom[ 1158]='h000007a8;  wr_data_rom[ 1158]='h00000000;
    rd_cycle[ 1159] = 1'b1;  wr_cycle[ 1159] = 1'b0;  addr_rom[ 1159]='h00000e2c;  wr_data_rom[ 1159]='h00000000;
    rd_cycle[ 1160] = 1'b0;  wr_cycle[ 1160] = 1'b1;  addr_rom[ 1160]='h0000062c;  wr_data_rom[ 1160]='h000007df;
    rd_cycle[ 1161] = 1'b1;  wr_cycle[ 1161] = 1'b0;  addr_rom[ 1161]='h000009b8;  wr_data_rom[ 1161]='h00000000;
    rd_cycle[ 1162] = 1'b1;  wr_cycle[ 1162] = 1'b0;  addr_rom[ 1162]='h00000d8c;  wr_data_rom[ 1162]='h00000000;
    rd_cycle[ 1163] = 1'b0;  wr_cycle[ 1163] = 1'b1;  addr_rom[ 1163]='h00000748;  wr_data_rom[ 1163]='h000003e0;
    rd_cycle[ 1164] = 1'b1;  wr_cycle[ 1164] = 1'b0;  addr_rom[ 1164]='h00000d88;  wr_data_rom[ 1164]='h00000000;
    rd_cycle[ 1165] = 1'b1;  wr_cycle[ 1165] = 1'b0;  addr_rom[ 1165]='h00000d30;  wr_data_rom[ 1165]='h00000000;
    rd_cycle[ 1166] = 1'b1;  wr_cycle[ 1166] = 1'b0;  addr_rom[ 1166]='h000009cc;  wr_data_rom[ 1166]='h00000000;
    rd_cycle[ 1167] = 1'b1;  wr_cycle[ 1167] = 1'b0;  addr_rom[ 1167]='h000003b4;  wr_data_rom[ 1167]='h00000000;
    rd_cycle[ 1168] = 1'b1;  wr_cycle[ 1168] = 1'b0;  addr_rom[ 1168]='h000003c0;  wr_data_rom[ 1168]='h00000000;
    rd_cycle[ 1169] = 1'b1;  wr_cycle[ 1169] = 1'b0;  addr_rom[ 1169]='h00000848;  wr_data_rom[ 1169]='h00000000;
    rd_cycle[ 1170] = 1'b1;  wr_cycle[ 1170] = 1'b0;  addr_rom[ 1170]='h000006dc;  wr_data_rom[ 1170]='h00000000;
    rd_cycle[ 1171] = 1'b1;  wr_cycle[ 1171] = 1'b0;  addr_rom[ 1171]='h000004e4;  wr_data_rom[ 1171]='h00000000;
    rd_cycle[ 1172] = 1'b0;  wr_cycle[ 1172] = 1'b1;  addr_rom[ 1172]='h00000088;  wr_data_rom[ 1172]='h00000d41;
    rd_cycle[ 1173] = 1'b0;  wr_cycle[ 1173] = 1'b1;  addr_rom[ 1173]='h000008b0;  wr_data_rom[ 1173]='h00000281;
    rd_cycle[ 1174] = 1'b1;  wr_cycle[ 1174] = 1'b0;  addr_rom[ 1174]='h00000e94;  wr_data_rom[ 1174]='h00000000;
    rd_cycle[ 1175] = 1'b1;  wr_cycle[ 1175] = 1'b0;  addr_rom[ 1175]='h00000ef8;  wr_data_rom[ 1175]='h00000000;
    rd_cycle[ 1176] = 1'b0;  wr_cycle[ 1176] = 1'b1;  addr_rom[ 1176]='h00000f1c;  wr_data_rom[ 1176]='h00000236;
    rd_cycle[ 1177] = 1'b1;  wr_cycle[ 1177] = 1'b0;  addr_rom[ 1177]='h000003f0;  wr_data_rom[ 1177]='h00000000;
    rd_cycle[ 1178] = 1'b1;  wr_cycle[ 1178] = 1'b0;  addr_rom[ 1178]='h00000b2c;  wr_data_rom[ 1178]='h00000000;
    rd_cycle[ 1179] = 1'b0;  wr_cycle[ 1179] = 1'b1;  addr_rom[ 1179]='h000005b0;  wr_data_rom[ 1179]='h00000753;
    rd_cycle[ 1180] = 1'b1;  wr_cycle[ 1180] = 1'b0;  addr_rom[ 1180]='h000006ac;  wr_data_rom[ 1180]='h00000000;
    rd_cycle[ 1181] = 1'b1;  wr_cycle[ 1181] = 1'b0;  addr_rom[ 1181]='h00000bac;  wr_data_rom[ 1181]='h00000000;
    rd_cycle[ 1182] = 1'b1;  wr_cycle[ 1182] = 1'b0;  addr_rom[ 1182]='h00000918;  wr_data_rom[ 1182]='h00000000;
    rd_cycle[ 1183] = 1'b0;  wr_cycle[ 1183] = 1'b1;  addr_rom[ 1183]='h00000450;  wr_data_rom[ 1183]='h00000f31;
    rd_cycle[ 1184] = 1'b0;  wr_cycle[ 1184] = 1'b1;  addr_rom[ 1184]='h00000cc4;  wr_data_rom[ 1184]='h00000ed4;
    rd_cycle[ 1185] = 1'b0;  wr_cycle[ 1185] = 1'b1;  addr_rom[ 1185]='h00000794;  wr_data_rom[ 1185]='h0000015a;
    rd_cycle[ 1186] = 1'b1;  wr_cycle[ 1186] = 1'b0;  addr_rom[ 1186]='h00000674;  wr_data_rom[ 1186]='h00000000;
    rd_cycle[ 1187] = 1'b1;  wr_cycle[ 1187] = 1'b0;  addr_rom[ 1187]='h00000bc8;  wr_data_rom[ 1187]='h00000000;
    rd_cycle[ 1188] = 1'b1;  wr_cycle[ 1188] = 1'b0;  addr_rom[ 1188]='h00000f5c;  wr_data_rom[ 1188]='h00000000;
    rd_cycle[ 1189] = 1'b1;  wr_cycle[ 1189] = 1'b0;  addr_rom[ 1189]='h00000bac;  wr_data_rom[ 1189]='h00000000;
    rd_cycle[ 1190] = 1'b0;  wr_cycle[ 1190] = 1'b1;  addr_rom[ 1190]='h000001e8;  wr_data_rom[ 1190]='h0000045f;
    rd_cycle[ 1191] = 1'b0;  wr_cycle[ 1191] = 1'b1;  addr_rom[ 1191]='h0000018c;  wr_data_rom[ 1191]='h000003d7;
    rd_cycle[ 1192] = 1'b0;  wr_cycle[ 1192] = 1'b1;  addr_rom[ 1192]='h00000040;  wr_data_rom[ 1192]='h00000081;
    rd_cycle[ 1193] = 1'b0;  wr_cycle[ 1193] = 1'b1;  addr_rom[ 1193]='h000004b4;  wr_data_rom[ 1193]='h00000457;
    rd_cycle[ 1194] = 1'b1;  wr_cycle[ 1194] = 1'b0;  addr_rom[ 1194]='h00000474;  wr_data_rom[ 1194]='h00000000;
    rd_cycle[ 1195] = 1'b0;  wr_cycle[ 1195] = 1'b1;  addr_rom[ 1195]='h00000418;  wr_data_rom[ 1195]='h00000ce3;
    rd_cycle[ 1196] = 1'b0;  wr_cycle[ 1196] = 1'b1;  addr_rom[ 1196]='h00000cf4;  wr_data_rom[ 1196]='h0000068a;
    rd_cycle[ 1197] = 1'b0;  wr_cycle[ 1197] = 1'b1;  addr_rom[ 1197]='h0000063c;  wr_data_rom[ 1197]='h000000a6;
    rd_cycle[ 1198] = 1'b1;  wr_cycle[ 1198] = 1'b0;  addr_rom[ 1198]='h00000ab8;  wr_data_rom[ 1198]='h00000000;
    rd_cycle[ 1199] = 1'b1;  wr_cycle[ 1199] = 1'b0;  addr_rom[ 1199]='h00000af4;  wr_data_rom[ 1199]='h00000000;
    rd_cycle[ 1200] = 1'b0;  wr_cycle[ 1200] = 1'b1;  addr_rom[ 1200]='h00000a14;  wr_data_rom[ 1200]='h00000a51;
    rd_cycle[ 1201] = 1'b1;  wr_cycle[ 1201] = 1'b0;  addr_rom[ 1201]='h00000220;  wr_data_rom[ 1201]='h00000000;
    rd_cycle[ 1202] = 1'b1;  wr_cycle[ 1202] = 1'b0;  addr_rom[ 1202]='h00000e84;  wr_data_rom[ 1202]='h00000000;
    rd_cycle[ 1203] = 1'b0;  wr_cycle[ 1203] = 1'b1;  addr_rom[ 1203]='h00000694;  wr_data_rom[ 1203]='h000005b7;
    rd_cycle[ 1204] = 1'b1;  wr_cycle[ 1204] = 1'b0;  addr_rom[ 1204]='h0000061c;  wr_data_rom[ 1204]='h00000000;
    rd_cycle[ 1205] = 1'b0;  wr_cycle[ 1205] = 1'b1;  addr_rom[ 1205]='h000002b0;  wr_data_rom[ 1205]='h000009d9;
    rd_cycle[ 1206] = 1'b1;  wr_cycle[ 1206] = 1'b0;  addr_rom[ 1206]='h00000a5c;  wr_data_rom[ 1206]='h00000000;
    rd_cycle[ 1207] = 1'b1;  wr_cycle[ 1207] = 1'b0;  addr_rom[ 1207]='h00000a70;  wr_data_rom[ 1207]='h00000000;
    rd_cycle[ 1208] = 1'b1;  wr_cycle[ 1208] = 1'b0;  addr_rom[ 1208]='h00000908;  wr_data_rom[ 1208]='h00000000;
    rd_cycle[ 1209] = 1'b1;  wr_cycle[ 1209] = 1'b0;  addr_rom[ 1209]='h000003f4;  wr_data_rom[ 1209]='h00000000;
    rd_cycle[ 1210] = 1'b1;  wr_cycle[ 1210] = 1'b0;  addr_rom[ 1210]='h00000ed8;  wr_data_rom[ 1210]='h00000000;
    rd_cycle[ 1211] = 1'b0;  wr_cycle[ 1211] = 1'b1;  addr_rom[ 1211]='h00000394;  wr_data_rom[ 1211]='h000007b2;
    rd_cycle[ 1212] = 1'b0;  wr_cycle[ 1212] = 1'b1;  addr_rom[ 1212]='h00000a0c;  wr_data_rom[ 1212]='h0000024f;
    rd_cycle[ 1213] = 1'b1;  wr_cycle[ 1213] = 1'b0;  addr_rom[ 1213]='h00000b5c;  wr_data_rom[ 1213]='h00000000;
    rd_cycle[ 1214] = 1'b0;  wr_cycle[ 1214] = 1'b1;  addr_rom[ 1214]='h000001dc;  wr_data_rom[ 1214]='h000005db;
    rd_cycle[ 1215] = 1'b1;  wr_cycle[ 1215] = 1'b0;  addr_rom[ 1215]='h00000218;  wr_data_rom[ 1215]='h00000000;
    rd_cycle[ 1216] = 1'b0;  wr_cycle[ 1216] = 1'b1;  addr_rom[ 1216]='h00000998;  wr_data_rom[ 1216]='h00000822;
    rd_cycle[ 1217] = 1'b0;  wr_cycle[ 1217] = 1'b1;  addr_rom[ 1217]='h00000bb4;  wr_data_rom[ 1217]='h00000ac3;
    rd_cycle[ 1218] = 1'b1;  wr_cycle[ 1218] = 1'b0;  addr_rom[ 1218]='h00000754;  wr_data_rom[ 1218]='h00000000;
    rd_cycle[ 1219] = 1'b1;  wr_cycle[ 1219] = 1'b0;  addr_rom[ 1219]='h00000d54;  wr_data_rom[ 1219]='h00000000;
    rd_cycle[ 1220] = 1'b1;  wr_cycle[ 1220] = 1'b0;  addr_rom[ 1220]='h0000073c;  wr_data_rom[ 1220]='h00000000;
    rd_cycle[ 1221] = 1'b1;  wr_cycle[ 1221] = 1'b0;  addr_rom[ 1221]='h000006d4;  wr_data_rom[ 1221]='h00000000;
    rd_cycle[ 1222] = 1'b0;  wr_cycle[ 1222] = 1'b1;  addr_rom[ 1222]='h00000b6c;  wr_data_rom[ 1222]='h000008e4;
    rd_cycle[ 1223] = 1'b1;  wr_cycle[ 1223] = 1'b0;  addr_rom[ 1223]='h00000310;  wr_data_rom[ 1223]='h00000000;
    rd_cycle[ 1224] = 1'b0;  wr_cycle[ 1224] = 1'b1;  addr_rom[ 1224]='h00000950;  wr_data_rom[ 1224]='h00000cc8;
    rd_cycle[ 1225] = 1'b1;  wr_cycle[ 1225] = 1'b0;  addr_rom[ 1225]='h000003f4;  wr_data_rom[ 1225]='h00000000;
    rd_cycle[ 1226] = 1'b1;  wr_cycle[ 1226] = 1'b0;  addr_rom[ 1226]='h00000120;  wr_data_rom[ 1226]='h00000000;
    rd_cycle[ 1227] = 1'b1;  wr_cycle[ 1227] = 1'b0;  addr_rom[ 1227]='h0000019c;  wr_data_rom[ 1227]='h00000000;
    rd_cycle[ 1228] = 1'b1;  wr_cycle[ 1228] = 1'b0;  addr_rom[ 1228]='h000002c4;  wr_data_rom[ 1228]='h00000000;
    rd_cycle[ 1229] = 1'b1;  wr_cycle[ 1229] = 1'b0;  addr_rom[ 1229]='h00000380;  wr_data_rom[ 1229]='h00000000;
    rd_cycle[ 1230] = 1'b0;  wr_cycle[ 1230] = 1'b1;  addr_rom[ 1230]='h000000f4;  wr_data_rom[ 1230]='h00000c76;
    rd_cycle[ 1231] = 1'b1;  wr_cycle[ 1231] = 1'b0;  addr_rom[ 1231]='h00000b4c;  wr_data_rom[ 1231]='h00000000;
    rd_cycle[ 1232] = 1'b1;  wr_cycle[ 1232] = 1'b0;  addr_rom[ 1232]='h00000348;  wr_data_rom[ 1232]='h00000000;
    rd_cycle[ 1233] = 1'b1;  wr_cycle[ 1233] = 1'b0;  addr_rom[ 1233]='h0000066c;  wr_data_rom[ 1233]='h00000000;
    rd_cycle[ 1234] = 1'b1;  wr_cycle[ 1234] = 1'b0;  addr_rom[ 1234]='h0000031c;  wr_data_rom[ 1234]='h00000000;
    rd_cycle[ 1235] = 1'b0;  wr_cycle[ 1235] = 1'b1;  addr_rom[ 1235]='h00000a58;  wr_data_rom[ 1235]='h00000bf1;
    rd_cycle[ 1236] = 1'b1;  wr_cycle[ 1236] = 1'b0;  addr_rom[ 1236]='h00000044;  wr_data_rom[ 1236]='h00000000;
    rd_cycle[ 1237] = 1'b1;  wr_cycle[ 1237] = 1'b0;  addr_rom[ 1237]='h00000e08;  wr_data_rom[ 1237]='h00000000;
    rd_cycle[ 1238] = 1'b1;  wr_cycle[ 1238] = 1'b0;  addr_rom[ 1238]='h0000023c;  wr_data_rom[ 1238]='h00000000;
    rd_cycle[ 1239] = 1'b1;  wr_cycle[ 1239] = 1'b0;  addr_rom[ 1239]='h00000e1c;  wr_data_rom[ 1239]='h00000000;
    rd_cycle[ 1240] = 1'b1;  wr_cycle[ 1240] = 1'b0;  addr_rom[ 1240]='h000000e0;  wr_data_rom[ 1240]='h00000000;
    rd_cycle[ 1241] = 1'b1;  wr_cycle[ 1241] = 1'b0;  addr_rom[ 1241]='h0000094c;  wr_data_rom[ 1241]='h00000000;
    rd_cycle[ 1242] = 1'b1;  wr_cycle[ 1242] = 1'b0;  addr_rom[ 1242]='h00000a64;  wr_data_rom[ 1242]='h00000000;
    rd_cycle[ 1243] = 1'b0;  wr_cycle[ 1243] = 1'b1;  addr_rom[ 1243]='h00000f40;  wr_data_rom[ 1243]='h00000078;
    rd_cycle[ 1244] = 1'b0;  wr_cycle[ 1244] = 1'b1;  addr_rom[ 1244]='h00000e68;  wr_data_rom[ 1244]='h00000e94;
    rd_cycle[ 1245] = 1'b1;  wr_cycle[ 1245] = 1'b0;  addr_rom[ 1245]='h000000c0;  wr_data_rom[ 1245]='h00000000;
    rd_cycle[ 1246] = 1'b0;  wr_cycle[ 1246] = 1'b1;  addr_rom[ 1246]='h00000b88;  wr_data_rom[ 1246]='h000003bc;
    rd_cycle[ 1247] = 1'b1;  wr_cycle[ 1247] = 1'b0;  addr_rom[ 1247]='h00000cf8;  wr_data_rom[ 1247]='h00000000;
    rd_cycle[ 1248] = 1'b1;  wr_cycle[ 1248] = 1'b0;  addr_rom[ 1248]='h00000310;  wr_data_rom[ 1248]='h00000000;
    rd_cycle[ 1249] = 1'b1;  wr_cycle[ 1249] = 1'b0;  addr_rom[ 1249]='h000000d4;  wr_data_rom[ 1249]='h00000000;
    rd_cycle[ 1250] = 1'b0;  wr_cycle[ 1250] = 1'b1;  addr_rom[ 1250]='h00000ac0;  wr_data_rom[ 1250]='h000006ea;
    rd_cycle[ 1251] = 1'b1;  wr_cycle[ 1251] = 1'b0;  addr_rom[ 1251]='h00000550;  wr_data_rom[ 1251]='h00000000;
    rd_cycle[ 1252] = 1'b1;  wr_cycle[ 1252] = 1'b0;  addr_rom[ 1252]='h000009b0;  wr_data_rom[ 1252]='h00000000;
    rd_cycle[ 1253] = 1'b1;  wr_cycle[ 1253] = 1'b0;  addr_rom[ 1253]='h00000d60;  wr_data_rom[ 1253]='h00000000;
    rd_cycle[ 1254] = 1'b1;  wr_cycle[ 1254] = 1'b0;  addr_rom[ 1254]='h00000460;  wr_data_rom[ 1254]='h00000000;
    rd_cycle[ 1255] = 1'b1;  wr_cycle[ 1255] = 1'b0;  addr_rom[ 1255]='h0000027c;  wr_data_rom[ 1255]='h00000000;
    rd_cycle[ 1256] = 1'b1;  wr_cycle[ 1256] = 1'b0;  addr_rom[ 1256]='h00000b24;  wr_data_rom[ 1256]='h00000000;
    rd_cycle[ 1257] = 1'b0;  wr_cycle[ 1257] = 1'b1;  addr_rom[ 1257]='h000001b0;  wr_data_rom[ 1257]='h00000b50;
    rd_cycle[ 1258] = 1'b0;  wr_cycle[ 1258] = 1'b1;  addr_rom[ 1258]='h000005a8;  wr_data_rom[ 1258]='h00000840;
    rd_cycle[ 1259] = 1'b1;  wr_cycle[ 1259] = 1'b0;  addr_rom[ 1259]='h00000b64;  wr_data_rom[ 1259]='h00000000;
    rd_cycle[ 1260] = 1'b1;  wr_cycle[ 1260] = 1'b0;  addr_rom[ 1260]='h00000a98;  wr_data_rom[ 1260]='h00000000;
    rd_cycle[ 1261] = 1'b0;  wr_cycle[ 1261] = 1'b1;  addr_rom[ 1261]='h00000ba8;  wr_data_rom[ 1261]='h00000eed;
    rd_cycle[ 1262] = 1'b0;  wr_cycle[ 1262] = 1'b1;  addr_rom[ 1262]='h00000ad8;  wr_data_rom[ 1262]='h00000bfd;
    rd_cycle[ 1263] = 1'b1;  wr_cycle[ 1263] = 1'b0;  addr_rom[ 1263]='h00000f70;  wr_data_rom[ 1263]='h00000000;
    rd_cycle[ 1264] = 1'b1;  wr_cycle[ 1264] = 1'b0;  addr_rom[ 1264]='h00000ae0;  wr_data_rom[ 1264]='h00000000;
    rd_cycle[ 1265] = 1'b1;  wr_cycle[ 1265] = 1'b0;  addr_rom[ 1265]='h00000a34;  wr_data_rom[ 1265]='h00000000;
    rd_cycle[ 1266] = 1'b0;  wr_cycle[ 1266] = 1'b1;  addr_rom[ 1266]='h00000778;  wr_data_rom[ 1266]='h00000d8e;
    rd_cycle[ 1267] = 1'b0;  wr_cycle[ 1267] = 1'b1;  addr_rom[ 1267]='h000007d4;  wr_data_rom[ 1267]='h0000053f;
    rd_cycle[ 1268] = 1'b1;  wr_cycle[ 1268] = 1'b0;  addr_rom[ 1268]='h000007cc;  wr_data_rom[ 1268]='h00000000;
    rd_cycle[ 1269] = 1'b0;  wr_cycle[ 1269] = 1'b1;  addr_rom[ 1269]='h000001dc;  wr_data_rom[ 1269]='h00000628;
    rd_cycle[ 1270] = 1'b0;  wr_cycle[ 1270] = 1'b1;  addr_rom[ 1270]='h00000f18;  wr_data_rom[ 1270]='h000005ea;
    rd_cycle[ 1271] = 1'b0;  wr_cycle[ 1271] = 1'b1;  addr_rom[ 1271]='h00000164;  wr_data_rom[ 1271]='h00000c7f;
    rd_cycle[ 1272] = 1'b0;  wr_cycle[ 1272] = 1'b1;  addr_rom[ 1272]='h00000bc4;  wr_data_rom[ 1272]='h00000516;
    rd_cycle[ 1273] = 1'b0;  wr_cycle[ 1273] = 1'b1;  addr_rom[ 1273]='h00000a34;  wr_data_rom[ 1273]='h0000034f;
    rd_cycle[ 1274] = 1'b0;  wr_cycle[ 1274] = 1'b1;  addr_rom[ 1274]='h00000f8c;  wr_data_rom[ 1274]='h00000236;
    rd_cycle[ 1275] = 1'b1;  wr_cycle[ 1275] = 1'b0;  addr_rom[ 1275]='h00000380;  wr_data_rom[ 1275]='h00000000;
    rd_cycle[ 1276] = 1'b1;  wr_cycle[ 1276] = 1'b0;  addr_rom[ 1276]='h000001ac;  wr_data_rom[ 1276]='h00000000;
    rd_cycle[ 1277] = 1'b0;  wr_cycle[ 1277] = 1'b1;  addr_rom[ 1277]='h00000af8;  wr_data_rom[ 1277]='h0000005d;
    rd_cycle[ 1278] = 1'b1;  wr_cycle[ 1278] = 1'b0;  addr_rom[ 1278]='h000002c0;  wr_data_rom[ 1278]='h00000000;
    rd_cycle[ 1279] = 1'b1;  wr_cycle[ 1279] = 1'b0;  addr_rom[ 1279]='h00000f90;  wr_data_rom[ 1279]='h00000000;
    rd_cycle[ 1280] = 1'b1;  wr_cycle[ 1280] = 1'b0;  addr_rom[ 1280]='h00000a8c;  wr_data_rom[ 1280]='h00000000;
    rd_cycle[ 1281] = 1'b1;  wr_cycle[ 1281] = 1'b0;  addr_rom[ 1281]='h00000794;  wr_data_rom[ 1281]='h00000000;
    rd_cycle[ 1282] = 1'b0;  wr_cycle[ 1282] = 1'b1;  addr_rom[ 1282]='h00000070;  wr_data_rom[ 1282]='h00000ab5;
    rd_cycle[ 1283] = 1'b1;  wr_cycle[ 1283] = 1'b0;  addr_rom[ 1283]='h0000080c;  wr_data_rom[ 1283]='h00000000;
    rd_cycle[ 1284] = 1'b0;  wr_cycle[ 1284] = 1'b1;  addr_rom[ 1284]='h00000264;  wr_data_rom[ 1284]='h00000d18;
    rd_cycle[ 1285] = 1'b0;  wr_cycle[ 1285] = 1'b1;  addr_rom[ 1285]='h000005b8;  wr_data_rom[ 1285]='h0000030b;
    rd_cycle[ 1286] = 1'b1;  wr_cycle[ 1286] = 1'b0;  addr_rom[ 1286]='h00000ed0;  wr_data_rom[ 1286]='h00000000;
    rd_cycle[ 1287] = 1'b1;  wr_cycle[ 1287] = 1'b0;  addr_rom[ 1287]='h00000260;  wr_data_rom[ 1287]='h00000000;
    rd_cycle[ 1288] = 1'b0;  wr_cycle[ 1288] = 1'b1;  addr_rom[ 1288]='h00000cfc;  wr_data_rom[ 1288]='h000000cd;
    rd_cycle[ 1289] = 1'b0;  wr_cycle[ 1289] = 1'b1;  addr_rom[ 1289]='h00000f94;  wr_data_rom[ 1289]='h00000609;
    rd_cycle[ 1290] = 1'b0;  wr_cycle[ 1290] = 1'b1;  addr_rom[ 1290]='h00000c6c;  wr_data_rom[ 1290]='h00000919;
    rd_cycle[ 1291] = 1'b1;  wr_cycle[ 1291] = 1'b0;  addr_rom[ 1291]='h00000d64;  wr_data_rom[ 1291]='h00000000;
    rd_cycle[ 1292] = 1'b0;  wr_cycle[ 1292] = 1'b1;  addr_rom[ 1292]='h00000d00;  wr_data_rom[ 1292]='h00000c9b;
    rd_cycle[ 1293] = 1'b1;  wr_cycle[ 1293] = 1'b0;  addr_rom[ 1293]='h00000474;  wr_data_rom[ 1293]='h00000000;
    rd_cycle[ 1294] = 1'b1;  wr_cycle[ 1294] = 1'b0;  addr_rom[ 1294]='h00000a84;  wr_data_rom[ 1294]='h00000000;
    rd_cycle[ 1295] = 1'b0;  wr_cycle[ 1295] = 1'b1;  addr_rom[ 1295]='h000003d0;  wr_data_rom[ 1295]='h00000539;
    rd_cycle[ 1296] = 1'b0;  wr_cycle[ 1296] = 1'b1;  addr_rom[ 1296]='h00000180;  wr_data_rom[ 1296]='h00000d00;
    rd_cycle[ 1297] = 1'b1;  wr_cycle[ 1297] = 1'b0;  addr_rom[ 1297]='h00000f4c;  wr_data_rom[ 1297]='h00000000;
    rd_cycle[ 1298] = 1'b0;  wr_cycle[ 1298] = 1'b1;  addr_rom[ 1298]='h000006b0;  wr_data_rom[ 1298]='h00000f62;
    rd_cycle[ 1299] = 1'b0;  wr_cycle[ 1299] = 1'b1;  addr_rom[ 1299]='h00000d40;  wr_data_rom[ 1299]='h00000972;
    rd_cycle[ 1300] = 1'b1;  wr_cycle[ 1300] = 1'b0;  addr_rom[ 1300]='h00000e68;  wr_data_rom[ 1300]='h00000000;
    rd_cycle[ 1301] = 1'b1;  wr_cycle[ 1301] = 1'b0;  addr_rom[ 1301]='h000005bc;  wr_data_rom[ 1301]='h00000000;
    rd_cycle[ 1302] = 1'b0;  wr_cycle[ 1302] = 1'b1;  addr_rom[ 1302]='h00000a24;  wr_data_rom[ 1302]='h00000c64;
    rd_cycle[ 1303] = 1'b0;  wr_cycle[ 1303] = 1'b1;  addr_rom[ 1303]='h00000258;  wr_data_rom[ 1303]='h000008f2;
    rd_cycle[ 1304] = 1'b0;  wr_cycle[ 1304] = 1'b1;  addr_rom[ 1304]='h0000058c;  wr_data_rom[ 1304]='h000006c7;
    rd_cycle[ 1305] = 1'b1;  wr_cycle[ 1305] = 1'b0;  addr_rom[ 1305]='h0000095c;  wr_data_rom[ 1305]='h00000000;
    rd_cycle[ 1306] = 1'b1;  wr_cycle[ 1306] = 1'b0;  addr_rom[ 1306]='h00000698;  wr_data_rom[ 1306]='h00000000;
    rd_cycle[ 1307] = 1'b1;  wr_cycle[ 1307] = 1'b0;  addr_rom[ 1307]='h00000630;  wr_data_rom[ 1307]='h00000000;
    rd_cycle[ 1308] = 1'b1;  wr_cycle[ 1308] = 1'b0;  addr_rom[ 1308]='h000001ac;  wr_data_rom[ 1308]='h00000000;
    rd_cycle[ 1309] = 1'b0;  wr_cycle[ 1309] = 1'b1;  addr_rom[ 1309]='h00000e68;  wr_data_rom[ 1309]='h00000cf3;
    rd_cycle[ 1310] = 1'b1;  wr_cycle[ 1310] = 1'b0;  addr_rom[ 1310]='h000009a4;  wr_data_rom[ 1310]='h00000000;
    rd_cycle[ 1311] = 1'b0;  wr_cycle[ 1311] = 1'b1;  addr_rom[ 1311]='h0000026c;  wr_data_rom[ 1311]='h00000854;
    rd_cycle[ 1312] = 1'b0;  wr_cycle[ 1312] = 1'b1;  addr_rom[ 1312]='h00000d4c;  wr_data_rom[ 1312]='h000008ba;
    rd_cycle[ 1313] = 1'b1;  wr_cycle[ 1313] = 1'b0;  addr_rom[ 1313]='h00000908;  wr_data_rom[ 1313]='h00000000;
    rd_cycle[ 1314] = 1'b1;  wr_cycle[ 1314] = 1'b0;  addr_rom[ 1314]='h00000594;  wr_data_rom[ 1314]='h00000000;
    rd_cycle[ 1315] = 1'b0;  wr_cycle[ 1315] = 1'b1;  addr_rom[ 1315]='h00000b58;  wr_data_rom[ 1315]='h000009a0;
    rd_cycle[ 1316] = 1'b0;  wr_cycle[ 1316] = 1'b1;  addr_rom[ 1316]='h00000360;  wr_data_rom[ 1316]='h00000d9d;
    rd_cycle[ 1317] = 1'b1;  wr_cycle[ 1317] = 1'b0;  addr_rom[ 1317]='h00000d84;  wr_data_rom[ 1317]='h00000000;
    rd_cycle[ 1318] = 1'b0;  wr_cycle[ 1318] = 1'b1;  addr_rom[ 1318]='h000000d8;  wr_data_rom[ 1318]='h0000058b;
    rd_cycle[ 1319] = 1'b1;  wr_cycle[ 1319] = 1'b0;  addr_rom[ 1319]='h00000e44;  wr_data_rom[ 1319]='h00000000;
    rd_cycle[ 1320] = 1'b0;  wr_cycle[ 1320] = 1'b1;  addr_rom[ 1320]='h00000538;  wr_data_rom[ 1320]='h00000065;
    rd_cycle[ 1321] = 1'b0;  wr_cycle[ 1321] = 1'b1;  addr_rom[ 1321]='h00000afc;  wr_data_rom[ 1321]='h00000865;
    rd_cycle[ 1322] = 1'b1;  wr_cycle[ 1322] = 1'b0;  addr_rom[ 1322]='h00000a20;  wr_data_rom[ 1322]='h00000000;
    rd_cycle[ 1323] = 1'b0;  wr_cycle[ 1323] = 1'b1;  addr_rom[ 1323]='h00000690;  wr_data_rom[ 1323]='h00000063;
    rd_cycle[ 1324] = 1'b1;  wr_cycle[ 1324] = 1'b0;  addr_rom[ 1324]='h000009c0;  wr_data_rom[ 1324]='h00000000;
    rd_cycle[ 1325] = 1'b0;  wr_cycle[ 1325] = 1'b1;  addr_rom[ 1325]='h000000a8;  wr_data_rom[ 1325]='h00000e32;
    rd_cycle[ 1326] = 1'b0;  wr_cycle[ 1326] = 1'b1;  addr_rom[ 1326]='h00000858;  wr_data_rom[ 1326]='h00000584;
    rd_cycle[ 1327] = 1'b0;  wr_cycle[ 1327] = 1'b1;  addr_rom[ 1327]='h0000053c;  wr_data_rom[ 1327]='h00000a90;
    rd_cycle[ 1328] = 1'b0;  wr_cycle[ 1328] = 1'b1;  addr_rom[ 1328]='h00000620;  wr_data_rom[ 1328]='h0000008c;
    rd_cycle[ 1329] = 1'b0;  wr_cycle[ 1329] = 1'b1;  addr_rom[ 1329]='h000007ec;  wr_data_rom[ 1329]='h000003f1;
    rd_cycle[ 1330] = 1'b0;  wr_cycle[ 1330] = 1'b1;  addr_rom[ 1330]='h0000010c;  wr_data_rom[ 1330]='h00000129;
    rd_cycle[ 1331] = 1'b0;  wr_cycle[ 1331] = 1'b1;  addr_rom[ 1331]='h00000424;  wr_data_rom[ 1331]='h00000028;
    rd_cycle[ 1332] = 1'b0;  wr_cycle[ 1332] = 1'b1;  addr_rom[ 1332]='h0000004c;  wr_data_rom[ 1332]='h000002de;
    rd_cycle[ 1333] = 1'b0;  wr_cycle[ 1333] = 1'b1;  addr_rom[ 1333]='h00000138;  wr_data_rom[ 1333]='h00000958;
    rd_cycle[ 1334] = 1'b1;  wr_cycle[ 1334] = 1'b0;  addr_rom[ 1334]='h00000158;  wr_data_rom[ 1334]='h00000000;
    rd_cycle[ 1335] = 1'b0;  wr_cycle[ 1335] = 1'b1;  addr_rom[ 1335]='h000007a8;  wr_data_rom[ 1335]='h000002e9;
    rd_cycle[ 1336] = 1'b1;  wr_cycle[ 1336] = 1'b0;  addr_rom[ 1336]='h000008f8;  wr_data_rom[ 1336]='h00000000;
    rd_cycle[ 1337] = 1'b0;  wr_cycle[ 1337] = 1'b1;  addr_rom[ 1337]='h00000d4c;  wr_data_rom[ 1337]='h00000186;
    rd_cycle[ 1338] = 1'b1;  wr_cycle[ 1338] = 1'b0;  addr_rom[ 1338]='h000001bc;  wr_data_rom[ 1338]='h00000000;
    rd_cycle[ 1339] = 1'b1;  wr_cycle[ 1339] = 1'b0;  addr_rom[ 1339]='h00000db0;  wr_data_rom[ 1339]='h00000000;
    rd_cycle[ 1340] = 1'b1;  wr_cycle[ 1340] = 1'b0;  addr_rom[ 1340]='h00000730;  wr_data_rom[ 1340]='h00000000;
    rd_cycle[ 1341] = 1'b0;  wr_cycle[ 1341] = 1'b1;  addr_rom[ 1341]='h0000001c;  wr_data_rom[ 1341]='h000007c0;
    rd_cycle[ 1342] = 1'b0;  wr_cycle[ 1342] = 1'b1;  addr_rom[ 1342]='h0000010c;  wr_data_rom[ 1342]='h0000083c;
    rd_cycle[ 1343] = 1'b1;  wr_cycle[ 1343] = 1'b0;  addr_rom[ 1343]='h00000a34;  wr_data_rom[ 1343]='h00000000;
    rd_cycle[ 1344] = 1'b0;  wr_cycle[ 1344] = 1'b1;  addr_rom[ 1344]='h000000c8;  wr_data_rom[ 1344]='h000006b6;
    rd_cycle[ 1345] = 1'b1;  wr_cycle[ 1345] = 1'b0;  addr_rom[ 1345]='h00000530;  wr_data_rom[ 1345]='h00000000;
    rd_cycle[ 1346] = 1'b1;  wr_cycle[ 1346] = 1'b0;  addr_rom[ 1346]='h00000744;  wr_data_rom[ 1346]='h00000000;
    rd_cycle[ 1347] = 1'b1;  wr_cycle[ 1347] = 1'b0;  addr_rom[ 1347]='h000002cc;  wr_data_rom[ 1347]='h00000000;
    rd_cycle[ 1348] = 1'b0;  wr_cycle[ 1348] = 1'b1;  addr_rom[ 1348]='h00000858;  wr_data_rom[ 1348]='h00000b40;
    rd_cycle[ 1349] = 1'b0;  wr_cycle[ 1349] = 1'b1;  addr_rom[ 1349]='h00000614;  wr_data_rom[ 1349]='h00000b64;
    rd_cycle[ 1350] = 1'b0;  wr_cycle[ 1350] = 1'b1;  addr_rom[ 1350]='h00000f40;  wr_data_rom[ 1350]='h0000039a;
    rd_cycle[ 1351] = 1'b0;  wr_cycle[ 1351] = 1'b1;  addr_rom[ 1351]='h000006bc;  wr_data_rom[ 1351]='h000006d8;
    rd_cycle[ 1352] = 1'b0;  wr_cycle[ 1352] = 1'b1;  addr_rom[ 1352]='h000001d0;  wr_data_rom[ 1352]='h000001ad;
    rd_cycle[ 1353] = 1'b1;  wr_cycle[ 1353] = 1'b0;  addr_rom[ 1353]='h00000a14;  wr_data_rom[ 1353]='h00000000;
    rd_cycle[ 1354] = 1'b0;  wr_cycle[ 1354] = 1'b1;  addr_rom[ 1354]='h000009a0;  wr_data_rom[ 1354]='h00000ddd;
    rd_cycle[ 1355] = 1'b1;  wr_cycle[ 1355] = 1'b0;  addr_rom[ 1355]='h0000058c;  wr_data_rom[ 1355]='h00000000;
    rd_cycle[ 1356] = 1'b1;  wr_cycle[ 1356] = 1'b0;  addr_rom[ 1356]='h00000984;  wr_data_rom[ 1356]='h00000000;
    rd_cycle[ 1357] = 1'b1;  wr_cycle[ 1357] = 1'b0;  addr_rom[ 1357]='h00000cd4;  wr_data_rom[ 1357]='h00000000;
    rd_cycle[ 1358] = 1'b0;  wr_cycle[ 1358] = 1'b1;  addr_rom[ 1358]='h000003e8;  wr_data_rom[ 1358]='h000007a1;
    rd_cycle[ 1359] = 1'b1;  wr_cycle[ 1359] = 1'b0;  addr_rom[ 1359]='h00000d58;  wr_data_rom[ 1359]='h00000000;
    rd_cycle[ 1360] = 1'b0;  wr_cycle[ 1360] = 1'b1;  addr_rom[ 1360]='h000004c0;  wr_data_rom[ 1360]='h00000cc0;
    rd_cycle[ 1361] = 1'b0;  wr_cycle[ 1361] = 1'b1;  addr_rom[ 1361]='h00000bfc;  wr_data_rom[ 1361]='h00000b6b;
    rd_cycle[ 1362] = 1'b1;  wr_cycle[ 1362] = 1'b0;  addr_rom[ 1362]='h000003e8;  wr_data_rom[ 1362]='h00000000;
    rd_cycle[ 1363] = 1'b1;  wr_cycle[ 1363] = 1'b0;  addr_rom[ 1363]='h00000460;  wr_data_rom[ 1363]='h00000000;
    rd_cycle[ 1364] = 1'b1;  wr_cycle[ 1364] = 1'b0;  addr_rom[ 1364]='h000002b8;  wr_data_rom[ 1364]='h00000000;
    rd_cycle[ 1365] = 1'b1;  wr_cycle[ 1365] = 1'b0;  addr_rom[ 1365]='h000006c8;  wr_data_rom[ 1365]='h00000000;
    rd_cycle[ 1366] = 1'b1;  wr_cycle[ 1366] = 1'b0;  addr_rom[ 1366]='h00000844;  wr_data_rom[ 1366]='h00000000;
    rd_cycle[ 1367] = 1'b0;  wr_cycle[ 1367] = 1'b1;  addr_rom[ 1367]='h00000dc0;  wr_data_rom[ 1367]='h0000053c;
    rd_cycle[ 1368] = 1'b1;  wr_cycle[ 1368] = 1'b0;  addr_rom[ 1368]='h00000464;  wr_data_rom[ 1368]='h00000000;
    rd_cycle[ 1369] = 1'b1;  wr_cycle[ 1369] = 1'b0;  addr_rom[ 1369]='h000000cc;  wr_data_rom[ 1369]='h00000000;
    rd_cycle[ 1370] = 1'b0;  wr_cycle[ 1370] = 1'b1;  addr_rom[ 1370]='h00000b48;  wr_data_rom[ 1370]='h00000e71;
    rd_cycle[ 1371] = 1'b0;  wr_cycle[ 1371] = 1'b1;  addr_rom[ 1371]='h00000050;  wr_data_rom[ 1371]='h00000d12;
    rd_cycle[ 1372] = 1'b1;  wr_cycle[ 1372] = 1'b0;  addr_rom[ 1372]='h00000e3c;  wr_data_rom[ 1372]='h00000000;
    rd_cycle[ 1373] = 1'b0;  wr_cycle[ 1373] = 1'b1;  addr_rom[ 1373]='h00000b28;  wr_data_rom[ 1373]='h0000063b;
    rd_cycle[ 1374] = 1'b1;  wr_cycle[ 1374] = 1'b0;  addr_rom[ 1374]='h000001fc;  wr_data_rom[ 1374]='h00000000;
    rd_cycle[ 1375] = 1'b1;  wr_cycle[ 1375] = 1'b0;  addr_rom[ 1375]='h000002d4;  wr_data_rom[ 1375]='h00000000;
    rd_cycle[ 1376] = 1'b0;  wr_cycle[ 1376] = 1'b1;  addr_rom[ 1376]='h000001f4;  wr_data_rom[ 1376]='h00000b86;
    rd_cycle[ 1377] = 1'b0;  wr_cycle[ 1377] = 1'b1;  addr_rom[ 1377]='h0000093c;  wr_data_rom[ 1377]='h000005aa;
    rd_cycle[ 1378] = 1'b0;  wr_cycle[ 1378] = 1'b1;  addr_rom[ 1378]='h00000838;  wr_data_rom[ 1378]='h0000092c;
    rd_cycle[ 1379] = 1'b1;  wr_cycle[ 1379] = 1'b0;  addr_rom[ 1379]='h000007ec;  wr_data_rom[ 1379]='h00000000;
    rd_cycle[ 1380] = 1'b0;  wr_cycle[ 1380] = 1'b1;  addr_rom[ 1380]='h000003b4;  wr_data_rom[ 1380]='h000006d2;
    rd_cycle[ 1381] = 1'b1;  wr_cycle[ 1381] = 1'b0;  addr_rom[ 1381]='h000008e4;  wr_data_rom[ 1381]='h00000000;
    rd_cycle[ 1382] = 1'b0;  wr_cycle[ 1382] = 1'b1;  addr_rom[ 1382]='h00000324;  wr_data_rom[ 1382]='h00000131;
    rd_cycle[ 1383] = 1'b0;  wr_cycle[ 1383] = 1'b1;  addr_rom[ 1383]='h00000668;  wr_data_rom[ 1383]='h00000b7c;
    rd_cycle[ 1384] = 1'b1;  wr_cycle[ 1384] = 1'b0;  addr_rom[ 1384]='h00000b8c;  wr_data_rom[ 1384]='h00000000;
    rd_cycle[ 1385] = 1'b1;  wr_cycle[ 1385] = 1'b0;  addr_rom[ 1385]='h00000850;  wr_data_rom[ 1385]='h00000000;
    rd_cycle[ 1386] = 1'b1;  wr_cycle[ 1386] = 1'b0;  addr_rom[ 1386]='h00000214;  wr_data_rom[ 1386]='h00000000;
    rd_cycle[ 1387] = 1'b1;  wr_cycle[ 1387] = 1'b0;  addr_rom[ 1387]='h00000178;  wr_data_rom[ 1387]='h00000000;
    rd_cycle[ 1388] = 1'b0;  wr_cycle[ 1388] = 1'b1;  addr_rom[ 1388]='h00000de0;  wr_data_rom[ 1388]='h00000ee6;
    rd_cycle[ 1389] = 1'b0;  wr_cycle[ 1389] = 1'b1;  addr_rom[ 1389]='h000003e4;  wr_data_rom[ 1389]='h00000b6d;
    rd_cycle[ 1390] = 1'b1;  wr_cycle[ 1390] = 1'b0;  addr_rom[ 1390]='h00000f70;  wr_data_rom[ 1390]='h00000000;
    rd_cycle[ 1391] = 1'b0;  wr_cycle[ 1391] = 1'b1;  addr_rom[ 1391]='h00000c78;  wr_data_rom[ 1391]='h0000015d;
    rd_cycle[ 1392] = 1'b0;  wr_cycle[ 1392] = 1'b1;  addr_rom[ 1392]='h00000e1c;  wr_data_rom[ 1392]='h00000401;
    rd_cycle[ 1393] = 1'b1;  wr_cycle[ 1393] = 1'b0;  addr_rom[ 1393]='h00000c7c;  wr_data_rom[ 1393]='h00000000;
    rd_cycle[ 1394] = 1'b1;  wr_cycle[ 1394] = 1'b0;  addr_rom[ 1394]='h000008b8;  wr_data_rom[ 1394]='h00000000;
    rd_cycle[ 1395] = 1'b0;  wr_cycle[ 1395] = 1'b1;  addr_rom[ 1395]='h00000498;  wr_data_rom[ 1395]='h00000a12;
    rd_cycle[ 1396] = 1'b1;  wr_cycle[ 1396] = 1'b0;  addr_rom[ 1396]='h00000828;  wr_data_rom[ 1396]='h00000000;
    rd_cycle[ 1397] = 1'b1;  wr_cycle[ 1397] = 1'b0;  addr_rom[ 1397]='h00000140;  wr_data_rom[ 1397]='h00000000;
    rd_cycle[ 1398] = 1'b1;  wr_cycle[ 1398] = 1'b0;  addr_rom[ 1398]='h00000a54;  wr_data_rom[ 1398]='h00000000;
    rd_cycle[ 1399] = 1'b1;  wr_cycle[ 1399] = 1'b0;  addr_rom[ 1399]='h0000050c;  wr_data_rom[ 1399]='h00000000;
    rd_cycle[ 1400] = 1'b0;  wr_cycle[ 1400] = 1'b1;  addr_rom[ 1400]='h000000c0;  wr_data_rom[ 1400]='h000007a0;
    rd_cycle[ 1401] = 1'b0;  wr_cycle[ 1401] = 1'b1;  addr_rom[ 1401]='h00000950;  wr_data_rom[ 1401]='h00000205;
    rd_cycle[ 1402] = 1'b1;  wr_cycle[ 1402] = 1'b0;  addr_rom[ 1402]='h000006b4;  wr_data_rom[ 1402]='h00000000;
    rd_cycle[ 1403] = 1'b0;  wr_cycle[ 1403] = 1'b1;  addr_rom[ 1403]='h00000688;  wr_data_rom[ 1403]='h00000f1f;
    rd_cycle[ 1404] = 1'b1;  wr_cycle[ 1404] = 1'b0;  addr_rom[ 1404]='h000002c0;  wr_data_rom[ 1404]='h00000000;
    rd_cycle[ 1405] = 1'b0;  wr_cycle[ 1405] = 1'b1;  addr_rom[ 1405]='h0000031c;  wr_data_rom[ 1405]='h00000cdf;
    rd_cycle[ 1406] = 1'b1;  wr_cycle[ 1406] = 1'b0;  addr_rom[ 1406]='h00000728;  wr_data_rom[ 1406]='h00000000;
    rd_cycle[ 1407] = 1'b1;  wr_cycle[ 1407] = 1'b0;  addr_rom[ 1407]='h000003f8;  wr_data_rom[ 1407]='h00000000;
    rd_cycle[ 1408] = 1'b1;  wr_cycle[ 1408] = 1'b0;  addr_rom[ 1408]='h0000052c;  wr_data_rom[ 1408]='h00000000;
    rd_cycle[ 1409] = 1'b0;  wr_cycle[ 1409] = 1'b1;  addr_rom[ 1409]='h00000a80;  wr_data_rom[ 1409]='h00000203;
    rd_cycle[ 1410] = 1'b1;  wr_cycle[ 1410] = 1'b0;  addr_rom[ 1410]='h00000a30;  wr_data_rom[ 1410]='h00000000;
    rd_cycle[ 1411] = 1'b1;  wr_cycle[ 1411] = 1'b0;  addr_rom[ 1411]='h00000a78;  wr_data_rom[ 1411]='h00000000;
    rd_cycle[ 1412] = 1'b0;  wr_cycle[ 1412] = 1'b1;  addr_rom[ 1412]='h000005bc;  wr_data_rom[ 1412]='h000004db;
    rd_cycle[ 1413] = 1'b0;  wr_cycle[ 1413] = 1'b1;  addr_rom[ 1413]='h0000090c;  wr_data_rom[ 1413]='h00000b0e;
    rd_cycle[ 1414] = 1'b0;  wr_cycle[ 1414] = 1'b1;  addr_rom[ 1414]='h00000008;  wr_data_rom[ 1414]='h00000e0f;
    rd_cycle[ 1415] = 1'b0;  wr_cycle[ 1415] = 1'b1;  addr_rom[ 1415]='h0000004c;  wr_data_rom[ 1415]='h00000202;
    rd_cycle[ 1416] = 1'b1;  wr_cycle[ 1416] = 1'b0;  addr_rom[ 1416]='h00000e08;  wr_data_rom[ 1416]='h00000000;
    rd_cycle[ 1417] = 1'b1;  wr_cycle[ 1417] = 1'b0;  addr_rom[ 1417]='h000002f0;  wr_data_rom[ 1417]='h00000000;
    rd_cycle[ 1418] = 1'b1;  wr_cycle[ 1418] = 1'b0;  addr_rom[ 1418]='h000003d8;  wr_data_rom[ 1418]='h00000000;
    rd_cycle[ 1419] = 1'b0;  wr_cycle[ 1419] = 1'b1;  addr_rom[ 1419]='h00000a8c;  wr_data_rom[ 1419]='h00000de8;
    rd_cycle[ 1420] = 1'b1;  wr_cycle[ 1420] = 1'b0;  addr_rom[ 1420]='h00000428;  wr_data_rom[ 1420]='h00000000;
    rd_cycle[ 1421] = 1'b1;  wr_cycle[ 1421] = 1'b0;  addr_rom[ 1421]='h000002a0;  wr_data_rom[ 1421]='h00000000;
    rd_cycle[ 1422] = 1'b1;  wr_cycle[ 1422] = 1'b0;  addr_rom[ 1422]='h000002b8;  wr_data_rom[ 1422]='h00000000;
    rd_cycle[ 1423] = 1'b1;  wr_cycle[ 1423] = 1'b0;  addr_rom[ 1423]='h00000490;  wr_data_rom[ 1423]='h00000000;
    rd_cycle[ 1424] = 1'b1;  wr_cycle[ 1424] = 1'b0;  addr_rom[ 1424]='h00000474;  wr_data_rom[ 1424]='h00000000;
    rd_cycle[ 1425] = 1'b0;  wr_cycle[ 1425] = 1'b1;  addr_rom[ 1425]='h00000b70;  wr_data_rom[ 1425]='h0000057f;
    rd_cycle[ 1426] = 1'b1;  wr_cycle[ 1426] = 1'b0;  addr_rom[ 1426]='h00000d78;  wr_data_rom[ 1426]='h00000000;
    rd_cycle[ 1427] = 1'b1;  wr_cycle[ 1427] = 1'b0;  addr_rom[ 1427]='h00000784;  wr_data_rom[ 1427]='h00000000;
    rd_cycle[ 1428] = 1'b1;  wr_cycle[ 1428] = 1'b0;  addr_rom[ 1428]='h00000810;  wr_data_rom[ 1428]='h00000000;
    rd_cycle[ 1429] = 1'b1;  wr_cycle[ 1429] = 1'b0;  addr_rom[ 1429]='h00000c7c;  wr_data_rom[ 1429]='h00000000;
    rd_cycle[ 1430] = 1'b1;  wr_cycle[ 1430] = 1'b0;  addr_rom[ 1430]='h00000270;  wr_data_rom[ 1430]='h00000000;
    rd_cycle[ 1431] = 1'b1;  wr_cycle[ 1431] = 1'b0;  addr_rom[ 1431]='h00000274;  wr_data_rom[ 1431]='h00000000;
    rd_cycle[ 1432] = 1'b1;  wr_cycle[ 1432] = 1'b0;  addr_rom[ 1432]='h000003d0;  wr_data_rom[ 1432]='h00000000;
    rd_cycle[ 1433] = 1'b0;  wr_cycle[ 1433] = 1'b1;  addr_rom[ 1433]='h00000398;  wr_data_rom[ 1433]='h00000215;
    rd_cycle[ 1434] = 1'b1;  wr_cycle[ 1434] = 1'b0;  addr_rom[ 1434]='h0000077c;  wr_data_rom[ 1434]='h00000000;
    rd_cycle[ 1435] = 1'b0;  wr_cycle[ 1435] = 1'b1;  addr_rom[ 1435]='h00000588;  wr_data_rom[ 1435]='h00000ae6;
    rd_cycle[ 1436] = 1'b1;  wr_cycle[ 1436] = 1'b0;  addr_rom[ 1436]='h00000a3c;  wr_data_rom[ 1436]='h00000000;
    rd_cycle[ 1437] = 1'b1;  wr_cycle[ 1437] = 1'b0;  addr_rom[ 1437]='h000003a0;  wr_data_rom[ 1437]='h00000000;
    rd_cycle[ 1438] = 1'b0;  wr_cycle[ 1438] = 1'b1;  addr_rom[ 1438]='h00000f4c;  wr_data_rom[ 1438]='h00000f48;
    rd_cycle[ 1439] = 1'b0;  wr_cycle[ 1439] = 1'b1;  addr_rom[ 1439]='h00000710;  wr_data_rom[ 1439]='h0000056d;
    rd_cycle[ 1440] = 1'b0;  wr_cycle[ 1440] = 1'b1;  addr_rom[ 1440]='h00000e78;  wr_data_rom[ 1440]='h000001b3;
    rd_cycle[ 1441] = 1'b1;  wr_cycle[ 1441] = 1'b0;  addr_rom[ 1441]='h0000049c;  wr_data_rom[ 1441]='h00000000;
    rd_cycle[ 1442] = 1'b0;  wr_cycle[ 1442] = 1'b1;  addr_rom[ 1442]='h000004cc;  wr_data_rom[ 1442]='h00000bb2;
    rd_cycle[ 1443] = 1'b1;  wr_cycle[ 1443] = 1'b0;  addr_rom[ 1443]='h0000030c;  wr_data_rom[ 1443]='h00000000;
    rd_cycle[ 1444] = 1'b0;  wr_cycle[ 1444] = 1'b1;  addr_rom[ 1444]='h0000081c;  wr_data_rom[ 1444]='h00000e87;
    rd_cycle[ 1445] = 1'b1;  wr_cycle[ 1445] = 1'b0;  addr_rom[ 1445]='h00000ce8;  wr_data_rom[ 1445]='h00000000;
    rd_cycle[ 1446] = 1'b1;  wr_cycle[ 1446] = 1'b0;  addr_rom[ 1446]='h00000a54;  wr_data_rom[ 1446]='h00000000;
    rd_cycle[ 1447] = 1'b0;  wr_cycle[ 1447] = 1'b1;  addr_rom[ 1447]='h0000012c;  wr_data_rom[ 1447]='h00000f99;
    rd_cycle[ 1448] = 1'b0;  wr_cycle[ 1448] = 1'b1;  addr_rom[ 1448]='h00000e38;  wr_data_rom[ 1448]='h00000186;
    rd_cycle[ 1449] = 1'b0;  wr_cycle[ 1449] = 1'b1;  addr_rom[ 1449]='h000002d8;  wr_data_rom[ 1449]='h000002bf;
    rd_cycle[ 1450] = 1'b0;  wr_cycle[ 1450] = 1'b1;  addr_rom[ 1450]='h0000078c;  wr_data_rom[ 1450]='h00000f67;
    rd_cycle[ 1451] = 1'b0;  wr_cycle[ 1451] = 1'b1;  addr_rom[ 1451]='h000004c8;  wr_data_rom[ 1451]='h00000027;
    rd_cycle[ 1452] = 1'b1;  wr_cycle[ 1452] = 1'b0;  addr_rom[ 1452]='h00000498;  wr_data_rom[ 1452]='h00000000;
    rd_cycle[ 1453] = 1'b0;  wr_cycle[ 1453] = 1'b1;  addr_rom[ 1453]='h00000784;  wr_data_rom[ 1453]='h000004cb;
    rd_cycle[ 1454] = 1'b0;  wr_cycle[ 1454] = 1'b1;  addr_rom[ 1454]='h00000cf4;  wr_data_rom[ 1454]='h00000b52;
    rd_cycle[ 1455] = 1'b0;  wr_cycle[ 1455] = 1'b1;  addr_rom[ 1455]='h00000350;  wr_data_rom[ 1455]='h00000307;
    rd_cycle[ 1456] = 1'b1;  wr_cycle[ 1456] = 1'b0;  addr_rom[ 1456]='h00000e5c;  wr_data_rom[ 1456]='h00000000;
    rd_cycle[ 1457] = 1'b1;  wr_cycle[ 1457] = 1'b0;  addr_rom[ 1457]='h00000e74;  wr_data_rom[ 1457]='h00000000;
    rd_cycle[ 1458] = 1'b1;  wr_cycle[ 1458] = 1'b0;  addr_rom[ 1458]='h00000994;  wr_data_rom[ 1458]='h00000000;
    rd_cycle[ 1459] = 1'b1;  wr_cycle[ 1459] = 1'b0;  addr_rom[ 1459]='h000006a4;  wr_data_rom[ 1459]='h00000000;
    rd_cycle[ 1460] = 1'b0;  wr_cycle[ 1460] = 1'b1;  addr_rom[ 1460]='h00000ca8;  wr_data_rom[ 1460]='h000000b5;
    rd_cycle[ 1461] = 1'b1;  wr_cycle[ 1461] = 1'b0;  addr_rom[ 1461]='h00000788;  wr_data_rom[ 1461]='h00000000;
    rd_cycle[ 1462] = 1'b1;  wr_cycle[ 1462] = 1'b0;  addr_rom[ 1462]='h00000b88;  wr_data_rom[ 1462]='h00000000;
    rd_cycle[ 1463] = 1'b0;  wr_cycle[ 1463] = 1'b1;  addr_rom[ 1463]='h00000734;  wr_data_rom[ 1463]='h000007c7;
    rd_cycle[ 1464] = 1'b0;  wr_cycle[ 1464] = 1'b1;  addr_rom[ 1464]='h00000078;  wr_data_rom[ 1464]='h0000038d;
    rd_cycle[ 1465] = 1'b0;  wr_cycle[ 1465] = 1'b1;  addr_rom[ 1465]='h00000cd0;  wr_data_rom[ 1465]='h00000487;
    rd_cycle[ 1466] = 1'b0;  wr_cycle[ 1466] = 1'b1;  addr_rom[ 1466]='h00000b0c;  wr_data_rom[ 1466]='h00000d59;
    rd_cycle[ 1467] = 1'b0;  wr_cycle[ 1467] = 1'b1;  addr_rom[ 1467]='h00000a7c;  wr_data_rom[ 1467]='h00000768;
    rd_cycle[ 1468] = 1'b0;  wr_cycle[ 1468] = 1'b1;  addr_rom[ 1468]='h000002d4;  wr_data_rom[ 1468]='h000007f9;
    rd_cycle[ 1469] = 1'b1;  wr_cycle[ 1469] = 1'b0;  addr_rom[ 1469]='h0000034c;  wr_data_rom[ 1469]='h00000000;
    rd_cycle[ 1470] = 1'b0;  wr_cycle[ 1470] = 1'b1;  addr_rom[ 1470]='h000007c8;  wr_data_rom[ 1470]='h00000d9f;
    rd_cycle[ 1471] = 1'b1;  wr_cycle[ 1471] = 1'b0;  addr_rom[ 1471]='h00000728;  wr_data_rom[ 1471]='h00000000;
    rd_cycle[ 1472] = 1'b1;  wr_cycle[ 1472] = 1'b0;  addr_rom[ 1472]='h00000090;  wr_data_rom[ 1472]='h00000000;
    rd_cycle[ 1473] = 1'b1;  wr_cycle[ 1473] = 1'b0;  addr_rom[ 1473]='h00000554;  wr_data_rom[ 1473]='h00000000;
    rd_cycle[ 1474] = 1'b0;  wr_cycle[ 1474] = 1'b1;  addr_rom[ 1474]='h00000684;  wr_data_rom[ 1474]='h00000341;
    rd_cycle[ 1475] = 1'b1;  wr_cycle[ 1475] = 1'b0;  addr_rom[ 1475]='h00000888;  wr_data_rom[ 1475]='h00000000;
    rd_cycle[ 1476] = 1'b1;  wr_cycle[ 1476] = 1'b0;  addr_rom[ 1476]='h00000254;  wr_data_rom[ 1476]='h00000000;
    rd_cycle[ 1477] = 1'b0;  wr_cycle[ 1477] = 1'b1;  addr_rom[ 1477]='h00000e1c;  wr_data_rom[ 1477]='h00000926;
    rd_cycle[ 1478] = 1'b1;  wr_cycle[ 1478] = 1'b0;  addr_rom[ 1478]='h000009f8;  wr_data_rom[ 1478]='h00000000;
    rd_cycle[ 1479] = 1'b1;  wr_cycle[ 1479] = 1'b0;  addr_rom[ 1479]='h00000738;  wr_data_rom[ 1479]='h00000000;
    rd_cycle[ 1480] = 1'b1;  wr_cycle[ 1480] = 1'b0;  addr_rom[ 1480]='h00000e1c;  wr_data_rom[ 1480]='h00000000;
    rd_cycle[ 1481] = 1'b0;  wr_cycle[ 1481] = 1'b1;  addr_rom[ 1481]='h00000610;  wr_data_rom[ 1481]='h000002f1;
    rd_cycle[ 1482] = 1'b0;  wr_cycle[ 1482] = 1'b1;  addr_rom[ 1482]='h000009b8;  wr_data_rom[ 1482]='h00000603;
    rd_cycle[ 1483] = 1'b0;  wr_cycle[ 1483] = 1'b1;  addr_rom[ 1483]='h000001fc;  wr_data_rom[ 1483]='h00000bac;
    rd_cycle[ 1484] = 1'b0;  wr_cycle[ 1484] = 1'b1;  addr_rom[ 1484]='h00000330;  wr_data_rom[ 1484]='h000005ba;
    rd_cycle[ 1485] = 1'b1;  wr_cycle[ 1485] = 1'b0;  addr_rom[ 1485]='h00000da0;  wr_data_rom[ 1485]='h00000000;
    rd_cycle[ 1486] = 1'b0;  wr_cycle[ 1486] = 1'b1;  addr_rom[ 1486]='h0000010c;  wr_data_rom[ 1486]='h00000c03;
    rd_cycle[ 1487] = 1'b1;  wr_cycle[ 1487] = 1'b0;  addr_rom[ 1487]='h00000cb8;  wr_data_rom[ 1487]='h00000000;
    rd_cycle[ 1488] = 1'b0;  wr_cycle[ 1488] = 1'b1;  addr_rom[ 1488]='h000007cc;  wr_data_rom[ 1488]='h00000709;
    rd_cycle[ 1489] = 1'b0;  wr_cycle[ 1489] = 1'b1;  addr_rom[ 1489]='h00000a84;  wr_data_rom[ 1489]='h00000a88;
    rd_cycle[ 1490] = 1'b1;  wr_cycle[ 1490] = 1'b0;  addr_rom[ 1490]='h00000f8c;  wr_data_rom[ 1490]='h00000000;
    rd_cycle[ 1491] = 1'b1;  wr_cycle[ 1491] = 1'b0;  addr_rom[ 1491]='h000000e0;  wr_data_rom[ 1491]='h00000000;
    rd_cycle[ 1492] = 1'b1;  wr_cycle[ 1492] = 1'b0;  addr_rom[ 1492]='h00000888;  wr_data_rom[ 1492]='h00000000;
    rd_cycle[ 1493] = 1'b0;  wr_cycle[ 1493] = 1'b1;  addr_rom[ 1493]='h000009f0;  wr_data_rom[ 1493]='h00000802;
    rd_cycle[ 1494] = 1'b0;  wr_cycle[ 1494] = 1'b1;  addr_rom[ 1494]='h000009e8;  wr_data_rom[ 1494]='h00000e5c;
    rd_cycle[ 1495] = 1'b0;  wr_cycle[ 1495] = 1'b1;  addr_rom[ 1495]='h00000864;  wr_data_rom[ 1495]='h00000e79;
    rd_cycle[ 1496] = 1'b1;  wr_cycle[ 1496] = 1'b0;  addr_rom[ 1496]='h000002ec;  wr_data_rom[ 1496]='h00000000;
    rd_cycle[ 1497] = 1'b0;  wr_cycle[ 1497] = 1'b1;  addr_rom[ 1497]='h00000f5c;  wr_data_rom[ 1497]='h000003f8;
    rd_cycle[ 1498] = 1'b1;  wr_cycle[ 1498] = 1'b0;  addr_rom[ 1498]='h00000530;  wr_data_rom[ 1498]='h00000000;
    rd_cycle[ 1499] = 1'b1;  wr_cycle[ 1499] = 1'b0;  addr_rom[ 1499]='h00000b58;  wr_data_rom[ 1499]='h00000000;
    rd_cycle[ 1500] = 1'b1;  wr_cycle[ 1500] = 1'b0;  addr_rom[ 1500]='h00000a34;  wr_data_rom[ 1500]='h00000000;
    rd_cycle[ 1501] = 1'b1;  wr_cycle[ 1501] = 1'b0;  addr_rom[ 1501]='h00000a78;  wr_data_rom[ 1501]='h00000000;
    rd_cycle[ 1502] = 1'b1;  wr_cycle[ 1502] = 1'b0;  addr_rom[ 1502]='h00000aac;  wr_data_rom[ 1502]='h00000000;
    rd_cycle[ 1503] = 1'b1;  wr_cycle[ 1503] = 1'b0;  addr_rom[ 1503]='h00000178;  wr_data_rom[ 1503]='h00000000;
    rd_cycle[ 1504] = 1'b1;  wr_cycle[ 1504] = 1'b0;  addr_rom[ 1504]='h00000ce0;  wr_data_rom[ 1504]='h00000000;
    rd_cycle[ 1505] = 1'b0;  wr_cycle[ 1505] = 1'b1;  addr_rom[ 1505]='h000002ac;  wr_data_rom[ 1505]='h00000a7a;
    rd_cycle[ 1506] = 1'b0;  wr_cycle[ 1506] = 1'b1;  addr_rom[ 1506]='h00000ba0;  wr_data_rom[ 1506]='h00000a98;
    rd_cycle[ 1507] = 1'b1;  wr_cycle[ 1507] = 1'b0;  addr_rom[ 1507]='h0000011c;  wr_data_rom[ 1507]='h00000000;
    rd_cycle[ 1508] = 1'b0;  wr_cycle[ 1508] = 1'b1;  addr_rom[ 1508]='h000004cc;  wr_data_rom[ 1508]='h00000e23;
    rd_cycle[ 1509] = 1'b1;  wr_cycle[ 1509] = 1'b0;  addr_rom[ 1509]='h00000850;  wr_data_rom[ 1509]='h00000000;
    rd_cycle[ 1510] = 1'b1;  wr_cycle[ 1510] = 1'b0;  addr_rom[ 1510]='h000005a0;  wr_data_rom[ 1510]='h00000000;
    rd_cycle[ 1511] = 1'b0;  wr_cycle[ 1511] = 1'b1;  addr_rom[ 1511]='h000007f8;  wr_data_rom[ 1511]='h000006a1;
    rd_cycle[ 1512] = 1'b0;  wr_cycle[ 1512] = 1'b1;  addr_rom[ 1512]='h00000648;  wr_data_rom[ 1512]='h000001f7;
    rd_cycle[ 1513] = 1'b0;  wr_cycle[ 1513] = 1'b1;  addr_rom[ 1513]='h000009f4;  wr_data_rom[ 1513]='h0000021b;
    rd_cycle[ 1514] = 1'b1;  wr_cycle[ 1514] = 1'b0;  addr_rom[ 1514]='h00000d6c;  wr_data_rom[ 1514]='h00000000;
    rd_cycle[ 1515] = 1'b1;  wr_cycle[ 1515] = 1'b0;  addr_rom[ 1515]='h0000039c;  wr_data_rom[ 1515]='h00000000;
    rd_cycle[ 1516] = 1'b1;  wr_cycle[ 1516] = 1'b0;  addr_rom[ 1516]='h000009c8;  wr_data_rom[ 1516]='h00000000;
    rd_cycle[ 1517] = 1'b1;  wr_cycle[ 1517] = 1'b0;  addr_rom[ 1517]='h000000bc;  wr_data_rom[ 1517]='h00000000;
    rd_cycle[ 1518] = 1'b1;  wr_cycle[ 1518] = 1'b0;  addr_rom[ 1518]='h000005f8;  wr_data_rom[ 1518]='h00000000;
    rd_cycle[ 1519] = 1'b1;  wr_cycle[ 1519] = 1'b0;  addr_rom[ 1519]='h00000ef8;  wr_data_rom[ 1519]='h00000000;
    rd_cycle[ 1520] = 1'b0;  wr_cycle[ 1520] = 1'b1;  addr_rom[ 1520]='h000001a8;  wr_data_rom[ 1520]='h000003e2;
    rd_cycle[ 1521] = 1'b0;  wr_cycle[ 1521] = 1'b1;  addr_rom[ 1521]='h00000994;  wr_data_rom[ 1521]='h000003f7;
    rd_cycle[ 1522] = 1'b1;  wr_cycle[ 1522] = 1'b0;  addr_rom[ 1522]='h000007dc;  wr_data_rom[ 1522]='h00000000;
    rd_cycle[ 1523] = 1'b0;  wr_cycle[ 1523] = 1'b1;  addr_rom[ 1523]='h0000076c;  wr_data_rom[ 1523]='h00000eb0;
    rd_cycle[ 1524] = 1'b1;  wr_cycle[ 1524] = 1'b0;  addr_rom[ 1524]='h00000eb0;  wr_data_rom[ 1524]='h00000000;
    rd_cycle[ 1525] = 1'b1;  wr_cycle[ 1525] = 1'b0;  addr_rom[ 1525]='h00000a28;  wr_data_rom[ 1525]='h00000000;
    rd_cycle[ 1526] = 1'b1;  wr_cycle[ 1526] = 1'b0;  addr_rom[ 1526]='h00000064;  wr_data_rom[ 1526]='h00000000;
    rd_cycle[ 1527] = 1'b0;  wr_cycle[ 1527] = 1'b1;  addr_rom[ 1527]='h00000b44;  wr_data_rom[ 1527]='h0000076f;
    rd_cycle[ 1528] = 1'b0;  wr_cycle[ 1528] = 1'b1;  addr_rom[ 1528]='h00000468;  wr_data_rom[ 1528]='h00000db6;
    rd_cycle[ 1529] = 1'b0;  wr_cycle[ 1529] = 1'b1;  addr_rom[ 1529]='h00000b04;  wr_data_rom[ 1529]='h00000bdf;
    rd_cycle[ 1530] = 1'b1;  wr_cycle[ 1530] = 1'b0;  addr_rom[ 1530]='h00000774;  wr_data_rom[ 1530]='h00000000;
    rd_cycle[ 1531] = 1'b1;  wr_cycle[ 1531] = 1'b0;  addr_rom[ 1531]='h00000c38;  wr_data_rom[ 1531]='h00000000;
    rd_cycle[ 1532] = 1'b1;  wr_cycle[ 1532] = 1'b0;  addr_rom[ 1532]='h000007cc;  wr_data_rom[ 1532]='h00000000;
    rd_cycle[ 1533] = 1'b1;  wr_cycle[ 1533] = 1'b0;  addr_rom[ 1533]='h00000d68;  wr_data_rom[ 1533]='h00000000;
    rd_cycle[ 1534] = 1'b1;  wr_cycle[ 1534] = 1'b0;  addr_rom[ 1534]='h00000224;  wr_data_rom[ 1534]='h00000000;
    rd_cycle[ 1535] = 1'b1;  wr_cycle[ 1535] = 1'b0;  addr_rom[ 1535]='h000007b8;  wr_data_rom[ 1535]='h00000000;
    rd_cycle[ 1536] = 1'b0;  wr_cycle[ 1536] = 1'b1;  addr_rom[ 1536]='h00000ae0;  wr_data_rom[ 1536]='h00000216;
    rd_cycle[ 1537] = 1'b1;  wr_cycle[ 1537] = 1'b0;  addr_rom[ 1537]='h00000704;  wr_data_rom[ 1537]='h00000000;
    rd_cycle[ 1538] = 1'b0;  wr_cycle[ 1538] = 1'b1;  addr_rom[ 1538]='h0000066c;  wr_data_rom[ 1538]='h00000ef0;
    rd_cycle[ 1539] = 1'b1;  wr_cycle[ 1539] = 1'b0;  addr_rom[ 1539]='h0000003c;  wr_data_rom[ 1539]='h00000000;
    rd_cycle[ 1540] = 1'b0;  wr_cycle[ 1540] = 1'b1;  addr_rom[ 1540]='h00000280;  wr_data_rom[ 1540]='h00000829;
    rd_cycle[ 1541] = 1'b1;  wr_cycle[ 1541] = 1'b0;  addr_rom[ 1541]='h00000e44;  wr_data_rom[ 1541]='h00000000;
    rd_cycle[ 1542] = 1'b0;  wr_cycle[ 1542] = 1'b1;  addr_rom[ 1542]='h00000b58;  wr_data_rom[ 1542]='h00000d11;
    rd_cycle[ 1543] = 1'b1;  wr_cycle[ 1543] = 1'b0;  addr_rom[ 1543]='h00000858;  wr_data_rom[ 1543]='h00000000;
    rd_cycle[ 1544] = 1'b1;  wr_cycle[ 1544] = 1'b0;  addr_rom[ 1544]='h000000ec;  wr_data_rom[ 1544]='h00000000;
    rd_cycle[ 1545] = 1'b1;  wr_cycle[ 1545] = 1'b0;  addr_rom[ 1545]='h0000016c;  wr_data_rom[ 1545]='h00000000;
    rd_cycle[ 1546] = 1'b0;  wr_cycle[ 1546] = 1'b1;  addr_rom[ 1546]='h000006e8;  wr_data_rom[ 1546]='h00000597;
    rd_cycle[ 1547] = 1'b1;  wr_cycle[ 1547] = 1'b0;  addr_rom[ 1547]='h00000b08;  wr_data_rom[ 1547]='h00000000;
    rd_cycle[ 1548] = 1'b1;  wr_cycle[ 1548] = 1'b0;  addr_rom[ 1548]='h000007dc;  wr_data_rom[ 1548]='h00000000;
    rd_cycle[ 1549] = 1'b1;  wr_cycle[ 1549] = 1'b0;  addr_rom[ 1549]='h000006ac;  wr_data_rom[ 1549]='h00000000;
    rd_cycle[ 1550] = 1'b1;  wr_cycle[ 1550] = 1'b0;  addr_rom[ 1550]='h0000093c;  wr_data_rom[ 1550]='h00000000;
    rd_cycle[ 1551] = 1'b1;  wr_cycle[ 1551] = 1'b0;  addr_rom[ 1551]='h000002ec;  wr_data_rom[ 1551]='h00000000;
    rd_cycle[ 1552] = 1'b0;  wr_cycle[ 1552] = 1'b1;  addr_rom[ 1552]='h00000cf0;  wr_data_rom[ 1552]='h000000f3;
    rd_cycle[ 1553] = 1'b0;  wr_cycle[ 1553] = 1'b1;  addr_rom[ 1553]='h000007e0;  wr_data_rom[ 1553]='h000007ff;
    rd_cycle[ 1554] = 1'b0;  wr_cycle[ 1554] = 1'b1;  addr_rom[ 1554]='h00000180;  wr_data_rom[ 1554]='h00000298;
    rd_cycle[ 1555] = 1'b1;  wr_cycle[ 1555] = 1'b0;  addr_rom[ 1555]='h000004e4;  wr_data_rom[ 1555]='h00000000;
    rd_cycle[ 1556] = 1'b1;  wr_cycle[ 1556] = 1'b0;  addr_rom[ 1556]='h00000aa8;  wr_data_rom[ 1556]='h00000000;
    rd_cycle[ 1557] = 1'b1;  wr_cycle[ 1557] = 1'b0;  addr_rom[ 1557]='h000000e0;  wr_data_rom[ 1557]='h00000000;
    rd_cycle[ 1558] = 1'b0;  wr_cycle[ 1558] = 1'b1;  addr_rom[ 1558]='h00000edc;  wr_data_rom[ 1558]='h000003c1;
    rd_cycle[ 1559] = 1'b1;  wr_cycle[ 1559] = 1'b0;  addr_rom[ 1559]='h00000568;  wr_data_rom[ 1559]='h00000000;
    rd_cycle[ 1560] = 1'b0;  wr_cycle[ 1560] = 1'b1;  addr_rom[ 1560]='h00000b10;  wr_data_rom[ 1560]='h0000029e;
    rd_cycle[ 1561] = 1'b1;  wr_cycle[ 1561] = 1'b0;  addr_rom[ 1561]='h00000544;  wr_data_rom[ 1561]='h00000000;
    rd_cycle[ 1562] = 1'b1;  wr_cycle[ 1562] = 1'b0;  addr_rom[ 1562]='h000003b8;  wr_data_rom[ 1562]='h00000000;
    rd_cycle[ 1563] = 1'b0;  wr_cycle[ 1563] = 1'b1;  addr_rom[ 1563]='h00000014;  wr_data_rom[ 1563]='h00000161;
    rd_cycle[ 1564] = 1'b1;  wr_cycle[ 1564] = 1'b0;  addr_rom[ 1564]='h00000470;  wr_data_rom[ 1564]='h00000000;
    rd_cycle[ 1565] = 1'b0;  wr_cycle[ 1565] = 1'b1;  addr_rom[ 1565]='h00000dc4;  wr_data_rom[ 1565]='h0000064a;
    rd_cycle[ 1566] = 1'b1;  wr_cycle[ 1566] = 1'b0;  addr_rom[ 1566]='h00000208;  wr_data_rom[ 1566]='h00000000;
    rd_cycle[ 1567] = 1'b1;  wr_cycle[ 1567] = 1'b0;  addr_rom[ 1567]='h0000004c;  wr_data_rom[ 1567]='h00000000;
    rd_cycle[ 1568] = 1'b0;  wr_cycle[ 1568] = 1'b1;  addr_rom[ 1568]='h00000060;  wr_data_rom[ 1568]='h000004bf;
    rd_cycle[ 1569] = 1'b1;  wr_cycle[ 1569] = 1'b0;  addr_rom[ 1569]='h000007fc;  wr_data_rom[ 1569]='h00000000;
    rd_cycle[ 1570] = 1'b1;  wr_cycle[ 1570] = 1'b0;  addr_rom[ 1570]='h000005b4;  wr_data_rom[ 1570]='h00000000;
    rd_cycle[ 1571] = 1'b1;  wr_cycle[ 1571] = 1'b0;  addr_rom[ 1571]='h00000ccc;  wr_data_rom[ 1571]='h00000000;
    rd_cycle[ 1572] = 1'b0;  wr_cycle[ 1572] = 1'b1;  addr_rom[ 1572]='h00000d38;  wr_data_rom[ 1572]='h00000a1d;
    rd_cycle[ 1573] = 1'b1;  wr_cycle[ 1573] = 1'b0;  addr_rom[ 1573]='h00000100;  wr_data_rom[ 1573]='h00000000;
    rd_cycle[ 1574] = 1'b1;  wr_cycle[ 1574] = 1'b0;  addr_rom[ 1574]='h00000f44;  wr_data_rom[ 1574]='h00000000;
    rd_cycle[ 1575] = 1'b1;  wr_cycle[ 1575] = 1'b0;  addr_rom[ 1575]='h00000d34;  wr_data_rom[ 1575]='h00000000;
    rd_cycle[ 1576] = 1'b0;  wr_cycle[ 1576] = 1'b1;  addr_rom[ 1576]='h00000cb0;  wr_data_rom[ 1576]='h00000747;
    rd_cycle[ 1577] = 1'b1;  wr_cycle[ 1577] = 1'b0;  addr_rom[ 1577]='h00000c34;  wr_data_rom[ 1577]='h00000000;
    rd_cycle[ 1578] = 1'b1;  wr_cycle[ 1578] = 1'b0;  addr_rom[ 1578]='h00000c34;  wr_data_rom[ 1578]='h00000000;
    rd_cycle[ 1579] = 1'b1;  wr_cycle[ 1579] = 1'b0;  addr_rom[ 1579]='h000008dc;  wr_data_rom[ 1579]='h00000000;
    rd_cycle[ 1580] = 1'b1;  wr_cycle[ 1580] = 1'b0;  addr_rom[ 1580]='h000005c8;  wr_data_rom[ 1580]='h00000000;
    rd_cycle[ 1581] = 1'b1;  wr_cycle[ 1581] = 1'b0;  addr_rom[ 1581]='h000006fc;  wr_data_rom[ 1581]='h00000000;
    rd_cycle[ 1582] = 1'b0;  wr_cycle[ 1582] = 1'b1;  addr_rom[ 1582]='h00000474;  wr_data_rom[ 1582]='h000006ff;
    rd_cycle[ 1583] = 1'b1;  wr_cycle[ 1583] = 1'b0;  addr_rom[ 1583]='h00000a28;  wr_data_rom[ 1583]='h00000000;
    rd_cycle[ 1584] = 1'b1;  wr_cycle[ 1584] = 1'b0;  addr_rom[ 1584]='h000000c4;  wr_data_rom[ 1584]='h00000000;
    rd_cycle[ 1585] = 1'b1;  wr_cycle[ 1585] = 1'b0;  addr_rom[ 1585]='h00000548;  wr_data_rom[ 1585]='h00000000;
    rd_cycle[ 1586] = 1'b1;  wr_cycle[ 1586] = 1'b0;  addr_rom[ 1586]='h000009b4;  wr_data_rom[ 1586]='h00000000;
    rd_cycle[ 1587] = 1'b1;  wr_cycle[ 1587] = 1'b0;  addr_rom[ 1587]='h00000690;  wr_data_rom[ 1587]='h00000000;
    rd_cycle[ 1588] = 1'b0;  wr_cycle[ 1588] = 1'b1;  addr_rom[ 1588]='h000007f0;  wr_data_rom[ 1588]='h00000f7d;
    rd_cycle[ 1589] = 1'b1;  wr_cycle[ 1589] = 1'b0;  addr_rom[ 1589]='h00000a94;  wr_data_rom[ 1589]='h00000000;
    rd_cycle[ 1590] = 1'b0;  wr_cycle[ 1590] = 1'b1;  addr_rom[ 1590]='h00000290;  wr_data_rom[ 1590]='h00000157;
    rd_cycle[ 1591] = 1'b0;  wr_cycle[ 1591] = 1'b1;  addr_rom[ 1591]='h00000a04;  wr_data_rom[ 1591]='h0000011f;
    rd_cycle[ 1592] = 1'b1;  wr_cycle[ 1592] = 1'b0;  addr_rom[ 1592]='h00000708;  wr_data_rom[ 1592]='h00000000;
    rd_cycle[ 1593] = 1'b0;  wr_cycle[ 1593] = 1'b1;  addr_rom[ 1593]='h00000144;  wr_data_rom[ 1593]='h00000606;
    rd_cycle[ 1594] = 1'b1;  wr_cycle[ 1594] = 1'b0;  addr_rom[ 1594]='h00000b90;  wr_data_rom[ 1594]='h00000000;
    rd_cycle[ 1595] = 1'b0;  wr_cycle[ 1595] = 1'b1;  addr_rom[ 1595]='h0000032c;  wr_data_rom[ 1595]='h00000a3e;
    rd_cycle[ 1596] = 1'b0;  wr_cycle[ 1596] = 1'b1;  addr_rom[ 1596]='h000005d0;  wr_data_rom[ 1596]='h00000972;
    rd_cycle[ 1597] = 1'b0;  wr_cycle[ 1597] = 1'b1;  addr_rom[ 1597]='h000001e0;  wr_data_rom[ 1597]='h00000c8d;
    rd_cycle[ 1598] = 1'b0;  wr_cycle[ 1598] = 1'b1;  addr_rom[ 1598]='h00000a20;  wr_data_rom[ 1598]='h00000bbc;
    rd_cycle[ 1599] = 1'b1;  wr_cycle[ 1599] = 1'b0;  addr_rom[ 1599]='h00000b28;  wr_data_rom[ 1599]='h00000000;
    rd_cycle[ 1600] = 1'b1;  wr_cycle[ 1600] = 1'b0;  addr_rom[ 1600]='h00000798;  wr_data_rom[ 1600]='h00000000;
    rd_cycle[ 1601] = 1'b0;  wr_cycle[ 1601] = 1'b1;  addr_rom[ 1601]='h00000d78;  wr_data_rom[ 1601]='h00000752;
    rd_cycle[ 1602] = 1'b1;  wr_cycle[ 1602] = 1'b0;  addr_rom[ 1602]='h00000430;  wr_data_rom[ 1602]='h00000000;
    rd_cycle[ 1603] = 1'b0;  wr_cycle[ 1603] = 1'b1;  addr_rom[ 1603]='h00000e3c;  wr_data_rom[ 1603]='h00000823;
    rd_cycle[ 1604] = 1'b0;  wr_cycle[ 1604] = 1'b1;  addr_rom[ 1604]='h00000538;  wr_data_rom[ 1604]='h00000ed2;
    rd_cycle[ 1605] = 1'b0;  wr_cycle[ 1605] = 1'b1;  addr_rom[ 1605]='h00000f58;  wr_data_rom[ 1605]='h00000802;
    rd_cycle[ 1606] = 1'b0;  wr_cycle[ 1606] = 1'b1;  addr_rom[ 1606]='h00000a5c;  wr_data_rom[ 1606]='h00000d04;
    rd_cycle[ 1607] = 1'b1;  wr_cycle[ 1607] = 1'b0;  addr_rom[ 1607]='h00000398;  wr_data_rom[ 1607]='h00000000;
    rd_cycle[ 1608] = 1'b0;  wr_cycle[ 1608] = 1'b1;  addr_rom[ 1608]='h000008a4;  wr_data_rom[ 1608]='h00000ed9;
    rd_cycle[ 1609] = 1'b1;  wr_cycle[ 1609] = 1'b0;  addr_rom[ 1609]='h00000264;  wr_data_rom[ 1609]='h00000000;
    rd_cycle[ 1610] = 1'b1;  wr_cycle[ 1610] = 1'b0;  addr_rom[ 1610]='h00000860;  wr_data_rom[ 1610]='h00000000;
    rd_cycle[ 1611] = 1'b1;  wr_cycle[ 1611] = 1'b0;  addr_rom[ 1611]='h00000e40;  wr_data_rom[ 1611]='h00000000;
    rd_cycle[ 1612] = 1'b1;  wr_cycle[ 1612] = 1'b0;  addr_rom[ 1612]='h00000d8c;  wr_data_rom[ 1612]='h00000000;
    rd_cycle[ 1613] = 1'b0;  wr_cycle[ 1613] = 1'b1;  addr_rom[ 1613]='h00000e54;  wr_data_rom[ 1613]='h00000515;
    rd_cycle[ 1614] = 1'b1;  wr_cycle[ 1614] = 1'b0;  addr_rom[ 1614]='h000009d0;  wr_data_rom[ 1614]='h00000000;
    rd_cycle[ 1615] = 1'b1;  wr_cycle[ 1615] = 1'b0;  addr_rom[ 1615]='h00000378;  wr_data_rom[ 1615]='h00000000;
    rd_cycle[ 1616] = 1'b1;  wr_cycle[ 1616] = 1'b0;  addr_rom[ 1616]='h00000f6c;  wr_data_rom[ 1616]='h00000000;
    rd_cycle[ 1617] = 1'b1;  wr_cycle[ 1617] = 1'b0;  addr_rom[ 1617]='h000008b4;  wr_data_rom[ 1617]='h00000000;
    rd_cycle[ 1618] = 1'b1;  wr_cycle[ 1618] = 1'b0;  addr_rom[ 1618]='h00000718;  wr_data_rom[ 1618]='h00000000;
    rd_cycle[ 1619] = 1'b0;  wr_cycle[ 1619] = 1'b1;  addr_rom[ 1619]='h000009c0;  wr_data_rom[ 1619]='h000002d5;
    rd_cycle[ 1620] = 1'b1;  wr_cycle[ 1620] = 1'b0;  addr_rom[ 1620]='h00000da4;  wr_data_rom[ 1620]='h00000000;
    rd_cycle[ 1621] = 1'b1;  wr_cycle[ 1621] = 1'b0;  addr_rom[ 1621]='h00000f30;  wr_data_rom[ 1621]='h00000000;
    rd_cycle[ 1622] = 1'b1;  wr_cycle[ 1622] = 1'b0;  addr_rom[ 1622]='h000007e8;  wr_data_rom[ 1622]='h00000000;
    rd_cycle[ 1623] = 1'b0;  wr_cycle[ 1623] = 1'b1;  addr_rom[ 1623]='h0000067c;  wr_data_rom[ 1623]='h00000910;
    rd_cycle[ 1624] = 1'b1;  wr_cycle[ 1624] = 1'b0;  addr_rom[ 1624]='h000007cc;  wr_data_rom[ 1624]='h00000000;
    rd_cycle[ 1625] = 1'b1;  wr_cycle[ 1625] = 1'b0;  addr_rom[ 1625]='h00000170;  wr_data_rom[ 1625]='h00000000;
    rd_cycle[ 1626] = 1'b1;  wr_cycle[ 1626] = 1'b0;  addr_rom[ 1626]='h00000aa4;  wr_data_rom[ 1626]='h00000000;
    rd_cycle[ 1627] = 1'b0;  wr_cycle[ 1627] = 1'b1;  addr_rom[ 1627]='h000008b4;  wr_data_rom[ 1627]='h00000185;
    rd_cycle[ 1628] = 1'b1;  wr_cycle[ 1628] = 1'b0;  addr_rom[ 1628]='h00000a4c;  wr_data_rom[ 1628]='h00000000;
    rd_cycle[ 1629] = 1'b0;  wr_cycle[ 1629] = 1'b1;  addr_rom[ 1629]='h0000025c;  wr_data_rom[ 1629]='h00000ea6;
    rd_cycle[ 1630] = 1'b1;  wr_cycle[ 1630] = 1'b0;  addr_rom[ 1630]='h00000560;  wr_data_rom[ 1630]='h00000000;
    rd_cycle[ 1631] = 1'b0;  wr_cycle[ 1631] = 1'b1;  addr_rom[ 1631]='h00000db8;  wr_data_rom[ 1631]='h00000d36;
    rd_cycle[ 1632] = 1'b1;  wr_cycle[ 1632] = 1'b0;  addr_rom[ 1632]='h00000254;  wr_data_rom[ 1632]='h00000000;
    rd_cycle[ 1633] = 1'b1;  wr_cycle[ 1633] = 1'b0;  addr_rom[ 1633]='h00000dac;  wr_data_rom[ 1633]='h00000000;
    rd_cycle[ 1634] = 1'b1;  wr_cycle[ 1634] = 1'b0;  addr_rom[ 1634]='h00000ae4;  wr_data_rom[ 1634]='h00000000;
    rd_cycle[ 1635] = 1'b0;  wr_cycle[ 1635] = 1'b1;  addr_rom[ 1635]='h000004a4;  wr_data_rom[ 1635]='h000003b3;
    rd_cycle[ 1636] = 1'b0;  wr_cycle[ 1636] = 1'b1;  addr_rom[ 1636]='h00000810;  wr_data_rom[ 1636]='h00000877;
    rd_cycle[ 1637] = 1'b1;  wr_cycle[ 1637] = 1'b0;  addr_rom[ 1637]='h00000814;  wr_data_rom[ 1637]='h00000000;
    rd_cycle[ 1638] = 1'b1;  wr_cycle[ 1638] = 1'b0;  addr_rom[ 1638]='h00000170;  wr_data_rom[ 1638]='h00000000;
    rd_cycle[ 1639] = 1'b0;  wr_cycle[ 1639] = 1'b1;  addr_rom[ 1639]='h00000f34;  wr_data_rom[ 1639]='h00000f6f;
    rd_cycle[ 1640] = 1'b0;  wr_cycle[ 1640] = 1'b1;  addr_rom[ 1640]='h000006cc;  wr_data_rom[ 1640]='h000003de;
    rd_cycle[ 1641] = 1'b1;  wr_cycle[ 1641] = 1'b0;  addr_rom[ 1641]='h00000ce0;  wr_data_rom[ 1641]='h00000000;
    rd_cycle[ 1642] = 1'b0;  wr_cycle[ 1642] = 1'b1;  addr_rom[ 1642]='h0000014c;  wr_data_rom[ 1642]='h0000090b;
    rd_cycle[ 1643] = 1'b1;  wr_cycle[ 1643] = 1'b0;  addr_rom[ 1643]='h000008b8;  wr_data_rom[ 1643]='h00000000;
    rd_cycle[ 1644] = 1'b1;  wr_cycle[ 1644] = 1'b0;  addr_rom[ 1644]='h00000e78;  wr_data_rom[ 1644]='h00000000;
    rd_cycle[ 1645] = 1'b0;  wr_cycle[ 1645] = 1'b1;  addr_rom[ 1645]='h00000260;  wr_data_rom[ 1645]='h00000c82;
    rd_cycle[ 1646] = 1'b0;  wr_cycle[ 1646] = 1'b1;  addr_rom[ 1646]='h00000f4c;  wr_data_rom[ 1646]='h0000067d;
    rd_cycle[ 1647] = 1'b1;  wr_cycle[ 1647] = 1'b0;  addr_rom[ 1647]='h00000464;  wr_data_rom[ 1647]='h00000000;
    rd_cycle[ 1648] = 1'b0;  wr_cycle[ 1648] = 1'b1;  addr_rom[ 1648]='h00000b8c;  wr_data_rom[ 1648]='h0000002c;
    rd_cycle[ 1649] = 1'b1;  wr_cycle[ 1649] = 1'b0;  addr_rom[ 1649]='h00000640;  wr_data_rom[ 1649]='h00000000;
    rd_cycle[ 1650] = 1'b0;  wr_cycle[ 1650] = 1'b1;  addr_rom[ 1650]='h00000be0;  wr_data_rom[ 1650]='h00000a31;
    rd_cycle[ 1651] = 1'b0;  wr_cycle[ 1651] = 1'b1;  addr_rom[ 1651]='h000000d4;  wr_data_rom[ 1651]='h00000e32;
    rd_cycle[ 1652] = 1'b0;  wr_cycle[ 1652] = 1'b1;  addr_rom[ 1652]='h00000b04;  wr_data_rom[ 1652]='h00000a00;
    rd_cycle[ 1653] = 1'b0;  wr_cycle[ 1653] = 1'b1;  addr_rom[ 1653]='h00000680;  wr_data_rom[ 1653]='h00000401;
    rd_cycle[ 1654] = 1'b1;  wr_cycle[ 1654] = 1'b0;  addr_rom[ 1654]='h00000068;  wr_data_rom[ 1654]='h00000000;
    rd_cycle[ 1655] = 1'b1;  wr_cycle[ 1655] = 1'b0;  addr_rom[ 1655]='h00000b1c;  wr_data_rom[ 1655]='h00000000;
    rd_cycle[ 1656] = 1'b1;  wr_cycle[ 1656] = 1'b0;  addr_rom[ 1656]='h000001dc;  wr_data_rom[ 1656]='h00000000;
    rd_cycle[ 1657] = 1'b1;  wr_cycle[ 1657] = 1'b0;  addr_rom[ 1657]='h00000d68;  wr_data_rom[ 1657]='h00000000;
    rd_cycle[ 1658] = 1'b1;  wr_cycle[ 1658] = 1'b0;  addr_rom[ 1658]='h00000910;  wr_data_rom[ 1658]='h00000000;
    rd_cycle[ 1659] = 1'b0;  wr_cycle[ 1659] = 1'b1;  addr_rom[ 1659]='h000006f4;  wr_data_rom[ 1659]='h0000070e;
    rd_cycle[ 1660] = 1'b0;  wr_cycle[ 1660] = 1'b1;  addr_rom[ 1660]='h000006d4;  wr_data_rom[ 1660]='h0000056b;
    rd_cycle[ 1661] = 1'b0;  wr_cycle[ 1661] = 1'b1;  addr_rom[ 1661]='h000009e8;  wr_data_rom[ 1661]='h0000053b;
    rd_cycle[ 1662] = 1'b1;  wr_cycle[ 1662] = 1'b0;  addr_rom[ 1662]='h00000290;  wr_data_rom[ 1662]='h00000000;
    rd_cycle[ 1663] = 1'b0;  wr_cycle[ 1663] = 1'b1;  addr_rom[ 1663]='h00000640;  wr_data_rom[ 1663]='h00000827;
    rd_cycle[ 1664] = 1'b1;  wr_cycle[ 1664] = 1'b0;  addr_rom[ 1664]='h00000474;  wr_data_rom[ 1664]='h00000000;
    rd_cycle[ 1665] = 1'b1;  wr_cycle[ 1665] = 1'b0;  addr_rom[ 1665]='h00000494;  wr_data_rom[ 1665]='h00000000;
    rd_cycle[ 1666] = 1'b1;  wr_cycle[ 1666] = 1'b0;  addr_rom[ 1666]='h00000df8;  wr_data_rom[ 1666]='h00000000;
    rd_cycle[ 1667] = 1'b0;  wr_cycle[ 1667] = 1'b1;  addr_rom[ 1667]='h00000100;  wr_data_rom[ 1667]='h00000ee8;
    rd_cycle[ 1668] = 1'b0;  wr_cycle[ 1668] = 1'b1;  addr_rom[ 1668]='h000004a8;  wr_data_rom[ 1668]='h0000097e;
    rd_cycle[ 1669] = 1'b0;  wr_cycle[ 1669] = 1'b1;  addr_rom[ 1669]='h00000654;  wr_data_rom[ 1669]='h00000f4c;
    rd_cycle[ 1670] = 1'b0;  wr_cycle[ 1670] = 1'b1;  addr_rom[ 1670]='h00000c4c;  wr_data_rom[ 1670]='h00000714;
    rd_cycle[ 1671] = 1'b0;  wr_cycle[ 1671] = 1'b1;  addr_rom[ 1671]='h0000093c;  wr_data_rom[ 1671]='h00000ded;
    rd_cycle[ 1672] = 1'b0;  wr_cycle[ 1672] = 1'b1;  addr_rom[ 1672]='h000005ec;  wr_data_rom[ 1672]='h00000718;
    rd_cycle[ 1673] = 1'b0;  wr_cycle[ 1673] = 1'b1;  addr_rom[ 1673]='h00000d5c;  wr_data_rom[ 1673]='h0000007f;
    rd_cycle[ 1674] = 1'b0;  wr_cycle[ 1674] = 1'b1;  addr_rom[ 1674]='h00000e28;  wr_data_rom[ 1674]='h0000007b;
    rd_cycle[ 1675] = 1'b1;  wr_cycle[ 1675] = 1'b0;  addr_rom[ 1675]='h000007a4;  wr_data_rom[ 1675]='h00000000;
    rd_cycle[ 1676] = 1'b0;  wr_cycle[ 1676] = 1'b1;  addr_rom[ 1676]='h00000818;  wr_data_rom[ 1676]='h00000e52;
    rd_cycle[ 1677] = 1'b1;  wr_cycle[ 1677] = 1'b0;  addr_rom[ 1677]='h000007f0;  wr_data_rom[ 1677]='h00000000;
    rd_cycle[ 1678] = 1'b1;  wr_cycle[ 1678] = 1'b0;  addr_rom[ 1678]='h00000ae0;  wr_data_rom[ 1678]='h00000000;
    rd_cycle[ 1679] = 1'b0;  wr_cycle[ 1679] = 1'b1;  addr_rom[ 1679]='h000004cc;  wr_data_rom[ 1679]='h0000068f;
    rd_cycle[ 1680] = 1'b0;  wr_cycle[ 1680] = 1'b1;  addr_rom[ 1680]='h00000f6c;  wr_data_rom[ 1680]='h00000bc0;
    rd_cycle[ 1681] = 1'b1;  wr_cycle[ 1681] = 1'b0;  addr_rom[ 1681]='h00000cc0;  wr_data_rom[ 1681]='h00000000;
    rd_cycle[ 1682] = 1'b1;  wr_cycle[ 1682] = 1'b0;  addr_rom[ 1682]='h000008dc;  wr_data_rom[ 1682]='h00000000;
    rd_cycle[ 1683] = 1'b0;  wr_cycle[ 1683] = 1'b1;  addr_rom[ 1683]='h00000630;  wr_data_rom[ 1683]='h00000066;
    rd_cycle[ 1684] = 1'b1;  wr_cycle[ 1684] = 1'b0;  addr_rom[ 1684]='h00000b2c;  wr_data_rom[ 1684]='h00000000;
    rd_cycle[ 1685] = 1'b0;  wr_cycle[ 1685] = 1'b1;  addr_rom[ 1685]='h000003d4;  wr_data_rom[ 1685]='h000008b2;
    rd_cycle[ 1686] = 1'b1;  wr_cycle[ 1686] = 1'b0;  addr_rom[ 1686]='h000006c4;  wr_data_rom[ 1686]='h00000000;
    rd_cycle[ 1687] = 1'b1;  wr_cycle[ 1687] = 1'b0;  addr_rom[ 1687]='h00000dbc;  wr_data_rom[ 1687]='h00000000;
    rd_cycle[ 1688] = 1'b1;  wr_cycle[ 1688] = 1'b0;  addr_rom[ 1688]='h00000620;  wr_data_rom[ 1688]='h00000000;
    rd_cycle[ 1689] = 1'b0;  wr_cycle[ 1689] = 1'b1;  addr_rom[ 1689]='h000005bc;  wr_data_rom[ 1689]='h0000008a;
    rd_cycle[ 1690] = 1'b0;  wr_cycle[ 1690] = 1'b1;  addr_rom[ 1690]='h00000020;  wr_data_rom[ 1690]='h00000519;
    rd_cycle[ 1691] = 1'b1;  wr_cycle[ 1691] = 1'b0;  addr_rom[ 1691]='h00000298;  wr_data_rom[ 1691]='h00000000;
    rd_cycle[ 1692] = 1'b1;  wr_cycle[ 1692] = 1'b0;  addr_rom[ 1692]='h000005f8;  wr_data_rom[ 1692]='h00000000;
    rd_cycle[ 1693] = 1'b1;  wr_cycle[ 1693] = 1'b0;  addr_rom[ 1693]='h00000138;  wr_data_rom[ 1693]='h00000000;
    rd_cycle[ 1694] = 1'b1;  wr_cycle[ 1694] = 1'b0;  addr_rom[ 1694]='h00000bd4;  wr_data_rom[ 1694]='h00000000;
    rd_cycle[ 1695] = 1'b0;  wr_cycle[ 1695] = 1'b1;  addr_rom[ 1695]='h00000874;  wr_data_rom[ 1695]='h0000052d;
    rd_cycle[ 1696] = 1'b0;  wr_cycle[ 1696] = 1'b1;  addr_rom[ 1696]='h00000140;  wr_data_rom[ 1696]='h00000b0b;
    rd_cycle[ 1697] = 1'b1;  wr_cycle[ 1697] = 1'b0;  addr_rom[ 1697]='h00000bcc;  wr_data_rom[ 1697]='h00000000;
    rd_cycle[ 1698] = 1'b0;  wr_cycle[ 1698] = 1'b1;  addr_rom[ 1698]='h00000e74;  wr_data_rom[ 1698]='h000007e5;
    rd_cycle[ 1699] = 1'b0;  wr_cycle[ 1699] = 1'b1;  addr_rom[ 1699]='h00000f48;  wr_data_rom[ 1699]='h000001c0;
    rd_cycle[ 1700] = 1'b1;  wr_cycle[ 1700] = 1'b0;  addr_rom[ 1700]='h0000057c;  wr_data_rom[ 1700]='h00000000;
    rd_cycle[ 1701] = 1'b0;  wr_cycle[ 1701] = 1'b1;  addr_rom[ 1701]='h000004c8;  wr_data_rom[ 1701]='h00000959;
    rd_cycle[ 1702] = 1'b0;  wr_cycle[ 1702] = 1'b1;  addr_rom[ 1702]='h00000750;  wr_data_rom[ 1702]='h00000571;
    rd_cycle[ 1703] = 1'b1;  wr_cycle[ 1703] = 1'b0;  addr_rom[ 1703]='h00000084;  wr_data_rom[ 1703]='h00000000;
    rd_cycle[ 1704] = 1'b0;  wr_cycle[ 1704] = 1'b1;  addr_rom[ 1704]='h00000c84;  wr_data_rom[ 1704]='h000003e8;
    rd_cycle[ 1705] = 1'b1;  wr_cycle[ 1705] = 1'b0;  addr_rom[ 1705]='h000006f4;  wr_data_rom[ 1705]='h00000000;
    rd_cycle[ 1706] = 1'b1;  wr_cycle[ 1706] = 1'b0;  addr_rom[ 1706]='h00000ae0;  wr_data_rom[ 1706]='h00000000;
    rd_cycle[ 1707] = 1'b0;  wr_cycle[ 1707] = 1'b1;  addr_rom[ 1707]='h00000c50;  wr_data_rom[ 1707]='h00000b3c;
    rd_cycle[ 1708] = 1'b0;  wr_cycle[ 1708] = 1'b1;  addr_rom[ 1708]='h00000de4;  wr_data_rom[ 1708]='h0000006f;
    rd_cycle[ 1709] = 1'b0;  wr_cycle[ 1709] = 1'b1;  addr_rom[ 1709]='h000003ac;  wr_data_rom[ 1709]='h00000eba;
    rd_cycle[ 1710] = 1'b0;  wr_cycle[ 1710] = 1'b1;  addr_rom[ 1710]='h000008b4;  wr_data_rom[ 1710]='h00000eec;
    rd_cycle[ 1711] = 1'b0;  wr_cycle[ 1711] = 1'b1;  addr_rom[ 1711]='h00000f50;  wr_data_rom[ 1711]='h00000640;
    rd_cycle[ 1712] = 1'b1;  wr_cycle[ 1712] = 1'b0;  addr_rom[ 1712]='h000000e0;  wr_data_rom[ 1712]='h00000000;
    rd_cycle[ 1713] = 1'b1;  wr_cycle[ 1713] = 1'b0;  addr_rom[ 1713]='h000000d8;  wr_data_rom[ 1713]='h00000000;
    rd_cycle[ 1714] = 1'b0;  wr_cycle[ 1714] = 1'b1;  addr_rom[ 1714]='h00000b58;  wr_data_rom[ 1714]='h0000010d;
    rd_cycle[ 1715] = 1'b1;  wr_cycle[ 1715] = 1'b0;  addr_rom[ 1715]='h00000030;  wr_data_rom[ 1715]='h00000000;
    rd_cycle[ 1716] = 1'b1;  wr_cycle[ 1716] = 1'b0;  addr_rom[ 1716]='h00000bb0;  wr_data_rom[ 1716]='h00000000;
    rd_cycle[ 1717] = 1'b1;  wr_cycle[ 1717] = 1'b0;  addr_rom[ 1717]='h000007fc;  wr_data_rom[ 1717]='h00000000;
    rd_cycle[ 1718] = 1'b0;  wr_cycle[ 1718] = 1'b1;  addr_rom[ 1718]='h00000b30;  wr_data_rom[ 1718]='h0000024e;
    rd_cycle[ 1719] = 1'b1;  wr_cycle[ 1719] = 1'b0;  addr_rom[ 1719]='h00000d7c;  wr_data_rom[ 1719]='h00000000;
    rd_cycle[ 1720] = 1'b0;  wr_cycle[ 1720] = 1'b1;  addr_rom[ 1720]='h00000d9c;  wr_data_rom[ 1720]='h00000d26;
    rd_cycle[ 1721] = 1'b1;  wr_cycle[ 1721] = 1'b0;  addr_rom[ 1721]='h00000f94;  wr_data_rom[ 1721]='h00000000;
    rd_cycle[ 1722] = 1'b1;  wr_cycle[ 1722] = 1'b0;  addr_rom[ 1722]='h0000047c;  wr_data_rom[ 1722]='h00000000;
    rd_cycle[ 1723] = 1'b0;  wr_cycle[ 1723] = 1'b1;  addr_rom[ 1723]='h00000f4c;  wr_data_rom[ 1723]='h00000d2e;
    rd_cycle[ 1724] = 1'b1;  wr_cycle[ 1724] = 1'b0;  addr_rom[ 1724]='h00000d00;  wr_data_rom[ 1724]='h00000000;
    rd_cycle[ 1725] = 1'b1;  wr_cycle[ 1725] = 1'b0;  addr_rom[ 1725]='h00000acc;  wr_data_rom[ 1725]='h00000000;
    rd_cycle[ 1726] = 1'b1;  wr_cycle[ 1726] = 1'b0;  addr_rom[ 1726]='h00000d74;  wr_data_rom[ 1726]='h00000000;
    rd_cycle[ 1727] = 1'b1;  wr_cycle[ 1727] = 1'b0;  addr_rom[ 1727]='h00000a40;  wr_data_rom[ 1727]='h00000000;
    rd_cycle[ 1728] = 1'b0;  wr_cycle[ 1728] = 1'b1;  addr_rom[ 1728]='h000003ac;  wr_data_rom[ 1728]='h00000b4a;
    rd_cycle[ 1729] = 1'b0;  wr_cycle[ 1729] = 1'b1;  addr_rom[ 1729]='h00000640;  wr_data_rom[ 1729]='h0000070c;
    rd_cycle[ 1730] = 1'b0;  wr_cycle[ 1730] = 1'b1;  addr_rom[ 1730]='h000004fc;  wr_data_rom[ 1730]='h00000f1f;
    rd_cycle[ 1731] = 1'b1;  wr_cycle[ 1731] = 1'b0;  addr_rom[ 1731]='h00000500;  wr_data_rom[ 1731]='h00000000;
    rd_cycle[ 1732] = 1'b0;  wr_cycle[ 1732] = 1'b1;  addr_rom[ 1732]='h00000610;  wr_data_rom[ 1732]='h000006c8;
    rd_cycle[ 1733] = 1'b1;  wr_cycle[ 1733] = 1'b0;  addr_rom[ 1733]='h00000e54;  wr_data_rom[ 1733]='h00000000;
    rd_cycle[ 1734] = 1'b0;  wr_cycle[ 1734] = 1'b1;  addr_rom[ 1734]='h00000ce4;  wr_data_rom[ 1734]='h000008f9;
    rd_cycle[ 1735] = 1'b0;  wr_cycle[ 1735] = 1'b1;  addr_rom[ 1735]='h00000960;  wr_data_rom[ 1735]='h00000910;
    rd_cycle[ 1736] = 1'b1;  wr_cycle[ 1736] = 1'b0;  addr_rom[ 1736]='h00000e00;  wr_data_rom[ 1736]='h00000000;
    rd_cycle[ 1737] = 1'b1;  wr_cycle[ 1737] = 1'b0;  addr_rom[ 1737]='h00000be8;  wr_data_rom[ 1737]='h00000000;
    rd_cycle[ 1738] = 1'b1;  wr_cycle[ 1738] = 1'b0;  addr_rom[ 1738]='h0000070c;  wr_data_rom[ 1738]='h00000000;
    rd_cycle[ 1739] = 1'b0;  wr_cycle[ 1739] = 1'b1;  addr_rom[ 1739]='h00000680;  wr_data_rom[ 1739]='h00000899;
    rd_cycle[ 1740] = 1'b0;  wr_cycle[ 1740] = 1'b1;  addr_rom[ 1740]='h00000254;  wr_data_rom[ 1740]='h00000057;
    rd_cycle[ 1741] = 1'b1;  wr_cycle[ 1741] = 1'b0;  addr_rom[ 1741]='h000009bc;  wr_data_rom[ 1741]='h00000000;
    rd_cycle[ 1742] = 1'b0;  wr_cycle[ 1742] = 1'b1;  addr_rom[ 1742]='h00000a5c;  wr_data_rom[ 1742]='h00000237;
    rd_cycle[ 1743] = 1'b1;  wr_cycle[ 1743] = 1'b0;  addr_rom[ 1743]='h000001b8;  wr_data_rom[ 1743]='h00000000;
    rd_cycle[ 1744] = 1'b1;  wr_cycle[ 1744] = 1'b0;  addr_rom[ 1744]='h00000b30;  wr_data_rom[ 1744]='h00000000;
    rd_cycle[ 1745] = 1'b1;  wr_cycle[ 1745] = 1'b0;  addr_rom[ 1745]='h00000254;  wr_data_rom[ 1745]='h00000000;
    rd_cycle[ 1746] = 1'b0;  wr_cycle[ 1746] = 1'b1;  addr_rom[ 1746]='h0000016c;  wr_data_rom[ 1746]='h00000c88;
    rd_cycle[ 1747] = 1'b1;  wr_cycle[ 1747] = 1'b0;  addr_rom[ 1747]='h00000190;  wr_data_rom[ 1747]='h00000000;
    rd_cycle[ 1748] = 1'b1;  wr_cycle[ 1748] = 1'b0;  addr_rom[ 1748]='h000000f4;  wr_data_rom[ 1748]='h00000000;
    rd_cycle[ 1749] = 1'b1;  wr_cycle[ 1749] = 1'b0;  addr_rom[ 1749]='h00000714;  wr_data_rom[ 1749]='h00000000;
    rd_cycle[ 1750] = 1'b0;  wr_cycle[ 1750] = 1'b1;  addr_rom[ 1750]='h000005cc;  wr_data_rom[ 1750]='h000005cd;
    rd_cycle[ 1751] = 1'b0;  wr_cycle[ 1751] = 1'b1;  addr_rom[ 1751]='h000003e8;  wr_data_rom[ 1751]='h00000578;
    rd_cycle[ 1752] = 1'b1;  wr_cycle[ 1752] = 1'b0;  addr_rom[ 1752]='h000001ec;  wr_data_rom[ 1752]='h00000000;
    rd_cycle[ 1753] = 1'b1;  wr_cycle[ 1753] = 1'b0;  addr_rom[ 1753]='h00000410;  wr_data_rom[ 1753]='h00000000;
    rd_cycle[ 1754] = 1'b0;  wr_cycle[ 1754] = 1'b1;  addr_rom[ 1754]='h00000d8c;  wr_data_rom[ 1754]='h0000008e;
    rd_cycle[ 1755] = 1'b1;  wr_cycle[ 1755] = 1'b0;  addr_rom[ 1755]='h000000f8;  wr_data_rom[ 1755]='h00000000;
    rd_cycle[ 1756] = 1'b0;  wr_cycle[ 1756] = 1'b1;  addr_rom[ 1756]='h000002dc;  wr_data_rom[ 1756]='h0000099a;
    rd_cycle[ 1757] = 1'b0;  wr_cycle[ 1757] = 1'b1;  addr_rom[ 1757]='h00000048;  wr_data_rom[ 1757]='h0000052d;
    rd_cycle[ 1758] = 1'b0;  wr_cycle[ 1758] = 1'b1;  addr_rom[ 1758]='h00000304;  wr_data_rom[ 1758]='h0000061f;
    rd_cycle[ 1759] = 1'b1;  wr_cycle[ 1759] = 1'b0;  addr_rom[ 1759]='h00000eec;  wr_data_rom[ 1759]='h00000000;
    rd_cycle[ 1760] = 1'b1;  wr_cycle[ 1760] = 1'b0;  addr_rom[ 1760]='h00000460;  wr_data_rom[ 1760]='h00000000;
    rd_cycle[ 1761] = 1'b0;  wr_cycle[ 1761] = 1'b1;  addr_rom[ 1761]='h00000198;  wr_data_rom[ 1761]='h0000071b;
    rd_cycle[ 1762] = 1'b0;  wr_cycle[ 1762] = 1'b1;  addr_rom[ 1762]='h00000584;  wr_data_rom[ 1762]='h00000add;
    rd_cycle[ 1763] = 1'b1;  wr_cycle[ 1763] = 1'b0;  addr_rom[ 1763]='h00000d40;  wr_data_rom[ 1763]='h00000000;
    rd_cycle[ 1764] = 1'b1;  wr_cycle[ 1764] = 1'b0;  addr_rom[ 1764]='h00000ed0;  wr_data_rom[ 1764]='h00000000;
    rd_cycle[ 1765] = 1'b1;  wr_cycle[ 1765] = 1'b0;  addr_rom[ 1765]='h000001e4;  wr_data_rom[ 1765]='h00000000;
    rd_cycle[ 1766] = 1'b0;  wr_cycle[ 1766] = 1'b1;  addr_rom[ 1766]='h000003bc;  wr_data_rom[ 1766]='h0000038d;
    rd_cycle[ 1767] = 1'b1;  wr_cycle[ 1767] = 1'b0;  addr_rom[ 1767]='h000001f8;  wr_data_rom[ 1767]='h00000000;
    rd_cycle[ 1768] = 1'b1;  wr_cycle[ 1768] = 1'b0;  addr_rom[ 1768]='h00000810;  wr_data_rom[ 1768]='h00000000;
    rd_cycle[ 1769] = 1'b1;  wr_cycle[ 1769] = 1'b0;  addr_rom[ 1769]='h00000824;  wr_data_rom[ 1769]='h00000000;
    rd_cycle[ 1770] = 1'b1;  wr_cycle[ 1770] = 1'b0;  addr_rom[ 1770]='h00000738;  wr_data_rom[ 1770]='h00000000;
    rd_cycle[ 1771] = 1'b1;  wr_cycle[ 1771] = 1'b0;  addr_rom[ 1771]='h00000d08;  wr_data_rom[ 1771]='h00000000;
    rd_cycle[ 1772] = 1'b1;  wr_cycle[ 1772] = 1'b0;  addr_rom[ 1772]='h00000ce4;  wr_data_rom[ 1772]='h00000000;
    rd_cycle[ 1773] = 1'b0;  wr_cycle[ 1773] = 1'b1;  addr_rom[ 1773]='h00000294;  wr_data_rom[ 1773]='h00000835;
    rd_cycle[ 1774] = 1'b1;  wr_cycle[ 1774] = 1'b0;  addr_rom[ 1774]='h00000ac8;  wr_data_rom[ 1774]='h00000000;
    rd_cycle[ 1775] = 1'b1;  wr_cycle[ 1775] = 1'b0;  addr_rom[ 1775]='h000009d0;  wr_data_rom[ 1775]='h00000000;
    rd_cycle[ 1776] = 1'b1;  wr_cycle[ 1776] = 1'b0;  addr_rom[ 1776]='h00000848;  wr_data_rom[ 1776]='h00000000;
    rd_cycle[ 1777] = 1'b0;  wr_cycle[ 1777] = 1'b1;  addr_rom[ 1777]='h00000abc;  wr_data_rom[ 1777]='h000004be;
    rd_cycle[ 1778] = 1'b1;  wr_cycle[ 1778] = 1'b0;  addr_rom[ 1778]='h00000d04;  wr_data_rom[ 1778]='h00000000;
    rd_cycle[ 1779] = 1'b1;  wr_cycle[ 1779] = 1'b0;  addr_rom[ 1779]='h00000078;  wr_data_rom[ 1779]='h00000000;
    rd_cycle[ 1780] = 1'b1;  wr_cycle[ 1780] = 1'b0;  addr_rom[ 1780]='h00000ec4;  wr_data_rom[ 1780]='h00000000;
    rd_cycle[ 1781] = 1'b1;  wr_cycle[ 1781] = 1'b0;  addr_rom[ 1781]='h00000174;  wr_data_rom[ 1781]='h00000000;
    rd_cycle[ 1782] = 1'b1;  wr_cycle[ 1782] = 1'b0;  addr_rom[ 1782]='h00000370;  wr_data_rom[ 1782]='h00000000;
    rd_cycle[ 1783] = 1'b0;  wr_cycle[ 1783] = 1'b1;  addr_rom[ 1783]='h000005c8;  wr_data_rom[ 1783]='h00000147;
    rd_cycle[ 1784] = 1'b0;  wr_cycle[ 1784] = 1'b1;  addr_rom[ 1784]='h00000140;  wr_data_rom[ 1784]='h0000094c;
    rd_cycle[ 1785] = 1'b1;  wr_cycle[ 1785] = 1'b0;  addr_rom[ 1785]='h00000e40;  wr_data_rom[ 1785]='h00000000;
    rd_cycle[ 1786] = 1'b1;  wr_cycle[ 1786] = 1'b0;  addr_rom[ 1786]='h000001a8;  wr_data_rom[ 1786]='h00000000;
    rd_cycle[ 1787] = 1'b1;  wr_cycle[ 1787] = 1'b0;  addr_rom[ 1787]='h00000c28;  wr_data_rom[ 1787]='h00000000;
    rd_cycle[ 1788] = 1'b1;  wr_cycle[ 1788] = 1'b0;  addr_rom[ 1788]='h00000324;  wr_data_rom[ 1788]='h00000000;
    rd_cycle[ 1789] = 1'b1;  wr_cycle[ 1789] = 1'b0;  addr_rom[ 1789]='h000007cc;  wr_data_rom[ 1789]='h00000000;
    rd_cycle[ 1790] = 1'b1;  wr_cycle[ 1790] = 1'b0;  addr_rom[ 1790]='h00000624;  wr_data_rom[ 1790]='h00000000;
    rd_cycle[ 1791] = 1'b0;  wr_cycle[ 1791] = 1'b1;  addr_rom[ 1791]='h000002e0;  wr_data_rom[ 1791]='h000009db;
    rd_cycle[ 1792] = 1'b1;  wr_cycle[ 1792] = 1'b0;  addr_rom[ 1792]='h00000a9c;  wr_data_rom[ 1792]='h00000000;
    rd_cycle[ 1793] = 1'b0;  wr_cycle[ 1793] = 1'b1;  addr_rom[ 1793]='h00000d10;  wr_data_rom[ 1793]='h00000eed;
    rd_cycle[ 1794] = 1'b0;  wr_cycle[ 1794] = 1'b1;  addr_rom[ 1794]='h000004ec;  wr_data_rom[ 1794]='h00000e57;
    rd_cycle[ 1795] = 1'b1;  wr_cycle[ 1795] = 1'b0;  addr_rom[ 1795]='h00000628;  wr_data_rom[ 1795]='h00000000;
    rd_cycle[ 1796] = 1'b1;  wr_cycle[ 1796] = 1'b0;  addr_rom[ 1796]='h000009f4;  wr_data_rom[ 1796]='h00000000;
    rd_cycle[ 1797] = 1'b1;  wr_cycle[ 1797] = 1'b0;  addr_rom[ 1797]='h00000704;  wr_data_rom[ 1797]='h00000000;
    rd_cycle[ 1798] = 1'b0;  wr_cycle[ 1798] = 1'b1;  addr_rom[ 1798]='h00000eec;  wr_data_rom[ 1798]='h00000111;
    rd_cycle[ 1799] = 1'b0;  wr_cycle[ 1799] = 1'b1;  addr_rom[ 1799]='h00000c18;  wr_data_rom[ 1799]='h00000e77;
    rd_cycle[ 1800] = 1'b1;  wr_cycle[ 1800] = 1'b0;  addr_rom[ 1800]='h000009d8;  wr_data_rom[ 1800]='h00000000;
    rd_cycle[ 1801] = 1'b0;  wr_cycle[ 1801] = 1'b1;  addr_rom[ 1801]='h00000c80;  wr_data_rom[ 1801]='h00000439;
    rd_cycle[ 1802] = 1'b0;  wr_cycle[ 1802] = 1'b1;  addr_rom[ 1802]='h00000520;  wr_data_rom[ 1802]='h00000603;
    rd_cycle[ 1803] = 1'b1;  wr_cycle[ 1803] = 1'b0;  addr_rom[ 1803]='h00000530;  wr_data_rom[ 1803]='h00000000;
    rd_cycle[ 1804] = 1'b0;  wr_cycle[ 1804] = 1'b1;  addr_rom[ 1804]='h00000124;  wr_data_rom[ 1804]='h000008cc;
    rd_cycle[ 1805] = 1'b0;  wr_cycle[ 1805] = 1'b1;  addr_rom[ 1805]='h00000aec;  wr_data_rom[ 1805]='h000005a0;
    rd_cycle[ 1806] = 1'b0;  wr_cycle[ 1806] = 1'b1;  addr_rom[ 1806]='h00000ad4;  wr_data_rom[ 1806]='h000001f2;
    rd_cycle[ 1807] = 1'b0;  wr_cycle[ 1807] = 1'b1;  addr_rom[ 1807]='h00000328;  wr_data_rom[ 1807]='h00000688;
    rd_cycle[ 1808] = 1'b1;  wr_cycle[ 1808] = 1'b0;  addr_rom[ 1808]='h000009a4;  wr_data_rom[ 1808]='h00000000;
    rd_cycle[ 1809] = 1'b0;  wr_cycle[ 1809] = 1'b1;  addr_rom[ 1809]='h0000009c;  wr_data_rom[ 1809]='h00000319;
    rd_cycle[ 1810] = 1'b1;  wr_cycle[ 1810] = 1'b0;  addr_rom[ 1810]='h00000d70;  wr_data_rom[ 1810]='h00000000;
    rd_cycle[ 1811] = 1'b0;  wr_cycle[ 1811] = 1'b1;  addr_rom[ 1811]='h00000a78;  wr_data_rom[ 1811]='h00000405;
    rd_cycle[ 1812] = 1'b1;  wr_cycle[ 1812] = 1'b0;  addr_rom[ 1812]='h00000e6c;  wr_data_rom[ 1812]='h00000000;
    rd_cycle[ 1813] = 1'b0;  wr_cycle[ 1813] = 1'b1;  addr_rom[ 1813]='h00000e18;  wr_data_rom[ 1813]='h00000bcf;
    rd_cycle[ 1814] = 1'b0;  wr_cycle[ 1814] = 1'b1;  addr_rom[ 1814]='h000005bc;  wr_data_rom[ 1814]='h00000465;
    rd_cycle[ 1815] = 1'b1;  wr_cycle[ 1815] = 1'b0;  addr_rom[ 1815]='h0000053c;  wr_data_rom[ 1815]='h00000000;
    rd_cycle[ 1816] = 1'b1;  wr_cycle[ 1816] = 1'b0;  addr_rom[ 1816]='h00000424;  wr_data_rom[ 1816]='h00000000;
    rd_cycle[ 1817] = 1'b0;  wr_cycle[ 1817] = 1'b1;  addr_rom[ 1817]='h00000698;  wr_data_rom[ 1817]='h000005de;
    rd_cycle[ 1818] = 1'b1;  wr_cycle[ 1818] = 1'b0;  addr_rom[ 1818]='h000004e8;  wr_data_rom[ 1818]='h00000000;
    rd_cycle[ 1819] = 1'b1;  wr_cycle[ 1819] = 1'b0;  addr_rom[ 1819]='h000001bc;  wr_data_rom[ 1819]='h00000000;
    rd_cycle[ 1820] = 1'b1;  wr_cycle[ 1820] = 1'b0;  addr_rom[ 1820]='h000007d0;  wr_data_rom[ 1820]='h00000000;
    rd_cycle[ 1821] = 1'b0;  wr_cycle[ 1821] = 1'b1;  addr_rom[ 1821]='h00000014;  wr_data_rom[ 1821]='h00000713;
    rd_cycle[ 1822] = 1'b1;  wr_cycle[ 1822] = 1'b0;  addr_rom[ 1822]='h000008a0;  wr_data_rom[ 1822]='h00000000;
    rd_cycle[ 1823] = 1'b0;  wr_cycle[ 1823] = 1'b1;  addr_rom[ 1823]='h0000021c;  wr_data_rom[ 1823]='h00000acc;
    rd_cycle[ 1824] = 1'b1;  wr_cycle[ 1824] = 1'b0;  addr_rom[ 1824]='h00000018;  wr_data_rom[ 1824]='h00000000;
    rd_cycle[ 1825] = 1'b1;  wr_cycle[ 1825] = 1'b0;  addr_rom[ 1825]='h000005d0;  wr_data_rom[ 1825]='h00000000;
    rd_cycle[ 1826] = 1'b1;  wr_cycle[ 1826] = 1'b0;  addr_rom[ 1826]='h000008dc;  wr_data_rom[ 1826]='h00000000;
    rd_cycle[ 1827] = 1'b1;  wr_cycle[ 1827] = 1'b0;  addr_rom[ 1827]='h000009b8;  wr_data_rom[ 1827]='h00000000;
    rd_cycle[ 1828] = 1'b0;  wr_cycle[ 1828] = 1'b1;  addr_rom[ 1828]='h00000900;  wr_data_rom[ 1828]='h0000039c;
    rd_cycle[ 1829] = 1'b1;  wr_cycle[ 1829] = 1'b0;  addr_rom[ 1829]='h00000758;  wr_data_rom[ 1829]='h00000000;
    rd_cycle[ 1830] = 1'b0;  wr_cycle[ 1830] = 1'b1;  addr_rom[ 1830]='h00000ebc;  wr_data_rom[ 1830]='h00000922;
    rd_cycle[ 1831] = 1'b0;  wr_cycle[ 1831] = 1'b1;  addr_rom[ 1831]='h00000210;  wr_data_rom[ 1831]='h00000915;
    rd_cycle[ 1832] = 1'b1;  wr_cycle[ 1832] = 1'b0;  addr_rom[ 1832]='h00000384;  wr_data_rom[ 1832]='h00000000;
    rd_cycle[ 1833] = 1'b1;  wr_cycle[ 1833] = 1'b0;  addr_rom[ 1833]='h000001a8;  wr_data_rom[ 1833]='h00000000;
    rd_cycle[ 1834] = 1'b1;  wr_cycle[ 1834] = 1'b0;  addr_rom[ 1834]='h00000220;  wr_data_rom[ 1834]='h00000000;
    rd_cycle[ 1835] = 1'b0;  wr_cycle[ 1835] = 1'b1;  addr_rom[ 1835]='h00000f08;  wr_data_rom[ 1835]='h00000d4a;
    rd_cycle[ 1836] = 1'b1;  wr_cycle[ 1836] = 1'b0;  addr_rom[ 1836]='h000005d4;  wr_data_rom[ 1836]='h00000000;
    rd_cycle[ 1837] = 1'b0;  wr_cycle[ 1837] = 1'b1;  addr_rom[ 1837]='h00000ce0;  wr_data_rom[ 1837]='h00000488;
    rd_cycle[ 1838] = 1'b0;  wr_cycle[ 1838] = 1'b1;  addr_rom[ 1838]='h000008f0;  wr_data_rom[ 1838]='h0000019f;
    rd_cycle[ 1839] = 1'b0;  wr_cycle[ 1839] = 1'b1;  addr_rom[ 1839]='h000003e4;  wr_data_rom[ 1839]='h00000c7c;
    rd_cycle[ 1840] = 1'b0;  wr_cycle[ 1840] = 1'b1;  addr_rom[ 1840]='h00000244;  wr_data_rom[ 1840]='h00000e13;
    rd_cycle[ 1841] = 1'b1;  wr_cycle[ 1841] = 1'b0;  addr_rom[ 1841]='h00000694;  wr_data_rom[ 1841]='h00000000;
    rd_cycle[ 1842] = 1'b1;  wr_cycle[ 1842] = 1'b0;  addr_rom[ 1842]='h00000e78;  wr_data_rom[ 1842]='h00000000;
    rd_cycle[ 1843] = 1'b1;  wr_cycle[ 1843] = 1'b0;  addr_rom[ 1843]='h000008cc;  wr_data_rom[ 1843]='h00000000;
    rd_cycle[ 1844] = 1'b0;  wr_cycle[ 1844] = 1'b1;  addr_rom[ 1844]='h0000025c;  wr_data_rom[ 1844]='h00000376;
    rd_cycle[ 1845] = 1'b1;  wr_cycle[ 1845] = 1'b0;  addr_rom[ 1845]='h00000b54;  wr_data_rom[ 1845]='h00000000;
    rd_cycle[ 1846] = 1'b0;  wr_cycle[ 1846] = 1'b1;  addr_rom[ 1846]='h00000940;  wr_data_rom[ 1846]='h00000ad4;
    rd_cycle[ 1847] = 1'b0;  wr_cycle[ 1847] = 1'b1;  addr_rom[ 1847]='h00000f2c;  wr_data_rom[ 1847]='h00000c6d;
    rd_cycle[ 1848] = 1'b0;  wr_cycle[ 1848] = 1'b1;  addr_rom[ 1848]='h00000474;  wr_data_rom[ 1848]='h00000cee;
    rd_cycle[ 1849] = 1'b0;  wr_cycle[ 1849] = 1'b1;  addr_rom[ 1849]='h00000c04;  wr_data_rom[ 1849]='h00000a2c;
    rd_cycle[ 1850] = 1'b0;  wr_cycle[ 1850] = 1'b1;  addr_rom[ 1850]='h00000880;  wr_data_rom[ 1850]='h00000f78;
    rd_cycle[ 1851] = 1'b0;  wr_cycle[ 1851] = 1'b1;  addr_rom[ 1851]='h00000a94;  wr_data_rom[ 1851]='h000007f3;
    rd_cycle[ 1852] = 1'b1;  wr_cycle[ 1852] = 1'b0;  addr_rom[ 1852]='h0000069c;  wr_data_rom[ 1852]='h00000000;
    rd_cycle[ 1853] = 1'b0;  wr_cycle[ 1853] = 1'b1;  addr_rom[ 1853]='h00000134;  wr_data_rom[ 1853]='h00000904;
    rd_cycle[ 1854] = 1'b1;  wr_cycle[ 1854] = 1'b0;  addr_rom[ 1854]='h000006bc;  wr_data_rom[ 1854]='h00000000;
    rd_cycle[ 1855] = 1'b0;  wr_cycle[ 1855] = 1'b1;  addr_rom[ 1855]='h000008b4;  wr_data_rom[ 1855]='h0000084d;
    rd_cycle[ 1856] = 1'b0;  wr_cycle[ 1856] = 1'b1;  addr_rom[ 1856]='h00000c9c;  wr_data_rom[ 1856]='h000001ca;
    rd_cycle[ 1857] = 1'b1;  wr_cycle[ 1857] = 1'b0;  addr_rom[ 1857]='h00000124;  wr_data_rom[ 1857]='h00000000;
    rd_cycle[ 1858] = 1'b1;  wr_cycle[ 1858] = 1'b0;  addr_rom[ 1858]='h00000328;  wr_data_rom[ 1858]='h00000000;
    rd_cycle[ 1859] = 1'b0;  wr_cycle[ 1859] = 1'b1;  addr_rom[ 1859]='h00000f44;  wr_data_rom[ 1859]='h00000951;
    rd_cycle[ 1860] = 1'b0;  wr_cycle[ 1860] = 1'b1;  addr_rom[ 1860]='h00000674;  wr_data_rom[ 1860]='h000008da;
    rd_cycle[ 1861] = 1'b1;  wr_cycle[ 1861] = 1'b0;  addr_rom[ 1861]='h00000cb4;  wr_data_rom[ 1861]='h00000000;
    rd_cycle[ 1862] = 1'b1;  wr_cycle[ 1862] = 1'b0;  addr_rom[ 1862]='h00000360;  wr_data_rom[ 1862]='h00000000;
    rd_cycle[ 1863] = 1'b1;  wr_cycle[ 1863] = 1'b0;  addr_rom[ 1863]='h00000930;  wr_data_rom[ 1863]='h00000000;
    rd_cycle[ 1864] = 1'b0;  wr_cycle[ 1864] = 1'b1;  addr_rom[ 1864]='h0000011c;  wr_data_rom[ 1864]='h00000255;
    rd_cycle[ 1865] = 1'b0;  wr_cycle[ 1865] = 1'b1;  addr_rom[ 1865]='h000008b0;  wr_data_rom[ 1865]='h000005c5;
    rd_cycle[ 1866] = 1'b1;  wr_cycle[ 1866] = 1'b0;  addr_rom[ 1866]='h000006c4;  wr_data_rom[ 1866]='h00000000;
    rd_cycle[ 1867] = 1'b1;  wr_cycle[ 1867] = 1'b0;  addr_rom[ 1867]='h00000e6c;  wr_data_rom[ 1867]='h00000000;
    rd_cycle[ 1868] = 1'b1;  wr_cycle[ 1868] = 1'b0;  addr_rom[ 1868]='h00000e20;  wr_data_rom[ 1868]='h00000000;
    rd_cycle[ 1869] = 1'b1;  wr_cycle[ 1869] = 1'b0;  addr_rom[ 1869]='h0000026c;  wr_data_rom[ 1869]='h00000000;
    rd_cycle[ 1870] = 1'b1;  wr_cycle[ 1870] = 1'b0;  addr_rom[ 1870]='h00000758;  wr_data_rom[ 1870]='h00000000;
    rd_cycle[ 1871] = 1'b1;  wr_cycle[ 1871] = 1'b0;  addr_rom[ 1871]='h00000b28;  wr_data_rom[ 1871]='h00000000;
    rd_cycle[ 1872] = 1'b1;  wr_cycle[ 1872] = 1'b0;  addr_rom[ 1872]='h00000de4;  wr_data_rom[ 1872]='h00000000;
    rd_cycle[ 1873] = 1'b1;  wr_cycle[ 1873] = 1'b0;  addr_rom[ 1873]='h000005c4;  wr_data_rom[ 1873]='h00000000;
    rd_cycle[ 1874] = 1'b1;  wr_cycle[ 1874] = 1'b0;  addr_rom[ 1874]='h00000cb4;  wr_data_rom[ 1874]='h00000000;
    rd_cycle[ 1875] = 1'b0;  wr_cycle[ 1875] = 1'b1;  addr_rom[ 1875]='h0000064c;  wr_data_rom[ 1875]='h00000c4a;
    rd_cycle[ 1876] = 1'b0;  wr_cycle[ 1876] = 1'b1;  addr_rom[ 1876]='h00000e58;  wr_data_rom[ 1876]='h000002d9;
    rd_cycle[ 1877] = 1'b0;  wr_cycle[ 1877] = 1'b1;  addr_rom[ 1877]='h000004a0;  wr_data_rom[ 1877]='h000000d6;
    rd_cycle[ 1878] = 1'b1;  wr_cycle[ 1878] = 1'b0;  addr_rom[ 1878]='h0000017c;  wr_data_rom[ 1878]='h00000000;
    rd_cycle[ 1879] = 1'b1;  wr_cycle[ 1879] = 1'b0;  addr_rom[ 1879]='h000002d0;  wr_data_rom[ 1879]='h00000000;
    rd_cycle[ 1880] = 1'b1;  wr_cycle[ 1880] = 1'b0;  addr_rom[ 1880]='h00000c28;  wr_data_rom[ 1880]='h00000000;
    rd_cycle[ 1881] = 1'b0;  wr_cycle[ 1881] = 1'b1;  addr_rom[ 1881]='h00000c20;  wr_data_rom[ 1881]='h000001b7;
    rd_cycle[ 1882] = 1'b0;  wr_cycle[ 1882] = 1'b1;  addr_rom[ 1882]='h00000d74;  wr_data_rom[ 1882]='h00000cd2;
    rd_cycle[ 1883] = 1'b0;  wr_cycle[ 1883] = 1'b1;  addr_rom[ 1883]='h00000550;  wr_data_rom[ 1883]='h00000be3;
    rd_cycle[ 1884] = 1'b1;  wr_cycle[ 1884] = 1'b0;  addr_rom[ 1884]='h000007ac;  wr_data_rom[ 1884]='h00000000;
    rd_cycle[ 1885] = 1'b0;  wr_cycle[ 1885] = 1'b1;  addr_rom[ 1885]='h00000064;  wr_data_rom[ 1885]='h00000385;
    rd_cycle[ 1886] = 1'b0;  wr_cycle[ 1886] = 1'b1;  addr_rom[ 1886]='h00000c78;  wr_data_rom[ 1886]='h00000d03;
    rd_cycle[ 1887] = 1'b0;  wr_cycle[ 1887] = 1'b1;  addr_rom[ 1887]='h000008f0;  wr_data_rom[ 1887]='h000004be;
    rd_cycle[ 1888] = 1'b1;  wr_cycle[ 1888] = 1'b0;  addr_rom[ 1888]='h0000046c;  wr_data_rom[ 1888]='h00000000;
    rd_cycle[ 1889] = 1'b0;  wr_cycle[ 1889] = 1'b1;  addr_rom[ 1889]='h0000021c;  wr_data_rom[ 1889]='h00000a22;
    rd_cycle[ 1890] = 1'b0;  wr_cycle[ 1890] = 1'b1;  addr_rom[ 1890]='h00000a64;  wr_data_rom[ 1890]='h00000cc3;
    rd_cycle[ 1891] = 1'b1;  wr_cycle[ 1891] = 1'b0;  addr_rom[ 1891]='h000006e8;  wr_data_rom[ 1891]='h00000000;
    rd_cycle[ 1892] = 1'b0;  wr_cycle[ 1892] = 1'b1;  addr_rom[ 1892]='h00000938;  wr_data_rom[ 1892]='h00000d0e;
    rd_cycle[ 1893] = 1'b1;  wr_cycle[ 1893] = 1'b0;  addr_rom[ 1893]='h00000c3c;  wr_data_rom[ 1893]='h00000000;
    rd_cycle[ 1894] = 1'b1;  wr_cycle[ 1894] = 1'b0;  addr_rom[ 1894]='h00000ec8;  wr_data_rom[ 1894]='h00000000;
    rd_cycle[ 1895] = 1'b1;  wr_cycle[ 1895] = 1'b0;  addr_rom[ 1895]='h00000408;  wr_data_rom[ 1895]='h00000000;
    rd_cycle[ 1896] = 1'b1;  wr_cycle[ 1896] = 1'b0;  addr_rom[ 1896]='h00000b50;  wr_data_rom[ 1896]='h00000000;
    rd_cycle[ 1897] = 1'b0;  wr_cycle[ 1897] = 1'b1;  addr_rom[ 1897]='h00000adc;  wr_data_rom[ 1897]='h000006bb;
    rd_cycle[ 1898] = 1'b1;  wr_cycle[ 1898] = 1'b0;  addr_rom[ 1898]='h00000b94;  wr_data_rom[ 1898]='h00000000;
    rd_cycle[ 1899] = 1'b1;  wr_cycle[ 1899] = 1'b0;  addr_rom[ 1899]='h00000ba0;  wr_data_rom[ 1899]='h00000000;
    rd_cycle[ 1900] = 1'b0;  wr_cycle[ 1900] = 1'b1;  addr_rom[ 1900]='h000003e4;  wr_data_rom[ 1900]='h00000e92;
    rd_cycle[ 1901] = 1'b0;  wr_cycle[ 1901] = 1'b1;  addr_rom[ 1901]='h00000ac0;  wr_data_rom[ 1901]='h000001f9;
    rd_cycle[ 1902] = 1'b1;  wr_cycle[ 1902] = 1'b0;  addr_rom[ 1902]='h00000b18;  wr_data_rom[ 1902]='h00000000;
    rd_cycle[ 1903] = 1'b1;  wr_cycle[ 1903] = 1'b0;  addr_rom[ 1903]='h00000e78;  wr_data_rom[ 1903]='h00000000;
    rd_cycle[ 1904] = 1'b0;  wr_cycle[ 1904] = 1'b1;  addr_rom[ 1904]='h00000240;  wr_data_rom[ 1904]='h000008db;
    rd_cycle[ 1905] = 1'b1;  wr_cycle[ 1905] = 1'b0;  addr_rom[ 1905]='h000000c0;  wr_data_rom[ 1905]='h00000000;
    rd_cycle[ 1906] = 1'b0;  wr_cycle[ 1906] = 1'b1;  addr_rom[ 1906]='h00000144;  wr_data_rom[ 1906]='h00000f99;
    rd_cycle[ 1907] = 1'b1;  wr_cycle[ 1907] = 1'b0;  addr_rom[ 1907]='h000004a0;  wr_data_rom[ 1907]='h00000000;
    rd_cycle[ 1908] = 1'b0;  wr_cycle[ 1908] = 1'b1;  addr_rom[ 1908]='h00000f50;  wr_data_rom[ 1908]='h0000058d;
    rd_cycle[ 1909] = 1'b1;  wr_cycle[ 1909] = 1'b0;  addr_rom[ 1909]='h00000a60;  wr_data_rom[ 1909]='h00000000;
    rd_cycle[ 1910] = 1'b1;  wr_cycle[ 1910] = 1'b0;  addr_rom[ 1910]='h000004cc;  wr_data_rom[ 1910]='h00000000;
    rd_cycle[ 1911] = 1'b0;  wr_cycle[ 1911] = 1'b1;  addr_rom[ 1911]='h00000940;  wr_data_rom[ 1911]='h000007ee;
    rd_cycle[ 1912] = 1'b0;  wr_cycle[ 1912] = 1'b1;  addr_rom[ 1912]='h00000a44;  wr_data_rom[ 1912]='h00000b90;
    rd_cycle[ 1913] = 1'b1;  wr_cycle[ 1913] = 1'b0;  addr_rom[ 1913]='h0000030c;  wr_data_rom[ 1913]='h00000000;
    rd_cycle[ 1914] = 1'b0;  wr_cycle[ 1914] = 1'b1;  addr_rom[ 1914]='h000005cc;  wr_data_rom[ 1914]='h00000f79;
    rd_cycle[ 1915] = 1'b1;  wr_cycle[ 1915] = 1'b0;  addr_rom[ 1915]='h0000039c;  wr_data_rom[ 1915]='h00000000;
    rd_cycle[ 1916] = 1'b1;  wr_cycle[ 1916] = 1'b0;  addr_rom[ 1916]='h00000e50;  wr_data_rom[ 1916]='h00000000;
    rd_cycle[ 1917] = 1'b1;  wr_cycle[ 1917] = 1'b0;  addr_rom[ 1917]='h00000f20;  wr_data_rom[ 1917]='h00000000;
    rd_cycle[ 1918] = 1'b1;  wr_cycle[ 1918] = 1'b0;  addr_rom[ 1918]='h00000720;  wr_data_rom[ 1918]='h00000000;
    rd_cycle[ 1919] = 1'b0;  wr_cycle[ 1919] = 1'b1;  addr_rom[ 1919]='h00000d34;  wr_data_rom[ 1919]='h00000065;
    rd_cycle[ 1920] = 1'b0;  wr_cycle[ 1920] = 1'b1;  addr_rom[ 1920]='h00000574;  wr_data_rom[ 1920]='h000007f0;
    rd_cycle[ 1921] = 1'b0;  wr_cycle[ 1921] = 1'b1;  addr_rom[ 1921]='h00000da4;  wr_data_rom[ 1921]='h00000e2c;
    rd_cycle[ 1922] = 1'b1;  wr_cycle[ 1922] = 1'b0;  addr_rom[ 1922]='h00000a20;  wr_data_rom[ 1922]='h00000000;
    rd_cycle[ 1923] = 1'b1;  wr_cycle[ 1923] = 1'b0;  addr_rom[ 1923]='h0000039c;  wr_data_rom[ 1923]='h00000000;
    rd_cycle[ 1924] = 1'b0;  wr_cycle[ 1924] = 1'b1;  addr_rom[ 1924]='h00000914;  wr_data_rom[ 1924]='h00000ef4;
    rd_cycle[ 1925] = 1'b0;  wr_cycle[ 1925] = 1'b1;  addr_rom[ 1925]='h00000d7c;  wr_data_rom[ 1925]='h000007db;
    rd_cycle[ 1926] = 1'b1;  wr_cycle[ 1926] = 1'b0;  addr_rom[ 1926]='h00000e20;  wr_data_rom[ 1926]='h00000000;
    rd_cycle[ 1927] = 1'b0;  wr_cycle[ 1927] = 1'b1;  addr_rom[ 1927]='h000006d8;  wr_data_rom[ 1927]='h000004aa;
    rd_cycle[ 1928] = 1'b1;  wr_cycle[ 1928] = 1'b0;  addr_rom[ 1928]='h000004cc;  wr_data_rom[ 1928]='h00000000;
    rd_cycle[ 1929] = 1'b1;  wr_cycle[ 1929] = 1'b0;  addr_rom[ 1929]='h00000a48;  wr_data_rom[ 1929]='h00000000;
    rd_cycle[ 1930] = 1'b0;  wr_cycle[ 1930] = 1'b1;  addr_rom[ 1930]='h00000d24;  wr_data_rom[ 1930]='h00000261;
    rd_cycle[ 1931] = 1'b0;  wr_cycle[ 1931] = 1'b1;  addr_rom[ 1931]='h00000454;  wr_data_rom[ 1931]='h00000390;
    rd_cycle[ 1932] = 1'b1;  wr_cycle[ 1932] = 1'b0;  addr_rom[ 1932]='h00000be4;  wr_data_rom[ 1932]='h00000000;
    rd_cycle[ 1933] = 1'b0;  wr_cycle[ 1933] = 1'b1;  addr_rom[ 1933]='h00000604;  wr_data_rom[ 1933]='h0000063e;
    rd_cycle[ 1934] = 1'b0;  wr_cycle[ 1934] = 1'b1;  addr_rom[ 1934]='h00000de4;  wr_data_rom[ 1934]='h00000102;
    rd_cycle[ 1935] = 1'b0;  wr_cycle[ 1935] = 1'b1;  addr_rom[ 1935]='h00000cfc;  wr_data_rom[ 1935]='h00000df2;
    rd_cycle[ 1936] = 1'b0;  wr_cycle[ 1936] = 1'b1;  addr_rom[ 1936]='h00000128;  wr_data_rom[ 1936]='h0000088b;
    rd_cycle[ 1937] = 1'b1;  wr_cycle[ 1937] = 1'b0;  addr_rom[ 1937]='h00000298;  wr_data_rom[ 1937]='h00000000;
    rd_cycle[ 1938] = 1'b1;  wr_cycle[ 1938] = 1'b0;  addr_rom[ 1938]='h00000a88;  wr_data_rom[ 1938]='h00000000;
    rd_cycle[ 1939] = 1'b1;  wr_cycle[ 1939] = 1'b0;  addr_rom[ 1939]='h000006c4;  wr_data_rom[ 1939]='h00000000;
    rd_cycle[ 1940] = 1'b1;  wr_cycle[ 1940] = 1'b0;  addr_rom[ 1940]='h00000790;  wr_data_rom[ 1940]='h00000000;
    rd_cycle[ 1941] = 1'b0;  wr_cycle[ 1941] = 1'b1;  addr_rom[ 1941]='h00000a78;  wr_data_rom[ 1941]='h00000714;
    rd_cycle[ 1942] = 1'b1;  wr_cycle[ 1942] = 1'b0;  addr_rom[ 1942]='h000006b4;  wr_data_rom[ 1942]='h00000000;
    rd_cycle[ 1943] = 1'b1;  wr_cycle[ 1943] = 1'b0;  addr_rom[ 1943]='h00000ee4;  wr_data_rom[ 1943]='h00000000;
    rd_cycle[ 1944] = 1'b1;  wr_cycle[ 1944] = 1'b0;  addr_rom[ 1944]='h000007d8;  wr_data_rom[ 1944]='h00000000;
    rd_cycle[ 1945] = 1'b1;  wr_cycle[ 1945] = 1'b0;  addr_rom[ 1945]='h00000ad0;  wr_data_rom[ 1945]='h00000000;
    rd_cycle[ 1946] = 1'b0;  wr_cycle[ 1946] = 1'b1;  addr_rom[ 1946]='h000003b4;  wr_data_rom[ 1946]='h00000220;
    rd_cycle[ 1947] = 1'b1;  wr_cycle[ 1947] = 1'b0;  addr_rom[ 1947]='h00000f74;  wr_data_rom[ 1947]='h00000000;
    rd_cycle[ 1948] = 1'b1;  wr_cycle[ 1948] = 1'b0;  addr_rom[ 1948]='h00000510;  wr_data_rom[ 1948]='h00000000;
    rd_cycle[ 1949] = 1'b0;  wr_cycle[ 1949] = 1'b1;  addr_rom[ 1949]='h00000b10;  wr_data_rom[ 1949]='h000008ea;
    rd_cycle[ 1950] = 1'b1;  wr_cycle[ 1950] = 1'b0;  addr_rom[ 1950]='h000000b0;  wr_data_rom[ 1950]='h00000000;
    rd_cycle[ 1951] = 1'b1;  wr_cycle[ 1951] = 1'b0;  addr_rom[ 1951]='h00000668;  wr_data_rom[ 1951]='h00000000;
    rd_cycle[ 1952] = 1'b1;  wr_cycle[ 1952] = 1'b0;  addr_rom[ 1952]='h00000ec0;  wr_data_rom[ 1952]='h00000000;
    rd_cycle[ 1953] = 1'b0;  wr_cycle[ 1953] = 1'b1;  addr_rom[ 1953]='h000001fc;  wr_data_rom[ 1953]='h00000e9b;
    rd_cycle[ 1954] = 1'b1;  wr_cycle[ 1954] = 1'b0;  addr_rom[ 1954]='h00000284;  wr_data_rom[ 1954]='h00000000;
    rd_cycle[ 1955] = 1'b1;  wr_cycle[ 1955] = 1'b0;  addr_rom[ 1955]='h00000bbc;  wr_data_rom[ 1955]='h00000000;
    rd_cycle[ 1956] = 1'b0;  wr_cycle[ 1956] = 1'b1;  addr_rom[ 1956]='h00000ed4;  wr_data_rom[ 1956]='h00000d94;
    rd_cycle[ 1957] = 1'b0;  wr_cycle[ 1957] = 1'b1;  addr_rom[ 1957]='h00000e50;  wr_data_rom[ 1957]='h00000511;
    rd_cycle[ 1958] = 1'b0;  wr_cycle[ 1958] = 1'b1;  addr_rom[ 1958]='h00000520;  wr_data_rom[ 1958]='h00000903;
    rd_cycle[ 1959] = 1'b0;  wr_cycle[ 1959] = 1'b1;  addr_rom[ 1959]='h00000edc;  wr_data_rom[ 1959]='h00000ef0;
    rd_cycle[ 1960] = 1'b0;  wr_cycle[ 1960] = 1'b1;  addr_rom[ 1960]='h00000120;  wr_data_rom[ 1960]='h00000cd5;
    rd_cycle[ 1961] = 1'b0;  wr_cycle[ 1961] = 1'b1;  addr_rom[ 1961]='h000003e0;  wr_data_rom[ 1961]='h00000628;
    rd_cycle[ 1962] = 1'b1;  wr_cycle[ 1962] = 1'b0;  addr_rom[ 1962]='h000005f8;  wr_data_rom[ 1962]='h00000000;
    rd_cycle[ 1963] = 1'b0;  wr_cycle[ 1963] = 1'b1;  addr_rom[ 1963]='h000003e8;  wr_data_rom[ 1963]='h000007a4;
    rd_cycle[ 1964] = 1'b0;  wr_cycle[ 1964] = 1'b1;  addr_rom[ 1964]='h00000014;  wr_data_rom[ 1964]='h00000a18;
    rd_cycle[ 1965] = 1'b0;  wr_cycle[ 1965] = 1'b1;  addr_rom[ 1965]='h00000a9c;  wr_data_rom[ 1965]='h00000c64;
    rd_cycle[ 1966] = 1'b0;  wr_cycle[ 1966] = 1'b1;  addr_rom[ 1966]='h00000614;  wr_data_rom[ 1966]='h0000099f;
    rd_cycle[ 1967] = 1'b0;  wr_cycle[ 1967] = 1'b1;  addr_rom[ 1967]='h00000d50;  wr_data_rom[ 1967]='h00000f93;
    rd_cycle[ 1968] = 1'b1;  wr_cycle[ 1968] = 1'b0;  addr_rom[ 1968]='h00000ee4;  wr_data_rom[ 1968]='h00000000;
    rd_cycle[ 1969] = 1'b0;  wr_cycle[ 1969] = 1'b1;  addr_rom[ 1969]='h00000b84;  wr_data_rom[ 1969]='h000004a8;
    rd_cycle[ 1970] = 1'b1;  wr_cycle[ 1970] = 1'b0;  addr_rom[ 1970]='h00000b40;  wr_data_rom[ 1970]='h00000000;
    rd_cycle[ 1971] = 1'b1;  wr_cycle[ 1971] = 1'b0;  addr_rom[ 1971]='h000002e8;  wr_data_rom[ 1971]='h00000000;
    rd_cycle[ 1972] = 1'b1;  wr_cycle[ 1972] = 1'b0;  addr_rom[ 1972]='h00000480;  wr_data_rom[ 1972]='h00000000;
    rd_cycle[ 1973] = 1'b0;  wr_cycle[ 1973] = 1'b1;  addr_rom[ 1973]='h000006b8;  wr_data_rom[ 1973]='h00000d83;
    rd_cycle[ 1974] = 1'b0;  wr_cycle[ 1974] = 1'b1;  addr_rom[ 1974]='h0000070c;  wr_data_rom[ 1974]='h000002e5;
    rd_cycle[ 1975] = 1'b0;  wr_cycle[ 1975] = 1'b1;  addr_rom[ 1975]='h00000648;  wr_data_rom[ 1975]='h000004b1;
    rd_cycle[ 1976] = 1'b0;  wr_cycle[ 1976] = 1'b1;  addr_rom[ 1976]='h00000da4;  wr_data_rom[ 1976]='h0000021e;
    rd_cycle[ 1977] = 1'b0;  wr_cycle[ 1977] = 1'b1;  addr_rom[ 1977]='h00000f88;  wr_data_rom[ 1977]='h00000b8c;
    rd_cycle[ 1978] = 1'b0;  wr_cycle[ 1978] = 1'b1;  addr_rom[ 1978]='h00000434;  wr_data_rom[ 1978]='h00000c13;
    rd_cycle[ 1979] = 1'b0;  wr_cycle[ 1979] = 1'b1;  addr_rom[ 1979]='h0000068c;  wr_data_rom[ 1979]='h00000741;
    rd_cycle[ 1980] = 1'b1;  wr_cycle[ 1980] = 1'b0;  addr_rom[ 1980]='h00000c30;  wr_data_rom[ 1980]='h00000000;
    rd_cycle[ 1981] = 1'b1;  wr_cycle[ 1981] = 1'b0;  addr_rom[ 1981]='h00000288;  wr_data_rom[ 1981]='h00000000;
    rd_cycle[ 1982] = 1'b0;  wr_cycle[ 1982] = 1'b1;  addr_rom[ 1982]='h00000f00;  wr_data_rom[ 1982]='h000000f0;
    rd_cycle[ 1983] = 1'b1;  wr_cycle[ 1983] = 1'b0;  addr_rom[ 1983]='h00000b8c;  wr_data_rom[ 1983]='h00000000;
    rd_cycle[ 1984] = 1'b0;  wr_cycle[ 1984] = 1'b1;  addr_rom[ 1984]='h00000f70;  wr_data_rom[ 1984]='h00000184;
    rd_cycle[ 1985] = 1'b1;  wr_cycle[ 1985] = 1'b0;  addr_rom[ 1985]='h00000d80;  wr_data_rom[ 1985]='h00000000;
    rd_cycle[ 1986] = 1'b1;  wr_cycle[ 1986] = 1'b0;  addr_rom[ 1986]='h00000ebc;  wr_data_rom[ 1986]='h00000000;
    rd_cycle[ 1987] = 1'b1;  wr_cycle[ 1987] = 1'b0;  addr_rom[ 1987]='h00000504;  wr_data_rom[ 1987]='h00000000;
    rd_cycle[ 1988] = 1'b1;  wr_cycle[ 1988] = 1'b0;  addr_rom[ 1988]='h000005fc;  wr_data_rom[ 1988]='h00000000;
    rd_cycle[ 1989] = 1'b1;  wr_cycle[ 1989] = 1'b0;  addr_rom[ 1989]='h0000035c;  wr_data_rom[ 1989]='h00000000;
    rd_cycle[ 1990] = 1'b1;  wr_cycle[ 1990] = 1'b0;  addr_rom[ 1990]='h000004fc;  wr_data_rom[ 1990]='h00000000;
    rd_cycle[ 1991] = 1'b0;  wr_cycle[ 1991] = 1'b1;  addr_rom[ 1991]='h00000d6c;  wr_data_rom[ 1991]='h00000d77;
    rd_cycle[ 1992] = 1'b0;  wr_cycle[ 1992] = 1'b1;  addr_rom[ 1992]='h0000040c;  wr_data_rom[ 1992]='h0000084d;
    rd_cycle[ 1993] = 1'b1;  wr_cycle[ 1993] = 1'b0;  addr_rom[ 1993]='h00000c20;  wr_data_rom[ 1993]='h00000000;
    rd_cycle[ 1994] = 1'b1;  wr_cycle[ 1994] = 1'b0;  addr_rom[ 1994]='h0000050c;  wr_data_rom[ 1994]='h00000000;
    rd_cycle[ 1995] = 1'b0;  wr_cycle[ 1995] = 1'b1;  addr_rom[ 1995]='h00000994;  wr_data_rom[ 1995]='h000003da;
    rd_cycle[ 1996] = 1'b1;  wr_cycle[ 1996] = 1'b0;  addr_rom[ 1996]='h0000006c;  wr_data_rom[ 1996]='h00000000;
    rd_cycle[ 1997] = 1'b1;  wr_cycle[ 1997] = 1'b0;  addr_rom[ 1997]='h00000444;  wr_data_rom[ 1997]='h00000000;
    rd_cycle[ 1998] = 1'b0;  wr_cycle[ 1998] = 1'b1;  addr_rom[ 1998]='h00000dec;  wr_data_rom[ 1998]='h0000041f;
    rd_cycle[ 1999] = 1'b0;  wr_cycle[ 1999] = 1'b1;  addr_rom[ 1999]='h00000e80;  wr_data_rom[ 1999]='h00000a34;
    rd_cycle[ 2000] = 1'b1;  wr_cycle[ 2000] = 1'b0;  addr_rom[ 2000]='h000001a8;  wr_data_rom[ 2000]='h00000000;
    rd_cycle[ 2001] = 1'b1;  wr_cycle[ 2001] = 1'b0;  addr_rom[ 2001]='h00000b38;  wr_data_rom[ 2001]='h00000000;
    rd_cycle[ 2002] = 1'b0;  wr_cycle[ 2002] = 1'b1;  addr_rom[ 2002]='h00000e84;  wr_data_rom[ 2002]='h00000381;
    rd_cycle[ 2003] = 1'b0;  wr_cycle[ 2003] = 1'b1;  addr_rom[ 2003]='h00000acc;  wr_data_rom[ 2003]='h000004c1;
    rd_cycle[ 2004] = 1'b0;  wr_cycle[ 2004] = 1'b1;  addr_rom[ 2004]='h00000468;  wr_data_rom[ 2004]='h00000e5d;
    rd_cycle[ 2005] = 1'b1;  wr_cycle[ 2005] = 1'b0;  addr_rom[ 2005]='h00000d88;  wr_data_rom[ 2005]='h00000000;
    rd_cycle[ 2006] = 1'b0;  wr_cycle[ 2006] = 1'b1;  addr_rom[ 2006]='h00000cd0;  wr_data_rom[ 2006]='h00000dd3;
    rd_cycle[ 2007] = 1'b0;  wr_cycle[ 2007] = 1'b1;  addr_rom[ 2007]='h000003e8;  wr_data_rom[ 2007]='h000008fc;
    rd_cycle[ 2008] = 1'b1;  wr_cycle[ 2008] = 1'b0;  addr_rom[ 2008]='h00000370;  wr_data_rom[ 2008]='h00000000;
    rd_cycle[ 2009] = 1'b1;  wr_cycle[ 2009] = 1'b0;  addr_rom[ 2009]='h000001d0;  wr_data_rom[ 2009]='h00000000;
    rd_cycle[ 2010] = 1'b1;  wr_cycle[ 2010] = 1'b0;  addr_rom[ 2010]='h00000c44;  wr_data_rom[ 2010]='h00000000;
    rd_cycle[ 2011] = 1'b0;  wr_cycle[ 2011] = 1'b1;  addr_rom[ 2011]='h00000718;  wr_data_rom[ 2011]='h0000049f;
    rd_cycle[ 2012] = 1'b1;  wr_cycle[ 2012] = 1'b0;  addr_rom[ 2012]='h00000290;  wr_data_rom[ 2012]='h00000000;
    rd_cycle[ 2013] = 1'b1;  wr_cycle[ 2013] = 1'b0;  addr_rom[ 2013]='h000006f8;  wr_data_rom[ 2013]='h00000000;
    rd_cycle[ 2014] = 1'b0;  wr_cycle[ 2014] = 1'b1;  addr_rom[ 2014]='h000006f0;  wr_data_rom[ 2014]='h000000d4;
    rd_cycle[ 2015] = 1'b0;  wr_cycle[ 2015] = 1'b1;  addr_rom[ 2015]='h00000754;  wr_data_rom[ 2015]='h00000ee4;
    rd_cycle[ 2016] = 1'b0;  wr_cycle[ 2016] = 1'b1;  addr_rom[ 2016]='h00000e28;  wr_data_rom[ 2016]='h00000945;
    rd_cycle[ 2017] = 1'b0;  wr_cycle[ 2017] = 1'b1;  addr_rom[ 2017]='h00000ebc;  wr_data_rom[ 2017]='h000001be;
    rd_cycle[ 2018] = 1'b1;  wr_cycle[ 2018] = 1'b0;  addr_rom[ 2018]='h00000b68;  wr_data_rom[ 2018]='h00000000;
    rd_cycle[ 2019] = 1'b0;  wr_cycle[ 2019] = 1'b1;  addr_rom[ 2019]='h00000c18;  wr_data_rom[ 2019]='h00000c78;
    rd_cycle[ 2020] = 1'b0;  wr_cycle[ 2020] = 1'b1;  addr_rom[ 2020]='h000004a0;  wr_data_rom[ 2020]='h00000de3;
    rd_cycle[ 2021] = 1'b0;  wr_cycle[ 2021] = 1'b1;  addr_rom[ 2021]='h000000a0;  wr_data_rom[ 2021]='h00000241;
    rd_cycle[ 2022] = 1'b0;  wr_cycle[ 2022] = 1'b1;  addr_rom[ 2022]='h00000c20;  wr_data_rom[ 2022]='h000003da;
    rd_cycle[ 2023] = 1'b0;  wr_cycle[ 2023] = 1'b1;  addr_rom[ 2023]='h000005e0;  wr_data_rom[ 2023]='h0000070e;
    rd_cycle[ 2024] = 1'b0;  wr_cycle[ 2024] = 1'b1;  addr_rom[ 2024]='h00000484;  wr_data_rom[ 2024]='h00000635;
    rd_cycle[ 2025] = 1'b1;  wr_cycle[ 2025] = 1'b0;  addr_rom[ 2025]='h000007a8;  wr_data_rom[ 2025]='h00000000;
    rd_cycle[ 2026] = 1'b1;  wr_cycle[ 2026] = 1'b0;  addr_rom[ 2026]='h00000068;  wr_data_rom[ 2026]='h00000000;
    rd_cycle[ 2027] = 1'b1;  wr_cycle[ 2027] = 1'b0;  addr_rom[ 2027]='h00000304;  wr_data_rom[ 2027]='h00000000;
    rd_cycle[ 2028] = 1'b0;  wr_cycle[ 2028] = 1'b1;  addr_rom[ 2028]='h00000c38;  wr_data_rom[ 2028]='h00000817;
    rd_cycle[ 2029] = 1'b0;  wr_cycle[ 2029] = 1'b1;  addr_rom[ 2029]='h00000c08;  wr_data_rom[ 2029]='h00000a3c;
    rd_cycle[ 2030] = 1'b0;  wr_cycle[ 2030] = 1'b1;  addr_rom[ 2030]='h00000a58;  wr_data_rom[ 2030]='h00000b5e;
    rd_cycle[ 2031] = 1'b0;  wr_cycle[ 2031] = 1'b1;  addr_rom[ 2031]='h00000494;  wr_data_rom[ 2031]='h000003d6;
    rd_cycle[ 2032] = 1'b1;  wr_cycle[ 2032] = 1'b0;  addr_rom[ 2032]='h00000ea0;  wr_data_rom[ 2032]='h00000000;
    rd_cycle[ 2033] = 1'b0;  wr_cycle[ 2033] = 1'b1;  addr_rom[ 2033]='h000004dc;  wr_data_rom[ 2033]='h000008e3;
    rd_cycle[ 2034] = 1'b0;  wr_cycle[ 2034] = 1'b1;  addr_rom[ 2034]='h0000020c;  wr_data_rom[ 2034]='h00000607;
    rd_cycle[ 2035] = 1'b0;  wr_cycle[ 2035] = 1'b1;  addr_rom[ 2035]='h0000076c;  wr_data_rom[ 2035]='h00000ac6;
    rd_cycle[ 2036] = 1'b0;  wr_cycle[ 2036] = 1'b1;  addr_rom[ 2036]='h0000091c;  wr_data_rom[ 2036]='h000001f7;
    rd_cycle[ 2037] = 1'b1;  wr_cycle[ 2037] = 1'b0;  addr_rom[ 2037]='h000004f4;  wr_data_rom[ 2037]='h00000000;
    rd_cycle[ 2038] = 1'b1;  wr_cycle[ 2038] = 1'b0;  addr_rom[ 2038]='h000000c0;  wr_data_rom[ 2038]='h00000000;
    rd_cycle[ 2039] = 1'b0;  wr_cycle[ 2039] = 1'b1;  addr_rom[ 2039]='h000003b0;  wr_data_rom[ 2039]='h00000e80;
    rd_cycle[ 2040] = 1'b0;  wr_cycle[ 2040] = 1'b1;  addr_rom[ 2040]='h000005f8;  wr_data_rom[ 2040]='h000009ef;
    rd_cycle[ 2041] = 1'b1;  wr_cycle[ 2041] = 1'b0;  addr_rom[ 2041]='h00000e90;  wr_data_rom[ 2041]='h00000000;
    rd_cycle[ 2042] = 1'b0;  wr_cycle[ 2042] = 1'b1;  addr_rom[ 2042]='h00000424;  wr_data_rom[ 2042]='h00000505;
    rd_cycle[ 2043] = 1'b1;  wr_cycle[ 2043] = 1'b0;  addr_rom[ 2043]='h00000804;  wr_data_rom[ 2043]='h00000000;
    rd_cycle[ 2044] = 1'b1;  wr_cycle[ 2044] = 1'b0;  addr_rom[ 2044]='h00000c5c;  wr_data_rom[ 2044]='h00000000;
    rd_cycle[ 2045] = 1'b1;  wr_cycle[ 2045] = 1'b0;  addr_rom[ 2045]='h00000278;  wr_data_rom[ 2045]='h00000000;
    rd_cycle[ 2046] = 1'b1;  wr_cycle[ 2046] = 1'b0;  addr_rom[ 2046]='h00000600;  wr_data_rom[ 2046]='h00000000;
    rd_cycle[ 2047] = 1'b0;  wr_cycle[ 2047] = 1'b1;  addr_rom[ 2047]='h00000944;  wr_data_rom[ 2047]='h00000206;
    rd_cycle[ 2048] = 1'b0;  wr_cycle[ 2048] = 1'b1;  addr_rom[ 2048]='h000006f8;  wr_data_rom[ 2048]='h00000707;
    rd_cycle[ 2049] = 1'b1;  wr_cycle[ 2049] = 1'b0;  addr_rom[ 2049]='h00000a40;  wr_data_rom[ 2049]='h00000000;
    rd_cycle[ 2050] = 1'b0;  wr_cycle[ 2050] = 1'b1;  addr_rom[ 2050]='h00000bb4;  wr_data_rom[ 2050]='h000008df;
    rd_cycle[ 2051] = 1'b0;  wr_cycle[ 2051] = 1'b1;  addr_rom[ 2051]='h00000f14;  wr_data_rom[ 2051]='h00000840;
    rd_cycle[ 2052] = 1'b0;  wr_cycle[ 2052] = 1'b1;  addr_rom[ 2052]='h000008c4;  wr_data_rom[ 2052]='h00000cd5;
    rd_cycle[ 2053] = 1'b0;  wr_cycle[ 2053] = 1'b1;  addr_rom[ 2053]='h00000bac;  wr_data_rom[ 2053]='h0000004f;
    rd_cycle[ 2054] = 1'b1;  wr_cycle[ 2054] = 1'b0;  addr_rom[ 2054]='h000001f8;  wr_data_rom[ 2054]='h00000000;
    rd_cycle[ 2055] = 1'b1;  wr_cycle[ 2055] = 1'b0;  addr_rom[ 2055]='h00000d90;  wr_data_rom[ 2055]='h00000000;
    rd_cycle[ 2056] = 1'b1;  wr_cycle[ 2056] = 1'b0;  addr_rom[ 2056]='h00000aa8;  wr_data_rom[ 2056]='h00000000;
    rd_cycle[ 2057] = 1'b0;  wr_cycle[ 2057] = 1'b1;  addr_rom[ 2057]='h000007a8;  wr_data_rom[ 2057]='h0000017c;
    rd_cycle[ 2058] = 1'b1;  wr_cycle[ 2058] = 1'b0;  addr_rom[ 2058]='h00000f44;  wr_data_rom[ 2058]='h00000000;
    rd_cycle[ 2059] = 1'b1;  wr_cycle[ 2059] = 1'b0;  addr_rom[ 2059]='h00000818;  wr_data_rom[ 2059]='h00000000;
    rd_cycle[ 2060] = 1'b1;  wr_cycle[ 2060] = 1'b0;  addr_rom[ 2060]='h00000a34;  wr_data_rom[ 2060]='h00000000;
    rd_cycle[ 2061] = 1'b0;  wr_cycle[ 2061] = 1'b1;  addr_rom[ 2061]='h00000b08;  wr_data_rom[ 2061]='h00000773;
    rd_cycle[ 2062] = 1'b1;  wr_cycle[ 2062] = 1'b0;  addr_rom[ 2062]='h000000a0;  wr_data_rom[ 2062]='h00000000;
    rd_cycle[ 2063] = 1'b0;  wr_cycle[ 2063] = 1'b1;  addr_rom[ 2063]='h00000780;  wr_data_rom[ 2063]='h00000704;
    rd_cycle[ 2064] = 1'b1;  wr_cycle[ 2064] = 1'b0;  addr_rom[ 2064]='h00000eb0;  wr_data_rom[ 2064]='h00000000;
    rd_cycle[ 2065] = 1'b1;  wr_cycle[ 2065] = 1'b0;  addr_rom[ 2065]='h00000164;  wr_data_rom[ 2065]='h00000000;
    rd_cycle[ 2066] = 1'b0;  wr_cycle[ 2066] = 1'b1;  addr_rom[ 2066]='h000001ac;  wr_data_rom[ 2066]='h000008b7;
    rd_cycle[ 2067] = 1'b0;  wr_cycle[ 2067] = 1'b1;  addr_rom[ 2067]='h00000008;  wr_data_rom[ 2067]='h00000f7e;
    rd_cycle[ 2068] = 1'b1;  wr_cycle[ 2068] = 1'b0;  addr_rom[ 2068]='h00000b4c;  wr_data_rom[ 2068]='h00000000;
    rd_cycle[ 2069] = 1'b1;  wr_cycle[ 2069] = 1'b0;  addr_rom[ 2069]='h00000268;  wr_data_rom[ 2069]='h00000000;
    rd_cycle[ 2070] = 1'b1;  wr_cycle[ 2070] = 1'b0;  addr_rom[ 2070]='h00000dc0;  wr_data_rom[ 2070]='h00000000;
    rd_cycle[ 2071] = 1'b0;  wr_cycle[ 2071] = 1'b1;  addr_rom[ 2071]='h00000a4c;  wr_data_rom[ 2071]='h0000020a;
    rd_cycle[ 2072] = 1'b0;  wr_cycle[ 2072] = 1'b1;  addr_rom[ 2072]='h00000a50;  wr_data_rom[ 2072]='h000007a0;
    rd_cycle[ 2073] = 1'b0;  wr_cycle[ 2073] = 1'b1;  addr_rom[ 2073]='h00000808;  wr_data_rom[ 2073]='h00000f97;
    rd_cycle[ 2074] = 1'b0;  wr_cycle[ 2074] = 1'b1;  addr_rom[ 2074]='h00000194;  wr_data_rom[ 2074]='h0000062e;
    rd_cycle[ 2075] = 1'b1;  wr_cycle[ 2075] = 1'b0;  addr_rom[ 2075]='h00000250;  wr_data_rom[ 2075]='h00000000;
    rd_cycle[ 2076] = 1'b1;  wr_cycle[ 2076] = 1'b0;  addr_rom[ 2076]='h000000c0;  wr_data_rom[ 2076]='h00000000;
    rd_cycle[ 2077] = 1'b1;  wr_cycle[ 2077] = 1'b0;  addr_rom[ 2077]='h00000824;  wr_data_rom[ 2077]='h00000000;
    rd_cycle[ 2078] = 1'b1;  wr_cycle[ 2078] = 1'b0;  addr_rom[ 2078]='h00000aac;  wr_data_rom[ 2078]='h00000000;
    rd_cycle[ 2079] = 1'b0;  wr_cycle[ 2079] = 1'b1;  addr_rom[ 2079]='h00000e84;  wr_data_rom[ 2079]='h0000099c;
    rd_cycle[ 2080] = 1'b0;  wr_cycle[ 2080] = 1'b1;  addr_rom[ 2080]='h00000cd0;  wr_data_rom[ 2080]='h000009bf;
    rd_cycle[ 2081] = 1'b0;  wr_cycle[ 2081] = 1'b1;  addr_rom[ 2081]='h00000410;  wr_data_rom[ 2081]='h00000f60;
    rd_cycle[ 2082] = 1'b1;  wr_cycle[ 2082] = 1'b0;  addr_rom[ 2082]='h00000224;  wr_data_rom[ 2082]='h00000000;
    rd_cycle[ 2083] = 1'b0;  wr_cycle[ 2083] = 1'b1;  addr_rom[ 2083]='h00000170;  wr_data_rom[ 2083]='h000009d8;
    rd_cycle[ 2084] = 1'b1;  wr_cycle[ 2084] = 1'b0;  addr_rom[ 2084]='h00000bfc;  wr_data_rom[ 2084]='h00000000;
    rd_cycle[ 2085] = 1'b1;  wr_cycle[ 2085] = 1'b0;  addr_rom[ 2085]='h000001f0;  wr_data_rom[ 2085]='h00000000;
    rd_cycle[ 2086] = 1'b0;  wr_cycle[ 2086] = 1'b1;  addr_rom[ 2086]='h000004f0;  wr_data_rom[ 2086]='h00000637;
    rd_cycle[ 2087] = 1'b0;  wr_cycle[ 2087] = 1'b1;  addr_rom[ 2087]='h0000054c;  wr_data_rom[ 2087]='h00000255;
    rd_cycle[ 2088] = 1'b1;  wr_cycle[ 2088] = 1'b0;  addr_rom[ 2088]='h00000178;  wr_data_rom[ 2088]='h00000000;
    rd_cycle[ 2089] = 1'b1;  wr_cycle[ 2089] = 1'b0;  addr_rom[ 2089]='h00000a3c;  wr_data_rom[ 2089]='h00000000;
    rd_cycle[ 2090] = 1'b0;  wr_cycle[ 2090] = 1'b1;  addr_rom[ 2090]='h00000c38;  wr_data_rom[ 2090]='h00000734;
    rd_cycle[ 2091] = 1'b0;  wr_cycle[ 2091] = 1'b1;  addr_rom[ 2091]='h00000c1c;  wr_data_rom[ 2091]='h000006db;
    rd_cycle[ 2092] = 1'b1;  wr_cycle[ 2092] = 1'b0;  addr_rom[ 2092]='h000008dc;  wr_data_rom[ 2092]='h00000000;
    rd_cycle[ 2093] = 1'b0;  wr_cycle[ 2093] = 1'b1;  addr_rom[ 2093]='h00000134;  wr_data_rom[ 2093]='h00000b3d;
    rd_cycle[ 2094] = 1'b0;  wr_cycle[ 2094] = 1'b1;  addr_rom[ 2094]='h00000910;  wr_data_rom[ 2094]='h000008b0;
    rd_cycle[ 2095] = 1'b1;  wr_cycle[ 2095] = 1'b0;  addr_rom[ 2095]='h000004ac;  wr_data_rom[ 2095]='h00000000;
    rd_cycle[ 2096] = 1'b0;  wr_cycle[ 2096] = 1'b1;  addr_rom[ 2096]='h00000ca0;  wr_data_rom[ 2096]='h00000111;
    rd_cycle[ 2097] = 1'b1;  wr_cycle[ 2097] = 1'b0;  addr_rom[ 2097]='h00000c78;  wr_data_rom[ 2097]='h00000000;
    rd_cycle[ 2098] = 1'b0;  wr_cycle[ 2098] = 1'b1;  addr_rom[ 2098]='h00000138;  wr_data_rom[ 2098]='h000008ad;
    rd_cycle[ 2099] = 1'b0;  wr_cycle[ 2099] = 1'b1;  addr_rom[ 2099]='h000003fc;  wr_data_rom[ 2099]='h00000431;
    rd_cycle[ 2100] = 1'b0;  wr_cycle[ 2100] = 1'b1;  addr_rom[ 2100]='h00000c2c;  wr_data_rom[ 2100]='h00000d53;
    rd_cycle[ 2101] = 1'b1;  wr_cycle[ 2101] = 1'b0;  addr_rom[ 2101]='h00000f04;  wr_data_rom[ 2101]='h00000000;
    rd_cycle[ 2102] = 1'b0;  wr_cycle[ 2102] = 1'b1;  addr_rom[ 2102]='h00000d14;  wr_data_rom[ 2102]='h00000acb;
    rd_cycle[ 2103] = 1'b1;  wr_cycle[ 2103] = 1'b0;  addr_rom[ 2103]='h00000b00;  wr_data_rom[ 2103]='h00000000;
    rd_cycle[ 2104] = 1'b0;  wr_cycle[ 2104] = 1'b1;  addr_rom[ 2104]='h00000144;  wr_data_rom[ 2104]='h00000ed0;
    rd_cycle[ 2105] = 1'b0;  wr_cycle[ 2105] = 1'b1;  addr_rom[ 2105]='h00000ba0;  wr_data_rom[ 2105]='h00000383;
    rd_cycle[ 2106] = 1'b0;  wr_cycle[ 2106] = 1'b1;  addr_rom[ 2106]='h00000628;  wr_data_rom[ 2106]='h00000c91;
    rd_cycle[ 2107] = 1'b1;  wr_cycle[ 2107] = 1'b0;  addr_rom[ 2107]='h000004ec;  wr_data_rom[ 2107]='h00000000;
    rd_cycle[ 2108] = 1'b0;  wr_cycle[ 2108] = 1'b1;  addr_rom[ 2108]='h0000070c;  wr_data_rom[ 2108]='h00000458;
    rd_cycle[ 2109] = 1'b1;  wr_cycle[ 2109] = 1'b0;  addr_rom[ 2109]='h00000f84;  wr_data_rom[ 2109]='h00000000;
    rd_cycle[ 2110] = 1'b1;  wr_cycle[ 2110] = 1'b0;  addr_rom[ 2110]='h0000011c;  wr_data_rom[ 2110]='h00000000;
    rd_cycle[ 2111] = 1'b1;  wr_cycle[ 2111] = 1'b0;  addr_rom[ 2111]='h00000900;  wr_data_rom[ 2111]='h00000000;
    rd_cycle[ 2112] = 1'b1;  wr_cycle[ 2112] = 1'b0;  addr_rom[ 2112]='h00000c40;  wr_data_rom[ 2112]='h00000000;
    rd_cycle[ 2113] = 1'b1;  wr_cycle[ 2113] = 1'b0;  addr_rom[ 2113]='h00000198;  wr_data_rom[ 2113]='h00000000;
    rd_cycle[ 2114] = 1'b0;  wr_cycle[ 2114] = 1'b1;  addr_rom[ 2114]='h00000c28;  wr_data_rom[ 2114]='h00000549;
    rd_cycle[ 2115] = 1'b0;  wr_cycle[ 2115] = 1'b1;  addr_rom[ 2115]='h0000044c;  wr_data_rom[ 2115]='h00000a3c;
    rd_cycle[ 2116] = 1'b0;  wr_cycle[ 2116] = 1'b1;  addr_rom[ 2116]='h00000a80;  wr_data_rom[ 2116]='h00000349;
    rd_cycle[ 2117] = 1'b0;  wr_cycle[ 2117] = 1'b1;  addr_rom[ 2117]='h00000c00;  wr_data_rom[ 2117]='h0000046a;
    rd_cycle[ 2118] = 1'b0;  wr_cycle[ 2118] = 1'b1;  addr_rom[ 2118]='h000007c0;  wr_data_rom[ 2118]='h000007a3;
    rd_cycle[ 2119] = 1'b0;  wr_cycle[ 2119] = 1'b1;  addr_rom[ 2119]='h00000818;  wr_data_rom[ 2119]='h000007f7;
    rd_cycle[ 2120] = 1'b0;  wr_cycle[ 2120] = 1'b1;  addr_rom[ 2120]='h00000220;  wr_data_rom[ 2120]='h000008bf;
    rd_cycle[ 2121] = 1'b0;  wr_cycle[ 2121] = 1'b1;  addr_rom[ 2121]='h000004a4;  wr_data_rom[ 2121]='h0000065e;
    rd_cycle[ 2122] = 1'b0;  wr_cycle[ 2122] = 1'b1;  addr_rom[ 2122]='h00000a84;  wr_data_rom[ 2122]='h00000959;
    rd_cycle[ 2123] = 1'b1;  wr_cycle[ 2123] = 1'b0;  addr_rom[ 2123]='h00000910;  wr_data_rom[ 2123]='h00000000;
    rd_cycle[ 2124] = 1'b0;  wr_cycle[ 2124] = 1'b1;  addr_rom[ 2124]='h00000340;  wr_data_rom[ 2124]='h00000dff;
    rd_cycle[ 2125] = 1'b0;  wr_cycle[ 2125] = 1'b1;  addr_rom[ 2125]='h0000033c;  wr_data_rom[ 2125]='h0000043e;
    rd_cycle[ 2126] = 1'b0;  wr_cycle[ 2126] = 1'b1;  addr_rom[ 2126]='h0000096c;  wr_data_rom[ 2126]='h0000059a;
    rd_cycle[ 2127] = 1'b0;  wr_cycle[ 2127] = 1'b1;  addr_rom[ 2127]='h00000ae0;  wr_data_rom[ 2127]='h00000357;
    rd_cycle[ 2128] = 1'b0;  wr_cycle[ 2128] = 1'b1;  addr_rom[ 2128]='h00000548;  wr_data_rom[ 2128]='h00000b44;
    rd_cycle[ 2129] = 1'b1;  wr_cycle[ 2129] = 1'b0;  addr_rom[ 2129]='h00000e14;  wr_data_rom[ 2129]='h00000000;
    rd_cycle[ 2130] = 1'b1;  wr_cycle[ 2130] = 1'b0;  addr_rom[ 2130]='h000008a0;  wr_data_rom[ 2130]='h00000000;
    rd_cycle[ 2131] = 1'b1;  wr_cycle[ 2131] = 1'b0;  addr_rom[ 2131]='h00000a50;  wr_data_rom[ 2131]='h00000000;
    rd_cycle[ 2132] = 1'b0;  wr_cycle[ 2132] = 1'b1;  addr_rom[ 2132]='h0000070c;  wr_data_rom[ 2132]='h000000c1;
    rd_cycle[ 2133] = 1'b0;  wr_cycle[ 2133] = 1'b1;  addr_rom[ 2133]='h00000418;  wr_data_rom[ 2133]='h0000053c;
    rd_cycle[ 2134] = 1'b0;  wr_cycle[ 2134] = 1'b1;  addr_rom[ 2134]='h00000944;  wr_data_rom[ 2134]='h000006fa;
    rd_cycle[ 2135] = 1'b0;  wr_cycle[ 2135] = 1'b1;  addr_rom[ 2135]='h00000924;  wr_data_rom[ 2135]='h00000a33;
    rd_cycle[ 2136] = 1'b0;  wr_cycle[ 2136] = 1'b1;  addr_rom[ 2136]='h00000104;  wr_data_rom[ 2136]='h000009fc;
    rd_cycle[ 2137] = 1'b0;  wr_cycle[ 2137] = 1'b1;  addr_rom[ 2137]='h00000b64;  wr_data_rom[ 2137]='h00000a61;
    rd_cycle[ 2138] = 1'b1;  wr_cycle[ 2138] = 1'b0;  addr_rom[ 2138]='h0000031c;  wr_data_rom[ 2138]='h00000000;
    rd_cycle[ 2139] = 1'b0;  wr_cycle[ 2139] = 1'b1;  addr_rom[ 2139]='h00000e44;  wr_data_rom[ 2139]='h0000098f;
    rd_cycle[ 2140] = 1'b0;  wr_cycle[ 2140] = 1'b1;  addr_rom[ 2140]='h000001d8;  wr_data_rom[ 2140]='h00000c08;
    rd_cycle[ 2141] = 1'b1;  wr_cycle[ 2141] = 1'b0;  addr_rom[ 2141]='h00000d3c;  wr_data_rom[ 2141]='h00000000;
    rd_cycle[ 2142] = 1'b1;  wr_cycle[ 2142] = 1'b0;  addr_rom[ 2142]='h000005a8;  wr_data_rom[ 2142]='h00000000;
    rd_cycle[ 2143] = 1'b0;  wr_cycle[ 2143] = 1'b1;  addr_rom[ 2143]='h000000ac;  wr_data_rom[ 2143]='h00000899;
    rd_cycle[ 2144] = 1'b0;  wr_cycle[ 2144] = 1'b1;  addr_rom[ 2144]='h00000304;  wr_data_rom[ 2144]='h00000d78;
    rd_cycle[ 2145] = 1'b0;  wr_cycle[ 2145] = 1'b1;  addr_rom[ 2145]='h00000490;  wr_data_rom[ 2145]='h000006d5;
    rd_cycle[ 2146] = 1'b1;  wr_cycle[ 2146] = 1'b0;  addr_rom[ 2146]='h00000a98;  wr_data_rom[ 2146]='h00000000;
    rd_cycle[ 2147] = 1'b1;  wr_cycle[ 2147] = 1'b0;  addr_rom[ 2147]='h00000c54;  wr_data_rom[ 2147]='h00000000;
    rd_cycle[ 2148] = 1'b1;  wr_cycle[ 2148] = 1'b0;  addr_rom[ 2148]='h00000510;  wr_data_rom[ 2148]='h00000000;
    rd_cycle[ 2149] = 1'b0;  wr_cycle[ 2149] = 1'b1;  addr_rom[ 2149]='h00000e30;  wr_data_rom[ 2149]='h00000005;
    rd_cycle[ 2150] = 1'b0;  wr_cycle[ 2150] = 1'b1;  addr_rom[ 2150]='h00000460;  wr_data_rom[ 2150]='h00000c9b;
    rd_cycle[ 2151] = 1'b1;  wr_cycle[ 2151] = 1'b0;  addr_rom[ 2151]='h00000aac;  wr_data_rom[ 2151]='h00000000;
    rd_cycle[ 2152] = 1'b1;  wr_cycle[ 2152] = 1'b0;  addr_rom[ 2152]='h00000860;  wr_data_rom[ 2152]='h00000000;
    rd_cycle[ 2153] = 1'b0;  wr_cycle[ 2153] = 1'b1;  addr_rom[ 2153]='h00000cc0;  wr_data_rom[ 2153]='h000004e4;
    rd_cycle[ 2154] = 1'b0;  wr_cycle[ 2154] = 1'b1;  addr_rom[ 2154]='h00000260;  wr_data_rom[ 2154]='h00000443;
    rd_cycle[ 2155] = 1'b0;  wr_cycle[ 2155] = 1'b1;  addr_rom[ 2155]='h000005d0;  wr_data_rom[ 2155]='h000001c5;
    rd_cycle[ 2156] = 1'b1;  wr_cycle[ 2156] = 1'b0;  addr_rom[ 2156]='h00000aa8;  wr_data_rom[ 2156]='h00000000;
    rd_cycle[ 2157] = 1'b0;  wr_cycle[ 2157] = 1'b1;  addr_rom[ 2157]='h00000f78;  wr_data_rom[ 2157]='h00000c84;
    rd_cycle[ 2158] = 1'b1;  wr_cycle[ 2158] = 1'b0;  addr_rom[ 2158]='h0000081c;  wr_data_rom[ 2158]='h00000000;
    rd_cycle[ 2159] = 1'b0;  wr_cycle[ 2159] = 1'b1;  addr_rom[ 2159]='h0000064c;  wr_data_rom[ 2159]='h0000052d;
    rd_cycle[ 2160] = 1'b0;  wr_cycle[ 2160] = 1'b1;  addr_rom[ 2160]='h000005ec;  wr_data_rom[ 2160]='h00000229;
    rd_cycle[ 2161] = 1'b0;  wr_cycle[ 2161] = 1'b1;  addr_rom[ 2161]='h00000e7c;  wr_data_rom[ 2161]='h0000047a;
    rd_cycle[ 2162] = 1'b1;  wr_cycle[ 2162] = 1'b0;  addr_rom[ 2162]='h00000f30;  wr_data_rom[ 2162]='h00000000;
    rd_cycle[ 2163] = 1'b0;  wr_cycle[ 2163] = 1'b1;  addr_rom[ 2163]='h00000694;  wr_data_rom[ 2163]='h000007e2;
    rd_cycle[ 2164] = 1'b0;  wr_cycle[ 2164] = 1'b1;  addr_rom[ 2164]='h00000af4;  wr_data_rom[ 2164]='h00000985;
    rd_cycle[ 2165] = 1'b0;  wr_cycle[ 2165] = 1'b1;  addr_rom[ 2165]='h00000c54;  wr_data_rom[ 2165]='h000004e2;
    rd_cycle[ 2166] = 1'b0;  wr_cycle[ 2166] = 1'b1;  addr_rom[ 2166]='h00000588;  wr_data_rom[ 2166]='h0000056a;
    rd_cycle[ 2167] = 1'b1;  wr_cycle[ 2167] = 1'b0;  addr_rom[ 2167]='h000002c8;  wr_data_rom[ 2167]='h00000000;
    rd_cycle[ 2168] = 1'b0;  wr_cycle[ 2168] = 1'b1;  addr_rom[ 2168]='h00000908;  wr_data_rom[ 2168]='h0000065e;
    rd_cycle[ 2169] = 1'b0;  wr_cycle[ 2169] = 1'b1;  addr_rom[ 2169]='h00000720;  wr_data_rom[ 2169]='h00000c10;
    rd_cycle[ 2170] = 1'b1;  wr_cycle[ 2170] = 1'b0;  addr_rom[ 2170]='h00000568;  wr_data_rom[ 2170]='h00000000;
    rd_cycle[ 2171] = 1'b1;  wr_cycle[ 2171] = 1'b0;  addr_rom[ 2171]='h00000290;  wr_data_rom[ 2171]='h00000000;
    rd_cycle[ 2172] = 1'b0;  wr_cycle[ 2172] = 1'b1;  addr_rom[ 2172]='h00000014;  wr_data_rom[ 2172]='h00000963;
    rd_cycle[ 2173] = 1'b1;  wr_cycle[ 2173] = 1'b0;  addr_rom[ 2173]='h00000660;  wr_data_rom[ 2173]='h00000000;
    rd_cycle[ 2174] = 1'b1;  wr_cycle[ 2174] = 1'b0;  addr_rom[ 2174]='h00000a80;  wr_data_rom[ 2174]='h00000000;
    rd_cycle[ 2175] = 1'b1;  wr_cycle[ 2175] = 1'b0;  addr_rom[ 2175]='h00000340;  wr_data_rom[ 2175]='h00000000;
    rd_cycle[ 2176] = 1'b0;  wr_cycle[ 2176] = 1'b1;  addr_rom[ 2176]='h00000a38;  wr_data_rom[ 2176]='h00000f17;
    rd_cycle[ 2177] = 1'b0;  wr_cycle[ 2177] = 1'b1;  addr_rom[ 2177]='h00000848;  wr_data_rom[ 2177]='h0000043d;
    rd_cycle[ 2178] = 1'b1;  wr_cycle[ 2178] = 1'b0;  addr_rom[ 2178]='h00000d30;  wr_data_rom[ 2178]='h00000000;
    rd_cycle[ 2179] = 1'b0;  wr_cycle[ 2179] = 1'b1;  addr_rom[ 2179]='h00000384;  wr_data_rom[ 2179]='h0000034c;
    rd_cycle[ 2180] = 1'b0;  wr_cycle[ 2180] = 1'b1;  addr_rom[ 2180]='h00000330;  wr_data_rom[ 2180]='h000007e3;
    rd_cycle[ 2181] = 1'b0;  wr_cycle[ 2181] = 1'b1;  addr_rom[ 2181]='h000000ac;  wr_data_rom[ 2181]='h000009a3;
    rd_cycle[ 2182] = 1'b0;  wr_cycle[ 2182] = 1'b1;  addr_rom[ 2182]='h000007c0;  wr_data_rom[ 2182]='h000005b2;
    rd_cycle[ 2183] = 1'b1;  wr_cycle[ 2183] = 1'b0;  addr_rom[ 2183]='h00000228;  wr_data_rom[ 2183]='h00000000;
    rd_cycle[ 2184] = 1'b0;  wr_cycle[ 2184] = 1'b1;  addr_rom[ 2184]='h000002a8;  wr_data_rom[ 2184]='h00000e3f;
    rd_cycle[ 2185] = 1'b1;  wr_cycle[ 2185] = 1'b0;  addr_rom[ 2185]='h000007c8;  wr_data_rom[ 2185]='h00000000;
    rd_cycle[ 2186] = 1'b0;  wr_cycle[ 2186] = 1'b1;  addr_rom[ 2186]='h0000049c;  wr_data_rom[ 2186]='h00000dcf;
    rd_cycle[ 2187] = 1'b0;  wr_cycle[ 2187] = 1'b1;  addr_rom[ 2187]='h00000604;  wr_data_rom[ 2187]='h00000839;
    rd_cycle[ 2188] = 1'b1;  wr_cycle[ 2188] = 1'b0;  addr_rom[ 2188]='h0000057c;  wr_data_rom[ 2188]='h00000000;
    rd_cycle[ 2189] = 1'b1;  wr_cycle[ 2189] = 1'b0;  addr_rom[ 2189]='h00000524;  wr_data_rom[ 2189]='h00000000;
    rd_cycle[ 2190] = 1'b1;  wr_cycle[ 2190] = 1'b0;  addr_rom[ 2190]='h00000df0;  wr_data_rom[ 2190]='h00000000;
    rd_cycle[ 2191] = 1'b0;  wr_cycle[ 2191] = 1'b1;  addr_rom[ 2191]='h0000019c;  wr_data_rom[ 2191]='h00000b3f;
    rd_cycle[ 2192] = 1'b0;  wr_cycle[ 2192] = 1'b1;  addr_rom[ 2192]='h00000110;  wr_data_rom[ 2192]='h00000da6;
    rd_cycle[ 2193] = 1'b0;  wr_cycle[ 2193] = 1'b1;  addr_rom[ 2193]='h00000b78;  wr_data_rom[ 2193]='h00000c58;
    rd_cycle[ 2194] = 1'b0;  wr_cycle[ 2194] = 1'b1;  addr_rom[ 2194]='h0000084c;  wr_data_rom[ 2194]='h000002de;
    rd_cycle[ 2195] = 1'b0;  wr_cycle[ 2195] = 1'b1;  addr_rom[ 2195]='h00000e80;  wr_data_rom[ 2195]='h0000014f;
    rd_cycle[ 2196] = 1'b0;  wr_cycle[ 2196] = 1'b1;  addr_rom[ 2196]='h00000458;  wr_data_rom[ 2196]='h000007e9;
    rd_cycle[ 2197] = 1'b1;  wr_cycle[ 2197] = 1'b0;  addr_rom[ 2197]='h00000424;  wr_data_rom[ 2197]='h00000000;
    rd_cycle[ 2198] = 1'b1;  wr_cycle[ 2198] = 1'b0;  addr_rom[ 2198]='h00000f6c;  wr_data_rom[ 2198]='h00000000;
    rd_cycle[ 2199] = 1'b0;  wr_cycle[ 2199] = 1'b1;  addr_rom[ 2199]='h00000614;  wr_data_rom[ 2199]='h00000421;
    rd_cycle[ 2200] = 1'b0;  wr_cycle[ 2200] = 1'b1;  addr_rom[ 2200]='h00000148;  wr_data_rom[ 2200]='h00000d87;
    rd_cycle[ 2201] = 1'b0;  wr_cycle[ 2201] = 1'b1;  addr_rom[ 2201]='h00000938;  wr_data_rom[ 2201]='h000008af;
    rd_cycle[ 2202] = 1'b1;  wr_cycle[ 2202] = 1'b0;  addr_rom[ 2202]='h00000120;  wr_data_rom[ 2202]='h00000000;
    rd_cycle[ 2203] = 1'b1;  wr_cycle[ 2203] = 1'b0;  addr_rom[ 2203]='h000005bc;  wr_data_rom[ 2203]='h00000000;
    rd_cycle[ 2204] = 1'b0;  wr_cycle[ 2204] = 1'b1;  addr_rom[ 2204]='h00000278;  wr_data_rom[ 2204]='h00000b35;
    rd_cycle[ 2205] = 1'b1;  wr_cycle[ 2205] = 1'b0;  addr_rom[ 2205]='h00000004;  wr_data_rom[ 2205]='h00000000;
    rd_cycle[ 2206] = 1'b0;  wr_cycle[ 2206] = 1'b1;  addr_rom[ 2206]='h00000ee4;  wr_data_rom[ 2206]='h0000091f;
    rd_cycle[ 2207] = 1'b0;  wr_cycle[ 2207] = 1'b1;  addr_rom[ 2207]='h00000af8;  wr_data_rom[ 2207]='h0000078e;
    rd_cycle[ 2208] = 1'b0;  wr_cycle[ 2208] = 1'b1;  addr_rom[ 2208]='h00000ee0;  wr_data_rom[ 2208]='h000003c8;
    rd_cycle[ 2209] = 1'b0;  wr_cycle[ 2209] = 1'b1;  addr_rom[ 2209]='h000005d8;  wr_data_rom[ 2209]='h00000552;
    rd_cycle[ 2210] = 1'b0;  wr_cycle[ 2210] = 1'b1;  addr_rom[ 2210]='h00000098;  wr_data_rom[ 2210]='h000007de;
    rd_cycle[ 2211] = 1'b0;  wr_cycle[ 2211] = 1'b1;  addr_rom[ 2211]='h00000208;  wr_data_rom[ 2211]='h00000a80;
    rd_cycle[ 2212] = 1'b1;  wr_cycle[ 2212] = 1'b0;  addr_rom[ 2212]='h00000654;  wr_data_rom[ 2212]='h00000000;
    rd_cycle[ 2213] = 1'b1;  wr_cycle[ 2213] = 1'b0;  addr_rom[ 2213]='h00000c18;  wr_data_rom[ 2213]='h00000000;
    rd_cycle[ 2214] = 1'b1;  wr_cycle[ 2214] = 1'b0;  addr_rom[ 2214]='h000001a4;  wr_data_rom[ 2214]='h00000000;
    rd_cycle[ 2215] = 1'b1;  wr_cycle[ 2215] = 1'b0;  addr_rom[ 2215]='h00000d08;  wr_data_rom[ 2215]='h00000000;
    rd_cycle[ 2216] = 1'b1;  wr_cycle[ 2216] = 1'b0;  addr_rom[ 2216]='h00000aac;  wr_data_rom[ 2216]='h00000000;
    rd_cycle[ 2217] = 1'b1;  wr_cycle[ 2217] = 1'b0;  addr_rom[ 2217]='h000000c4;  wr_data_rom[ 2217]='h00000000;
    rd_cycle[ 2218] = 1'b1;  wr_cycle[ 2218] = 1'b0;  addr_rom[ 2218]='h00000ec0;  wr_data_rom[ 2218]='h00000000;
    rd_cycle[ 2219] = 1'b0;  wr_cycle[ 2219] = 1'b1;  addr_rom[ 2219]='h00000600;  wr_data_rom[ 2219]='h00000e9d;
    rd_cycle[ 2220] = 1'b1;  wr_cycle[ 2220] = 1'b0;  addr_rom[ 2220]='h000007c8;  wr_data_rom[ 2220]='h00000000;
    rd_cycle[ 2221] = 1'b0;  wr_cycle[ 2221] = 1'b1;  addr_rom[ 2221]='h0000028c;  wr_data_rom[ 2221]='h00000a86;
    rd_cycle[ 2222] = 1'b1;  wr_cycle[ 2222] = 1'b0;  addr_rom[ 2222]='h0000054c;  wr_data_rom[ 2222]='h00000000;
    rd_cycle[ 2223] = 1'b0;  wr_cycle[ 2223] = 1'b1;  addr_rom[ 2223]='h0000009c;  wr_data_rom[ 2223]='h000001ff;
    rd_cycle[ 2224] = 1'b1;  wr_cycle[ 2224] = 1'b0;  addr_rom[ 2224]='h0000061c;  wr_data_rom[ 2224]='h00000000;
    rd_cycle[ 2225] = 1'b0;  wr_cycle[ 2225] = 1'b1;  addr_rom[ 2225]='h00000910;  wr_data_rom[ 2225]='h00000ee5;
    rd_cycle[ 2226] = 1'b0;  wr_cycle[ 2226] = 1'b1;  addr_rom[ 2226]='h00000e6c;  wr_data_rom[ 2226]='h00000d92;
    rd_cycle[ 2227] = 1'b1;  wr_cycle[ 2227] = 1'b0;  addr_rom[ 2227]='h000009d4;  wr_data_rom[ 2227]='h00000000;
    rd_cycle[ 2228] = 1'b1;  wr_cycle[ 2228] = 1'b0;  addr_rom[ 2228]='h00000920;  wr_data_rom[ 2228]='h00000000;
    rd_cycle[ 2229] = 1'b0;  wr_cycle[ 2229] = 1'b1;  addr_rom[ 2229]='h00000f2c;  wr_data_rom[ 2229]='h0000006f;
    rd_cycle[ 2230] = 1'b0;  wr_cycle[ 2230] = 1'b1;  addr_rom[ 2230]='h000004d8;  wr_data_rom[ 2230]='h00000edf;
    rd_cycle[ 2231] = 1'b1;  wr_cycle[ 2231] = 1'b0;  addr_rom[ 2231]='h0000098c;  wr_data_rom[ 2231]='h00000000;
    rd_cycle[ 2232] = 1'b0;  wr_cycle[ 2232] = 1'b1;  addr_rom[ 2232]='h00000670;  wr_data_rom[ 2232]='h00000a80;
    rd_cycle[ 2233] = 1'b1;  wr_cycle[ 2233] = 1'b0;  addr_rom[ 2233]='h00000550;  wr_data_rom[ 2233]='h00000000;
    rd_cycle[ 2234] = 1'b0;  wr_cycle[ 2234] = 1'b1;  addr_rom[ 2234]='h00000bd4;  wr_data_rom[ 2234]='h000003be;
    rd_cycle[ 2235] = 1'b0;  wr_cycle[ 2235] = 1'b1;  addr_rom[ 2235]='h0000096c;  wr_data_rom[ 2235]='h00000168;
    rd_cycle[ 2236] = 1'b0;  wr_cycle[ 2236] = 1'b1;  addr_rom[ 2236]='h00000d20;  wr_data_rom[ 2236]='h00000c0b;
    rd_cycle[ 2237] = 1'b1;  wr_cycle[ 2237] = 1'b0;  addr_rom[ 2237]='h00000b08;  wr_data_rom[ 2237]='h00000000;
    rd_cycle[ 2238] = 1'b1;  wr_cycle[ 2238] = 1'b0;  addr_rom[ 2238]='h00000334;  wr_data_rom[ 2238]='h00000000;
    rd_cycle[ 2239] = 1'b0;  wr_cycle[ 2239] = 1'b1;  addr_rom[ 2239]='h00000284;  wr_data_rom[ 2239]='h00000ce3;
    rd_cycle[ 2240] = 1'b0;  wr_cycle[ 2240] = 1'b1;  addr_rom[ 2240]='h000003f0;  wr_data_rom[ 2240]='h000005c0;
    rd_cycle[ 2241] = 1'b0;  wr_cycle[ 2241] = 1'b1;  addr_rom[ 2241]='h000005b8;  wr_data_rom[ 2241]='h00000820;
    rd_cycle[ 2242] = 1'b1;  wr_cycle[ 2242] = 1'b0;  addr_rom[ 2242]='h000009a4;  wr_data_rom[ 2242]='h00000000;
    rd_cycle[ 2243] = 1'b1;  wr_cycle[ 2243] = 1'b0;  addr_rom[ 2243]='h00000178;  wr_data_rom[ 2243]='h00000000;
    rd_cycle[ 2244] = 1'b0;  wr_cycle[ 2244] = 1'b1;  addr_rom[ 2244]='h00000c44;  wr_data_rom[ 2244]='h00000649;
    rd_cycle[ 2245] = 1'b0;  wr_cycle[ 2245] = 1'b1;  addr_rom[ 2245]='h0000097c;  wr_data_rom[ 2245]='h00000786;
    rd_cycle[ 2246] = 1'b0;  wr_cycle[ 2246] = 1'b1;  addr_rom[ 2246]='h00000ca8;  wr_data_rom[ 2246]='h000007b3;
    rd_cycle[ 2247] = 1'b1;  wr_cycle[ 2247] = 1'b0;  addr_rom[ 2247]='h00000f48;  wr_data_rom[ 2247]='h00000000;
    rd_cycle[ 2248] = 1'b0;  wr_cycle[ 2248] = 1'b1;  addr_rom[ 2248]='h00000ae0;  wr_data_rom[ 2248]='h00000d64;
    rd_cycle[ 2249] = 1'b0;  wr_cycle[ 2249] = 1'b1;  addr_rom[ 2249]='h00000c64;  wr_data_rom[ 2249]='h000007c0;
    rd_cycle[ 2250] = 1'b0;  wr_cycle[ 2250] = 1'b1;  addr_rom[ 2250]='h0000024c;  wr_data_rom[ 2250]='h00000f13;
    rd_cycle[ 2251] = 1'b1;  wr_cycle[ 2251] = 1'b0;  addr_rom[ 2251]='h00000660;  wr_data_rom[ 2251]='h00000000;
    rd_cycle[ 2252] = 1'b0;  wr_cycle[ 2252] = 1'b1;  addr_rom[ 2252]='h0000061c;  wr_data_rom[ 2252]='h00000ecc;
    rd_cycle[ 2253] = 1'b1;  wr_cycle[ 2253] = 1'b0;  addr_rom[ 2253]='h00000c24;  wr_data_rom[ 2253]='h00000000;
    rd_cycle[ 2254] = 1'b0;  wr_cycle[ 2254] = 1'b1;  addr_rom[ 2254]='h000004d0;  wr_data_rom[ 2254]='h00000c44;
    rd_cycle[ 2255] = 1'b0;  wr_cycle[ 2255] = 1'b1;  addr_rom[ 2255]='h0000079c;  wr_data_rom[ 2255]='h00000a5e;
    rd_cycle[ 2256] = 1'b1;  wr_cycle[ 2256] = 1'b0;  addr_rom[ 2256]='h0000049c;  wr_data_rom[ 2256]='h00000000;
    rd_cycle[ 2257] = 1'b0;  wr_cycle[ 2257] = 1'b1;  addr_rom[ 2257]='h00000b14;  wr_data_rom[ 2257]='h00000de9;
    rd_cycle[ 2258] = 1'b1;  wr_cycle[ 2258] = 1'b0;  addr_rom[ 2258]='h00000834;  wr_data_rom[ 2258]='h00000000;
    rd_cycle[ 2259] = 1'b0;  wr_cycle[ 2259] = 1'b1;  addr_rom[ 2259]='h00000dc4;  wr_data_rom[ 2259]='h0000081b;
    rd_cycle[ 2260] = 1'b0;  wr_cycle[ 2260] = 1'b1;  addr_rom[ 2260]='h00000724;  wr_data_rom[ 2260]='h0000034d;
    rd_cycle[ 2261] = 1'b1;  wr_cycle[ 2261] = 1'b0;  addr_rom[ 2261]='h00000a30;  wr_data_rom[ 2261]='h00000000;
    rd_cycle[ 2262] = 1'b0;  wr_cycle[ 2262] = 1'b1;  addr_rom[ 2262]='h00000ca4;  wr_data_rom[ 2262]='h00000335;
    rd_cycle[ 2263] = 1'b1;  wr_cycle[ 2263] = 1'b0;  addr_rom[ 2263]='h000006bc;  wr_data_rom[ 2263]='h00000000;
    rd_cycle[ 2264] = 1'b0;  wr_cycle[ 2264] = 1'b1;  addr_rom[ 2264]='h000007c0;  wr_data_rom[ 2264]='h0000035b;
    rd_cycle[ 2265] = 1'b1;  wr_cycle[ 2265] = 1'b0;  addr_rom[ 2265]='h00000610;  wr_data_rom[ 2265]='h00000000;
    rd_cycle[ 2266] = 1'b1;  wr_cycle[ 2266] = 1'b0;  addr_rom[ 2266]='h0000034c;  wr_data_rom[ 2266]='h00000000;
    rd_cycle[ 2267] = 1'b1;  wr_cycle[ 2267] = 1'b0;  addr_rom[ 2267]='h00000f6c;  wr_data_rom[ 2267]='h00000000;
    rd_cycle[ 2268] = 1'b0;  wr_cycle[ 2268] = 1'b1;  addr_rom[ 2268]='h00000a24;  wr_data_rom[ 2268]='h00000b72;
    rd_cycle[ 2269] = 1'b0;  wr_cycle[ 2269] = 1'b1;  addr_rom[ 2269]='h00000134;  wr_data_rom[ 2269]='h00000b7c;
    rd_cycle[ 2270] = 1'b1;  wr_cycle[ 2270] = 1'b0;  addr_rom[ 2270]='h00000974;  wr_data_rom[ 2270]='h00000000;
    rd_cycle[ 2271] = 1'b1;  wr_cycle[ 2271] = 1'b0;  addr_rom[ 2271]='h000007d0;  wr_data_rom[ 2271]='h00000000;
    rd_cycle[ 2272] = 1'b1;  wr_cycle[ 2272] = 1'b0;  addr_rom[ 2272]='h00000bf8;  wr_data_rom[ 2272]='h00000000;
    rd_cycle[ 2273] = 1'b1;  wr_cycle[ 2273] = 1'b0;  addr_rom[ 2273]='h00000c2c;  wr_data_rom[ 2273]='h00000000;
    rd_cycle[ 2274] = 1'b0;  wr_cycle[ 2274] = 1'b1;  addr_rom[ 2274]='h000005c8;  wr_data_rom[ 2274]='h0000055d;
    rd_cycle[ 2275] = 1'b1;  wr_cycle[ 2275] = 1'b0;  addr_rom[ 2275]='h00000e74;  wr_data_rom[ 2275]='h00000000;
    rd_cycle[ 2276] = 1'b0;  wr_cycle[ 2276] = 1'b1;  addr_rom[ 2276]='h00000eb8;  wr_data_rom[ 2276]='h000005d0;
    rd_cycle[ 2277] = 1'b0;  wr_cycle[ 2277] = 1'b1;  addr_rom[ 2277]='h000001e8;  wr_data_rom[ 2277]='h000007b8;
    rd_cycle[ 2278] = 1'b1;  wr_cycle[ 2278] = 1'b0;  addr_rom[ 2278]='h0000091c;  wr_data_rom[ 2278]='h00000000;
    rd_cycle[ 2279] = 1'b0;  wr_cycle[ 2279] = 1'b1;  addr_rom[ 2279]='h000008f0;  wr_data_rom[ 2279]='h00000b45;
    rd_cycle[ 2280] = 1'b0;  wr_cycle[ 2280] = 1'b1;  addr_rom[ 2280]='h00000f34;  wr_data_rom[ 2280]='h000002f1;
    rd_cycle[ 2281] = 1'b1;  wr_cycle[ 2281] = 1'b0;  addr_rom[ 2281]='h0000058c;  wr_data_rom[ 2281]='h00000000;
    rd_cycle[ 2282] = 1'b0;  wr_cycle[ 2282] = 1'b1;  addr_rom[ 2282]='h000000d4;  wr_data_rom[ 2282]='h00000f70;
    rd_cycle[ 2283] = 1'b1;  wr_cycle[ 2283] = 1'b0;  addr_rom[ 2283]='h000004c8;  wr_data_rom[ 2283]='h00000000;
    rd_cycle[ 2284] = 1'b0;  wr_cycle[ 2284] = 1'b1;  addr_rom[ 2284]='h00000458;  wr_data_rom[ 2284]='h00000429;
    rd_cycle[ 2285] = 1'b0;  wr_cycle[ 2285] = 1'b1;  addr_rom[ 2285]='h00000b9c;  wr_data_rom[ 2285]='h00000082;
    rd_cycle[ 2286] = 1'b0;  wr_cycle[ 2286] = 1'b1;  addr_rom[ 2286]='h00000d00;  wr_data_rom[ 2286]='h00000e91;
    rd_cycle[ 2287] = 1'b1;  wr_cycle[ 2287] = 1'b0;  addr_rom[ 2287]='h00000344;  wr_data_rom[ 2287]='h00000000;
    rd_cycle[ 2288] = 1'b1;  wr_cycle[ 2288] = 1'b0;  addr_rom[ 2288]='h0000038c;  wr_data_rom[ 2288]='h00000000;
    rd_cycle[ 2289] = 1'b0;  wr_cycle[ 2289] = 1'b1;  addr_rom[ 2289]='h00000be4;  wr_data_rom[ 2289]='h00000900;
    rd_cycle[ 2290] = 1'b0;  wr_cycle[ 2290] = 1'b1;  addr_rom[ 2290]='h00000744;  wr_data_rom[ 2290]='h000003bf;
    rd_cycle[ 2291] = 1'b0;  wr_cycle[ 2291] = 1'b1;  addr_rom[ 2291]='h00000e60;  wr_data_rom[ 2291]='h00000d68;
    rd_cycle[ 2292] = 1'b0;  wr_cycle[ 2292] = 1'b1;  addr_rom[ 2292]='h0000011c;  wr_data_rom[ 2292]='h0000061b;
    rd_cycle[ 2293] = 1'b1;  wr_cycle[ 2293] = 1'b0;  addr_rom[ 2293]='h00000d2c;  wr_data_rom[ 2293]='h00000000;
    rd_cycle[ 2294] = 1'b1;  wr_cycle[ 2294] = 1'b0;  addr_rom[ 2294]='h00000778;  wr_data_rom[ 2294]='h00000000;
    rd_cycle[ 2295] = 1'b1;  wr_cycle[ 2295] = 1'b0;  addr_rom[ 2295]='h00000b1c;  wr_data_rom[ 2295]='h00000000;
    rd_cycle[ 2296] = 1'b1;  wr_cycle[ 2296] = 1'b0;  addr_rom[ 2296]='h00000c8c;  wr_data_rom[ 2296]='h00000000;
    rd_cycle[ 2297] = 1'b1;  wr_cycle[ 2297] = 1'b0;  addr_rom[ 2297]='h00000938;  wr_data_rom[ 2297]='h00000000;
    rd_cycle[ 2298] = 1'b0;  wr_cycle[ 2298] = 1'b1;  addr_rom[ 2298]='h00000c24;  wr_data_rom[ 2298]='h000001c6;
    rd_cycle[ 2299] = 1'b1;  wr_cycle[ 2299] = 1'b0;  addr_rom[ 2299]='h00000e70;  wr_data_rom[ 2299]='h00000000;
    rd_cycle[ 2300] = 1'b1;  wr_cycle[ 2300] = 1'b0;  addr_rom[ 2300]='h00000d1c;  wr_data_rom[ 2300]='h00000000;
    rd_cycle[ 2301] = 1'b1;  wr_cycle[ 2301] = 1'b0;  addr_rom[ 2301]='h00000a74;  wr_data_rom[ 2301]='h00000000;
    rd_cycle[ 2302] = 1'b1;  wr_cycle[ 2302] = 1'b0;  addr_rom[ 2302]='h00000d48;  wr_data_rom[ 2302]='h00000000;
    rd_cycle[ 2303] = 1'b0;  wr_cycle[ 2303] = 1'b1;  addr_rom[ 2303]='h00000cb4;  wr_data_rom[ 2303]='h00000c61;
    rd_cycle[ 2304] = 1'b1;  wr_cycle[ 2304] = 1'b0;  addr_rom[ 2304]='h00000d14;  wr_data_rom[ 2304]='h00000000;
    rd_cycle[ 2305] = 1'b0;  wr_cycle[ 2305] = 1'b1;  addr_rom[ 2305]='h00000e58;  wr_data_rom[ 2305]='h000007ab;
    rd_cycle[ 2306] = 1'b1;  wr_cycle[ 2306] = 1'b0;  addr_rom[ 2306]='h00000714;  wr_data_rom[ 2306]='h00000000;
    rd_cycle[ 2307] = 1'b0;  wr_cycle[ 2307] = 1'b1;  addr_rom[ 2307]='h000007d8;  wr_data_rom[ 2307]='h00000618;
    rd_cycle[ 2308] = 1'b0;  wr_cycle[ 2308] = 1'b1;  addr_rom[ 2308]='h00000854;  wr_data_rom[ 2308]='h0000049e;
    rd_cycle[ 2309] = 1'b0;  wr_cycle[ 2309] = 1'b1;  addr_rom[ 2309]='h00000a7c;  wr_data_rom[ 2309]='h0000075b;
    rd_cycle[ 2310] = 1'b1;  wr_cycle[ 2310] = 1'b0;  addr_rom[ 2310]='h00000a68;  wr_data_rom[ 2310]='h00000000;
    rd_cycle[ 2311] = 1'b1;  wr_cycle[ 2311] = 1'b0;  addr_rom[ 2311]='h00000540;  wr_data_rom[ 2311]='h00000000;
    rd_cycle[ 2312] = 1'b0;  wr_cycle[ 2312] = 1'b1;  addr_rom[ 2312]='h000006e8;  wr_data_rom[ 2312]='h00000421;
    rd_cycle[ 2313] = 1'b1;  wr_cycle[ 2313] = 1'b0;  addr_rom[ 2313]='h00000e10;  wr_data_rom[ 2313]='h00000000;
    rd_cycle[ 2314] = 1'b1;  wr_cycle[ 2314] = 1'b0;  addr_rom[ 2314]='h00000c34;  wr_data_rom[ 2314]='h00000000;
    rd_cycle[ 2315] = 1'b0;  wr_cycle[ 2315] = 1'b1;  addr_rom[ 2315]='h00000658;  wr_data_rom[ 2315]='h00000309;
    rd_cycle[ 2316] = 1'b0;  wr_cycle[ 2316] = 1'b1;  addr_rom[ 2316]='h000006f0;  wr_data_rom[ 2316]='h000006db;
    rd_cycle[ 2317] = 1'b0;  wr_cycle[ 2317] = 1'b1;  addr_rom[ 2317]='h000008f8;  wr_data_rom[ 2317]='h0000017b;
    rd_cycle[ 2318] = 1'b0;  wr_cycle[ 2318] = 1'b1;  addr_rom[ 2318]='h000004f8;  wr_data_rom[ 2318]='h00000e69;
    rd_cycle[ 2319] = 1'b1;  wr_cycle[ 2319] = 1'b0;  addr_rom[ 2319]='h000001cc;  wr_data_rom[ 2319]='h00000000;
    rd_cycle[ 2320] = 1'b0;  wr_cycle[ 2320] = 1'b1;  addr_rom[ 2320]='h00000a04;  wr_data_rom[ 2320]='h00000a9a;
    rd_cycle[ 2321] = 1'b1;  wr_cycle[ 2321] = 1'b0;  addr_rom[ 2321]='h00000f1c;  wr_data_rom[ 2321]='h00000000;
    rd_cycle[ 2322] = 1'b1;  wr_cycle[ 2322] = 1'b0;  addr_rom[ 2322]='h000008b8;  wr_data_rom[ 2322]='h00000000;
    rd_cycle[ 2323] = 1'b0;  wr_cycle[ 2323] = 1'b1;  addr_rom[ 2323]='h00000344;  wr_data_rom[ 2323]='h000002b5;
    rd_cycle[ 2324] = 1'b0;  wr_cycle[ 2324] = 1'b1;  addr_rom[ 2324]='h00000da4;  wr_data_rom[ 2324]='h00000034;
    rd_cycle[ 2325] = 1'b1;  wr_cycle[ 2325] = 1'b0;  addr_rom[ 2325]='h000001b0;  wr_data_rom[ 2325]='h00000000;
    rd_cycle[ 2326] = 1'b0;  wr_cycle[ 2326] = 1'b1;  addr_rom[ 2326]='h00000ce8;  wr_data_rom[ 2326]='h000009fb;
    rd_cycle[ 2327] = 1'b1;  wr_cycle[ 2327] = 1'b0;  addr_rom[ 2327]='h00000930;  wr_data_rom[ 2327]='h00000000;
    rd_cycle[ 2328] = 1'b0;  wr_cycle[ 2328] = 1'b1;  addr_rom[ 2328]='h000009e4;  wr_data_rom[ 2328]='h000006dd;
    rd_cycle[ 2329] = 1'b0;  wr_cycle[ 2329] = 1'b1;  addr_rom[ 2329]='h000005a8;  wr_data_rom[ 2329]='h00000af9;
    rd_cycle[ 2330] = 1'b1;  wr_cycle[ 2330] = 1'b0;  addr_rom[ 2330]='h00000f6c;  wr_data_rom[ 2330]='h00000000;
    rd_cycle[ 2331] = 1'b1;  wr_cycle[ 2331] = 1'b0;  addr_rom[ 2331]='h00000bc8;  wr_data_rom[ 2331]='h00000000;
    rd_cycle[ 2332] = 1'b1;  wr_cycle[ 2332] = 1'b0;  addr_rom[ 2332]='h0000034c;  wr_data_rom[ 2332]='h00000000;
    rd_cycle[ 2333] = 1'b1;  wr_cycle[ 2333] = 1'b0;  addr_rom[ 2333]='h000008d8;  wr_data_rom[ 2333]='h00000000;
    rd_cycle[ 2334] = 1'b0;  wr_cycle[ 2334] = 1'b1;  addr_rom[ 2334]='h000001ec;  wr_data_rom[ 2334]='h00000d64;
    rd_cycle[ 2335] = 1'b1;  wr_cycle[ 2335] = 1'b0;  addr_rom[ 2335]='h00000c68;  wr_data_rom[ 2335]='h00000000;
    rd_cycle[ 2336] = 1'b1;  wr_cycle[ 2336] = 1'b0;  addr_rom[ 2336]='h00000124;  wr_data_rom[ 2336]='h00000000;
    rd_cycle[ 2337] = 1'b0;  wr_cycle[ 2337] = 1'b1;  addr_rom[ 2337]='h00000504;  wr_data_rom[ 2337]='h0000070f;
    rd_cycle[ 2338] = 1'b1;  wr_cycle[ 2338] = 1'b0;  addr_rom[ 2338]='h00000a3c;  wr_data_rom[ 2338]='h00000000;
    rd_cycle[ 2339] = 1'b1;  wr_cycle[ 2339] = 1'b0;  addr_rom[ 2339]='h00000624;  wr_data_rom[ 2339]='h00000000;
    rd_cycle[ 2340] = 1'b0;  wr_cycle[ 2340] = 1'b1;  addr_rom[ 2340]='h00000494;  wr_data_rom[ 2340]='h00000180;
    rd_cycle[ 2341] = 1'b1;  wr_cycle[ 2341] = 1'b0;  addr_rom[ 2341]='h0000072c;  wr_data_rom[ 2341]='h00000000;
    rd_cycle[ 2342] = 1'b1;  wr_cycle[ 2342] = 1'b0;  addr_rom[ 2342]='h00000ecc;  wr_data_rom[ 2342]='h00000000;
    rd_cycle[ 2343] = 1'b1;  wr_cycle[ 2343] = 1'b0;  addr_rom[ 2343]='h00000a34;  wr_data_rom[ 2343]='h00000000;
    rd_cycle[ 2344] = 1'b1;  wr_cycle[ 2344] = 1'b0;  addr_rom[ 2344]='h00000954;  wr_data_rom[ 2344]='h00000000;
    rd_cycle[ 2345] = 1'b0;  wr_cycle[ 2345] = 1'b1;  addr_rom[ 2345]='h0000038c;  wr_data_rom[ 2345]='h00000076;
    rd_cycle[ 2346] = 1'b1;  wr_cycle[ 2346] = 1'b0;  addr_rom[ 2346]='h00000130;  wr_data_rom[ 2346]='h00000000;
    rd_cycle[ 2347] = 1'b0;  wr_cycle[ 2347] = 1'b1;  addr_rom[ 2347]='h000001a0;  wr_data_rom[ 2347]='h000003dd;
    rd_cycle[ 2348] = 1'b1;  wr_cycle[ 2348] = 1'b0;  addr_rom[ 2348]='h000001c8;  wr_data_rom[ 2348]='h00000000;
    rd_cycle[ 2349] = 1'b0;  wr_cycle[ 2349] = 1'b1;  addr_rom[ 2349]='h00000cfc;  wr_data_rom[ 2349]='h00000a24;
    rd_cycle[ 2350] = 1'b1;  wr_cycle[ 2350] = 1'b0;  addr_rom[ 2350]='h00000120;  wr_data_rom[ 2350]='h00000000;
    rd_cycle[ 2351] = 1'b1;  wr_cycle[ 2351] = 1'b0;  addr_rom[ 2351]='h000009c0;  wr_data_rom[ 2351]='h00000000;
    rd_cycle[ 2352] = 1'b1;  wr_cycle[ 2352] = 1'b0;  addr_rom[ 2352]='h00000d64;  wr_data_rom[ 2352]='h00000000;
    rd_cycle[ 2353] = 1'b1;  wr_cycle[ 2353] = 1'b0;  addr_rom[ 2353]='h000005e4;  wr_data_rom[ 2353]='h00000000;
    rd_cycle[ 2354] = 1'b1;  wr_cycle[ 2354] = 1'b0;  addr_rom[ 2354]='h000006b8;  wr_data_rom[ 2354]='h00000000;
    rd_cycle[ 2355] = 1'b0;  wr_cycle[ 2355] = 1'b1;  addr_rom[ 2355]='h000006d4;  wr_data_rom[ 2355]='h0000064d;
    rd_cycle[ 2356] = 1'b0;  wr_cycle[ 2356] = 1'b1;  addr_rom[ 2356]='h0000052c;  wr_data_rom[ 2356]='h00000579;
    rd_cycle[ 2357] = 1'b1;  wr_cycle[ 2357] = 1'b0;  addr_rom[ 2357]='h00000f58;  wr_data_rom[ 2357]='h00000000;
    rd_cycle[ 2358] = 1'b0;  wr_cycle[ 2358] = 1'b1;  addr_rom[ 2358]='h000007b4;  wr_data_rom[ 2358]='h000007c3;
    rd_cycle[ 2359] = 1'b1;  wr_cycle[ 2359] = 1'b0;  addr_rom[ 2359]='h000008d8;  wr_data_rom[ 2359]='h00000000;
    rd_cycle[ 2360] = 1'b0;  wr_cycle[ 2360] = 1'b1;  addr_rom[ 2360]='h00000224;  wr_data_rom[ 2360]='h000000d6;
    rd_cycle[ 2361] = 1'b0;  wr_cycle[ 2361] = 1'b1;  addr_rom[ 2361]='h00000a40;  wr_data_rom[ 2361]='h000008c0;
    rd_cycle[ 2362] = 1'b0;  wr_cycle[ 2362] = 1'b1;  addr_rom[ 2362]='h00000d0c;  wr_data_rom[ 2362]='h00000d51;
    rd_cycle[ 2363] = 1'b1;  wr_cycle[ 2363] = 1'b0;  addr_rom[ 2363]='h000008e0;  wr_data_rom[ 2363]='h00000000;
    rd_cycle[ 2364] = 1'b1;  wr_cycle[ 2364] = 1'b0;  addr_rom[ 2364]='h000004f0;  wr_data_rom[ 2364]='h00000000;
    rd_cycle[ 2365] = 1'b1;  wr_cycle[ 2365] = 1'b0;  addr_rom[ 2365]='h000007e4;  wr_data_rom[ 2365]='h00000000;
    rd_cycle[ 2366] = 1'b1;  wr_cycle[ 2366] = 1'b0;  addr_rom[ 2366]='h000005e0;  wr_data_rom[ 2366]='h00000000;
    rd_cycle[ 2367] = 1'b1;  wr_cycle[ 2367] = 1'b0;  addr_rom[ 2367]='h00000b34;  wr_data_rom[ 2367]='h00000000;
    rd_cycle[ 2368] = 1'b0;  wr_cycle[ 2368] = 1'b1;  addr_rom[ 2368]='h000005bc;  wr_data_rom[ 2368]='h00000700;
    rd_cycle[ 2369] = 1'b1;  wr_cycle[ 2369] = 1'b0;  addr_rom[ 2369]='h00000e94;  wr_data_rom[ 2369]='h00000000;
    rd_cycle[ 2370] = 1'b1;  wr_cycle[ 2370] = 1'b0;  addr_rom[ 2370]='h000002b0;  wr_data_rom[ 2370]='h00000000;
    rd_cycle[ 2371] = 1'b0;  wr_cycle[ 2371] = 1'b1;  addr_rom[ 2371]='h000004e8;  wr_data_rom[ 2371]='h0000000a;
    rd_cycle[ 2372] = 1'b1;  wr_cycle[ 2372] = 1'b0;  addr_rom[ 2372]='h000000e8;  wr_data_rom[ 2372]='h00000000;
    rd_cycle[ 2373] = 1'b0;  wr_cycle[ 2373] = 1'b1;  addr_rom[ 2373]='h00000998;  wr_data_rom[ 2373]='h00000670;
    rd_cycle[ 2374] = 1'b0;  wr_cycle[ 2374] = 1'b1;  addr_rom[ 2374]='h00000374;  wr_data_rom[ 2374]='h000009e6;
    rd_cycle[ 2375] = 1'b1;  wr_cycle[ 2375] = 1'b0;  addr_rom[ 2375]='h000000ec;  wr_data_rom[ 2375]='h00000000;
    rd_cycle[ 2376] = 1'b1;  wr_cycle[ 2376] = 1'b0;  addr_rom[ 2376]='h00000a70;  wr_data_rom[ 2376]='h00000000;
    rd_cycle[ 2377] = 1'b1;  wr_cycle[ 2377] = 1'b0;  addr_rom[ 2377]='h0000036c;  wr_data_rom[ 2377]='h00000000;
    rd_cycle[ 2378] = 1'b1;  wr_cycle[ 2378] = 1'b0;  addr_rom[ 2378]='h00000984;  wr_data_rom[ 2378]='h00000000;
    rd_cycle[ 2379] = 1'b0;  wr_cycle[ 2379] = 1'b1;  addr_rom[ 2379]='h00000778;  wr_data_rom[ 2379]='h000005a5;
    rd_cycle[ 2380] = 1'b1;  wr_cycle[ 2380] = 1'b0;  addr_rom[ 2380]='h00000bd4;  wr_data_rom[ 2380]='h00000000;
    rd_cycle[ 2381] = 1'b1;  wr_cycle[ 2381] = 1'b0;  addr_rom[ 2381]='h000000bc;  wr_data_rom[ 2381]='h00000000;
    rd_cycle[ 2382] = 1'b0;  wr_cycle[ 2382] = 1'b1;  addr_rom[ 2382]='h00000a34;  wr_data_rom[ 2382]='h000004ec;
    rd_cycle[ 2383] = 1'b1;  wr_cycle[ 2383] = 1'b0;  addr_rom[ 2383]='h000002e0;  wr_data_rom[ 2383]='h00000000;
    rd_cycle[ 2384] = 1'b1;  wr_cycle[ 2384] = 1'b0;  addr_rom[ 2384]='h00000898;  wr_data_rom[ 2384]='h00000000;
    rd_cycle[ 2385] = 1'b0;  wr_cycle[ 2385] = 1'b1;  addr_rom[ 2385]='h000007e4;  wr_data_rom[ 2385]='h00000852;
    rd_cycle[ 2386] = 1'b0;  wr_cycle[ 2386] = 1'b1;  addr_rom[ 2386]='h00000e98;  wr_data_rom[ 2386]='h0000058f;
    rd_cycle[ 2387] = 1'b0;  wr_cycle[ 2387] = 1'b1;  addr_rom[ 2387]='h00000388;  wr_data_rom[ 2387]='h00000124;
    rd_cycle[ 2388] = 1'b1;  wr_cycle[ 2388] = 1'b0;  addr_rom[ 2388]='h00000bd0;  wr_data_rom[ 2388]='h00000000;
    rd_cycle[ 2389] = 1'b0;  wr_cycle[ 2389] = 1'b1;  addr_rom[ 2389]='h00000374;  wr_data_rom[ 2389]='h00000cd8;
    rd_cycle[ 2390] = 1'b0;  wr_cycle[ 2390] = 1'b1;  addr_rom[ 2390]='h000002e4;  wr_data_rom[ 2390]='h00000c79;
    rd_cycle[ 2391] = 1'b0;  wr_cycle[ 2391] = 1'b1;  addr_rom[ 2391]='h00000330;  wr_data_rom[ 2391]='h00000cbc;
    rd_cycle[ 2392] = 1'b1;  wr_cycle[ 2392] = 1'b0;  addr_rom[ 2392]='h00000260;  wr_data_rom[ 2392]='h00000000;
    rd_cycle[ 2393] = 1'b1;  wr_cycle[ 2393] = 1'b0;  addr_rom[ 2393]='h000003e8;  wr_data_rom[ 2393]='h00000000;
    rd_cycle[ 2394] = 1'b0;  wr_cycle[ 2394] = 1'b1;  addr_rom[ 2394]='h00000020;  wr_data_rom[ 2394]='h00000503;
    rd_cycle[ 2395] = 1'b1;  wr_cycle[ 2395] = 1'b0;  addr_rom[ 2395]='h00000c3c;  wr_data_rom[ 2395]='h00000000;
    rd_cycle[ 2396] = 1'b1;  wr_cycle[ 2396] = 1'b0;  addr_rom[ 2396]='h00000f74;  wr_data_rom[ 2396]='h00000000;
    rd_cycle[ 2397] = 1'b1;  wr_cycle[ 2397] = 1'b0;  addr_rom[ 2397]='h00000ba0;  wr_data_rom[ 2397]='h00000000;
    rd_cycle[ 2398] = 1'b1;  wr_cycle[ 2398] = 1'b0;  addr_rom[ 2398]='h00000650;  wr_data_rom[ 2398]='h00000000;
    rd_cycle[ 2399] = 1'b1;  wr_cycle[ 2399] = 1'b0;  addr_rom[ 2399]='h00000700;  wr_data_rom[ 2399]='h00000000;
    rd_cycle[ 2400] = 1'b0;  wr_cycle[ 2400] = 1'b1;  addr_rom[ 2400]='h00000648;  wr_data_rom[ 2400]='h000005c7;
    rd_cycle[ 2401] = 1'b0;  wr_cycle[ 2401] = 1'b1;  addr_rom[ 2401]='h000003ec;  wr_data_rom[ 2401]='h0000048c;
    rd_cycle[ 2402] = 1'b1;  wr_cycle[ 2402] = 1'b0;  addr_rom[ 2402]='h00000374;  wr_data_rom[ 2402]='h00000000;
    rd_cycle[ 2403] = 1'b0;  wr_cycle[ 2403] = 1'b1;  addr_rom[ 2403]='h0000004c;  wr_data_rom[ 2403]='h000000d2;
    rd_cycle[ 2404] = 1'b1;  wr_cycle[ 2404] = 1'b0;  addr_rom[ 2404]='h00000340;  wr_data_rom[ 2404]='h00000000;
    rd_cycle[ 2405] = 1'b1;  wr_cycle[ 2405] = 1'b0;  addr_rom[ 2405]='h00000c18;  wr_data_rom[ 2405]='h00000000;
    rd_cycle[ 2406] = 1'b0;  wr_cycle[ 2406] = 1'b1;  addr_rom[ 2406]='h0000020c;  wr_data_rom[ 2406]='h000009c1;
    rd_cycle[ 2407] = 1'b0;  wr_cycle[ 2407] = 1'b1;  addr_rom[ 2407]='h00000a40;  wr_data_rom[ 2407]='h00000792;
    rd_cycle[ 2408] = 1'b1;  wr_cycle[ 2408] = 1'b0;  addr_rom[ 2408]='h00000df4;  wr_data_rom[ 2408]='h00000000;
    rd_cycle[ 2409] = 1'b1;  wr_cycle[ 2409] = 1'b0;  addr_rom[ 2409]='h00000a70;  wr_data_rom[ 2409]='h00000000;
    rd_cycle[ 2410] = 1'b0;  wr_cycle[ 2410] = 1'b1;  addr_rom[ 2410]='h000009d4;  wr_data_rom[ 2410]='h00000839;
    rd_cycle[ 2411] = 1'b1;  wr_cycle[ 2411] = 1'b0;  addr_rom[ 2411]='h000003e8;  wr_data_rom[ 2411]='h00000000;
    rd_cycle[ 2412] = 1'b1;  wr_cycle[ 2412] = 1'b0;  addr_rom[ 2412]='h00000360;  wr_data_rom[ 2412]='h00000000;
    rd_cycle[ 2413] = 1'b1;  wr_cycle[ 2413] = 1'b0;  addr_rom[ 2413]='h00000234;  wr_data_rom[ 2413]='h00000000;
    rd_cycle[ 2414] = 1'b0;  wr_cycle[ 2414] = 1'b1;  addr_rom[ 2414]='h00000094;  wr_data_rom[ 2414]='h000006e6;
    rd_cycle[ 2415] = 1'b1;  wr_cycle[ 2415] = 1'b0;  addr_rom[ 2415]='h0000008c;  wr_data_rom[ 2415]='h00000000;
    rd_cycle[ 2416] = 1'b1;  wr_cycle[ 2416] = 1'b0;  addr_rom[ 2416]='h0000085c;  wr_data_rom[ 2416]='h00000000;
    rd_cycle[ 2417] = 1'b1;  wr_cycle[ 2417] = 1'b0;  addr_rom[ 2417]='h00000544;  wr_data_rom[ 2417]='h00000000;
    rd_cycle[ 2418] = 1'b1;  wr_cycle[ 2418] = 1'b0;  addr_rom[ 2418]='h0000085c;  wr_data_rom[ 2418]='h00000000;
    rd_cycle[ 2419] = 1'b1;  wr_cycle[ 2419] = 1'b0;  addr_rom[ 2419]='h00000d34;  wr_data_rom[ 2419]='h00000000;
    rd_cycle[ 2420] = 1'b0;  wr_cycle[ 2420] = 1'b1;  addr_rom[ 2420]='h000001c8;  wr_data_rom[ 2420]='h00000bf1;
    rd_cycle[ 2421] = 1'b0;  wr_cycle[ 2421] = 1'b1;  addr_rom[ 2421]='h00000454;  wr_data_rom[ 2421]='h0000075b;
    rd_cycle[ 2422] = 1'b1;  wr_cycle[ 2422] = 1'b0;  addr_rom[ 2422]='h000003d8;  wr_data_rom[ 2422]='h00000000;
    rd_cycle[ 2423] = 1'b1;  wr_cycle[ 2423] = 1'b0;  addr_rom[ 2423]='h00000724;  wr_data_rom[ 2423]='h00000000;
    rd_cycle[ 2424] = 1'b0;  wr_cycle[ 2424] = 1'b1;  addr_rom[ 2424]='h000004f8;  wr_data_rom[ 2424]='h00000e2b;
    rd_cycle[ 2425] = 1'b0;  wr_cycle[ 2425] = 1'b1;  addr_rom[ 2425]='h00000174;  wr_data_rom[ 2425]='h00000129;
    rd_cycle[ 2426] = 1'b0;  wr_cycle[ 2426] = 1'b1;  addr_rom[ 2426]='h00000740;  wr_data_rom[ 2426]='h0000006f;
    rd_cycle[ 2427] = 1'b1;  wr_cycle[ 2427] = 1'b0;  addr_rom[ 2427]='h00000808;  wr_data_rom[ 2427]='h00000000;
    rd_cycle[ 2428] = 1'b0;  wr_cycle[ 2428] = 1'b1;  addr_rom[ 2428]='h00000610;  wr_data_rom[ 2428]='h000001c6;
    rd_cycle[ 2429] = 1'b0;  wr_cycle[ 2429] = 1'b1;  addr_rom[ 2429]='h00000d40;  wr_data_rom[ 2429]='h00000711;
    rd_cycle[ 2430] = 1'b1;  wr_cycle[ 2430] = 1'b0;  addr_rom[ 2430]='h00000a34;  wr_data_rom[ 2430]='h00000000;
    rd_cycle[ 2431] = 1'b1;  wr_cycle[ 2431] = 1'b0;  addr_rom[ 2431]='h000007d4;  wr_data_rom[ 2431]='h00000000;
    rd_cycle[ 2432] = 1'b0;  wr_cycle[ 2432] = 1'b1;  addr_rom[ 2432]='h00000e54;  wr_data_rom[ 2432]='h000003bf;
    rd_cycle[ 2433] = 1'b1;  wr_cycle[ 2433] = 1'b0;  addr_rom[ 2433]='h00000300;  wr_data_rom[ 2433]='h00000000;
    rd_cycle[ 2434] = 1'b1;  wr_cycle[ 2434] = 1'b0;  addr_rom[ 2434]='h00000eb8;  wr_data_rom[ 2434]='h00000000;
    rd_cycle[ 2435] = 1'b0;  wr_cycle[ 2435] = 1'b1;  addr_rom[ 2435]='h000002c8;  wr_data_rom[ 2435]='h00000a50;
    rd_cycle[ 2436] = 1'b1;  wr_cycle[ 2436] = 1'b0;  addr_rom[ 2436]='h00000334;  wr_data_rom[ 2436]='h00000000;
    rd_cycle[ 2437] = 1'b0;  wr_cycle[ 2437] = 1'b1;  addr_rom[ 2437]='h0000093c;  wr_data_rom[ 2437]='h000005c3;
    rd_cycle[ 2438] = 1'b0;  wr_cycle[ 2438] = 1'b1;  addr_rom[ 2438]='h000003bc;  wr_data_rom[ 2438]='h0000093c;
    rd_cycle[ 2439] = 1'b0;  wr_cycle[ 2439] = 1'b1;  addr_rom[ 2439]='h00000094;  wr_data_rom[ 2439]='h00000e17;
    rd_cycle[ 2440] = 1'b1;  wr_cycle[ 2440] = 1'b0;  addr_rom[ 2440]='h00000c18;  wr_data_rom[ 2440]='h00000000;
    rd_cycle[ 2441] = 1'b0;  wr_cycle[ 2441] = 1'b1;  addr_rom[ 2441]='h00000058;  wr_data_rom[ 2441]='h00000d40;
    rd_cycle[ 2442] = 1'b1;  wr_cycle[ 2442] = 1'b0;  addr_rom[ 2442]='h000007b4;  wr_data_rom[ 2442]='h00000000;
    rd_cycle[ 2443] = 1'b1;  wr_cycle[ 2443] = 1'b0;  addr_rom[ 2443]='h00000848;  wr_data_rom[ 2443]='h00000000;
    rd_cycle[ 2444] = 1'b1;  wr_cycle[ 2444] = 1'b0;  addr_rom[ 2444]='h00000b88;  wr_data_rom[ 2444]='h00000000;
    rd_cycle[ 2445] = 1'b0;  wr_cycle[ 2445] = 1'b1;  addr_rom[ 2445]='h00000454;  wr_data_rom[ 2445]='h00000a4d;
    rd_cycle[ 2446] = 1'b1;  wr_cycle[ 2446] = 1'b0;  addr_rom[ 2446]='h00000404;  wr_data_rom[ 2446]='h00000000;
    rd_cycle[ 2447] = 1'b1;  wr_cycle[ 2447] = 1'b0;  addr_rom[ 2447]='h00000c68;  wr_data_rom[ 2447]='h00000000;
    rd_cycle[ 2448] = 1'b1;  wr_cycle[ 2448] = 1'b0;  addr_rom[ 2448]='h000002ac;  wr_data_rom[ 2448]='h00000000;
    rd_cycle[ 2449] = 1'b0;  wr_cycle[ 2449] = 1'b1;  addr_rom[ 2449]='h00000dc4;  wr_data_rom[ 2449]='h00000d5c;
    rd_cycle[ 2450] = 1'b1;  wr_cycle[ 2450] = 1'b0;  addr_rom[ 2450]='h00000f28;  wr_data_rom[ 2450]='h00000000;
    rd_cycle[ 2451] = 1'b1;  wr_cycle[ 2451] = 1'b0;  addr_rom[ 2451]='h00000b9c;  wr_data_rom[ 2451]='h00000000;
    rd_cycle[ 2452] = 1'b0;  wr_cycle[ 2452] = 1'b1;  addr_rom[ 2452]='h00000218;  wr_data_rom[ 2452]='h00000134;
    rd_cycle[ 2453] = 1'b1;  wr_cycle[ 2453] = 1'b0;  addr_rom[ 2453]='h00000900;  wr_data_rom[ 2453]='h00000000;
    rd_cycle[ 2454] = 1'b0;  wr_cycle[ 2454] = 1'b1;  addr_rom[ 2454]='h00000e50;  wr_data_rom[ 2454]='h0000000c;
    rd_cycle[ 2455] = 1'b0;  wr_cycle[ 2455] = 1'b1;  addr_rom[ 2455]='h00000c04;  wr_data_rom[ 2455]='h00000246;
    rd_cycle[ 2456] = 1'b1;  wr_cycle[ 2456] = 1'b0;  addr_rom[ 2456]='h0000097c;  wr_data_rom[ 2456]='h00000000;
    rd_cycle[ 2457] = 1'b1;  wr_cycle[ 2457] = 1'b0;  addr_rom[ 2457]='h000006d4;  wr_data_rom[ 2457]='h00000000;
    rd_cycle[ 2458] = 1'b1;  wr_cycle[ 2458] = 1'b0;  addr_rom[ 2458]='h00000de4;  wr_data_rom[ 2458]='h00000000;
    rd_cycle[ 2459] = 1'b1;  wr_cycle[ 2459] = 1'b0;  addr_rom[ 2459]='h00000a40;  wr_data_rom[ 2459]='h00000000;
    rd_cycle[ 2460] = 1'b0;  wr_cycle[ 2460] = 1'b1;  addr_rom[ 2460]='h000002cc;  wr_data_rom[ 2460]='h00000a4b;
    rd_cycle[ 2461] = 1'b0;  wr_cycle[ 2461] = 1'b1;  addr_rom[ 2461]='h000007e0;  wr_data_rom[ 2461]='h00000768;
    rd_cycle[ 2462] = 1'b1;  wr_cycle[ 2462] = 1'b0;  addr_rom[ 2462]='h00000aa0;  wr_data_rom[ 2462]='h00000000;
    rd_cycle[ 2463] = 1'b1;  wr_cycle[ 2463] = 1'b0;  addr_rom[ 2463]='h00000954;  wr_data_rom[ 2463]='h00000000;
    rd_cycle[ 2464] = 1'b0;  wr_cycle[ 2464] = 1'b1;  addr_rom[ 2464]='h000003e8;  wr_data_rom[ 2464]='h000006e3;
    rd_cycle[ 2465] = 1'b0;  wr_cycle[ 2465] = 1'b1;  addr_rom[ 2465]='h00000a50;  wr_data_rom[ 2465]='h000002eb;
    rd_cycle[ 2466] = 1'b1;  wr_cycle[ 2466] = 1'b0;  addr_rom[ 2466]='h00000820;  wr_data_rom[ 2466]='h00000000;
    rd_cycle[ 2467] = 1'b1;  wr_cycle[ 2467] = 1'b0;  addr_rom[ 2467]='h000000c8;  wr_data_rom[ 2467]='h00000000;
    rd_cycle[ 2468] = 1'b0;  wr_cycle[ 2468] = 1'b1;  addr_rom[ 2468]='h00000500;  wr_data_rom[ 2468]='h000001b7;
    rd_cycle[ 2469] = 1'b1;  wr_cycle[ 2469] = 1'b0;  addr_rom[ 2469]='h000006f0;  wr_data_rom[ 2469]='h00000000;
    rd_cycle[ 2470] = 1'b0;  wr_cycle[ 2470] = 1'b1;  addr_rom[ 2470]='h00000c18;  wr_data_rom[ 2470]='h000000c6;
    rd_cycle[ 2471] = 1'b0;  wr_cycle[ 2471] = 1'b1;  addr_rom[ 2471]='h000002a0;  wr_data_rom[ 2471]='h00000918;
    rd_cycle[ 2472] = 1'b1;  wr_cycle[ 2472] = 1'b0;  addr_rom[ 2472]='h0000032c;  wr_data_rom[ 2472]='h00000000;
    rd_cycle[ 2473] = 1'b0;  wr_cycle[ 2473] = 1'b1;  addr_rom[ 2473]='h00000d20;  wr_data_rom[ 2473]='h00000e8a;
    rd_cycle[ 2474] = 1'b0;  wr_cycle[ 2474] = 1'b1;  addr_rom[ 2474]='h000002ec;  wr_data_rom[ 2474]='h000007cf;
    rd_cycle[ 2475] = 1'b0;  wr_cycle[ 2475] = 1'b1;  addr_rom[ 2475]='h000006c0;  wr_data_rom[ 2475]='h00000e02;
    rd_cycle[ 2476] = 1'b1;  wr_cycle[ 2476] = 1'b0;  addr_rom[ 2476]='h000004fc;  wr_data_rom[ 2476]='h00000000;
    rd_cycle[ 2477] = 1'b0;  wr_cycle[ 2477] = 1'b1;  addr_rom[ 2477]='h000002e0;  wr_data_rom[ 2477]='h0000080e;
    rd_cycle[ 2478] = 1'b1;  wr_cycle[ 2478] = 1'b0;  addr_rom[ 2478]='h000008a4;  wr_data_rom[ 2478]='h00000000;
    rd_cycle[ 2479] = 1'b1;  wr_cycle[ 2479] = 1'b0;  addr_rom[ 2479]='h000006c0;  wr_data_rom[ 2479]='h00000000;
    rd_cycle[ 2480] = 1'b0;  wr_cycle[ 2480] = 1'b1;  addr_rom[ 2480]='h000000a4;  wr_data_rom[ 2480]='h00000623;
    rd_cycle[ 2481] = 1'b1;  wr_cycle[ 2481] = 1'b0;  addr_rom[ 2481]='h000000f4;  wr_data_rom[ 2481]='h00000000;
    rd_cycle[ 2482] = 1'b1;  wr_cycle[ 2482] = 1'b0;  addr_rom[ 2482]='h0000034c;  wr_data_rom[ 2482]='h00000000;
    rd_cycle[ 2483] = 1'b0;  wr_cycle[ 2483] = 1'b1;  addr_rom[ 2483]='h000002d4;  wr_data_rom[ 2483]='h0000084d;
    rd_cycle[ 2484] = 1'b0;  wr_cycle[ 2484] = 1'b1;  addr_rom[ 2484]='h000007d0;  wr_data_rom[ 2484]='h000007f7;
    rd_cycle[ 2485] = 1'b0;  wr_cycle[ 2485] = 1'b1;  addr_rom[ 2485]='h00000894;  wr_data_rom[ 2485]='h00000bd6;
    rd_cycle[ 2486] = 1'b1;  wr_cycle[ 2486] = 1'b0;  addr_rom[ 2486]='h00000e10;  wr_data_rom[ 2486]='h00000000;
    rd_cycle[ 2487] = 1'b1;  wr_cycle[ 2487] = 1'b0;  addr_rom[ 2487]='h000006ec;  wr_data_rom[ 2487]='h00000000;
    rd_cycle[ 2488] = 1'b0;  wr_cycle[ 2488] = 1'b1;  addr_rom[ 2488]='h00000c04;  wr_data_rom[ 2488]='h000009f2;
    rd_cycle[ 2489] = 1'b1;  wr_cycle[ 2489] = 1'b0;  addr_rom[ 2489]='h00000d70;  wr_data_rom[ 2489]='h00000000;
    rd_cycle[ 2490] = 1'b1;  wr_cycle[ 2490] = 1'b0;  addr_rom[ 2490]='h000003f4;  wr_data_rom[ 2490]='h00000000;
    rd_cycle[ 2491] = 1'b1;  wr_cycle[ 2491] = 1'b0;  addr_rom[ 2491]='h0000000c;  wr_data_rom[ 2491]='h00000000;
    rd_cycle[ 2492] = 1'b0;  wr_cycle[ 2492] = 1'b1;  addr_rom[ 2492]='h000004a8;  wr_data_rom[ 2492]='h00000620;
    rd_cycle[ 2493] = 1'b1;  wr_cycle[ 2493] = 1'b0;  addr_rom[ 2493]='h000005e4;  wr_data_rom[ 2493]='h00000000;
    rd_cycle[ 2494] = 1'b1;  wr_cycle[ 2494] = 1'b0;  addr_rom[ 2494]='h00000b2c;  wr_data_rom[ 2494]='h00000000;
    rd_cycle[ 2495] = 1'b0;  wr_cycle[ 2495] = 1'b1;  addr_rom[ 2495]='h00000534;  wr_data_rom[ 2495]='h0000049e;
    rd_cycle[ 2496] = 1'b1;  wr_cycle[ 2496] = 1'b0;  addr_rom[ 2496]='h00000580;  wr_data_rom[ 2496]='h00000000;
    rd_cycle[ 2497] = 1'b0;  wr_cycle[ 2497] = 1'b1;  addr_rom[ 2497]='h0000095c;  wr_data_rom[ 2497]='h00000b2e;
    rd_cycle[ 2498] = 1'b0;  wr_cycle[ 2498] = 1'b1;  addr_rom[ 2498]='h00000d78;  wr_data_rom[ 2498]='h00000474;
    rd_cycle[ 2499] = 1'b1;  wr_cycle[ 2499] = 1'b0;  addr_rom[ 2499]='h000001bc;  wr_data_rom[ 2499]='h00000000;
    rd_cycle[ 2500] = 1'b1;  wr_cycle[ 2500] = 1'b0;  addr_rom[ 2500]='h00000664;  wr_data_rom[ 2500]='h00000000;
    rd_cycle[ 2501] = 1'b1;  wr_cycle[ 2501] = 1'b0;  addr_rom[ 2501]='h00000794;  wr_data_rom[ 2501]='h00000000;
    rd_cycle[ 2502] = 1'b0;  wr_cycle[ 2502] = 1'b1;  addr_rom[ 2502]='h00000910;  wr_data_rom[ 2502]='h00000302;
    rd_cycle[ 2503] = 1'b1;  wr_cycle[ 2503] = 1'b0;  addr_rom[ 2503]='h00000de4;  wr_data_rom[ 2503]='h00000000;
    rd_cycle[ 2504] = 1'b1;  wr_cycle[ 2504] = 1'b0;  addr_rom[ 2504]='h0000027c;  wr_data_rom[ 2504]='h00000000;
    rd_cycle[ 2505] = 1'b0;  wr_cycle[ 2505] = 1'b1;  addr_rom[ 2505]='h00000a90;  wr_data_rom[ 2505]='h00000107;
    rd_cycle[ 2506] = 1'b1;  wr_cycle[ 2506] = 1'b0;  addr_rom[ 2506]='h000001f4;  wr_data_rom[ 2506]='h00000000;
    rd_cycle[ 2507] = 1'b1;  wr_cycle[ 2507] = 1'b0;  addr_rom[ 2507]='h00000f2c;  wr_data_rom[ 2507]='h00000000;
    rd_cycle[ 2508] = 1'b0;  wr_cycle[ 2508] = 1'b1;  addr_rom[ 2508]='h00000330;  wr_data_rom[ 2508]='h0000051c;
    rd_cycle[ 2509] = 1'b1;  wr_cycle[ 2509] = 1'b0;  addr_rom[ 2509]='h000001f8;  wr_data_rom[ 2509]='h00000000;
    rd_cycle[ 2510] = 1'b0;  wr_cycle[ 2510] = 1'b1;  addr_rom[ 2510]='h00000274;  wr_data_rom[ 2510]='h00000a37;
    rd_cycle[ 2511] = 1'b0;  wr_cycle[ 2511] = 1'b1;  addr_rom[ 2511]='h0000036c;  wr_data_rom[ 2511]='h00000719;
    rd_cycle[ 2512] = 1'b0;  wr_cycle[ 2512] = 1'b1;  addr_rom[ 2512]='h000002c4;  wr_data_rom[ 2512]='h00000ce5;
    rd_cycle[ 2513] = 1'b0;  wr_cycle[ 2513] = 1'b1;  addr_rom[ 2513]='h00000174;  wr_data_rom[ 2513]='h000005ac;
    rd_cycle[ 2514] = 1'b1;  wr_cycle[ 2514] = 1'b0;  addr_rom[ 2514]='h000004f4;  wr_data_rom[ 2514]='h00000000;
    rd_cycle[ 2515] = 1'b1;  wr_cycle[ 2515] = 1'b0;  addr_rom[ 2515]='h000008c4;  wr_data_rom[ 2515]='h00000000;
    rd_cycle[ 2516] = 1'b1;  wr_cycle[ 2516] = 1'b0;  addr_rom[ 2516]='h00000764;  wr_data_rom[ 2516]='h00000000;
    rd_cycle[ 2517] = 1'b0;  wr_cycle[ 2517] = 1'b1;  addr_rom[ 2517]='h000004ec;  wr_data_rom[ 2517]='h00000b5c;
    rd_cycle[ 2518] = 1'b0;  wr_cycle[ 2518] = 1'b1;  addr_rom[ 2518]='h000001ec;  wr_data_rom[ 2518]='h00000758;
    rd_cycle[ 2519] = 1'b1;  wr_cycle[ 2519] = 1'b0;  addr_rom[ 2519]='h0000013c;  wr_data_rom[ 2519]='h00000000;
    rd_cycle[ 2520] = 1'b0;  wr_cycle[ 2520] = 1'b1;  addr_rom[ 2520]='h0000032c;  wr_data_rom[ 2520]='h00000080;
    rd_cycle[ 2521] = 1'b1;  wr_cycle[ 2521] = 1'b0;  addr_rom[ 2521]='h00000370;  wr_data_rom[ 2521]='h00000000;
    rd_cycle[ 2522] = 1'b0;  wr_cycle[ 2522] = 1'b1;  addr_rom[ 2522]='h000001b0;  wr_data_rom[ 2522]='h000008f5;
    rd_cycle[ 2523] = 1'b1;  wr_cycle[ 2523] = 1'b0;  addr_rom[ 2523]='h00000f90;  wr_data_rom[ 2523]='h00000000;
    rd_cycle[ 2524] = 1'b1;  wr_cycle[ 2524] = 1'b0;  addr_rom[ 2524]='h000006c8;  wr_data_rom[ 2524]='h00000000;
    rd_cycle[ 2525] = 1'b0;  wr_cycle[ 2525] = 1'b1;  addr_rom[ 2525]='h000009a0;  wr_data_rom[ 2525]='h000007a9;
    rd_cycle[ 2526] = 1'b1;  wr_cycle[ 2526] = 1'b0;  addr_rom[ 2526]='h0000081c;  wr_data_rom[ 2526]='h00000000;
    rd_cycle[ 2527] = 1'b1;  wr_cycle[ 2527] = 1'b0;  addr_rom[ 2527]='h00000620;  wr_data_rom[ 2527]='h00000000;
    rd_cycle[ 2528] = 1'b1;  wr_cycle[ 2528] = 1'b0;  addr_rom[ 2528]='h00000d9c;  wr_data_rom[ 2528]='h00000000;
    rd_cycle[ 2529] = 1'b1;  wr_cycle[ 2529] = 1'b0;  addr_rom[ 2529]='h00000f78;  wr_data_rom[ 2529]='h00000000;
    rd_cycle[ 2530] = 1'b1;  wr_cycle[ 2530] = 1'b0;  addr_rom[ 2530]='h00000140;  wr_data_rom[ 2530]='h00000000;
    rd_cycle[ 2531] = 1'b1;  wr_cycle[ 2531] = 1'b0;  addr_rom[ 2531]='h00000094;  wr_data_rom[ 2531]='h00000000;
    rd_cycle[ 2532] = 1'b0;  wr_cycle[ 2532] = 1'b1;  addr_rom[ 2532]='h00000bf0;  wr_data_rom[ 2532]='h0000008c;
    rd_cycle[ 2533] = 1'b0;  wr_cycle[ 2533] = 1'b1;  addr_rom[ 2533]='h00000328;  wr_data_rom[ 2533]='h00000dc4;
    rd_cycle[ 2534] = 1'b1;  wr_cycle[ 2534] = 1'b0;  addr_rom[ 2534]='h000001f4;  wr_data_rom[ 2534]='h00000000;
    rd_cycle[ 2535] = 1'b0;  wr_cycle[ 2535] = 1'b1;  addr_rom[ 2535]='h0000084c;  wr_data_rom[ 2535]='h0000025c;
    rd_cycle[ 2536] = 1'b0;  wr_cycle[ 2536] = 1'b1;  addr_rom[ 2536]='h00000808;  wr_data_rom[ 2536]='h0000072a;
    rd_cycle[ 2537] = 1'b0;  wr_cycle[ 2537] = 1'b1;  addr_rom[ 2537]='h00000214;  wr_data_rom[ 2537]='h000006f1;
    rd_cycle[ 2538] = 1'b1;  wr_cycle[ 2538] = 1'b0;  addr_rom[ 2538]='h00000eb8;  wr_data_rom[ 2538]='h00000000;
    rd_cycle[ 2539] = 1'b1;  wr_cycle[ 2539] = 1'b0;  addr_rom[ 2539]='h00000a10;  wr_data_rom[ 2539]='h00000000;
    rd_cycle[ 2540] = 1'b1;  wr_cycle[ 2540] = 1'b0;  addr_rom[ 2540]='h000009e0;  wr_data_rom[ 2540]='h00000000;
    rd_cycle[ 2541] = 1'b0;  wr_cycle[ 2541] = 1'b1;  addr_rom[ 2541]='h00000bcc;  wr_data_rom[ 2541]='h00000f85;
    rd_cycle[ 2542] = 1'b1;  wr_cycle[ 2542] = 1'b0;  addr_rom[ 2542]='h000004e4;  wr_data_rom[ 2542]='h00000000;
    rd_cycle[ 2543] = 1'b1;  wr_cycle[ 2543] = 1'b0;  addr_rom[ 2543]='h00000478;  wr_data_rom[ 2543]='h00000000;
    rd_cycle[ 2544] = 1'b0;  wr_cycle[ 2544] = 1'b1;  addr_rom[ 2544]='h00000b38;  wr_data_rom[ 2544]='h00000350;
    rd_cycle[ 2545] = 1'b0;  wr_cycle[ 2545] = 1'b1;  addr_rom[ 2545]='h00000078;  wr_data_rom[ 2545]='h000000cf;
    rd_cycle[ 2546] = 1'b1;  wr_cycle[ 2546] = 1'b0;  addr_rom[ 2546]='h00000398;  wr_data_rom[ 2546]='h00000000;
    rd_cycle[ 2547] = 1'b1;  wr_cycle[ 2547] = 1'b0;  addr_rom[ 2547]='h000007e4;  wr_data_rom[ 2547]='h00000000;
    rd_cycle[ 2548] = 1'b1;  wr_cycle[ 2548] = 1'b0;  addr_rom[ 2548]='h00000240;  wr_data_rom[ 2548]='h00000000;
    rd_cycle[ 2549] = 1'b1;  wr_cycle[ 2549] = 1'b0;  addr_rom[ 2549]='h000008e0;  wr_data_rom[ 2549]='h00000000;
    rd_cycle[ 2550] = 1'b1;  wr_cycle[ 2550] = 1'b0;  addr_rom[ 2550]='h00000930;  wr_data_rom[ 2550]='h00000000;
    rd_cycle[ 2551] = 1'b1;  wr_cycle[ 2551] = 1'b0;  addr_rom[ 2551]='h00000cf0;  wr_data_rom[ 2551]='h00000000;
    rd_cycle[ 2552] = 1'b1;  wr_cycle[ 2552] = 1'b0;  addr_rom[ 2552]='h00000a24;  wr_data_rom[ 2552]='h00000000;
    rd_cycle[ 2553] = 1'b1;  wr_cycle[ 2553] = 1'b0;  addr_rom[ 2553]='h0000019c;  wr_data_rom[ 2553]='h00000000;
    rd_cycle[ 2554] = 1'b1;  wr_cycle[ 2554] = 1'b0;  addr_rom[ 2554]='h00000b7c;  wr_data_rom[ 2554]='h00000000;
    rd_cycle[ 2555] = 1'b1;  wr_cycle[ 2555] = 1'b0;  addr_rom[ 2555]='h0000098c;  wr_data_rom[ 2555]='h00000000;
    rd_cycle[ 2556] = 1'b1;  wr_cycle[ 2556] = 1'b0;  addr_rom[ 2556]='h000005ec;  wr_data_rom[ 2556]='h00000000;
    rd_cycle[ 2557] = 1'b1;  wr_cycle[ 2557] = 1'b0;  addr_rom[ 2557]='h000004bc;  wr_data_rom[ 2557]='h00000000;
    rd_cycle[ 2558] = 1'b1;  wr_cycle[ 2558] = 1'b0;  addr_rom[ 2558]='h00000b5c;  wr_data_rom[ 2558]='h00000000;
    rd_cycle[ 2559] = 1'b1;  wr_cycle[ 2559] = 1'b0;  addr_rom[ 2559]='h000003f8;  wr_data_rom[ 2559]='h00000000;
    rd_cycle[ 2560] = 1'b0;  wr_cycle[ 2560] = 1'b1;  addr_rom[ 2560]='h00000598;  wr_data_rom[ 2560]='h00000acc;
    rd_cycle[ 2561] = 1'b1;  wr_cycle[ 2561] = 1'b0;  addr_rom[ 2561]='h000008d4;  wr_data_rom[ 2561]='h00000000;
    rd_cycle[ 2562] = 1'b0;  wr_cycle[ 2562] = 1'b1;  addr_rom[ 2562]='h00000cec;  wr_data_rom[ 2562]='h00000a7c;
    rd_cycle[ 2563] = 1'b1;  wr_cycle[ 2563] = 1'b0;  addr_rom[ 2563]='h00000a08;  wr_data_rom[ 2563]='h00000000;
    rd_cycle[ 2564] = 1'b0;  wr_cycle[ 2564] = 1'b1;  addr_rom[ 2564]='h000009a8;  wr_data_rom[ 2564]='h00000ccd;
    rd_cycle[ 2565] = 1'b1;  wr_cycle[ 2565] = 1'b0;  addr_rom[ 2565]='h0000016c;  wr_data_rom[ 2565]='h00000000;
    rd_cycle[ 2566] = 1'b1;  wr_cycle[ 2566] = 1'b0;  addr_rom[ 2566]='h0000079c;  wr_data_rom[ 2566]='h00000000;
    rd_cycle[ 2567] = 1'b0;  wr_cycle[ 2567] = 1'b1;  addr_rom[ 2567]='h00000778;  wr_data_rom[ 2567]='h000006ae;
    rd_cycle[ 2568] = 1'b1;  wr_cycle[ 2568] = 1'b0;  addr_rom[ 2568]='h00000bc0;  wr_data_rom[ 2568]='h00000000;
    rd_cycle[ 2569] = 1'b0;  wr_cycle[ 2569] = 1'b1;  addr_rom[ 2569]='h00000eb0;  wr_data_rom[ 2569]='h00000a83;
    rd_cycle[ 2570] = 1'b0;  wr_cycle[ 2570] = 1'b1;  addr_rom[ 2570]='h00000814;  wr_data_rom[ 2570]='h00000782;
    rd_cycle[ 2571] = 1'b0;  wr_cycle[ 2571] = 1'b1;  addr_rom[ 2571]='h00000298;  wr_data_rom[ 2571]='h00000983;
    rd_cycle[ 2572] = 1'b1;  wr_cycle[ 2572] = 1'b0;  addr_rom[ 2572]='h00000c78;  wr_data_rom[ 2572]='h00000000;
    rd_cycle[ 2573] = 1'b0;  wr_cycle[ 2573] = 1'b1;  addr_rom[ 2573]='h000003b0;  wr_data_rom[ 2573]='h000007f6;
    rd_cycle[ 2574] = 1'b1;  wr_cycle[ 2574] = 1'b0;  addr_rom[ 2574]='h0000088c;  wr_data_rom[ 2574]='h00000000;
    rd_cycle[ 2575] = 1'b0;  wr_cycle[ 2575] = 1'b1;  addr_rom[ 2575]='h00000cc0;  wr_data_rom[ 2575]='h00000c69;
    rd_cycle[ 2576] = 1'b0;  wr_cycle[ 2576] = 1'b1;  addr_rom[ 2576]='h00000578;  wr_data_rom[ 2576]='h00000a01;
    rd_cycle[ 2577] = 1'b1;  wr_cycle[ 2577] = 1'b0;  addr_rom[ 2577]='h00000228;  wr_data_rom[ 2577]='h00000000;
    rd_cycle[ 2578] = 1'b0;  wr_cycle[ 2578] = 1'b1;  addr_rom[ 2578]='h0000097c;  wr_data_rom[ 2578]='h00000adc;
    rd_cycle[ 2579] = 1'b1;  wr_cycle[ 2579] = 1'b0;  addr_rom[ 2579]='h00000a34;  wr_data_rom[ 2579]='h00000000;
    rd_cycle[ 2580] = 1'b1;  wr_cycle[ 2580] = 1'b0;  addr_rom[ 2580]='h00000784;  wr_data_rom[ 2580]='h00000000;
    rd_cycle[ 2581] = 1'b0;  wr_cycle[ 2581] = 1'b1;  addr_rom[ 2581]='h00000cb0;  wr_data_rom[ 2581]='h00000c7a;
    rd_cycle[ 2582] = 1'b0;  wr_cycle[ 2582] = 1'b1;  addr_rom[ 2582]='h00000bcc;  wr_data_rom[ 2582]='h0000069d;
    rd_cycle[ 2583] = 1'b0;  wr_cycle[ 2583] = 1'b1;  addr_rom[ 2583]='h00000b08;  wr_data_rom[ 2583]='h00000a70;
    rd_cycle[ 2584] = 1'b1;  wr_cycle[ 2584] = 1'b0;  addr_rom[ 2584]='h000001f0;  wr_data_rom[ 2584]='h00000000;
    rd_cycle[ 2585] = 1'b0;  wr_cycle[ 2585] = 1'b1;  addr_rom[ 2585]='h00000878;  wr_data_rom[ 2585]='h00000f97;
    rd_cycle[ 2586] = 1'b0;  wr_cycle[ 2586] = 1'b1;  addr_rom[ 2586]='h00000e34;  wr_data_rom[ 2586]='h00000d2e;
    rd_cycle[ 2587] = 1'b1;  wr_cycle[ 2587] = 1'b0;  addr_rom[ 2587]='h00000614;  wr_data_rom[ 2587]='h00000000;
    rd_cycle[ 2588] = 1'b0;  wr_cycle[ 2588] = 1'b1;  addr_rom[ 2588]='h000000fc;  wr_data_rom[ 2588]='h00000378;
    rd_cycle[ 2589] = 1'b1;  wr_cycle[ 2589] = 1'b0;  addr_rom[ 2589]='h00000514;  wr_data_rom[ 2589]='h00000000;
    rd_cycle[ 2590] = 1'b0;  wr_cycle[ 2590] = 1'b1;  addr_rom[ 2590]='h00000300;  wr_data_rom[ 2590]='h00000f0c;
    rd_cycle[ 2591] = 1'b1;  wr_cycle[ 2591] = 1'b0;  addr_rom[ 2591]='h00000cc8;  wr_data_rom[ 2591]='h00000000;
    rd_cycle[ 2592] = 1'b0;  wr_cycle[ 2592] = 1'b1;  addr_rom[ 2592]='h000005e4;  wr_data_rom[ 2592]='h000005be;
    rd_cycle[ 2593] = 1'b0;  wr_cycle[ 2593] = 1'b1;  addr_rom[ 2593]='h00000d3c;  wr_data_rom[ 2593]='h00000144;
    rd_cycle[ 2594] = 1'b0;  wr_cycle[ 2594] = 1'b1;  addr_rom[ 2594]='h00000124;  wr_data_rom[ 2594]='h00000d39;
    rd_cycle[ 2595] = 1'b0;  wr_cycle[ 2595] = 1'b1;  addr_rom[ 2595]='h00000e7c;  wr_data_rom[ 2595]='h0000093c;
    rd_cycle[ 2596] = 1'b0;  wr_cycle[ 2596] = 1'b1;  addr_rom[ 2596]='h00000a00;  wr_data_rom[ 2596]='h00000c3c;
    rd_cycle[ 2597] = 1'b1;  wr_cycle[ 2597] = 1'b0;  addr_rom[ 2597]='h00000f7c;  wr_data_rom[ 2597]='h00000000;
    rd_cycle[ 2598] = 1'b1;  wr_cycle[ 2598] = 1'b0;  addr_rom[ 2598]='h0000091c;  wr_data_rom[ 2598]='h00000000;
    rd_cycle[ 2599] = 1'b0;  wr_cycle[ 2599] = 1'b1;  addr_rom[ 2599]='h00000220;  wr_data_rom[ 2599]='h00000d3d;
    rd_cycle[ 2600] = 1'b1;  wr_cycle[ 2600] = 1'b0;  addr_rom[ 2600]='h00000c40;  wr_data_rom[ 2600]='h00000000;
    rd_cycle[ 2601] = 1'b1;  wr_cycle[ 2601] = 1'b0;  addr_rom[ 2601]='h00000c78;  wr_data_rom[ 2601]='h00000000;
    rd_cycle[ 2602] = 1'b0;  wr_cycle[ 2602] = 1'b1;  addr_rom[ 2602]='h0000018c;  wr_data_rom[ 2602]='h000006ad;
    rd_cycle[ 2603] = 1'b1;  wr_cycle[ 2603] = 1'b0;  addr_rom[ 2603]='h00000bf4;  wr_data_rom[ 2603]='h00000000;
    rd_cycle[ 2604] = 1'b1;  wr_cycle[ 2604] = 1'b0;  addr_rom[ 2604]='h00000d84;  wr_data_rom[ 2604]='h00000000;
    rd_cycle[ 2605] = 1'b1;  wr_cycle[ 2605] = 1'b0;  addr_rom[ 2605]='h000002c0;  wr_data_rom[ 2605]='h00000000;
    rd_cycle[ 2606] = 1'b1;  wr_cycle[ 2606] = 1'b0;  addr_rom[ 2606]='h00000c24;  wr_data_rom[ 2606]='h00000000;
    rd_cycle[ 2607] = 1'b0;  wr_cycle[ 2607] = 1'b1;  addr_rom[ 2607]='h00000b14;  wr_data_rom[ 2607]='h00000cab;
    rd_cycle[ 2608] = 1'b0;  wr_cycle[ 2608] = 1'b1;  addr_rom[ 2608]='h00000b00;  wr_data_rom[ 2608]='h000003cd;
    rd_cycle[ 2609] = 1'b0;  wr_cycle[ 2609] = 1'b1;  addr_rom[ 2609]='h00000f68;  wr_data_rom[ 2609]='h00000b8e;
    rd_cycle[ 2610] = 1'b0;  wr_cycle[ 2610] = 1'b1;  addr_rom[ 2610]='h000003c8;  wr_data_rom[ 2610]='h00000d2c;
    rd_cycle[ 2611] = 1'b1;  wr_cycle[ 2611] = 1'b0;  addr_rom[ 2611]='h00000a1c;  wr_data_rom[ 2611]='h00000000;
    rd_cycle[ 2612] = 1'b1;  wr_cycle[ 2612] = 1'b0;  addr_rom[ 2612]='h000005f0;  wr_data_rom[ 2612]='h00000000;
    rd_cycle[ 2613] = 1'b0;  wr_cycle[ 2613] = 1'b1;  addr_rom[ 2613]='h000003a4;  wr_data_rom[ 2613]='h00000b7d;
    rd_cycle[ 2614] = 1'b0;  wr_cycle[ 2614] = 1'b1;  addr_rom[ 2614]='h00000070;  wr_data_rom[ 2614]='h000008ce;
    rd_cycle[ 2615] = 1'b1;  wr_cycle[ 2615] = 1'b0;  addr_rom[ 2615]='h000000bc;  wr_data_rom[ 2615]='h00000000;
    rd_cycle[ 2616] = 1'b0;  wr_cycle[ 2616] = 1'b1;  addr_rom[ 2616]='h000001e8;  wr_data_rom[ 2616]='h0000035e;
    rd_cycle[ 2617] = 1'b0;  wr_cycle[ 2617] = 1'b1;  addr_rom[ 2617]='h0000021c;  wr_data_rom[ 2617]='h000005e5;
    rd_cycle[ 2618] = 1'b0;  wr_cycle[ 2618] = 1'b1;  addr_rom[ 2618]='h00000978;  wr_data_rom[ 2618]='h00000ae1;
    rd_cycle[ 2619] = 1'b0;  wr_cycle[ 2619] = 1'b1;  addr_rom[ 2619]='h00000220;  wr_data_rom[ 2619]='h00000d69;
    rd_cycle[ 2620] = 1'b1;  wr_cycle[ 2620] = 1'b0;  addr_rom[ 2620]='h0000074c;  wr_data_rom[ 2620]='h00000000;
    rd_cycle[ 2621] = 1'b0;  wr_cycle[ 2621] = 1'b1;  addr_rom[ 2621]='h00000d9c;  wr_data_rom[ 2621]='h00000338;
    rd_cycle[ 2622] = 1'b1;  wr_cycle[ 2622] = 1'b0;  addr_rom[ 2622]='h00000df8;  wr_data_rom[ 2622]='h00000000;
    rd_cycle[ 2623] = 1'b1;  wr_cycle[ 2623] = 1'b0;  addr_rom[ 2623]='h00000068;  wr_data_rom[ 2623]='h00000000;
    rd_cycle[ 2624] = 1'b0;  wr_cycle[ 2624] = 1'b1;  addr_rom[ 2624]='h000001e8;  wr_data_rom[ 2624]='h00000316;
    rd_cycle[ 2625] = 1'b1;  wr_cycle[ 2625] = 1'b0;  addr_rom[ 2625]='h000001b0;  wr_data_rom[ 2625]='h00000000;
    rd_cycle[ 2626] = 1'b1;  wr_cycle[ 2626] = 1'b0;  addr_rom[ 2626]='h00000b54;  wr_data_rom[ 2626]='h00000000;
    rd_cycle[ 2627] = 1'b1;  wr_cycle[ 2627] = 1'b0;  addr_rom[ 2627]='h0000058c;  wr_data_rom[ 2627]='h00000000;
    rd_cycle[ 2628] = 1'b1;  wr_cycle[ 2628] = 1'b0;  addr_rom[ 2628]='h00000ec8;  wr_data_rom[ 2628]='h00000000;
    rd_cycle[ 2629] = 1'b1;  wr_cycle[ 2629] = 1'b0;  addr_rom[ 2629]='h00000c20;  wr_data_rom[ 2629]='h00000000;
    rd_cycle[ 2630] = 1'b0;  wr_cycle[ 2630] = 1'b1;  addr_rom[ 2630]='h00000c0c;  wr_data_rom[ 2630]='h000008fb;
    rd_cycle[ 2631] = 1'b0;  wr_cycle[ 2631] = 1'b1;  addr_rom[ 2631]='h00000974;  wr_data_rom[ 2631]='h00000357;
    rd_cycle[ 2632] = 1'b1;  wr_cycle[ 2632] = 1'b0;  addr_rom[ 2632]='h00000c88;  wr_data_rom[ 2632]='h00000000;
    rd_cycle[ 2633] = 1'b1;  wr_cycle[ 2633] = 1'b0;  addr_rom[ 2633]='h000007d8;  wr_data_rom[ 2633]='h00000000;
    rd_cycle[ 2634] = 1'b0;  wr_cycle[ 2634] = 1'b1;  addr_rom[ 2634]='h00000b40;  wr_data_rom[ 2634]='h000008d5;
    rd_cycle[ 2635] = 1'b0;  wr_cycle[ 2635] = 1'b1;  addr_rom[ 2635]='h00000860;  wr_data_rom[ 2635]='h00000842;
    rd_cycle[ 2636] = 1'b1;  wr_cycle[ 2636] = 1'b0;  addr_rom[ 2636]='h000004d4;  wr_data_rom[ 2636]='h00000000;
    rd_cycle[ 2637] = 1'b0;  wr_cycle[ 2637] = 1'b1;  addr_rom[ 2637]='h00000114;  wr_data_rom[ 2637]='h000006d8;
    rd_cycle[ 2638] = 1'b0;  wr_cycle[ 2638] = 1'b1;  addr_rom[ 2638]='h00000b18;  wr_data_rom[ 2638]='h00000edd;
    rd_cycle[ 2639] = 1'b1;  wr_cycle[ 2639] = 1'b0;  addr_rom[ 2639]='h00000f30;  wr_data_rom[ 2639]='h00000000;
    rd_cycle[ 2640] = 1'b0;  wr_cycle[ 2640] = 1'b1;  addr_rom[ 2640]='h0000051c;  wr_data_rom[ 2640]='h00000958;
    rd_cycle[ 2641] = 1'b1;  wr_cycle[ 2641] = 1'b0;  addr_rom[ 2641]='h00000450;  wr_data_rom[ 2641]='h00000000;
    rd_cycle[ 2642] = 1'b0;  wr_cycle[ 2642] = 1'b1;  addr_rom[ 2642]='h000005c0;  wr_data_rom[ 2642]='h00000507;
    rd_cycle[ 2643] = 1'b1;  wr_cycle[ 2643] = 1'b0;  addr_rom[ 2643]='h00000560;  wr_data_rom[ 2643]='h00000000;
    rd_cycle[ 2644] = 1'b0;  wr_cycle[ 2644] = 1'b1;  addr_rom[ 2644]='h00000ecc;  wr_data_rom[ 2644]='h00000c5a;
    rd_cycle[ 2645] = 1'b0;  wr_cycle[ 2645] = 1'b1;  addr_rom[ 2645]='h00000318;  wr_data_rom[ 2645]='h000006b8;
    rd_cycle[ 2646] = 1'b0;  wr_cycle[ 2646] = 1'b1;  addr_rom[ 2646]='h00000930;  wr_data_rom[ 2646]='h0000027c;
    rd_cycle[ 2647] = 1'b0;  wr_cycle[ 2647] = 1'b1;  addr_rom[ 2647]='h00000eac;  wr_data_rom[ 2647]='h00000eac;
    rd_cycle[ 2648] = 1'b1;  wr_cycle[ 2648] = 1'b0;  addr_rom[ 2648]='h00000680;  wr_data_rom[ 2648]='h00000000;
    rd_cycle[ 2649] = 1'b1;  wr_cycle[ 2649] = 1'b0;  addr_rom[ 2649]='h00000f10;  wr_data_rom[ 2649]='h00000000;
    rd_cycle[ 2650] = 1'b0;  wr_cycle[ 2650] = 1'b1;  addr_rom[ 2650]='h000002d8;  wr_data_rom[ 2650]='h00000d95;
    rd_cycle[ 2651] = 1'b0;  wr_cycle[ 2651] = 1'b1;  addr_rom[ 2651]='h00000dd8;  wr_data_rom[ 2651]='h000002cf;
    rd_cycle[ 2652] = 1'b0;  wr_cycle[ 2652] = 1'b1;  addr_rom[ 2652]='h00000ea8;  wr_data_rom[ 2652]='h00000330;
    rd_cycle[ 2653] = 1'b1;  wr_cycle[ 2653] = 1'b0;  addr_rom[ 2653]='h0000009c;  wr_data_rom[ 2653]='h00000000;
    rd_cycle[ 2654] = 1'b1;  wr_cycle[ 2654] = 1'b0;  addr_rom[ 2654]='h00000924;  wr_data_rom[ 2654]='h00000000;
    rd_cycle[ 2655] = 1'b0;  wr_cycle[ 2655] = 1'b1;  addr_rom[ 2655]='h00000a38;  wr_data_rom[ 2655]='h00000f60;
    rd_cycle[ 2656] = 1'b1;  wr_cycle[ 2656] = 1'b0;  addr_rom[ 2656]='h00000278;  wr_data_rom[ 2656]='h00000000;
    rd_cycle[ 2657] = 1'b1;  wr_cycle[ 2657] = 1'b0;  addr_rom[ 2657]='h00000db4;  wr_data_rom[ 2657]='h00000000;
    rd_cycle[ 2658] = 1'b1;  wr_cycle[ 2658] = 1'b0;  addr_rom[ 2658]='h00000c08;  wr_data_rom[ 2658]='h00000000;
    rd_cycle[ 2659] = 1'b0;  wr_cycle[ 2659] = 1'b1;  addr_rom[ 2659]='h00000878;  wr_data_rom[ 2659]='h000000c5;
    rd_cycle[ 2660] = 1'b0;  wr_cycle[ 2660] = 1'b1;  addr_rom[ 2660]='h000000c4;  wr_data_rom[ 2660]='h00000e31;
    rd_cycle[ 2661] = 1'b0;  wr_cycle[ 2661] = 1'b1;  addr_rom[ 2661]='h000007d8;  wr_data_rom[ 2661]='h00000ab1;
    rd_cycle[ 2662] = 1'b1;  wr_cycle[ 2662] = 1'b0;  addr_rom[ 2662]='h000001e0;  wr_data_rom[ 2662]='h00000000;
    rd_cycle[ 2663] = 1'b0;  wr_cycle[ 2663] = 1'b1;  addr_rom[ 2663]='h000009a8;  wr_data_rom[ 2663]='h00000a5a;
    rd_cycle[ 2664] = 1'b1;  wr_cycle[ 2664] = 1'b0;  addr_rom[ 2664]='h00000894;  wr_data_rom[ 2664]='h00000000;
    rd_cycle[ 2665] = 1'b0;  wr_cycle[ 2665] = 1'b1;  addr_rom[ 2665]='h000005ec;  wr_data_rom[ 2665]='h00000452;
    rd_cycle[ 2666] = 1'b1;  wr_cycle[ 2666] = 1'b0;  addr_rom[ 2666]='h00000834;  wr_data_rom[ 2666]='h00000000;
    rd_cycle[ 2667] = 1'b1;  wr_cycle[ 2667] = 1'b0;  addr_rom[ 2667]='h000000d8;  wr_data_rom[ 2667]='h00000000;
    rd_cycle[ 2668] = 1'b0;  wr_cycle[ 2668] = 1'b1;  addr_rom[ 2668]='h000008a0;  wr_data_rom[ 2668]='h00000961;
    rd_cycle[ 2669] = 1'b1;  wr_cycle[ 2669] = 1'b0;  addr_rom[ 2669]='h00000438;  wr_data_rom[ 2669]='h00000000;
    rd_cycle[ 2670] = 1'b0;  wr_cycle[ 2670] = 1'b1;  addr_rom[ 2670]='h00000ec4;  wr_data_rom[ 2670]='h0000023f;
    rd_cycle[ 2671] = 1'b1;  wr_cycle[ 2671] = 1'b0;  addr_rom[ 2671]='h00000110;  wr_data_rom[ 2671]='h00000000;
    rd_cycle[ 2672] = 1'b0;  wr_cycle[ 2672] = 1'b1;  addr_rom[ 2672]='h00000e14;  wr_data_rom[ 2672]='h000006bf;
    rd_cycle[ 2673] = 1'b1;  wr_cycle[ 2673] = 1'b0;  addr_rom[ 2673]='h00000a58;  wr_data_rom[ 2673]='h00000000;
    rd_cycle[ 2674] = 1'b0;  wr_cycle[ 2674] = 1'b1;  addr_rom[ 2674]='h00000c7c;  wr_data_rom[ 2674]='h00000965;
    rd_cycle[ 2675] = 1'b0;  wr_cycle[ 2675] = 1'b1;  addr_rom[ 2675]='h00000efc;  wr_data_rom[ 2675]='h000006bc;
    rd_cycle[ 2676] = 1'b1;  wr_cycle[ 2676] = 1'b0;  addr_rom[ 2676]='h00000528;  wr_data_rom[ 2676]='h00000000;
    rd_cycle[ 2677] = 1'b0;  wr_cycle[ 2677] = 1'b1;  addr_rom[ 2677]='h00000bfc;  wr_data_rom[ 2677]='h000004f8;
    rd_cycle[ 2678] = 1'b0;  wr_cycle[ 2678] = 1'b1;  addr_rom[ 2678]='h00000c4c;  wr_data_rom[ 2678]='h00000cd7;
    rd_cycle[ 2679] = 1'b0;  wr_cycle[ 2679] = 1'b1;  addr_rom[ 2679]='h00000624;  wr_data_rom[ 2679]='h00000088;
    rd_cycle[ 2680] = 1'b1;  wr_cycle[ 2680] = 1'b0;  addr_rom[ 2680]='h00000420;  wr_data_rom[ 2680]='h00000000;
    rd_cycle[ 2681] = 1'b1;  wr_cycle[ 2681] = 1'b0;  addr_rom[ 2681]='h00000600;  wr_data_rom[ 2681]='h00000000;
    rd_cycle[ 2682] = 1'b1;  wr_cycle[ 2682] = 1'b0;  addr_rom[ 2682]='h00000ee8;  wr_data_rom[ 2682]='h00000000;
    rd_cycle[ 2683] = 1'b0;  wr_cycle[ 2683] = 1'b1;  addr_rom[ 2683]='h0000042c;  wr_data_rom[ 2683]='h00000f59;
    rd_cycle[ 2684] = 1'b0;  wr_cycle[ 2684] = 1'b1;  addr_rom[ 2684]='h00000028;  wr_data_rom[ 2684]='h0000090a;
    rd_cycle[ 2685] = 1'b1;  wr_cycle[ 2685] = 1'b0;  addr_rom[ 2685]='h00000b54;  wr_data_rom[ 2685]='h00000000;
    rd_cycle[ 2686] = 1'b1;  wr_cycle[ 2686] = 1'b0;  addr_rom[ 2686]='h00000d10;  wr_data_rom[ 2686]='h00000000;
    rd_cycle[ 2687] = 1'b0;  wr_cycle[ 2687] = 1'b1;  addr_rom[ 2687]='h000009a8;  wr_data_rom[ 2687]='h00000338;
    rd_cycle[ 2688] = 1'b0;  wr_cycle[ 2688] = 1'b1;  addr_rom[ 2688]='h00000d0c;  wr_data_rom[ 2688]='h000007bd;
    rd_cycle[ 2689] = 1'b1;  wr_cycle[ 2689] = 1'b0;  addr_rom[ 2689]='h000001a8;  wr_data_rom[ 2689]='h00000000;
    rd_cycle[ 2690] = 1'b0;  wr_cycle[ 2690] = 1'b1;  addr_rom[ 2690]='h0000082c;  wr_data_rom[ 2690]='h000000af;
    rd_cycle[ 2691] = 1'b1;  wr_cycle[ 2691] = 1'b0;  addr_rom[ 2691]='h00000f40;  wr_data_rom[ 2691]='h00000000;
    rd_cycle[ 2692] = 1'b1;  wr_cycle[ 2692] = 1'b0;  addr_rom[ 2692]='h00000544;  wr_data_rom[ 2692]='h00000000;
    rd_cycle[ 2693] = 1'b0;  wr_cycle[ 2693] = 1'b1;  addr_rom[ 2693]='h00000488;  wr_data_rom[ 2693]='h0000077a;
    rd_cycle[ 2694] = 1'b0;  wr_cycle[ 2694] = 1'b1;  addr_rom[ 2694]='h0000049c;  wr_data_rom[ 2694]='h00000b27;
    rd_cycle[ 2695] = 1'b0;  wr_cycle[ 2695] = 1'b1;  addr_rom[ 2695]='h00000b8c;  wr_data_rom[ 2695]='h000003a1;
    rd_cycle[ 2696] = 1'b0;  wr_cycle[ 2696] = 1'b1;  addr_rom[ 2696]='h000005bc;  wr_data_rom[ 2696]='h00000e65;
    rd_cycle[ 2697] = 1'b0;  wr_cycle[ 2697] = 1'b1;  addr_rom[ 2697]='h00000abc;  wr_data_rom[ 2697]='h000006c5;
    rd_cycle[ 2698] = 1'b0;  wr_cycle[ 2698] = 1'b1;  addr_rom[ 2698]='h00000348;  wr_data_rom[ 2698]='h000008dd;
    rd_cycle[ 2699] = 1'b1;  wr_cycle[ 2699] = 1'b0;  addr_rom[ 2699]='h000005ac;  wr_data_rom[ 2699]='h00000000;
    rd_cycle[ 2700] = 1'b1;  wr_cycle[ 2700] = 1'b0;  addr_rom[ 2700]='h000009cc;  wr_data_rom[ 2700]='h00000000;
    rd_cycle[ 2701] = 1'b1;  wr_cycle[ 2701] = 1'b0;  addr_rom[ 2701]='h00000cc8;  wr_data_rom[ 2701]='h00000000;
    rd_cycle[ 2702] = 1'b1;  wr_cycle[ 2702] = 1'b0;  addr_rom[ 2702]='h00000dec;  wr_data_rom[ 2702]='h00000000;
    rd_cycle[ 2703] = 1'b0;  wr_cycle[ 2703] = 1'b1;  addr_rom[ 2703]='h00000e4c;  wr_data_rom[ 2703]='h00000414;
    rd_cycle[ 2704] = 1'b0;  wr_cycle[ 2704] = 1'b1;  addr_rom[ 2704]='h00000218;  wr_data_rom[ 2704]='h00000476;
    rd_cycle[ 2705] = 1'b0;  wr_cycle[ 2705] = 1'b1;  addr_rom[ 2705]='h00000a78;  wr_data_rom[ 2705]='h00000e1c;
    rd_cycle[ 2706] = 1'b1;  wr_cycle[ 2706] = 1'b0;  addr_rom[ 2706]='h000000cc;  wr_data_rom[ 2706]='h00000000;
    rd_cycle[ 2707] = 1'b0;  wr_cycle[ 2707] = 1'b1;  addr_rom[ 2707]='h000005ec;  wr_data_rom[ 2707]='h00000378;
    rd_cycle[ 2708] = 1'b1;  wr_cycle[ 2708] = 1'b0;  addr_rom[ 2708]='h00000a34;  wr_data_rom[ 2708]='h00000000;
    rd_cycle[ 2709] = 1'b1;  wr_cycle[ 2709] = 1'b0;  addr_rom[ 2709]='h00000ee4;  wr_data_rom[ 2709]='h00000000;
    rd_cycle[ 2710] = 1'b0;  wr_cycle[ 2710] = 1'b1;  addr_rom[ 2710]='h0000041c;  wr_data_rom[ 2710]='h00000d52;
    rd_cycle[ 2711] = 1'b0;  wr_cycle[ 2711] = 1'b1;  addr_rom[ 2711]='h000007e8;  wr_data_rom[ 2711]='h00000079;
    rd_cycle[ 2712] = 1'b0;  wr_cycle[ 2712] = 1'b1;  addr_rom[ 2712]='h00000494;  wr_data_rom[ 2712]='h00000c15;
    rd_cycle[ 2713] = 1'b1;  wr_cycle[ 2713] = 1'b0;  addr_rom[ 2713]='h00000550;  wr_data_rom[ 2713]='h00000000;
    rd_cycle[ 2714] = 1'b1;  wr_cycle[ 2714] = 1'b0;  addr_rom[ 2714]='h000004e4;  wr_data_rom[ 2714]='h00000000;
    rd_cycle[ 2715] = 1'b0;  wr_cycle[ 2715] = 1'b1;  addr_rom[ 2715]='h00000088;  wr_data_rom[ 2715]='h000006e4;
    rd_cycle[ 2716] = 1'b1;  wr_cycle[ 2716] = 1'b0;  addr_rom[ 2716]='h00000bec;  wr_data_rom[ 2716]='h00000000;
    rd_cycle[ 2717] = 1'b0;  wr_cycle[ 2717] = 1'b1;  addr_rom[ 2717]='h0000060c;  wr_data_rom[ 2717]='h000000b0;
    rd_cycle[ 2718] = 1'b1;  wr_cycle[ 2718] = 1'b0;  addr_rom[ 2718]='h00000918;  wr_data_rom[ 2718]='h00000000;
    rd_cycle[ 2719] = 1'b0;  wr_cycle[ 2719] = 1'b1;  addr_rom[ 2719]='h0000084c;  wr_data_rom[ 2719]='h00000d4f;
    rd_cycle[ 2720] = 1'b1;  wr_cycle[ 2720] = 1'b0;  addr_rom[ 2720]='h00000270;  wr_data_rom[ 2720]='h00000000;
    rd_cycle[ 2721] = 1'b0;  wr_cycle[ 2721] = 1'b1;  addr_rom[ 2721]='h000004fc;  wr_data_rom[ 2721]='h00000f40;
    rd_cycle[ 2722] = 1'b0;  wr_cycle[ 2722] = 1'b1;  addr_rom[ 2722]='h0000044c;  wr_data_rom[ 2722]='h00000017;
    rd_cycle[ 2723] = 1'b0;  wr_cycle[ 2723] = 1'b1;  addr_rom[ 2723]='h00000c48;  wr_data_rom[ 2723]='h00000747;
    rd_cycle[ 2724] = 1'b0;  wr_cycle[ 2724] = 1'b1;  addr_rom[ 2724]='h000003dc;  wr_data_rom[ 2724]='h00000711;
    rd_cycle[ 2725] = 1'b0;  wr_cycle[ 2725] = 1'b1;  addr_rom[ 2725]='h00000f98;  wr_data_rom[ 2725]='h0000076b;
    rd_cycle[ 2726] = 1'b0;  wr_cycle[ 2726] = 1'b1;  addr_rom[ 2726]='h00000a78;  wr_data_rom[ 2726]='h0000096b;
    rd_cycle[ 2727] = 1'b1;  wr_cycle[ 2727] = 1'b0;  addr_rom[ 2727]='h00000bac;  wr_data_rom[ 2727]='h00000000;
    rd_cycle[ 2728] = 1'b0;  wr_cycle[ 2728] = 1'b1;  addr_rom[ 2728]='h00000e7c;  wr_data_rom[ 2728]='h00000069;
    rd_cycle[ 2729] = 1'b0;  wr_cycle[ 2729] = 1'b1;  addr_rom[ 2729]='h00000048;  wr_data_rom[ 2729]='h0000041c;
    rd_cycle[ 2730] = 1'b1;  wr_cycle[ 2730] = 1'b0;  addr_rom[ 2730]='h00000788;  wr_data_rom[ 2730]='h00000000;
    rd_cycle[ 2731] = 1'b1;  wr_cycle[ 2731] = 1'b0;  addr_rom[ 2731]='h00000150;  wr_data_rom[ 2731]='h00000000;
    rd_cycle[ 2732] = 1'b1;  wr_cycle[ 2732] = 1'b0;  addr_rom[ 2732]='h00000a90;  wr_data_rom[ 2732]='h00000000;
    rd_cycle[ 2733] = 1'b1;  wr_cycle[ 2733] = 1'b0;  addr_rom[ 2733]='h0000078c;  wr_data_rom[ 2733]='h00000000;
    rd_cycle[ 2734] = 1'b1;  wr_cycle[ 2734] = 1'b0;  addr_rom[ 2734]='h00000664;  wr_data_rom[ 2734]='h00000000;
    rd_cycle[ 2735] = 1'b1;  wr_cycle[ 2735] = 1'b0;  addr_rom[ 2735]='h00000648;  wr_data_rom[ 2735]='h00000000;
    rd_cycle[ 2736] = 1'b1;  wr_cycle[ 2736] = 1'b0;  addr_rom[ 2736]='h0000000c;  wr_data_rom[ 2736]='h00000000;
    rd_cycle[ 2737] = 1'b1;  wr_cycle[ 2737] = 1'b0;  addr_rom[ 2737]='h000001ec;  wr_data_rom[ 2737]='h00000000;
    rd_cycle[ 2738] = 1'b1;  wr_cycle[ 2738] = 1'b0;  addr_rom[ 2738]='h00000130;  wr_data_rom[ 2738]='h00000000;
    rd_cycle[ 2739] = 1'b1;  wr_cycle[ 2739] = 1'b0;  addr_rom[ 2739]='h00000b58;  wr_data_rom[ 2739]='h00000000;
    rd_cycle[ 2740] = 1'b1;  wr_cycle[ 2740] = 1'b0;  addr_rom[ 2740]='h00000d10;  wr_data_rom[ 2740]='h00000000;
    rd_cycle[ 2741] = 1'b1;  wr_cycle[ 2741] = 1'b0;  addr_rom[ 2741]='h000005dc;  wr_data_rom[ 2741]='h00000000;
    rd_cycle[ 2742] = 1'b1;  wr_cycle[ 2742] = 1'b0;  addr_rom[ 2742]='h00000bb8;  wr_data_rom[ 2742]='h00000000;
    rd_cycle[ 2743] = 1'b0;  wr_cycle[ 2743] = 1'b1;  addr_rom[ 2743]='h00000b48;  wr_data_rom[ 2743]='h000003fc;
    rd_cycle[ 2744] = 1'b1;  wr_cycle[ 2744] = 1'b0;  addr_rom[ 2744]='h000002dc;  wr_data_rom[ 2744]='h00000000;
    rd_cycle[ 2745] = 1'b1;  wr_cycle[ 2745] = 1'b0;  addr_rom[ 2745]='h00000d4c;  wr_data_rom[ 2745]='h00000000;
    rd_cycle[ 2746] = 1'b0;  wr_cycle[ 2746] = 1'b1;  addr_rom[ 2746]='h00000d74;  wr_data_rom[ 2746]='h00000a12;
    rd_cycle[ 2747] = 1'b0;  wr_cycle[ 2747] = 1'b1;  addr_rom[ 2747]='h00000304;  wr_data_rom[ 2747]='h00000f8d;
    rd_cycle[ 2748] = 1'b1;  wr_cycle[ 2748] = 1'b0;  addr_rom[ 2748]='h00000b08;  wr_data_rom[ 2748]='h00000000;
    rd_cycle[ 2749] = 1'b1;  wr_cycle[ 2749] = 1'b0;  addr_rom[ 2749]='h00000454;  wr_data_rom[ 2749]='h00000000;
    rd_cycle[ 2750] = 1'b0;  wr_cycle[ 2750] = 1'b1;  addr_rom[ 2750]='h00000b74;  wr_data_rom[ 2750]='h00000eb3;
    rd_cycle[ 2751] = 1'b1;  wr_cycle[ 2751] = 1'b0;  addr_rom[ 2751]='h00000454;  wr_data_rom[ 2751]='h00000000;
    rd_cycle[ 2752] = 1'b0;  wr_cycle[ 2752] = 1'b1;  addr_rom[ 2752]='h00000328;  wr_data_rom[ 2752]='h00000338;
    rd_cycle[ 2753] = 1'b1;  wr_cycle[ 2753] = 1'b0;  addr_rom[ 2753]='h00000e90;  wr_data_rom[ 2753]='h00000000;
    rd_cycle[ 2754] = 1'b0;  wr_cycle[ 2754] = 1'b1;  addr_rom[ 2754]='h00000884;  wr_data_rom[ 2754]='h00000678;
    rd_cycle[ 2755] = 1'b1;  wr_cycle[ 2755] = 1'b0;  addr_rom[ 2755]='h0000032c;  wr_data_rom[ 2755]='h00000000;
    rd_cycle[ 2756] = 1'b0;  wr_cycle[ 2756] = 1'b1;  addr_rom[ 2756]='h000008a4;  wr_data_rom[ 2756]='h000002cd;
    rd_cycle[ 2757] = 1'b1;  wr_cycle[ 2757] = 1'b0;  addr_rom[ 2757]='h000004e8;  wr_data_rom[ 2757]='h00000000;
    rd_cycle[ 2758] = 1'b0;  wr_cycle[ 2758] = 1'b1;  addr_rom[ 2758]='h00000590;  wr_data_rom[ 2758]='h0000090b;
    rd_cycle[ 2759] = 1'b0;  wr_cycle[ 2759] = 1'b1;  addr_rom[ 2759]='h00000160;  wr_data_rom[ 2759]='h00000a79;
    rd_cycle[ 2760] = 1'b1;  wr_cycle[ 2760] = 1'b0;  addr_rom[ 2760]='h00000b58;  wr_data_rom[ 2760]='h00000000;
    rd_cycle[ 2761] = 1'b0;  wr_cycle[ 2761] = 1'b1;  addr_rom[ 2761]='h00000f9c;  wr_data_rom[ 2761]='h00000e29;
    rd_cycle[ 2762] = 1'b1;  wr_cycle[ 2762] = 1'b0;  addr_rom[ 2762]='h00000dc0;  wr_data_rom[ 2762]='h00000000;
    rd_cycle[ 2763] = 1'b0;  wr_cycle[ 2763] = 1'b1;  addr_rom[ 2763]='h000006f4;  wr_data_rom[ 2763]='h0000020a;
    rd_cycle[ 2764] = 1'b0;  wr_cycle[ 2764] = 1'b1;  addr_rom[ 2764]='h0000047c;  wr_data_rom[ 2764]='h00000000;
    rd_cycle[ 2765] = 1'b0;  wr_cycle[ 2765] = 1'b1;  addr_rom[ 2765]='h00000d74;  wr_data_rom[ 2765]='h00000c5e;
    rd_cycle[ 2766] = 1'b0;  wr_cycle[ 2766] = 1'b1;  addr_rom[ 2766]='h00000760;  wr_data_rom[ 2766]='h00000d17;
    rd_cycle[ 2767] = 1'b0;  wr_cycle[ 2767] = 1'b1;  addr_rom[ 2767]='h00000718;  wr_data_rom[ 2767]='h00000080;
    rd_cycle[ 2768] = 1'b1;  wr_cycle[ 2768] = 1'b0;  addr_rom[ 2768]='h00000ec8;  wr_data_rom[ 2768]='h00000000;
    rd_cycle[ 2769] = 1'b1;  wr_cycle[ 2769] = 1'b0;  addr_rom[ 2769]='h00000900;  wr_data_rom[ 2769]='h00000000;
    rd_cycle[ 2770] = 1'b1;  wr_cycle[ 2770] = 1'b0;  addr_rom[ 2770]='h000005d4;  wr_data_rom[ 2770]='h00000000;
    rd_cycle[ 2771] = 1'b0;  wr_cycle[ 2771] = 1'b1;  addr_rom[ 2771]='h00000d0c;  wr_data_rom[ 2771]='h0000076b;
    rd_cycle[ 2772] = 1'b0;  wr_cycle[ 2772] = 1'b1;  addr_rom[ 2772]='h00000438;  wr_data_rom[ 2772]='h00000ab0;
    rd_cycle[ 2773] = 1'b1;  wr_cycle[ 2773] = 1'b0;  addr_rom[ 2773]='h00000ab4;  wr_data_rom[ 2773]='h00000000;
    rd_cycle[ 2774] = 1'b1;  wr_cycle[ 2774] = 1'b0;  addr_rom[ 2774]='h00000abc;  wr_data_rom[ 2774]='h00000000;
    rd_cycle[ 2775] = 1'b1;  wr_cycle[ 2775] = 1'b0;  addr_rom[ 2775]='h00000520;  wr_data_rom[ 2775]='h00000000;
    rd_cycle[ 2776] = 1'b0;  wr_cycle[ 2776] = 1'b1;  addr_rom[ 2776]='h000005e8;  wr_data_rom[ 2776]='h00000f82;
    rd_cycle[ 2777] = 1'b1;  wr_cycle[ 2777] = 1'b0;  addr_rom[ 2777]='h00000f98;  wr_data_rom[ 2777]='h00000000;
    rd_cycle[ 2778] = 1'b1;  wr_cycle[ 2778] = 1'b0;  addr_rom[ 2778]='h00000b94;  wr_data_rom[ 2778]='h00000000;
    rd_cycle[ 2779] = 1'b0;  wr_cycle[ 2779] = 1'b1;  addr_rom[ 2779]='h00000d70;  wr_data_rom[ 2779]='h0000097a;
    rd_cycle[ 2780] = 1'b0;  wr_cycle[ 2780] = 1'b1;  addr_rom[ 2780]='h0000009c;  wr_data_rom[ 2780]='h00000867;
    rd_cycle[ 2781] = 1'b1;  wr_cycle[ 2781] = 1'b0;  addr_rom[ 2781]='h00000d00;  wr_data_rom[ 2781]='h00000000;
    rd_cycle[ 2782] = 1'b0;  wr_cycle[ 2782] = 1'b1;  addr_rom[ 2782]='h00000148;  wr_data_rom[ 2782]='h000002c4;
    rd_cycle[ 2783] = 1'b1;  wr_cycle[ 2783] = 1'b0;  addr_rom[ 2783]='h00000d00;  wr_data_rom[ 2783]='h00000000;
    rd_cycle[ 2784] = 1'b0;  wr_cycle[ 2784] = 1'b1;  addr_rom[ 2784]='h00000348;  wr_data_rom[ 2784]='h0000074f;
    rd_cycle[ 2785] = 1'b1;  wr_cycle[ 2785] = 1'b0;  addr_rom[ 2785]='h000009d0;  wr_data_rom[ 2785]='h00000000;
    rd_cycle[ 2786] = 1'b1;  wr_cycle[ 2786] = 1'b0;  addr_rom[ 2786]='h00000e60;  wr_data_rom[ 2786]='h00000000;
    rd_cycle[ 2787] = 1'b1;  wr_cycle[ 2787] = 1'b0;  addr_rom[ 2787]='h00000024;  wr_data_rom[ 2787]='h00000000;
    rd_cycle[ 2788] = 1'b0;  wr_cycle[ 2788] = 1'b1;  addr_rom[ 2788]='h000000a8;  wr_data_rom[ 2788]='h00000257;
    rd_cycle[ 2789] = 1'b0;  wr_cycle[ 2789] = 1'b1;  addr_rom[ 2789]='h00000684;  wr_data_rom[ 2789]='h00000b94;
    rd_cycle[ 2790] = 1'b0;  wr_cycle[ 2790] = 1'b1;  addr_rom[ 2790]='h00000040;  wr_data_rom[ 2790]='h0000031f;
    rd_cycle[ 2791] = 1'b1;  wr_cycle[ 2791] = 1'b0;  addr_rom[ 2791]='h00000914;  wr_data_rom[ 2791]='h00000000;
    rd_cycle[ 2792] = 1'b0;  wr_cycle[ 2792] = 1'b1;  addr_rom[ 2792]='h00000448;  wr_data_rom[ 2792]='h0000055f;
    rd_cycle[ 2793] = 1'b0;  wr_cycle[ 2793] = 1'b1;  addr_rom[ 2793]='h00000970;  wr_data_rom[ 2793]='h00000e46;
    rd_cycle[ 2794] = 1'b1;  wr_cycle[ 2794] = 1'b0;  addr_rom[ 2794]='h00000ef8;  wr_data_rom[ 2794]='h00000000;
    rd_cycle[ 2795] = 1'b0;  wr_cycle[ 2795] = 1'b1;  addr_rom[ 2795]='h0000064c;  wr_data_rom[ 2795]='h0000042c;
    rd_cycle[ 2796] = 1'b1;  wr_cycle[ 2796] = 1'b0;  addr_rom[ 2796]='h000006a4;  wr_data_rom[ 2796]='h00000000;
    rd_cycle[ 2797] = 1'b1;  wr_cycle[ 2797] = 1'b0;  addr_rom[ 2797]='h000007b8;  wr_data_rom[ 2797]='h00000000;
    rd_cycle[ 2798] = 1'b1;  wr_cycle[ 2798] = 1'b0;  addr_rom[ 2798]='h0000088c;  wr_data_rom[ 2798]='h00000000;
    rd_cycle[ 2799] = 1'b1;  wr_cycle[ 2799] = 1'b0;  addr_rom[ 2799]='h000008e0;  wr_data_rom[ 2799]='h00000000;
    rd_cycle[ 2800] = 1'b0;  wr_cycle[ 2800] = 1'b1;  addr_rom[ 2800]='h000000a4;  wr_data_rom[ 2800]='h00000108;
    rd_cycle[ 2801] = 1'b1;  wr_cycle[ 2801] = 1'b0;  addr_rom[ 2801]='h0000083c;  wr_data_rom[ 2801]='h00000000;
    rd_cycle[ 2802] = 1'b1;  wr_cycle[ 2802] = 1'b0;  addr_rom[ 2802]='h00000374;  wr_data_rom[ 2802]='h00000000;
    rd_cycle[ 2803] = 1'b0;  wr_cycle[ 2803] = 1'b1;  addr_rom[ 2803]='h00000454;  wr_data_rom[ 2803]='h0000018f;
    rd_cycle[ 2804] = 1'b1;  wr_cycle[ 2804] = 1'b0;  addr_rom[ 2804]='h000006bc;  wr_data_rom[ 2804]='h00000000;
    rd_cycle[ 2805] = 1'b1;  wr_cycle[ 2805] = 1'b0;  addr_rom[ 2805]='h00000958;  wr_data_rom[ 2805]='h00000000;
    rd_cycle[ 2806] = 1'b1;  wr_cycle[ 2806] = 1'b0;  addr_rom[ 2806]='h000007b8;  wr_data_rom[ 2806]='h00000000;
    rd_cycle[ 2807] = 1'b0;  wr_cycle[ 2807] = 1'b1;  addr_rom[ 2807]='h000007d4;  wr_data_rom[ 2807]='h00000683;
    rd_cycle[ 2808] = 1'b0;  wr_cycle[ 2808] = 1'b1;  addr_rom[ 2808]='h00000770;  wr_data_rom[ 2808]='h00000be4;
    rd_cycle[ 2809] = 1'b1;  wr_cycle[ 2809] = 1'b0;  addr_rom[ 2809]='h000000b0;  wr_data_rom[ 2809]='h00000000;
    rd_cycle[ 2810] = 1'b1;  wr_cycle[ 2810] = 1'b0;  addr_rom[ 2810]='h00000458;  wr_data_rom[ 2810]='h00000000;
    rd_cycle[ 2811] = 1'b0;  wr_cycle[ 2811] = 1'b1;  addr_rom[ 2811]='h0000045c;  wr_data_rom[ 2811]='h000006c8;
    rd_cycle[ 2812] = 1'b0;  wr_cycle[ 2812] = 1'b1;  addr_rom[ 2812]='h00000500;  wr_data_rom[ 2812]='h00000123;
    rd_cycle[ 2813] = 1'b0;  wr_cycle[ 2813] = 1'b1;  addr_rom[ 2813]='h00000828;  wr_data_rom[ 2813]='h00000778;
    rd_cycle[ 2814] = 1'b0;  wr_cycle[ 2814] = 1'b1;  addr_rom[ 2814]='h00000c98;  wr_data_rom[ 2814]='h00000856;
    rd_cycle[ 2815] = 1'b0;  wr_cycle[ 2815] = 1'b1;  addr_rom[ 2815]='h00000054;  wr_data_rom[ 2815]='h00000946;
    rd_cycle[ 2816] = 1'b1;  wr_cycle[ 2816] = 1'b0;  addr_rom[ 2816]='h00000244;  wr_data_rom[ 2816]='h00000000;
    rd_cycle[ 2817] = 1'b0;  wr_cycle[ 2817] = 1'b1;  addr_rom[ 2817]='h00000960;  wr_data_rom[ 2817]='h00000a86;
    rd_cycle[ 2818] = 1'b0;  wr_cycle[ 2818] = 1'b1;  addr_rom[ 2818]='h00000580;  wr_data_rom[ 2818]='h00000554;
    rd_cycle[ 2819] = 1'b1;  wr_cycle[ 2819] = 1'b0;  addr_rom[ 2819]='h00000d68;  wr_data_rom[ 2819]='h00000000;
    rd_cycle[ 2820] = 1'b0;  wr_cycle[ 2820] = 1'b1;  addr_rom[ 2820]='h0000026c;  wr_data_rom[ 2820]='h00000b54;
    rd_cycle[ 2821] = 1'b1;  wr_cycle[ 2821] = 1'b0;  addr_rom[ 2821]='h00000a64;  wr_data_rom[ 2821]='h00000000;
    rd_cycle[ 2822] = 1'b0;  wr_cycle[ 2822] = 1'b1;  addr_rom[ 2822]='h00000420;  wr_data_rom[ 2822]='h00000cab;
    rd_cycle[ 2823] = 1'b0;  wr_cycle[ 2823] = 1'b1;  addr_rom[ 2823]='h00000d54;  wr_data_rom[ 2823]='h00000d8a;
    rd_cycle[ 2824] = 1'b1;  wr_cycle[ 2824] = 1'b0;  addr_rom[ 2824]='h00000d58;  wr_data_rom[ 2824]='h00000000;
    rd_cycle[ 2825] = 1'b0;  wr_cycle[ 2825] = 1'b1;  addr_rom[ 2825]='h00000e9c;  wr_data_rom[ 2825]='h00000b58;
    rd_cycle[ 2826] = 1'b0;  wr_cycle[ 2826] = 1'b1;  addr_rom[ 2826]='h000009bc;  wr_data_rom[ 2826]='h000005f4;
    rd_cycle[ 2827] = 1'b0;  wr_cycle[ 2827] = 1'b1;  addr_rom[ 2827]='h0000005c;  wr_data_rom[ 2827]='h000009f8;
    rd_cycle[ 2828] = 1'b0;  wr_cycle[ 2828] = 1'b1;  addr_rom[ 2828]='h00000c14;  wr_data_rom[ 2828]='h00000049;
    rd_cycle[ 2829] = 1'b1;  wr_cycle[ 2829] = 1'b0;  addr_rom[ 2829]='h0000060c;  wr_data_rom[ 2829]='h00000000;
    rd_cycle[ 2830] = 1'b1;  wr_cycle[ 2830] = 1'b0;  addr_rom[ 2830]='h00000864;  wr_data_rom[ 2830]='h00000000;
    rd_cycle[ 2831] = 1'b0;  wr_cycle[ 2831] = 1'b1;  addr_rom[ 2831]='h000004d0;  wr_data_rom[ 2831]='h000006bf;
    rd_cycle[ 2832] = 1'b1;  wr_cycle[ 2832] = 1'b0;  addr_rom[ 2832]='h00000648;  wr_data_rom[ 2832]='h00000000;
    rd_cycle[ 2833] = 1'b1;  wr_cycle[ 2833] = 1'b0;  addr_rom[ 2833]='h00000c58;  wr_data_rom[ 2833]='h00000000;
    rd_cycle[ 2834] = 1'b0;  wr_cycle[ 2834] = 1'b1;  addr_rom[ 2834]='h00000f84;  wr_data_rom[ 2834]='h0000049c;
    rd_cycle[ 2835] = 1'b1;  wr_cycle[ 2835] = 1'b0;  addr_rom[ 2835]='h00000c38;  wr_data_rom[ 2835]='h00000000;
    rd_cycle[ 2836] = 1'b1;  wr_cycle[ 2836] = 1'b0;  addr_rom[ 2836]='h00000d18;  wr_data_rom[ 2836]='h00000000;
    rd_cycle[ 2837] = 1'b1;  wr_cycle[ 2837] = 1'b0;  addr_rom[ 2837]='h0000050c;  wr_data_rom[ 2837]='h00000000;
    rd_cycle[ 2838] = 1'b0;  wr_cycle[ 2838] = 1'b1;  addr_rom[ 2838]='h00000b44;  wr_data_rom[ 2838]='h00000230;
    rd_cycle[ 2839] = 1'b1;  wr_cycle[ 2839] = 1'b0;  addr_rom[ 2839]='h00000ef4;  wr_data_rom[ 2839]='h00000000;
    rd_cycle[ 2840] = 1'b1;  wr_cycle[ 2840] = 1'b0;  addr_rom[ 2840]='h00000544;  wr_data_rom[ 2840]='h00000000;
    rd_cycle[ 2841] = 1'b0;  wr_cycle[ 2841] = 1'b1;  addr_rom[ 2841]='h000005a4;  wr_data_rom[ 2841]='h00000169;
    rd_cycle[ 2842] = 1'b1;  wr_cycle[ 2842] = 1'b0;  addr_rom[ 2842]='h00000018;  wr_data_rom[ 2842]='h00000000;
    rd_cycle[ 2843] = 1'b1;  wr_cycle[ 2843] = 1'b0;  addr_rom[ 2843]='h00000f14;  wr_data_rom[ 2843]='h00000000;
    rd_cycle[ 2844] = 1'b0;  wr_cycle[ 2844] = 1'b1;  addr_rom[ 2844]='h00000ba8;  wr_data_rom[ 2844]='h000006a0;
    rd_cycle[ 2845] = 1'b0;  wr_cycle[ 2845] = 1'b1;  addr_rom[ 2845]='h000000b8;  wr_data_rom[ 2845]='h000004b8;
    rd_cycle[ 2846] = 1'b0;  wr_cycle[ 2846] = 1'b1;  addr_rom[ 2846]='h00000610;  wr_data_rom[ 2846]='h0000036c;
    rd_cycle[ 2847] = 1'b0;  wr_cycle[ 2847] = 1'b1;  addr_rom[ 2847]='h00000c98;  wr_data_rom[ 2847]='h00000110;
    rd_cycle[ 2848] = 1'b0;  wr_cycle[ 2848] = 1'b1;  addr_rom[ 2848]='h00000160;  wr_data_rom[ 2848]='h00000ddd;
    rd_cycle[ 2849] = 1'b0;  wr_cycle[ 2849] = 1'b1;  addr_rom[ 2849]='h00000d0c;  wr_data_rom[ 2849]='h000002e4;
    rd_cycle[ 2850] = 1'b0;  wr_cycle[ 2850] = 1'b1;  addr_rom[ 2850]='h00000f28;  wr_data_rom[ 2850]='h00000c19;
    rd_cycle[ 2851] = 1'b0;  wr_cycle[ 2851] = 1'b1;  addr_rom[ 2851]='h00000504;  wr_data_rom[ 2851]='h00000f2b;
    rd_cycle[ 2852] = 1'b1;  wr_cycle[ 2852] = 1'b0;  addr_rom[ 2852]='h00000b18;  wr_data_rom[ 2852]='h00000000;
    rd_cycle[ 2853] = 1'b0;  wr_cycle[ 2853] = 1'b1;  addr_rom[ 2853]='h00000534;  wr_data_rom[ 2853]='h00000f94;
    rd_cycle[ 2854] = 1'b0;  wr_cycle[ 2854] = 1'b1;  addr_rom[ 2854]='h000003dc;  wr_data_rom[ 2854]='h00000653;
    rd_cycle[ 2855] = 1'b0;  wr_cycle[ 2855] = 1'b1;  addr_rom[ 2855]='h000007b0;  wr_data_rom[ 2855]='h0000094b;
    rd_cycle[ 2856] = 1'b1;  wr_cycle[ 2856] = 1'b0;  addr_rom[ 2856]='h00000e58;  wr_data_rom[ 2856]='h00000000;
    rd_cycle[ 2857] = 1'b0;  wr_cycle[ 2857] = 1'b1;  addr_rom[ 2857]='h00000e58;  wr_data_rom[ 2857]='h00000c0a;
    rd_cycle[ 2858] = 1'b1;  wr_cycle[ 2858] = 1'b0;  addr_rom[ 2858]='h000001f8;  wr_data_rom[ 2858]='h00000000;
    rd_cycle[ 2859] = 1'b1;  wr_cycle[ 2859] = 1'b0;  addr_rom[ 2859]='h00000dbc;  wr_data_rom[ 2859]='h00000000;
    rd_cycle[ 2860] = 1'b1;  wr_cycle[ 2860] = 1'b0;  addr_rom[ 2860]='h00000998;  wr_data_rom[ 2860]='h00000000;
    rd_cycle[ 2861] = 1'b0;  wr_cycle[ 2861] = 1'b1;  addr_rom[ 2861]='h00000abc;  wr_data_rom[ 2861]='h000001f0;
    rd_cycle[ 2862] = 1'b0;  wr_cycle[ 2862] = 1'b1;  addr_rom[ 2862]='h000006cc;  wr_data_rom[ 2862]='h00000243;
    rd_cycle[ 2863] = 1'b1;  wr_cycle[ 2863] = 1'b0;  addr_rom[ 2863]='h000004a8;  wr_data_rom[ 2863]='h00000000;
    rd_cycle[ 2864] = 1'b0;  wr_cycle[ 2864] = 1'b1;  addr_rom[ 2864]='h00000bf0;  wr_data_rom[ 2864]='h0000084f;
    rd_cycle[ 2865] = 1'b1;  wr_cycle[ 2865] = 1'b0;  addr_rom[ 2865]='h000003a0;  wr_data_rom[ 2865]='h00000000;
    rd_cycle[ 2866] = 1'b0;  wr_cycle[ 2866] = 1'b1;  addr_rom[ 2866]='h00000900;  wr_data_rom[ 2866]='h00000a61;
    rd_cycle[ 2867] = 1'b1;  wr_cycle[ 2867] = 1'b0;  addr_rom[ 2867]='h00000634;  wr_data_rom[ 2867]='h00000000;
    rd_cycle[ 2868] = 1'b1;  wr_cycle[ 2868] = 1'b0;  addr_rom[ 2868]='h00000874;  wr_data_rom[ 2868]='h00000000;
    rd_cycle[ 2869] = 1'b0;  wr_cycle[ 2869] = 1'b1;  addr_rom[ 2869]='h000007bc;  wr_data_rom[ 2869]='h00000d59;
    rd_cycle[ 2870] = 1'b1;  wr_cycle[ 2870] = 1'b0;  addr_rom[ 2870]='h00000028;  wr_data_rom[ 2870]='h00000000;
    rd_cycle[ 2871] = 1'b0;  wr_cycle[ 2871] = 1'b1;  addr_rom[ 2871]='h000003cc;  wr_data_rom[ 2871]='h00000907;
    rd_cycle[ 2872] = 1'b1;  wr_cycle[ 2872] = 1'b0;  addr_rom[ 2872]='h00000534;  wr_data_rom[ 2872]='h00000000;
    rd_cycle[ 2873] = 1'b0;  wr_cycle[ 2873] = 1'b1;  addr_rom[ 2873]='h0000054c;  wr_data_rom[ 2873]='h0000092d;
    rd_cycle[ 2874] = 1'b1;  wr_cycle[ 2874] = 1'b0;  addr_rom[ 2874]='h00000538;  wr_data_rom[ 2874]='h00000000;
    rd_cycle[ 2875] = 1'b1;  wr_cycle[ 2875] = 1'b0;  addr_rom[ 2875]='h00000f64;  wr_data_rom[ 2875]='h00000000;
    rd_cycle[ 2876] = 1'b1;  wr_cycle[ 2876] = 1'b0;  addr_rom[ 2876]='h000001d4;  wr_data_rom[ 2876]='h00000000;
    rd_cycle[ 2877] = 1'b1;  wr_cycle[ 2877] = 1'b0;  addr_rom[ 2877]='h00000cac;  wr_data_rom[ 2877]='h00000000;
    rd_cycle[ 2878] = 1'b0;  wr_cycle[ 2878] = 1'b1;  addr_rom[ 2878]='h0000039c;  wr_data_rom[ 2878]='h0000039c;
    rd_cycle[ 2879] = 1'b1;  wr_cycle[ 2879] = 1'b0;  addr_rom[ 2879]='h00000920;  wr_data_rom[ 2879]='h00000000;
    rd_cycle[ 2880] = 1'b0;  wr_cycle[ 2880] = 1'b1;  addr_rom[ 2880]='h00000bb0;  wr_data_rom[ 2880]='h000001f6;
    rd_cycle[ 2881] = 1'b1;  wr_cycle[ 2881] = 1'b0;  addr_rom[ 2881]='h00000cf0;  wr_data_rom[ 2881]='h00000000;
    rd_cycle[ 2882] = 1'b1;  wr_cycle[ 2882] = 1'b0;  addr_rom[ 2882]='h000001d8;  wr_data_rom[ 2882]='h00000000;
    rd_cycle[ 2883] = 1'b0;  wr_cycle[ 2883] = 1'b1;  addr_rom[ 2883]='h00000a9c;  wr_data_rom[ 2883]='h00000c4b;
    rd_cycle[ 2884] = 1'b0;  wr_cycle[ 2884] = 1'b1;  addr_rom[ 2884]='h000003a0;  wr_data_rom[ 2884]='h00000e02;
    rd_cycle[ 2885] = 1'b0;  wr_cycle[ 2885] = 1'b1;  addr_rom[ 2885]='h00000f64;  wr_data_rom[ 2885]='h00000a48;
    rd_cycle[ 2886] = 1'b1;  wr_cycle[ 2886] = 1'b0;  addr_rom[ 2886]='h00000964;  wr_data_rom[ 2886]='h00000000;
    rd_cycle[ 2887] = 1'b1;  wr_cycle[ 2887] = 1'b0;  addr_rom[ 2887]='h00000f94;  wr_data_rom[ 2887]='h00000000;
    rd_cycle[ 2888] = 1'b1;  wr_cycle[ 2888] = 1'b0;  addr_rom[ 2888]='h00000d90;  wr_data_rom[ 2888]='h00000000;
    rd_cycle[ 2889] = 1'b1;  wr_cycle[ 2889] = 1'b0;  addr_rom[ 2889]='h00000dc8;  wr_data_rom[ 2889]='h00000000;
    rd_cycle[ 2890] = 1'b1;  wr_cycle[ 2890] = 1'b0;  addr_rom[ 2890]='h000002ac;  wr_data_rom[ 2890]='h00000000;
    rd_cycle[ 2891] = 1'b0;  wr_cycle[ 2891] = 1'b1;  addr_rom[ 2891]='h00000598;  wr_data_rom[ 2891]='h0000079e;
    rd_cycle[ 2892] = 1'b1;  wr_cycle[ 2892] = 1'b0;  addr_rom[ 2892]='h00000d34;  wr_data_rom[ 2892]='h00000000;
    rd_cycle[ 2893] = 1'b0;  wr_cycle[ 2893] = 1'b1;  addr_rom[ 2893]='h000007e4;  wr_data_rom[ 2893]='h000005ad;
    rd_cycle[ 2894] = 1'b0;  wr_cycle[ 2894] = 1'b1;  addr_rom[ 2894]='h00000ad4;  wr_data_rom[ 2894]='h00000836;
    rd_cycle[ 2895] = 1'b1;  wr_cycle[ 2895] = 1'b0;  addr_rom[ 2895]='h00000874;  wr_data_rom[ 2895]='h00000000;
    rd_cycle[ 2896] = 1'b1;  wr_cycle[ 2896] = 1'b0;  addr_rom[ 2896]='h00000f00;  wr_data_rom[ 2896]='h00000000;
    rd_cycle[ 2897] = 1'b1;  wr_cycle[ 2897] = 1'b0;  addr_rom[ 2897]='h000009d8;  wr_data_rom[ 2897]='h00000000;
    rd_cycle[ 2898] = 1'b0;  wr_cycle[ 2898] = 1'b1;  addr_rom[ 2898]='h000008a8;  wr_data_rom[ 2898]='h00000d42;
    rd_cycle[ 2899] = 1'b1;  wr_cycle[ 2899] = 1'b0;  addr_rom[ 2899]='h00000944;  wr_data_rom[ 2899]='h00000000;
    rd_cycle[ 2900] = 1'b1;  wr_cycle[ 2900] = 1'b0;  addr_rom[ 2900]='h00000698;  wr_data_rom[ 2900]='h00000000;
    rd_cycle[ 2901] = 1'b1;  wr_cycle[ 2901] = 1'b0;  addr_rom[ 2901]='h00000d58;  wr_data_rom[ 2901]='h00000000;
    rd_cycle[ 2902] = 1'b1;  wr_cycle[ 2902] = 1'b0;  addr_rom[ 2902]='h00000498;  wr_data_rom[ 2902]='h00000000;
    rd_cycle[ 2903] = 1'b1;  wr_cycle[ 2903] = 1'b0;  addr_rom[ 2903]='h000002c4;  wr_data_rom[ 2903]='h00000000;
    rd_cycle[ 2904] = 1'b1;  wr_cycle[ 2904] = 1'b0;  addr_rom[ 2904]='h0000091c;  wr_data_rom[ 2904]='h00000000;
    rd_cycle[ 2905] = 1'b0;  wr_cycle[ 2905] = 1'b1;  addr_rom[ 2905]='h000007f8;  wr_data_rom[ 2905]='h00000b7e;
    rd_cycle[ 2906] = 1'b0;  wr_cycle[ 2906] = 1'b1;  addr_rom[ 2906]='h00000944;  wr_data_rom[ 2906]='h00000884;
    rd_cycle[ 2907] = 1'b1;  wr_cycle[ 2907] = 1'b0;  addr_rom[ 2907]='h00000db8;  wr_data_rom[ 2907]='h00000000;
    rd_cycle[ 2908] = 1'b1;  wr_cycle[ 2908] = 1'b0;  addr_rom[ 2908]='h00000f64;  wr_data_rom[ 2908]='h00000000;
    rd_cycle[ 2909] = 1'b1;  wr_cycle[ 2909] = 1'b0;  addr_rom[ 2909]='h000007f8;  wr_data_rom[ 2909]='h00000000;
    rd_cycle[ 2910] = 1'b1;  wr_cycle[ 2910] = 1'b0;  addr_rom[ 2910]='h00000df0;  wr_data_rom[ 2910]='h00000000;
    rd_cycle[ 2911] = 1'b1;  wr_cycle[ 2911] = 1'b0;  addr_rom[ 2911]='h000009fc;  wr_data_rom[ 2911]='h00000000;
    rd_cycle[ 2912] = 1'b1;  wr_cycle[ 2912] = 1'b0;  addr_rom[ 2912]='h00000ca8;  wr_data_rom[ 2912]='h00000000;
    rd_cycle[ 2913] = 1'b0;  wr_cycle[ 2913] = 1'b1;  addr_rom[ 2913]='h00000f8c;  wr_data_rom[ 2913]='h00000a0e;
    rd_cycle[ 2914] = 1'b0;  wr_cycle[ 2914] = 1'b1;  addr_rom[ 2914]='h00000c7c;  wr_data_rom[ 2914]='h000007c3;
    rd_cycle[ 2915] = 1'b1;  wr_cycle[ 2915] = 1'b0;  addr_rom[ 2915]='h00000910;  wr_data_rom[ 2915]='h00000000;
    rd_cycle[ 2916] = 1'b1;  wr_cycle[ 2916] = 1'b0;  addr_rom[ 2916]='h00000860;  wr_data_rom[ 2916]='h00000000;
    rd_cycle[ 2917] = 1'b0;  wr_cycle[ 2917] = 1'b1;  addr_rom[ 2917]='h000005e8;  wr_data_rom[ 2917]='h00000cec;
    rd_cycle[ 2918] = 1'b1;  wr_cycle[ 2918] = 1'b0;  addr_rom[ 2918]='h00000ef4;  wr_data_rom[ 2918]='h00000000;
    rd_cycle[ 2919] = 1'b0;  wr_cycle[ 2919] = 1'b1;  addr_rom[ 2919]='h0000005c;  wr_data_rom[ 2919]='h00000e7a;
    rd_cycle[ 2920] = 1'b1;  wr_cycle[ 2920] = 1'b0;  addr_rom[ 2920]='h000001d4;  wr_data_rom[ 2920]='h00000000;
    rd_cycle[ 2921] = 1'b0;  wr_cycle[ 2921] = 1'b1;  addr_rom[ 2921]='h00000db8;  wr_data_rom[ 2921]='h000004a0;
    rd_cycle[ 2922] = 1'b1;  wr_cycle[ 2922] = 1'b0;  addr_rom[ 2922]='h000001a4;  wr_data_rom[ 2922]='h00000000;
    rd_cycle[ 2923] = 1'b1;  wr_cycle[ 2923] = 1'b0;  addr_rom[ 2923]='h00000d2c;  wr_data_rom[ 2923]='h00000000;
    rd_cycle[ 2924] = 1'b1;  wr_cycle[ 2924] = 1'b0;  addr_rom[ 2924]='h000005d0;  wr_data_rom[ 2924]='h00000000;
    rd_cycle[ 2925] = 1'b1;  wr_cycle[ 2925] = 1'b0;  addr_rom[ 2925]='h0000035c;  wr_data_rom[ 2925]='h00000000;
    rd_cycle[ 2926] = 1'b0;  wr_cycle[ 2926] = 1'b1;  addr_rom[ 2926]='h00000ba4;  wr_data_rom[ 2926]='h00000882;
    rd_cycle[ 2927] = 1'b0;  wr_cycle[ 2927] = 1'b1;  addr_rom[ 2927]='h00000ef0;  wr_data_rom[ 2927]='h00000c51;
    rd_cycle[ 2928] = 1'b0;  wr_cycle[ 2928] = 1'b1;  addr_rom[ 2928]='h000006c8;  wr_data_rom[ 2928]='h00000a62;
    rd_cycle[ 2929] = 1'b0;  wr_cycle[ 2929] = 1'b1;  addr_rom[ 2929]='h000004b8;  wr_data_rom[ 2929]='h00000496;
    rd_cycle[ 2930] = 1'b1;  wr_cycle[ 2930] = 1'b0;  addr_rom[ 2930]='h00000574;  wr_data_rom[ 2930]='h00000000;
    rd_cycle[ 2931] = 1'b1;  wr_cycle[ 2931] = 1'b0;  addr_rom[ 2931]='h000009a4;  wr_data_rom[ 2931]='h00000000;
    rd_cycle[ 2932] = 1'b1;  wr_cycle[ 2932] = 1'b0;  addr_rom[ 2932]='h000001d4;  wr_data_rom[ 2932]='h00000000;
    rd_cycle[ 2933] = 1'b0;  wr_cycle[ 2933] = 1'b1;  addr_rom[ 2933]='h00000dc0;  wr_data_rom[ 2933]='h000002cd;
    rd_cycle[ 2934] = 1'b0;  wr_cycle[ 2934] = 1'b1;  addr_rom[ 2934]='h00000ee0;  wr_data_rom[ 2934]='h00000453;
    rd_cycle[ 2935] = 1'b0;  wr_cycle[ 2935] = 1'b1;  addr_rom[ 2935]='h00000dbc;  wr_data_rom[ 2935]='h00000a42;
    rd_cycle[ 2936] = 1'b1;  wr_cycle[ 2936] = 1'b0;  addr_rom[ 2936]='h00000008;  wr_data_rom[ 2936]='h00000000;
    rd_cycle[ 2937] = 1'b1;  wr_cycle[ 2937] = 1'b0;  addr_rom[ 2937]='h00000be8;  wr_data_rom[ 2937]='h00000000;
    rd_cycle[ 2938] = 1'b0;  wr_cycle[ 2938] = 1'b1;  addr_rom[ 2938]='h00000378;  wr_data_rom[ 2938]='h00000195;
    rd_cycle[ 2939] = 1'b0;  wr_cycle[ 2939] = 1'b1;  addr_rom[ 2939]='h00000e30;  wr_data_rom[ 2939]='h0000032b;
    rd_cycle[ 2940] = 1'b0;  wr_cycle[ 2940] = 1'b1;  addr_rom[ 2940]='h00000408;  wr_data_rom[ 2940]='h00000614;
    rd_cycle[ 2941] = 1'b1;  wr_cycle[ 2941] = 1'b0;  addr_rom[ 2941]='h00000034;  wr_data_rom[ 2941]='h00000000;
    rd_cycle[ 2942] = 1'b1;  wr_cycle[ 2942] = 1'b0;  addr_rom[ 2942]='h00000a64;  wr_data_rom[ 2942]='h00000000;
    rd_cycle[ 2943] = 1'b1;  wr_cycle[ 2943] = 1'b0;  addr_rom[ 2943]='h00000400;  wr_data_rom[ 2943]='h00000000;
    rd_cycle[ 2944] = 1'b1;  wr_cycle[ 2944] = 1'b0;  addr_rom[ 2944]='h0000018c;  wr_data_rom[ 2944]='h00000000;
    rd_cycle[ 2945] = 1'b0;  wr_cycle[ 2945] = 1'b1;  addr_rom[ 2945]='h0000028c;  wr_data_rom[ 2945]='h0000038f;
    rd_cycle[ 2946] = 1'b0;  wr_cycle[ 2946] = 1'b1;  addr_rom[ 2946]='h00000384;  wr_data_rom[ 2946]='h00000212;
    rd_cycle[ 2947] = 1'b1;  wr_cycle[ 2947] = 1'b0;  addr_rom[ 2947]='h00000150;  wr_data_rom[ 2947]='h00000000;
    rd_cycle[ 2948] = 1'b0;  wr_cycle[ 2948] = 1'b1;  addr_rom[ 2948]='h000003b4;  wr_data_rom[ 2948]='h000008fc;
    rd_cycle[ 2949] = 1'b1;  wr_cycle[ 2949] = 1'b0;  addr_rom[ 2949]='h00000254;  wr_data_rom[ 2949]='h00000000;
    rd_cycle[ 2950] = 1'b0;  wr_cycle[ 2950] = 1'b1;  addr_rom[ 2950]='h00000d80;  wr_data_rom[ 2950]='h0000058c;
    rd_cycle[ 2951] = 1'b1;  wr_cycle[ 2951] = 1'b0;  addr_rom[ 2951]='h00000198;  wr_data_rom[ 2951]='h00000000;
    rd_cycle[ 2952] = 1'b0;  wr_cycle[ 2952] = 1'b1;  addr_rom[ 2952]='h0000074c;  wr_data_rom[ 2952]='h00000d4c;
    rd_cycle[ 2953] = 1'b0;  wr_cycle[ 2953] = 1'b1;  addr_rom[ 2953]='h00000374;  wr_data_rom[ 2953]='h00000d7d;
    rd_cycle[ 2954] = 1'b0;  wr_cycle[ 2954] = 1'b1;  addr_rom[ 2954]='h000004e4;  wr_data_rom[ 2954]='h00000521;
    rd_cycle[ 2955] = 1'b1;  wr_cycle[ 2955] = 1'b0;  addr_rom[ 2955]='h0000049c;  wr_data_rom[ 2955]='h00000000;
    rd_cycle[ 2956] = 1'b0;  wr_cycle[ 2956] = 1'b1;  addr_rom[ 2956]='h000006e4;  wr_data_rom[ 2956]='h00000143;
    rd_cycle[ 2957] = 1'b0;  wr_cycle[ 2957] = 1'b1;  addr_rom[ 2957]='h00000d00;  wr_data_rom[ 2957]='h0000095b;
    rd_cycle[ 2958] = 1'b1;  wr_cycle[ 2958] = 1'b0;  addr_rom[ 2958]='h000001e8;  wr_data_rom[ 2958]='h00000000;
    rd_cycle[ 2959] = 1'b1;  wr_cycle[ 2959] = 1'b0;  addr_rom[ 2959]='h00000abc;  wr_data_rom[ 2959]='h00000000;
    rd_cycle[ 2960] = 1'b0;  wr_cycle[ 2960] = 1'b1;  addr_rom[ 2960]='h00000df4;  wr_data_rom[ 2960]='h000003c0;
    rd_cycle[ 2961] = 1'b1;  wr_cycle[ 2961] = 1'b0;  addr_rom[ 2961]='h00000328;  wr_data_rom[ 2961]='h00000000;
    rd_cycle[ 2962] = 1'b1;  wr_cycle[ 2962] = 1'b0;  addr_rom[ 2962]='h00000f30;  wr_data_rom[ 2962]='h00000000;
    rd_cycle[ 2963] = 1'b1;  wr_cycle[ 2963] = 1'b0;  addr_rom[ 2963]='h00000ee0;  wr_data_rom[ 2963]='h00000000;
    rd_cycle[ 2964] = 1'b0;  wr_cycle[ 2964] = 1'b1;  addr_rom[ 2964]='h000004a0;  wr_data_rom[ 2964]='h00000b12;
    rd_cycle[ 2965] = 1'b0;  wr_cycle[ 2965] = 1'b1;  addr_rom[ 2965]='h00000764;  wr_data_rom[ 2965]='h00000911;
    rd_cycle[ 2966] = 1'b0;  wr_cycle[ 2966] = 1'b1;  addr_rom[ 2966]='h00000424;  wr_data_rom[ 2966]='h00000de1;
    rd_cycle[ 2967] = 1'b0;  wr_cycle[ 2967] = 1'b1;  addr_rom[ 2967]='h00000a94;  wr_data_rom[ 2967]='h00000eb7;
    rd_cycle[ 2968] = 1'b1;  wr_cycle[ 2968] = 1'b0;  addr_rom[ 2968]='h00000b14;  wr_data_rom[ 2968]='h00000000;
    rd_cycle[ 2969] = 1'b1;  wr_cycle[ 2969] = 1'b0;  addr_rom[ 2969]='h0000031c;  wr_data_rom[ 2969]='h00000000;
    rd_cycle[ 2970] = 1'b0;  wr_cycle[ 2970] = 1'b1;  addr_rom[ 2970]='h00000adc;  wr_data_rom[ 2970]='h000007cd;
    rd_cycle[ 2971] = 1'b1;  wr_cycle[ 2971] = 1'b0;  addr_rom[ 2971]='h00000d20;  wr_data_rom[ 2971]='h00000000;
    rd_cycle[ 2972] = 1'b0;  wr_cycle[ 2972] = 1'b1;  addr_rom[ 2972]='h000009e4;  wr_data_rom[ 2972]='h00000a4f;
    rd_cycle[ 2973] = 1'b0;  wr_cycle[ 2973] = 1'b1;  addr_rom[ 2973]='h00000418;  wr_data_rom[ 2973]='h00000e48;
    rd_cycle[ 2974] = 1'b0;  wr_cycle[ 2974] = 1'b1;  addr_rom[ 2974]='h00000c10;  wr_data_rom[ 2974]='h00000189;
    rd_cycle[ 2975] = 1'b0;  wr_cycle[ 2975] = 1'b1;  addr_rom[ 2975]='h00000c18;  wr_data_rom[ 2975]='h000009ad;
    rd_cycle[ 2976] = 1'b0;  wr_cycle[ 2976] = 1'b1;  addr_rom[ 2976]='h00000960;  wr_data_rom[ 2976]='h00000c9a;
    rd_cycle[ 2977] = 1'b0;  wr_cycle[ 2977] = 1'b1;  addr_rom[ 2977]='h00000e08;  wr_data_rom[ 2977]='h0000037b;
    rd_cycle[ 2978] = 1'b0;  wr_cycle[ 2978] = 1'b1;  addr_rom[ 2978]='h00000788;  wr_data_rom[ 2978]='h000004b1;
    rd_cycle[ 2979] = 1'b0;  wr_cycle[ 2979] = 1'b1;  addr_rom[ 2979]='h00000090;  wr_data_rom[ 2979]='h00000cca;
    rd_cycle[ 2980] = 1'b0;  wr_cycle[ 2980] = 1'b1;  addr_rom[ 2980]='h00000cf8;  wr_data_rom[ 2980]='h00000946;
    rd_cycle[ 2981] = 1'b1;  wr_cycle[ 2981] = 1'b0;  addr_rom[ 2981]='h00000784;  wr_data_rom[ 2981]='h00000000;
    rd_cycle[ 2982] = 1'b1;  wr_cycle[ 2982] = 1'b0;  addr_rom[ 2982]='h000002e0;  wr_data_rom[ 2982]='h00000000;
    rd_cycle[ 2983] = 1'b0;  wr_cycle[ 2983] = 1'b1;  addr_rom[ 2983]='h00000df0;  wr_data_rom[ 2983]='h00000cef;
    rd_cycle[ 2984] = 1'b0;  wr_cycle[ 2984] = 1'b1;  addr_rom[ 2984]='h00000bd0;  wr_data_rom[ 2984]='h000000ad;
    rd_cycle[ 2985] = 1'b0;  wr_cycle[ 2985] = 1'b1;  addr_rom[ 2985]='h000006e4;  wr_data_rom[ 2985]='h00000c0a;
    rd_cycle[ 2986] = 1'b1;  wr_cycle[ 2986] = 1'b0;  addr_rom[ 2986]='h00000504;  wr_data_rom[ 2986]='h00000000;
    rd_cycle[ 2987] = 1'b0;  wr_cycle[ 2987] = 1'b1;  addr_rom[ 2987]='h0000085c;  wr_data_rom[ 2987]='h00000e2f;
    rd_cycle[ 2988] = 1'b0;  wr_cycle[ 2988] = 1'b1;  addr_rom[ 2988]='h00000098;  wr_data_rom[ 2988]='h00000bb1;
    rd_cycle[ 2989] = 1'b1;  wr_cycle[ 2989] = 1'b0;  addr_rom[ 2989]='h00000b00;  wr_data_rom[ 2989]='h00000000;
    rd_cycle[ 2990] = 1'b1;  wr_cycle[ 2990] = 1'b0;  addr_rom[ 2990]='h00000e20;  wr_data_rom[ 2990]='h00000000;
    rd_cycle[ 2991] = 1'b1;  wr_cycle[ 2991] = 1'b0;  addr_rom[ 2991]='h000005d8;  wr_data_rom[ 2991]='h00000000;
    rd_cycle[ 2992] = 1'b0;  wr_cycle[ 2992] = 1'b1;  addr_rom[ 2992]='h000003e4;  wr_data_rom[ 2992]='h0000088a;
    rd_cycle[ 2993] = 1'b1;  wr_cycle[ 2993] = 1'b0;  addr_rom[ 2993]='h00000e30;  wr_data_rom[ 2993]='h00000000;
    rd_cycle[ 2994] = 1'b0;  wr_cycle[ 2994] = 1'b1;  addr_rom[ 2994]='h00000eb0;  wr_data_rom[ 2994]='h0000060f;
    rd_cycle[ 2995] = 1'b1;  wr_cycle[ 2995] = 1'b0;  addr_rom[ 2995]='h00000c00;  wr_data_rom[ 2995]='h00000000;
    rd_cycle[ 2996] = 1'b0;  wr_cycle[ 2996] = 1'b1;  addr_rom[ 2996]='h0000027c;  wr_data_rom[ 2996]='h00000f8a;
    rd_cycle[ 2997] = 1'b1;  wr_cycle[ 2997] = 1'b0;  addr_rom[ 2997]='h00000478;  wr_data_rom[ 2997]='h00000000;
    rd_cycle[ 2998] = 1'b1;  wr_cycle[ 2998] = 1'b0;  addr_rom[ 2998]='h00000794;  wr_data_rom[ 2998]='h00000000;
    rd_cycle[ 2999] = 1'b0;  wr_cycle[ 2999] = 1'b1;  addr_rom[ 2999]='h000001d4;  wr_data_rom[ 2999]='h000004b6;
    rd_cycle[ 3000] = 1'b0;  wr_cycle[ 3000] = 1'b1;  addr_rom[ 3000]='h00000ac4;  wr_data_rom[ 3000]='h000007f6;
    rd_cycle[ 3001] = 1'b0;  wr_cycle[ 3001] = 1'b1;  addr_rom[ 3001]='h000004b8;  wr_data_rom[ 3001]='h000001b1;
    rd_cycle[ 3002] = 1'b1;  wr_cycle[ 3002] = 1'b0;  addr_rom[ 3002]='h0000008c;  wr_data_rom[ 3002]='h00000000;
    rd_cycle[ 3003] = 1'b0;  wr_cycle[ 3003] = 1'b1;  addr_rom[ 3003]='h00000830;  wr_data_rom[ 3003]='h000003c3;
    rd_cycle[ 3004] = 1'b0;  wr_cycle[ 3004] = 1'b1;  addr_rom[ 3004]='h00000d68;  wr_data_rom[ 3004]='h00000d6e;
    rd_cycle[ 3005] = 1'b0;  wr_cycle[ 3005] = 1'b1;  addr_rom[ 3005]='h000005fc;  wr_data_rom[ 3005]='h00000199;
    rd_cycle[ 3006] = 1'b1;  wr_cycle[ 3006] = 1'b0;  addr_rom[ 3006]='h00000340;  wr_data_rom[ 3006]='h00000000;
    rd_cycle[ 3007] = 1'b1;  wr_cycle[ 3007] = 1'b0;  addr_rom[ 3007]='h0000032c;  wr_data_rom[ 3007]='h00000000;
    rd_cycle[ 3008] = 1'b1;  wr_cycle[ 3008] = 1'b0;  addr_rom[ 3008]='h00000638;  wr_data_rom[ 3008]='h00000000;
    rd_cycle[ 3009] = 1'b0;  wr_cycle[ 3009] = 1'b1;  addr_rom[ 3009]='h00000c94;  wr_data_rom[ 3009]='h000004bc;
    rd_cycle[ 3010] = 1'b0;  wr_cycle[ 3010] = 1'b1;  addr_rom[ 3010]='h000007d0;  wr_data_rom[ 3010]='h00000566;
    rd_cycle[ 3011] = 1'b1;  wr_cycle[ 3011] = 1'b0;  addr_rom[ 3011]='h00000f84;  wr_data_rom[ 3011]='h00000000;
    rd_cycle[ 3012] = 1'b0;  wr_cycle[ 3012] = 1'b1;  addr_rom[ 3012]='h00000cf4;  wr_data_rom[ 3012]='h00000cb5;
    rd_cycle[ 3013] = 1'b1;  wr_cycle[ 3013] = 1'b0;  addr_rom[ 3013]='h000009c0;  wr_data_rom[ 3013]='h00000000;
    rd_cycle[ 3014] = 1'b0;  wr_cycle[ 3014] = 1'b1;  addr_rom[ 3014]='h00000b74;  wr_data_rom[ 3014]='h00000133;
    rd_cycle[ 3015] = 1'b1;  wr_cycle[ 3015] = 1'b0;  addr_rom[ 3015]='h000002c0;  wr_data_rom[ 3015]='h00000000;
    rd_cycle[ 3016] = 1'b0;  wr_cycle[ 3016] = 1'b1;  addr_rom[ 3016]='h00000b24;  wr_data_rom[ 3016]='h00000f83;
    rd_cycle[ 3017] = 1'b1;  wr_cycle[ 3017] = 1'b0;  addr_rom[ 3017]='h00000b08;  wr_data_rom[ 3017]='h00000000;
    rd_cycle[ 3018] = 1'b1;  wr_cycle[ 3018] = 1'b0;  addr_rom[ 3018]='h00000ec0;  wr_data_rom[ 3018]='h00000000;
    rd_cycle[ 3019] = 1'b0;  wr_cycle[ 3019] = 1'b1;  addr_rom[ 3019]='h00000208;  wr_data_rom[ 3019]='h00000bcd;
    rd_cycle[ 3020] = 1'b0;  wr_cycle[ 3020] = 1'b1;  addr_rom[ 3020]='h00000748;  wr_data_rom[ 3020]='h00000f59;
    rd_cycle[ 3021] = 1'b1;  wr_cycle[ 3021] = 1'b0;  addr_rom[ 3021]='h00000034;  wr_data_rom[ 3021]='h00000000;
    rd_cycle[ 3022] = 1'b0;  wr_cycle[ 3022] = 1'b1;  addr_rom[ 3022]='h00000888;  wr_data_rom[ 3022]='h00000b85;
    rd_cycle[ 3023] = 1'b1;  wr_cycle[ 3023] = 1'b0;  addr_rom[ 3023]='h00000aa4;  wr_data_rom[ 3023]='h00000000;
    rd_cycle[ 3024] = 1'b0;  wr_cycle[ 3024] = 1'b1;  addr_rom[ 3024]='h000009e0;  wr_data_rom[ 3024]='h00000257;
    rd_cycle[ 3025] = 1'b0;  wr_cycle[ 3025] = 1'b1;  addr_rom[ 3025]='h000002d8;  wr_data_rom[ 3025]='h00000c56;
    rd_cycle[ 3026] = 1'b1;  wr_cycle[ 3026] = 1'b0;  addr_rom[ 3026]='h00000dcc;  wr_data_rom[ 3026]='h00000000;
    rd_cycle[ 3027] = 1'b1;  wr_cycle[ 3027] = 1'b0;  addr_rom[ 3027]='h0000011c;  wr_data_rom[ 3027]='h00000000;
    rd_cycle[ 3028] = 1'b1;  wr_cycle[ 3028] = 1'b0;  addr_rom[ 3028]='h00000890;  wr_data_rom[ 3028]='h00000000;
    rd_cycle[ 3029] = 1'b1;  wr_cycle[ 3029] = 1'b0;  addr_rom[ 3029]='h00000f10;  wr_data_rom[ 3029]='h00000000;
    rd_cycle[ 3030] = 1'b0;  wr_cycle[ 3030] = 1'b1;  addr_rom[ 3030]='h00000b78;  wr_data_rom[ 3030]='h00000072;
    rd_cycle[ 3031] = 1'b0;  wr_cycle[ 3031] = 1'b1;  addr_rom[ 3031]='h00000bb8;  wr_data_rom[ 3031]='h0000073b;
    rd_cycle[ 3032] = 1'b1;  wr_cycle[ 3032] = 1'b0;  addr_rom[ 3032]='h00000608;  wr_data_rom[ 3032]='h00000000;
    rd_cycle[ 3033] = 1'b1;  wr_cycle[ 3033] = 1'b0;  addr_rom[ 3033]='h00000254;  wr_data_rom[ 3033]='h00000000;
    rd_cycle[ 3034] = 1'b1;  wr_cycle[ 3034] = 1'b0;  addr_rom[ 3034]='h0000032c;  wr_data_rom[ 3034]='h00000000;
    rd_cycle[ 3035] = 1'b0;  wr_cycle[ 3035] = 1'b1;  addr_rom[ 3035]='h000005ac;  wr_data_rom[ 3035]='h00000142;
    rd_cycle[ 3036] = 1'b0;  wr_cycle[ 3036] = 1'b1;  addr_rom[ 3036]='h00000e64;  wr_data_rom[ 3036]='h000009a4;
    rd_cycle[ 3037] = 1'b0;  wr_cycle[ 3037] = 1'b1;  addr_rom[ 3037]='h00000aa0;  wr_data_rom[ 3037]='h000000f2;
    rd_cycle[ 3038] = 1'b0;  wr_cycle[ 3038] = 1'b1;  addr_rom[ 3038]='h00000320;  wr_data_rom[ 3038]='h00000f3f;
    rd_cycle[ 3039] = 1'b0;  wr_cycle[ 3039] = 1'b1;  addr_rom[ 3039]='h00000298;  wr_data_rom[ 3039]='h00000207;
    rd_cycle[ 3040] = 1'b1;  wr_cycle[ 3040] = 1'b0;  addr_rom[ 3040]='h000004a8;  wr_data_rom[ 3040]='h00000000;
    rd_cycle[ 3041] = 1'b1;  wr_cycle[ 3041] = 1'b0;  addr_rom[ 3041]='h00000a84;  wr_data_rom[ 3041]='h00000000;
    rd_cycle[ 3042] = 1'b0;  wr_cycle[ 3042] = 1'b1;  addr_rom[ 3042]='h000000e0;  wr_data_rom[ 3042]='h00000c56;
    rd_cycle[ 3043] = 1'b0;  wr_cycle[ 3043] = 1'b1;  addr_rom[ 3043]='h00000be8;  wr_data_rom[ 3043]='h00000860;
    rd_cycle[ 3044] = 1'b1;  wr_cycle[ 3044] = 1'b0;  addr_rom[ 3044]='h000007f4;  wr_data_rom[ 3044]='h00000000;
    rd_cycle[ 3045] = 1'b1;  wr_cycle[ 3045] = 1'b0;  addr_rom[ 3045]='h0000005c;  wr_data_rom[ 3045]='h00000000;
    rd_cycle[ 3046] = 1'b1;  wr_cycle[ 3046] = 1'b0;  addr_rom[ 3046]='h0000052c;  wr_data_rom[ 3046]='h00000000;
    rd_cycle[ 3047] = 1'b1;  wr_cycle[ 3047] = 1'b0;  addr_rom[ 3047]='h00000a4c;  wr_data_rom[ 3047]='h00000000;
    rd_cycle[ 3048] = 1'b0;  wr_cycle[ 3048] = 1'b1;  addr_rom[ 3048]='h00000138;  wr_data_rom[ 3048]='h00000e15;
    rd_cycle[ 3049] = 1'b1;  wr_cycle[ 3049] = 1'b0;  addr_rom[ 3049]='h00000274;  wr_data_rom[ 3049]='h00000000;
    rd_cycle[ 3050] = 1'b0;  wr_cycle[ 3050] = 1'b1;  addr_rom[ 3050]='h00000d3c;  wr_data_rom[ 3050]='h00000306;
    rd_cycle[ 3051] = 1'b0;  wr_cycle[ 3051] = 1'b1;  addr_rom[ 3051]='h00000854;  wr_data_rom[ 3051]='h00000b36;
    rd_cycle[ 3052] = 1'b0;  wr_cycle[ 3052] = 1'b1;  addr_rom[ 3052]='h00000d64;  wr_data_rom[ 3052]='h00000eac;
    rd_cycle[ 3053] = 1'b1;  wr_cycle[ 3053] = 1'b0;  addr_rom[ 3053]='h00000380;  wr_data_rom[ 3053]='h00000000;
    rd_cycle[ 3054] = 1'b0;  wr_cycle[ 3054] = 1'b1;  addr_rom[ 3054]='h0000053c;  wr_data_rom[ 3054]='h00000a61;
    rd_cycle[ 3055] = 1'b0;  wr_cycle[ 3055] = 1'b1;  addr_rom[ 3055]='h00000eac;  wr_data_rom[ 3055]='h00000280;
    rd_cycle[ 3056] = 1'b0;  wr_cycle[ 3056] = 1'b1;  addr_rom[ 3056]='h000000e0;  wr_data_rom[ 3056]='h0000039e;
    rd_cycle[ 3057] = 1'b1;  wr_cycle[ 3057] = 1'b0;  addr_rom[ 3057]='h00000784;  wr_data_rom[ 3057]='h00000000;
    rd_cycle[ 3058] = 1'b1;  wr_cycle[ 3058] = 1'b0;  addr_rom[ 3058]='h00000a34;  wr_data_rom[ 3058]='h00000000;
    rd_cycle[ 3059] = 1'b1;  wr_cycle[ 3059] = 1'b0;  addr_rom[ 3059]='h00000a04;  wr_data_rom[ 3059]='h00000000;
    rd_cycle[ 3060] = 1'b1;  wr_cycle[ 3060] = 1'b0;  addr_rom[ 3060]='h00000a5c;  wr_data_rom[ 3060]='h00000000;
    rd_cycle[ 3061] = 1'b1;  wr_cycle[ 3061] = 1'b0;  addr_rom[ 3061]='h0000083c;  wr_data_rom[ 3061]='h00000000;
    rd_cycle[ 3062] = 1'b1;  wr_cycle[ 3062] = 1'b0;  addr_rom[ 3062]='h00000830;  wr_data_rom[ 3062]='h00000000;
    rd_cycle[ 3063] = 1'b1;  wr_cycle[ 3063] = 1'b0;  addr_rom[ 3063]='h000007e8;  wr_data_rom[ 3063]='h00000000;
    rd_cycle[ 3064] = 1'b0;  wr_cycle[ 3064] = 1'b1;  addr_rom[ 3064]='h00000dc0;  wr_data_rom[ 3064]='h00000065;
    rd_cycle[ 3065] = 1'b0;  wr_cycle[ 3065] = 1'b1;  addr_rom[ 3065]='h00000ee4;  wr_data_rom[ 3065]='h000006b5;
    rd_cycle[ 3066] = 1'b1;  wr_cycle[ 3066] = 1'b0;  addr_rom[ 3066]='h000006a0;  wr_data_rom[ 3066]='h00000000;
    rd_cycle[ 3067] = 1'b0;  wr_cycle[ 3067] = 1'b1;  addr_rom[ 3067]='h00000474;  wr_data_rom[ 3067]='h00000283;
    rd_cycle[ 3068] = 1'b0;  wr_cycle[ 3068] = 1'b1;  addr_rom[ 3068]='h00000f20;  wr_data_rom[ 3068]='h00000e64;
    rd_cycle[ 3069] = 1'b0;  wr_cycle[ 3069] = 1'b1;  addr_rom[ 3069]='h00000a1c;  wr_data_rom[ 3069]='h00000672;
    rd_cycle[ 3070] = 1'b0;  wr_cycle[ 3070] = 1'b1;  addr_rom[ 3070]='h00000acc;  wr_data_rom[ 3070]='h000002ca;
    rd_cycle[ 3071] = 1'b1;  wr_cycle[ 3071] = 1'b0;  addr_rom[ 3071]='h00000f04;  wr_data_rom[ 3071]='h00000000;
    rd_cycle[ 3072] = 1'b0;  wr_cycle[ 3072] = 1'b1;  addr_rom[ 3072]='h0000049c;  wr_data_rom[ 3072]='h00000ad4;
    rd_cycle[ 3073] = 1'b1;  wr_cycle[ 3073] = 1'b0;  addr_rom[ 3073]='h00000eb4;  wr_data_rom[ 3073]='h00000000;
    rd_cycle[ 3074] = 1'b0;  wr_cycle[ 3074] = 1'b1;  addr_rom[ 3074]='h00000550;  wr_data_rom[ 3074]='h00000551;
    rd_cycle[ 3075] = 1'b1;  wr_cycle[ 3075] = 1'b0;  addr_rom[ 3075]='h00000734;  wr_data_rom[ 3075]='h00000000;
    rd_cycle[ 3076] = 1'b1;  wr_cycle[ 3076] = 1'b0;  addr_rom[ 3076]='h00000414;  wr_data_rom[ 3076]='h00000000;
    rd_cycle[ 3077] = 1'b1;  wr_cycle[ 3077] = 1'b0;  addr_rom[ 3077]='h0000029c;  wr_data_rom[ 3077]='h00000000;
    rd_cycle[ 3078] = 1'b0;  wr_cycle[ 3078] = 1'b1;  addr_rom[ 3078]='h0000014c;  wr_data_rom[ 3078]='h00000267;
    rd_cycle[ 3079] = 1'b0;  wr_cycle[ 3079] = 1'b1;  addr_rom[ 3079]='h00000ea4;  wr_data_rom[ 3079]='h00000907;
    rd_cycle[ 3080] = 1'b1;  wr_cycle[ 3080] = 1'b0;  addr_rom[ 3080]='h0000070c;  wr_data_rom[ 3080]='h00000000;
    rd_cycle[ 3081] = 1'b0;  wr_cycle[ 3081] = 1'b1;  addr_rom[ 3081]='h00000af8;  wr_data_rom[ 3081]='h00000f14;
    rd_cycle[ 3082] = 1'b1;  wr_cycle[ 3082] = 1'b0;  addr_rom[ 3082]='h00000600;  wr_data_rom[ 3082]='h00000000;
    rd_cycle[ 3083] = 1'b1;  wr_cycle[ 3083] = 1'b0;  addr_rom[ 3083]='h00000418;  wr_data_rom[ 3083]='h00000000;
    rd_cycle[ 3084] = 1'b1;  wr_cycle[ 3084] = 1'b0;  addr_rom[ 3084]='h00000b80;  wr_data_rom[ 3084]='h00000000;
    rd_cycle[ 3085] = 1'b0;  wr_cycle[ 3085] = 1'b1;  addr_rom[ 3085]='h00000eb8;  wr_data_rom[ 3085]='h00000317;
    rd_cycle[ 3086] = 1'b1;  wr_cycle[ 3086] = 1'b0;  addr_rom[ 3086]='h000009bc;  wr_data_rom[ 3086]='h00000000;
    rd_cycle[ 3087] = 1'b1;  wr_cycle[ 3087] = 1'b0;  addr_rom[ 3087]='h00000c1c;  wr_data_rom[ 3087]='h00000000;
    rd_cycle[ 3088] = 1'b0;  wr_cycle[ 3088] = 1'b1;  addr_rom[ 3088]='h00000778;  wr_data_rom[ 3088]='h00000bf4;
    rd_cycle[ 3089] = 1'b1;  wr_cycle[ 3089] = 1'b0;  addr_rom[ 3089]='h000008c0;  wr_data_rom[ 3089]='h00000000;
    rd_cycle[ 3090] = 1'b1;  wr_cycle[ 3090] = 1'b0;  addr_rom[ 3090]='h00000074;  wr_data_rom[ 3090]='h00000000;
    rd_cycle[ 3091] = 1'b0;  wr_cycle[ 3091] = 1'b1;  addr_rom[ 3091]='h00000048;  wr_data_rom[ 3091]='h00000335;
    rd_cycle[ 3092] = 1'b1;  wr_cycle[ 3092] = 1'b0;  addr_rom[ 3092]='h000008d0;  wr_data_rom[ 3092]='h00000000;
    rd_cycle[ 3093] = 1'b1;  wr_cycle[ 3093] = 1'b0;  addr_rom[ 3093]='h00000404;  wr_data_rom[ 3093]='h00000000;
    rd_cycle[ 3094] = 1'b0;  wr_cycle[ 3094] = 1'b1;  addr_rom[ 3094]='h00000c48;  wr_data_rom[ 3094]='h000001bf;
    rd_cycle[ 3095] = 1'b0;  wr_cycle[ 3095] = 1'b1;  addr_rom[ 3095]='h000005f4;  wr_data_rom[ 3095]='h000000f7;
    rd_cycle[ 3096] = 1'b1;  wr_cycle[ 3096] = 1'b0;  addr_rom[ 3096]='h000008ac;  wr_data_rom[ 3096]='h00000000;
    rd_cycle[ 3097] = 1'b1;  wr_cycle[ 3097] = 1'b0;  addr_rom[ 3097]='h000006f0;  wr_data_rom[ 3097]='h00000000;
    rd_cycle[ 3098] = 1'b0;  wr_cycle[ 3098] = 1'b1;  addr_rom[ 3098]='h000006e0;  wr_data_rom[ 3098]='h00000917;
    rd_cycle[ 3099] = 1'b1;  wr_cycle[ 3099] = 1'b0;  addr_rom[ 3099]='h00000854;  wr_data_rom[ 3099]='h00000000;
    rd_cycle[ 3100] = 1'b1;  wr_cycle[ 3100] = 1'b0;  addr_rom[ 3100]='h00000b54;  wr_data_rom[ 3100]='h00000000;
    rd_cycle[ 3101] = 1'b1;  wr_cycle[ 3101] = 1'b0;  addr_rom[ 3101]='h00000f64;  wr_data_rom[ 3101]='h00000000;
    rd_cycle[ 3102] = 1'b1;  wr_cycle[ 3102] = 1'b0;  addr_rom[ 3102]='h00000c08;  wr_data_rom[ 3102]='h00000000;
    rd_cycle[ 3103] = 1'b0;  wr_cycle[ 3103] = 1'b1;  addr_rom[ 3103]='h00000dc8;  wr_data_rom[ 3103]='h00000051;
    rd_cycle[ 3104] = 1'b0;  wr_cycle[ 3104] = 1'b1;  addr_rom[ 3104]='h000001e8;  wr_data_rom[ 3104]='h00000f7f;
    rd_cycle[ 3105] = 1'b1;  wr_cycle[ 3105] = 1'b0;  addr_rom[ 3105]='h00000ac8;  wr_data_rom[ 3105]='h00000000;
    rd_cycle[ 3106] = 1'b0;  wr_cycle[ 3106] = 1'b1;  addr_rom[ 3106]='h00000664;  wr_data_rom[ 3106]='h00000e85;
    rd_cycle[ 3107] = 1'b0;  wr_cycle[ 3107] = 1'b1;  addr_rom[ 3107]='h00000738;  wr_data_rom[ 3107]='h0000048a;
    rd_cycle[ 3108] = 1'b1;  wr_cycle[ 3108] = 1'b0;  addr_rom[ 3108]='h000001d0;  wr_data_rom[ 3108]='h00000000;
    rd_cycle[ 3109] = 1'b0;  wr_cycle[ 3109] = 1'b1;  addr_rom[ 3109]='h00000d78;  wr_data_rom[ 3109]='h0000069a;
    rd_cycle[ 3110] = 1'b0;  wr_cycle[ 3110] = 1'b1;  addr_rom[ 3110]='h00000be4;  wr_data_rom[ 3110]='h00000f14;
    rd_cycle[ 3111] = 1'b1;  wr_cycle[ 3111] = 1'b0;  addr_rom[ 3111]='h000003b8;  wr_data_rom[ 3111]='h00000000;
    rd_cycle[ 3112] = 1'b1;  wr_cycle[ 3112] = 1'b0;  addr_rom[ 3112]='h0000042c;  wr_data_rom[ 3112]='h00000000;
    rd_cycle[ 3113] = 1'b0;  wr_cycle[ 3113] = 1'b1;  addr_rom[ 3113]='h00000ed8;  wr_data_rom[ 3113]='h00000cc8;
    rd_cycle[ 3114] = 1'b0;  wr_cycle[ 3114] = 1'b1;  addr_rom[ 3114]='h00000714;  wr_data_rom[ 3114]='h00000324;
    rd_cycle[ 3115] = 1'b0;  wr_cycle[ 3115] = 1'b1;  addr_rom[ 3115]='h000006d8;  wr_data_rom[ 3115]='h00000295;
    rd_cycle[ 3116] = 1'b0;  wr_cycle[ 3116] = 1'b1;  addr_rom[ 3116]='h00000d28;  wr_data_rom[ 3116]='h000005c4;
    rd_cycle[ 3117] = 1'b1;  wr_cycle[ 3117] = 1'b0;  addr_rom[ 3117]='h00000918;  wr_data_rom[ 3117]='h00000000;
    rd_cycle[ 3118] = 1'b0;  wr_cycle[ 3118] = 1'b1;  addr_rom[ 3118]='h000006e0;  wr_data_rom[ 3118]='h00000b8a;
    rd_cycle[ 3119] = 1'b1;  wr_cycle[ 3119] = 1'b0;  addr_rom[ 3119]='h000000a8;  wr_data_rom[ 3119]='h00000000;
    rd_cycle[ 3120] = 1'b1;  wr_cycle[ 3120] = 1'b0;  addr_rom[ 3120]='h00000264;  wr_data_rom[ 3120]='h00000000;
    rd_cycle[ 3121] = 1'b1;  wr_cycle[ 3121] = 1'b0;  addr_rom[ 3121]='h00000258;  wr_data_rom[ 3121]='h00000000;
    rd_cycle[ 3122] = 1'b0;  wr_cycle[ 3122] = 1'b1;  addr_rom[ 3122]='h00000adc;  wr_data_rom[ 3122]='h00000493;
    rd_cycle[ 3123] = 1'b1;  wr_cycle[ 3123] = 1'b0;  addr_rom[ 3123]='h000008c0;  wr_data_rom[ 3123]='h00000000;
    rd_cycle[ 3124] = 1'b1;  wr_cycle[ 3124] = 1'b0;  addr_rom[ 3124]='h00000b88;  wr_data_rom[ 3124]='h00000000;
    rd_cycle[ 3125] = 1'b0;  wr_cycle[ 3125] = 1'b1;  addr_rom[ 3125]='h00000d94;  wr_data_rom[ 3125]='h00000118;
    rd_cycle[ 3126] = 1'b1;  wr_cycle[ 3126] = 1'b0;  addr_rom[ 3126]='h00000da4;  wr_data_rom[ 3126]='h00000000;
    rd_cycle[ 3127] = 1'b1;  wr_cycle[ 3127] = 1'b0;  addr_rom[ 3127]='h00000ddc;  wr_data_rom[ 3127]='h00000000;
    rd_cycle[ 3128] = 1'b0;  wr_cycle[ 3128] = 1'b1;  addr_rom[ 3128]='h00000444;  wr_data_rom[ 3128]='h00000690;
    rd_cycle[ 3129] = 1'b1;  wr_cycle[ 3129] = 1'b0;  addr_rom[ 3129]='h00000590;  wr_data_rom[ 3129]='h00000000;
    rd_cycle[ 3130] = 1'b1;  wr_cycle[ 3130] = 1'b0;  addr_rom[ 3130]='h000000dc;  wr_data_rom[ 3130]='h00000000;
    rd_cycle[ 3131] = 1'b1;  wr_cycle[ 3131] = 1'b0;  addr_rom[ 3131]='h0000027c;  wr_data_rom[ 3131]='h00000000;
    rd_cycle[ 3132] = 1'b1;  wr_cycle[ 3132] = 1'b0;  addr_rom[ 3132]='h00000da0;  wr_data_rom[ 3132]='h00000000;
    rd_cycle[ 3133] = 1'b0;  wr_cycle[ 3133] = 1'b1;  addr_rom[ 3133]='h0000072c;  wr_data_rom[ 3133]='h0000016c;
    rd_cycle[ 3134] = 1'b1;  wr_cycle[ 3134] = 1'b0;  addr_rom[ 3134]='h00000d18;  wr_data_rom[ 3134]='h00000000;
    rd_cycle[ 3135] = 1'b1;  wr_cycle[ 3135] = 1'b0;  addr_rom[ 3135]='h000009b8;  wr_data_rom[ 3135]='h00000000;
    rd_cycle[ 3136] = 1'b0;  wr_cycle[ 3136] = 1'b1;  addr_rom[ 3136]='h00000ee0;  wr_data_rom[ 3136]='h000008a3;
    rd_cycle[ 3137] = 1'b1;  wr_cycle[ 3137] = 1'b0;  addr_rom[ 3137]='h00000578;  wr_data_rom[ 3137]='h00000000;
    rd_cycle[ 3138] = 1'b0;  wr_cycle[ 3138] = 1'b1;  addr_rom[ 3138]='h00000398;  wr_data_rom[ 3138]='h00000501;
    rd_cycle[ 3139] = 1'b0;  wr_cycle[ 3139] = 1'b1;  addr_rom[ 3139]='h000005b0;  wr_data_rom[ 3139]='h000006a1;
    rd_cycle[ 3140] = 1'b0;  wr_cycle[ 3140] = 1'b1;  addr_rom[ 3140]='h0000081c;  wr_data_rom[ 3140]='h00000187;
    rd_cycle[ 3141] = 1'b0;  wr_cycle[ 3141] = 1'b1;  addr_rom[ 3141]='h00000f40;  wr_data_rom[ 3141]='h00000e88;
    rd_cycle[ 3142] = 1'b1;  wr_cycle[ 3142] = 1'b0;  addr_rom[ 3142]='h000002b0;  wr_data_rom[ 3142]='h00000000;
    rd_cycle[ 3143] = 1'b0;  wr_cycle[ 3143] = 1'b1;  addr_rom[ 3143]='h000002b8;  wr_data_rom[ 3143]='h000008cf;
    rd_cycle[ 3144] = 1'b0;  wr_cycle[ 3144] = 1'b1;  addr_rom[ 3144]='h0000028c;  wr_data_rom[ 3144]='h00000e7a;
    rd_cycle[ 3145] = 1'b1;  wr_cycle[ 3145] = 1'b0;  addr_rom[ 3145]='h00000e08;  wr_data_rom[ 3145]='h00000000;
    rd_cycle[ 3146] = 1'b1;  wr_cycle[ 3146] = 1'b0;  addr_rom[ 3146]='h0000067c;  wr_data_rom[ 3146]='h00000000;
    rd_cycle[ 3147] = 1'b1;  wr_cycle[ 3147] = 1'b0;  addr_rom[ 3147]='h00000120;  wr_data_rom[ 3147]='h00000000;
    rd_cycle[ 3148] = 1'b1;  wr_cycle[ 3148] = 1'b0;  addr_rom[ 3148]='h00000c7c;  wr_data_rom[ 3148]='h00000000;
    rd_cycle[ 3149] = 1'b0;  wr_cycle[ 3149] = 1'b1;  addr_rom[ 3149]='h000009f0;  wr_data_rom[ 3149]='h00000932;
    rd_cycle[ 3150] = 1'b0;  wr_cycle[ 3150] = 1'b1;  addr_rom[ 3150]='h00000d34;  wr_data_rom[ 3150]='h00000c44;
    rd_cycle[ 3151] = 1'b0;  wr_cycle[ 3151] = 1'b1;  addr_rom[ 3151]='h00000e0c;  wr_data_rom[ 3151]='h0000011e;
    rd_cycle[ 3152] = 1'b0;  wr_cycle[ 3152] = 1'b1;  addr_rom[ 3152]='h00000e70;  wr_data_rom[ 3152]='h000003fb;
    rd_cycle[ 3153] = 1'b0;  wr_cycle[ 3153] = 1'b1;  addr_rom[ 3153]='h00000bfc;  wr_data_rom[ 3153]='h00000ef3;
    rd_cycle[ 3154] = 1'b0;  wr_cycle[ 3154] = 1'b1;  addr_rom[ 3154]='h000008d0;  wr_data_rom[ 3154]='h00000d99;
    rd_cycle[ 3155] = 1'b1;  wr_cycle[ 3155] = 1'b0;  addr_rom[ 3155]='h00000688;  wr_data_rom[ 3155]='h00000000;
    rd_cycle[ 3156] = 1'b0;  wr_cycle[ 3156] = 1'b1;  addr_rom[ 3156]='h00000a2c;  wr_data_rom[ 3156]='h0000030f;
    rd_cycle[ 3157] = 1'b1;  wr_cycle[ 3157] = 1'b0;  addr_rom[ 3157]='h00000204;  wr_data_rom[ 3157]='h00000000;
    rd_cycle[ 3158] = 1'b1;  wr_cycle[ 3158] = 1'b0;  addr_rom[ 3158]='h00000a00;  wr_data_rom[ 3158]='h00000000;
    rd_cycle[ 3159] = 1'b0;  wr_cycle[ 3159] = 1'b1;  addr_rom[ 3159]='h000001c8;  wr_data_rom[ 3159]='h000008c2;
    rd_cycle[ 3160] = 1'b0;  wr_cycle[ 3160] = 1'b1;  addr_rom[ 3160]='h00000c84;  wr_data_rom[ 3160]='h00000657;
    rd_cycle[ 3161] = 1'b1;  wr_cycle[ 3161] = 1'b0;  addr_rom[ 3161]='h00000828;  wr_data_rom[ 3161]='h00000000;
    rd_cycle[ 3162] = 1'b0;  wr_cycle[ 3162] = 1'b1;  addr_rom[ 3162]='h0000009c;  wr_data_rom[ 3162]='h00000e24;
    rd_cycle[ 3163] = 1'b1;  wr_cycle[ 3163] = 1'b0;  addr_rom[ 3163]='h00000d50;  wr_data_rom[ 3163]='h00000000;
    rd_cycle[ 3164] = 1'b0;  wr_cycle[ 3164] = 1'b1;  addr_rom[ 3164]='h0000034c;  wr_data_rom[ 3164]='h00000bf7;
    rd_cycle[ 3165] = 1'b0;  wr_cycle[ 3165] = 1'b1;  addr_rom[ 3165]='h00000150;  wr_data_rom[ 3165]='h00000411;
    rd_cycle[ 3166] = 1'b1;  wr_cycle[ 3166] = 1'b0;  addr_rom[ 3166]='h00000ea4;  wr_data_rom[ 3166]='h00000000;
    rd_cycle[ 3167] = 1'b0;  wr_cycle[ 3167] = 1'b1;  addr_rom[ 3167]='h00000748;  wr_data_rom[ 3167]='h000007d4;
    rd_cycle[ 3168] = 1'b0;  wr_cycle[ 3168] = 1'b1;  addr_rom[ 3168]='h00000148;  wr_data_rom[ 3168]='h00000e88;
    rd_cycle[ 3169] = 1'b0;  wr_cycle[ 3169] = 1'b1;  addr_rom[ 3169]='h00000d20;  wr_data_rom[ 3169]='h000001b5;
    rd_cycle[ 3170] = 1'b1;  wr_cycle[ 3170] = 1'b0;  addr_rom[ 3170]='h00000f74;  wr_data_rom[ 3170]='h00000000;
    rd_cycle[ 3171] = 1'b1;  wr_cycle[ 3171] = 1'b0;  addr_rom[ 3171]='h00000208;  wr_data_rom[ 3171]='h00000000;
    rd_cycle[ 3172] = 1'b0;  wr_cycle[ 3172] = 1'b1;  addr_rom[ 3172]='h00000910;  wr_data_rom[ 3172]='h00000d7f;
    rd_cycle[ 3173] = 1'b1;  wr_cycle[ 3173] = 1'b0;  addr_rom[ 3173]='h000008b0;  wr_data_rom[ 3173]='h00000000;
    rd_cycle[ 3174] = 1'b0;  wr_cycle[ 3174] = 1'b1;  addr_rom[ 3174]='h00000f08;  wr_data_rom[ 3174]='h0000012f;
    rd_cycle[ 3175] = 1'b1;  wr_cycle[ 3175] = 1'b0;  addr_rom[ 3175]='h00000e60;  wr_data_rom[ 3175]='h00000000;
    rd_cycle[ 3176] = 1'b0;  wr_cycle[ 3176] = 1'b1;  addr_rom[ 3176]='h000002dc;  wr_data_rom[ 3176]='h000002cf;
    rd_cycle[ 3177] = 1'b1;  wr_cycle[ 3177] = 1'b0;  addr_rom[ 3177]='h00000bf4;  wr_data_rom[ 3177]='h00000000;
    rd_cycle[ 3178] = 1'b1;  wr_cycle[ 3178] = 1'b0;  addr_rom[ 3178]='h00000410;  wr_data_rom[ 3178]='h00000000;
    rd_cycle[ 3179] = 1'b0;  wr_cycle[ 3179] = 1'b1;  addr_rom[ 3179]='h00000b2c;  wr_data_rom[ 3179]='h00000d93;
    rd_cycle[ 3180] = 1'b1;  wr_cycle[ 3180] = 1'b0;  addr_rom[ 3180]='h00000168;  wr_data_rom[ 3180]='h00000000;
    rd_cycle[ 3181] = 1'b0;  wr_cycle[ 3181] = 1'b1;  addr_rom[ 3181]='h000006d0;  wr_data_rom[ 3181]='h000000cc;
    rd_cycle[ 3182] = 1'b0;  wr_cycle[ 3182] = 1'b1;  addr_rom[ 3182]='h00000c2c;  wr_data_rom[ 3182]='h000002f3;
    rd_cycle[ 3183] = 1'b0;  wr_cycle[ 3183] = 1'b1;  addr_rom[ 3183]='h00000514;  wr_data_rom[ 3183]='h00000c33;
    rd_cycle[ 3184] = 1'b1;  wr_cycle[ 3184] = 1'b0;  addr_rom[ 3184]='h00000708;  wr_data_rom[ 3184]='h00000000;
    rd_cycle[ 3185] = 1'b1;  wr_cycle[ 3185] = 1'b0;  addr_rom[ 3185]='h00000ad0;  wr_data_rom[ 3185]='h00000000;
    rd_cycle[ 3186] = 1'b1;  wr_cycle[ 3186] = 1'b0;  addr_rom[ 3186]='h00000d2c;  wr_data_rom[ 3186]='h00000000;
    rd_cycle[ 3187] = 1'b1;  wr_cycle[ 3187] = 1'b0;  addr_rom[ 3187]='h00000334;  wr_data_rom[ 3187]='h00000000;
    rd_cycle[ 3188] = 1'b1;  wr_cycle[ 3188] = 1'b0;  addr_rom[ 3188]='h00000628;  wr_data_rom[ 3188]='h00000000;
    rd_cycle[ 3189] = 1'b0;  wr_cycle[ 3189] = 1'b1;  addr_rom[ 3189]='h00000f4c;  wr_data_rom[ 3189]='h0000040a;
    rd_cycle[ 3190] = 1'b0;  wr_cycle[ 3190] = 1'b1;  addr_rom[ 3190]='h000002b4;  wr_data_rom[ 3190]='h000007de;
    rd_cycle[ 3191] = 1'b1;  wr_cycle[ 3191] = 1'b0;  addr_rom[ 3191]='h0000060c;  wr_data_rom[ 3191]='h00000000;
    rd_cycle[ 3192] = 1'b0;  wr_cycle[ 3192] = 1'b1;  addr_rom[ 3192]='h00000684;  wr_data_rom[ 3192]='h000007f7;
    rd_cycle[ 3193] = 1'b0;  wr_cycle[ 3193] = 1'b1;  addr_rom[ 3193]='h00000590;  wr_data_rom[ 3193]='h00000540;
    rd_cycle[ 3194] = 1'b0;  wr_cycle[ 3194] = 1'b1;  addr_rom[ 3194]='h00000544;  wr_data_rom[ 3194]='h000002cc;
    rd_cycle[ 3195] = 1'b0;  wr_cycle[ 3195] = 1'b1;  addr_rom[ 3195]='h00000bdc;  wr_data_rom[ 3195]='h00000c40;
    rd_cycle[ 3196] = 1'b1;  wr_cycle[ 3196] = 1'b0;  addr_rom[ 3196]='h00000a20;  wr_data_rom[ 3196]='h00000000;
    rd_cycle[ 3197] = 1'b1;  wr_cycle[ 3197] = 1'b0;  addr_rom[ 3197]='h00000bdc;  wr_data_rom[ 3197]='h00000000;
    rd_cycle[ 3198] = 1'b0;  wr_cycle[ 3198] = 1'b1;  addr_rom[ 3198]='h0000030c;  wr_data_rom[ 3198]='h00000e3a;
    rd_cycle[ 3199] = 1'b0;  wr_cycle[ 3199] = 1'b1;  addr_rom[ 3199]='h00000828;  wr_data_rom[ 3199]='h00000541;
    rd_cycle[ 3200] = 1'b0;  wr_cycle[ 3200] = 1'b1;  addr_rom[ 3200]='h00000b20;  wr_data_rom[ 3200]='h00000219;
    rd_cycle[ 3201] = 1'b1;  wr_cycle[ 3201] = 1'b0;  addr_rom[ 3201]='h00000148;  wr_data_rom[ 3201]='h00000000;
    rd_cycle[ 3202] = 1'b1;  wr_cycle[ 3202] = 1'b0;  addr_rom[ 3202]='h000005a4;  wr_data_rom[ 3202]='h00000000;
    rd_cycle[ 3203] = 1'b0;  wr_cycle[ 3203] = 1'b1;  addr_rom[ 3203]='h000005bc;  wr_data_rom[ 3203]='h0000023a;
    rd_cycle[ 3204] = 1'b0;  wr_cycle[ 3204] = 1'b1;  addr_rom[ 3204]='h000006f4;  wr_data_rom[ 3204]='h00000568;
    rd_cycle[ 3205] = 1'b1;  wr_cycle[ 3205] = 1'b0;  addr_rom[ 3205]='h00000764;  wr_data_rom[ 3205]='h00000000;
    rd_cycle[ 3206] = 1'b0;  wr_cycle[ 3206] = 1'b1;  addr_rom[ 3206]='h00000b0c;  wr_data_rom[ 3206]='h00000a0c;
    rd_cycle[ 3207] = 1'b1;  wr_cycle[ 3207] = 1'b0;  addr_rom[ 3207]='h000001b4;  wr_data_rom[ 3207]='h00000000;
    rd_cycle[ 3208] = 1'b0;  wr_cycle[ 3208] = 1'b1;  addr_rom[ 3208]='h00000f10;  wr_data_rom[ 3208]='h00000b62;
    rd_cycle[ 3209] = 1'b1;  wr_cycle[ 3209] = 1'b0;  addr_rom[ 3209]='h00000494;  wr_data_rom[ 3209]='h00000000;
    rd_cycle[ 3210] = 1'b0;  wr_cycle[ 3210] = 1'b1;  addr_rom[ 3210]='h00000048;  wr_data_rom[ 3210]='h00000c3b;
    rd_cycle[ 3211] = 1'b0;  wr_cycle[ 3211] = 1'b1;  addr_rom[ 3211]='h00000124;  wr_data_rom[ 3211]='h000001a3;
    rd_cycle[ 3212] = 1'b0;  wr_cycle[ 3212] = 1'b1;  addr_rom[ 3212]='h000008b8;  wr_data_rom[ 3212]='h00000552;
    rd_cycle[ 3213] = 1'b1;  wr_cycle[ 3213] = 1'b0;  addr_rom[ 3213]='h00000d68;  wr_data_rom[ 3213]='h00000000;
    rd_cycle[ 3214] = 1'b1;  wr_cycle[ 3214] = 1'b0;  addr_rom[ 3214]='h000001ac;  wr_data_rom[ 3214]='h00000000;
    rd_cycle[ 3215] = 1'b1;  wr_cycle[ 3215] = 1'b0;  addr_rom[ 3215]='h000003c0;  wr_data_rom[ 3215]='h00000000;
    rd_cycle[ 3216] = 1'b0;  wr_cycle[ 3216] = 1'b1;  addr_rom[ 3216]='h000003bc;  wr_data_rom[ 3216]='h00000080;
    rd_cycle[ 3217] = 1'b0;  wr_cycle[ 3217] = 1'b1;  addr_rom[ 3217]='h000006b8;  wr_data_rom[ 3217]='h00000f1d;
    rd_cycle[ 3218] = 1'b0;  wr_cycle[ 3218] = 1'b1;  addr_rom[ 3218]='h0000047c;  wr_data_rom[ 3218]='h000003c6;
    rd_cycle[ 3219] = 1'b0;  wr_cycle[ 3219] = 1'b1;  addr_rom[ 3219]='h00000478;  wr_data_rom[ 3219]='h00000f90;
    rd_cycle[ 3220] = 1'b1;  wr_cycle[ 3220] = 1'b0;  addr_rom[ 3220]='h00000b04;  wr_data_rom[ 3220]='h00000000;
    rd_cycle[ 3221] = 1'b0;  wr_cycle[ 3221] = 1'b1;  addr_rom[ 3221]='h0000020c;  wr_data_rom[ 3221]='h000007c8;
    rd_cycle[ 3222] = 1'b0;  wr_cycle[ 3222] = 1'b1;  addr_rom[ 3222]='h00000d7c;  wr_data_rom[ 3222]='h000000e9;
    rd_cycle[ 3223] = 1'b1;  wr_cycle[ 3223] = 1'b0;  addr_rom[ 3223]='h0000072c;  wr_data_rom[ 3223]='h00000000;
    rd_cycle[ 3224] = 1'b1;  wr_cycle[ 3224] = 1'b0;  addr_rom[ 3224]='h00000708;  wr_data_rom[ 3224]='h00000000;
    rd_cycle[ 3225] = 1'b0;  wr_cycle[ 3225] = 1'b1;  addr_rom[ 3225]='h00000188;  wr_data_rom[ 3225]='h00000d4a;
    rd_cycle[ 3226] = 1'b0;  wr_cycle[ 3226] = 1'b1;  addr_rom[ 3226]='h00000700;  wr_data_rom[ 3226]='h00000b4e;
    rd_cycle[ 3227] = 1'b1;  wr_cycle[ 3227] = 1'b0;  addr_rom[ 3227]='h000001c0;  wr_data_rom[ 3227]='h00000000;
    rd_cycle[ 3228] = 1'b1;  wr_cycle[ 3228] = 1'b0;  addr_rom[ 3228]='h00000828;  wr_data_rom[ 3228]='h00000000;
    rd_cycle[ 3229] = 1'b0;  wr_cycle[ 3229] = 1'b1;  addr_rom[ 3229]='h00000f44;  wr_data_rom[ 3229]='h00000b7a;
    rd_cycle[ 3230] = 1'b0;  wr_cycle[ 3230] = 1'b1;  addr_rom[ 3230]='h0000023c;  wr_data_rom[ 3230]='h00000d23;
    rd_cycle[ 3231] = 1'b0;  wr_cycle[ 3231] = 1'b1;  addr_rom[ 3231]='h00000e2c;  wr_data_rom[ 3231]='h000009b9;
    rd_cycle[ 3232] = 1'b1;  wr_cycle[ 3232] = 1'b0;  addr_rom[ 3232]='h00000178;  wr_data_rom[ 3232]='h00000000;
    rd_cycle[ 3233] = 1'b0;  wr_cycle[ 3233] = 1'b1;  addr_rom[ 3233]='h000001d8;  wr_data_rom[ 3233]='h000007fd;
    rd_cycle[ 3234] = 1'b1;  wr_cycle[ 3234] = 1'b0;  addr_rom[ 3234]='h00000a68;  wr_data_rom[ 3234]='h00000000;
    rd_cycle[ 3235] = 1'b1;  wr_cycle[ 3235] = 1'b0;  addr_rom[ 3235]='h00000f90;  wr_data_rom[ 3235]='h00000000;
    rd_cycle[ 3236] = 1'b1;  wr_cycle[ 3236] = 1'b0;  addr_rom[ 3236]='h00000324;  wr_data_rom[ 3236]='h00000000;
    rd_cycle[ 3237] = 1'b0;  wr_cycle[ 3237] = 1'b1;  addr_rom[ 3237]='h000009b8;  wr_data_rom[ 3237]='h00000a50;
    rd_cycle[ 3238] = 1'b0;  wr_cycle[ 3238] = 1'b1;  addr_rom[ 3238]='h000009a8;  wr_data_rom[ 3238]='h00000233;
    rd_cycle[ 3239] = 1'b1;  wr_cycle[ 3239] = 1'b0;  addr_rom[ 3239]='h00000934;  wr_data_rom[ 3239]='h00000000;
    rd_cycle[ 3240] = 1'b1;  wr_cycle[ 3240] = 1'b0;  addr_rom[ 3240]='h00000af0;  wr_data_rom[ 3240]='h00000000;
    rd_cycle[ 3241] = 1'b1;  wr_cycle[ 3241] = 1'b0;  addr_rom[ 3241]='h0000020c;  wr_data_rom[ 3241]='h00000000;
    rd_cycle[ 3242] = 1'b1;  wr_cycle[ 3242] = 1'b0;  addr_rom[ 3242]='h00000128;  wr_data_rom[ 3242]='h00000000;
    rd_cycle[ 3243] = 1'b1;  wr_cycle[ 3243] = 1'b0;  addr_rom[ 3243]='h00000920;  wr_data_rom[ 3243]='h00000000;
    rd_cycle[ 3244] = 1'b1;  wr_cycle[ 3244] = 1'b0;  addr_rom[ 3244]='h000002c0;  wr_data_rom[ 3244]='h00000000;
    rd_cycle[ 3245] = 1'b0;  wr_cycle[ 3245] = 1'b1;  addr_rom[ 3245]='h00000db0;  wr_data_rom[ 3245]='h000002dc;
    rd_cycle[ 3246] = 1'b0;  wr_cycle[ 3246] = 1'b1;  addr_rom[ 3246]='h00000088;  wr_data_rom[ 3246]='h00000a79;
    rd_cycle[ 3247] = 1'b1;  wr_cycle[ 3247] = 1'b0;  addr_rom[ 3247]='h00000338;  wr_data_rom[ 3247]='h00000000;
    rd_cycle[ 3248] = 1'b1;  wr_cycle[ 3248] = 1'b0;  addr_rom[ 3248]='h00000b28;  wr_data_rom[ 3248]='h00000000;
    rd_cycle[ 3249] = 1'b1;  wr_cycle[ 3249] = 1'b0;  addr_rom[ 3249]='h00000634;  wr_data_rom[ 3249]='h00000000;
    rd_cycle[ 3250] = 1'b1;  wr_cycle[ 3250] = 1'b0;  addr_rom[ 3250]='h00000598;  wr_data_rom[ 3250]='h00000000;
    rd_cycle[ 3251] = 1'b0;  wr_cycle[ 3251] = 1'b1;  addr_rom[ 3251]='h0000080c;  wr_data_rom[ 3251]='h00000969;
    rd_cycle[ 3252] = 1'b0;  wr_cycle[ 3252] = 1'b1;  addr_rom[ 3252]='h00000944;  wr_data_rom[ 3252]='h00000dd3;
    rd_cycle[ 3253] = 1'b0;  wr_cycle[ 3253] = 1'b1;  addr_rom[ 3253]='h00000258;  wr_data_rom[ 3253]='h00000670;
    rd_cycle[ 3254] = 1'b0;  wr_cycle[ 3254] = 1'b1;  addr_rom[ 3254]='h00000b24;  wr_data_rom[ 3254]='h00000652;
    rd_cycle[ 3255] = 1'b0;  wr_cycle[ 3255] = 1'b1;  addr_rom[ 3255]='h00000cc0;  wr_data_rom[ 3255]='h000008aa;
    rd_cycle[ 3256] = 1'b1;  wr_cycle[ 3256] = 1'b0;  addr_rom[ 3256]='h00000c7c;  wr_data_rom[ 3256]='h00000000;
    rd_cycle[ 3257] = 1'b0;  wr_cycle[ 3257] = 1'b1;  addr_rom[ 3257]='h00000714;  wr_data_rom[ 3257]='h00000cad;
    rd_cycle[ 3258] = 1'b1;  wr_cycle[ 3258] = 1'b0;  addr_rom[ 3258]='h00000b64;  wr_data_rom[ 3258]='h00000000;
    rd_cycle[ 3259] = 1'b0;  wr_cycle[ 3259] = 1'b1;  addr_rom[ 3259]='h00000738;  wr_data_rom[ 3259]='h00000af2;
    rd_cycle[ 3260] = 1'b0;  wr_cycle[ 3260] = 1'b1;  addr_rom[ 3260]='h0000073c;  wr_data_rom[ 3260]='h00000414;
    rd_cycle[ 3261] = 1'b1;  wr_cycle[ 3261] = 1'b0;  addr_rom[ 3261]='h00000f14;  wr_data_rom[ 3261]='h00000000;
    rd_cycle[ 3262] = 1'b0;  wr_cycle[ 3262] = 1'b1;  addr_rom[ 3262]='h00000d80;  wr_data_rom[ 3262]='h00000b0b;
    rd_cycle[ 3263] = 1'b0;  wr_cycle[ 3263] = 1'b1;  addr_rom[ 3263]='h00000f2c;  wr_data_rom[ 3263]='h0000056a;
    rd_cycle[ 3264] = 1'b0;  wr_cycle[ 3264] = 1'b1;  addr_rom[ 3264]='h00000514;  wr_data_rom[ 3264]='h00000d8e;
    rd_cycle[ 3265] = 1'b1;  wr_cycle[ 3265] = 1'b0;  addr_rom[ 3265]='h000000e4;  wr_data_rom[ 3265]='h00000000;
    rd_cycle[ 3266] = 1'b0;  wr_cycle[ 3266] = 1'b1;  addr_rom[ 3266]='h00000bfc;  wr_data_rom[ 3266]='h00000a99;
    rd_cycle[ 3267] = 1'b0;  wr_cycle[ 3267] = 1'b1;  addr_rom[ 3267]='h000000d0;  wr_data_rom[ 3267]='h00000607;
    rd_cycle[ 3268] = 1'b1;  wr_cycle[ 3268] = 1'b0;  addr_rom[ 3268]='h000003a8;  wr_data_rom[ 3268]='h00000000;
    rd_cycle[ 3269] = 1'b0;  wr_cycle[ 3269] = 1'b1;  addr_rom[ 3269]='h000006bc;  wr_data_rom[ 3269]='h000007f0;
    rd_cycle[ 3270] = 1'b1;  wr_cycle[ 3270] = 1'b0;  addr_rom[ 3270]='h00000ac4;  wr_data_rom[ 3270]='h00000000;
    rd_cycle[ 3271] = 1'b1;  wr_cycle[ 3271] = 1'b0;  addr_rom[ 3271]='h0000086c;  wr_data_rom[ 3271]='h00000000;
    rd_cycle[ 3272] = 1'b1;  wr_cycle[ 3272] = 1'b0;  addr_rom[ 3272]='h0000089c;  wr_data_rom[ 3272]='h00000000;
    rd_cycle[ 3273] = 1'b1;  wr_cycle[ 3273] = 1'b0;  addr_rom[ 3273]='h00000ec4;  wr_data_rom[ 3273]='h00000000;
    rd_cycle[ 3274] = 1'b1;  wr_cycle[ 3274] = 1'b0;  addr_rom[ 3274]='h00000c1c;  wr_data_rom[ 3274]='h00000000;
    rd_cycle[ 3275] = 1'b1;  wr_cycle[ 3275] = 1'b0;  addr_rom[ 3275]='h00000b34;  wr_data_rom[ 3275]='h00000000;
    rd_cycle[ 3276] = 1'b0;  wr_cycle[ 3276] = 1'b1;  addr_rom[ 3276]='h00000d6c;  wr_data_rom[ 3276]='h00000a57;
    rd_cycle[ 3277] = 1'b1;  wr_cycle[ 3277] = 1'b0;  addr_rom[ 3277]='h000009f8;  wr_data_rom[ 3277]='h00000000;
    rd_cycle[ 3278] = 1'b0;  wr_cycle[ 3278] = 1'b1;  addr_rom[ 3278]='h00000630;  wr_data_rom[ 3278]='h00000f93;
    rd_cycle[ 3279] = 1'b0;  wr_cycle[ 3279] = 1'b1;  addr_rom[ 3279]='h000000c4;  wr_data_rom[ 3279]='h000000ba;
    rd_cycle[ 3280] = 1'b1;  wr_cycle[ 3280] = 1'b0;  addr_rom[ 3280]='h00000558;  wr_data_rom[ 3280]='h00000000;
    rd_cycle[ 3281] = 1'b0;  wr_cycle[ 3281] = 1'b1;  addr_rom[ 3281]='h000001e8;  wr_data_rom[ 3281]='h00000a1e;
    rd_cycle[ 3282] = 1'b0;  wr_cycle[ 3282] = 1'b1;  addr_rom[ 3282]='h00000344;  wr_data_rom[ 3282]='h0000027e;
    rd_cycle[ 3283] = 1'b0;  wr_cycle[ 3283] = 1'b1;  addr_rom[ 3283]='h00000bb4;  wr_data_rom[ 3283]='h00000886;
    rd_cycle[ 3284] = 1'b1;  wr_cycle[ 3284] = 1'b0;  addr_rom[ 3284]='h00000ec0;  wr_data_rom[ 3284]='h00000000;
    rd_cycle[ 3285] = 1'b1;  wr_cycle[ 3285] = 1'b0;  addr_rom[ 3285]='h00000c74;  wr_data_rom[ 3285]='h00000000;
    rd_cycle[ 3286] = 1'b1;  wr_cycle[ 3286] = 1'b0;  addr_rom[ 3286]='h000009b0;  wr_data_rom[ 3286]='h00000000;
    rd_cycle[ 3287] = 1'b0;  wr_cycle[ 3287] = 1'b1;  addr_rom[ 3287]='h00000c98;  wr_data_rom[ 3287]='h0000035b;
    rd_cycle[ 3288] = 1'b0;  wr_cycle[ 3288] = 1'b1;  addr_rom[ 3288]='h00000ad0;  wr_data_rom[ 3288]='h000005d0;
    rd_cycle[ 3289] = 1'b0;  wr_cycle[ 3289] = 1'b1;  addr_rom[ 3289]='h00000880;  wr_data_rom[ 3289]='h00000786;
    rd_cycle[ 3290] = 1'b1;  wr_cycle[ 3290] = 1'b0;  addr_rom[ 3290]='h000005b0;  wr_data_rom[ 3290]='h00000000;
    rd_cycle[ 3291] = 1'b1;  wr_cycle[ 3291] = 1'b0;  addr_rom[ 3291]='h00000d4c;  wr_data_rom[ 3291]='h00000000;
    rd_cycle[ 3292] = 1'b0;  wr_cycle[ 3292] = 1'b1;  addr_rom[ 3292]='h00000200;  wr_data_rom[ 3292]='h00000884;
    rd_cycle[ 3293] = 1'b0;  wr_cycle[ 3293] = 1'b1;  addr_rom[ 3293]='h0000011c;  wr_data_rom[ 3293]='h00000af3;
    rd_cycle[ 3294] = 1'b0;  wr_cycle[ 3294] = 1'b1;  addr_rom[ 3294]='h000004e4;  wr_data_rom[ 3294]='h00000243;
    rd_cycle[ 3295] = 1'b0;  wr_cycle[ 3295] = 1'b1;  addr_rom[ 3295]='h000001a8;  wr_data_rom[ 3295]='h00000203;
    rd_cycle[ 3296] = 1'b1;  wr_cycle[ 3296] = 1'b0;  addr_rom[ 3296]='h00000820;  wr_data_rom[ 3296]='h00000000;
    rd_cycle[ 3297] = 1'b1;  wr_cycle[ 3297] = 1'b0;  addr_rom[ 3297]='h00000930;  wr_data_rom[ 3297]='h00000000;
    rd_cycle[ 3298] = 1'b1;  wr_cycle[ 3298] = 1'b0;  addr_rom[ 3298]='h00000f5c;  wr_data_rom[ 3298]='h00000000;
    rd_cycle[ 3299] = 1'b1;  wr_cycle[ 3299] = 1'b0;  addr_rom[ 3299]='h00000b88;  wr_data_rom[ 3299]='h00000000;
    rd_cycle[ 3300] = 1'b0;  wr_cycle[ 3300] = 1'b1;  addr_rom[ 3300]='h00000f64;  wr_data_rom[ 3300]='h00000a16;
    rd_cycle[ 3301] = 1'b1;  wr_cycle[ 3301] = 1'b0;  addr_rom[ 3301]='h00000d48;  wr_data_rom[ 3301]='h00000000;
    rd_cycle[ 3302] = 1'b0;  wr_cycle[ 3302] = 1'b1;  addr_rom[ 3302]='h00000a8c;  wr_data_rom[ 3302]='h00000f6b;
    rd_cycle[ 3303] = 1'b1;  wr_cycle[ 3303] = 1'b0;  addr_rom[ 3303]='h000001c4;  wr_data_rom[ 3303]='h00000000;
    rd_cycle[ 3304] = 1'b1;  wr_cycle[ 3304] = 1'b0;  addr_rom[ 3304]='h00000f44;  wr_data_rom[ 3304]='h00000000;
    rd_cycle[ 3305] = 1'b1;  wr_cycle[ 3305] = 1'b0;  addr_rom[ 3305]='h00000474;  wr_data_rom[ 3305]='h00000000;
    rd_cycle[ 3306] = 1'b0;  wr_cycle[ 3306] = 1'b1;  addr_rom[ 3306]='h00000e24;  wr_data_rom[ 3306]='h00000686;
    rd_cycle[ 3307] = 1'b0;  wr_cycle[ 3307] = 1'b1;  addr_rom[ 3307]='h00000888;  wr_data_rom[ 3307]='h00000e65;
    rd_cycle[ 3308] = 1'b1;  wr_cycle[ 3308] = 1'b0;  addr_rom[ 3308]='h00000cc8;  wr_data_rom[ 3308]='h00000000;
    rd_cycle[ 3309] = 1'b0;  wr_cycle[ 3309] = 1'b1;  addr_rom[ 3309]='h0000054c;  wr_data_rom[ 3309]='h000005c6;
    rd_cycle[ 3310] = 1'b0;  wr_cycle[ 3310] = 1'b1;  addr_rom[ 3310]='h00000b94;  wr_data_rom[ 3310]='h0000000f;
    rd_cycle[ 3311] = 1'b0;  wr_cycle[ 3311] = 1'b1;  addr_rom[ 3311]='h00000808;  wr_data_rom[ 3311]='h00000b0c;
    rd_cycle[ 3312] = 1'b1;  wr_cycle[ 3312] = 1'b0;  addr_rom[ 3312]='h00000558;  wr_data_rom[ 3312]='h00000000;
    rd_cycle[ 3313] = 1'b1;  wr_cycle[ 3313] = 1'b0;  addr_rom[ 3313]='h00000824;  wr_data_rom[ 3313]='h00000000;
    rd_cycle[ 3314] = 1'b0;  wr_cycle[ 3314] = 1'b1;  addr_rom[ 3314]='h00000f38;  wr_data_rom[ 3314]='h0000062c;
    rd_cycle[ 3315] = 1'b1;  wr_cycle[ 3315] = 1'b0;  addr_rom[ 3315]='h0000095c;  wr_data_rom[ 3315]='h00000000;
    rd_cycle[ 3316] = 1'b0;  wr_cycle[ 3316] = 1'b1;  addr_rom[ 3316]='h00000bd0;  wr_data_rom[ 3316]='h00000d51;
    rd_cycle[ 3317] = 1'b1;  wr_cycle[ 3317] = 1'b0;  addr_rom[ 3317]='h00000e4c;  wr_data_rom[ 3317]='h00000000;
    rd_cycle[ 3318] = 1'b0;  wr_cycle[ 3318] = 1'b1;  addr_rom[ 3318]='h000004e0;  wr_data_rom[ 3318]='h000008fd;
    rd_cycle[ 3319] = 1'b0;  wr_cycle[ 3319] = 1'b1;  addr_rom[ 3319]='h00000df8;  wr_data_rom[ 3319]='h00000ca7;
    rd_cycle[ 3320] = 1'b0;  wr_cycle[ 3320] = 1'b1;  addr_rom[ 3320]='h00000e28;  wr_data_rom[ 3320]='h000008e5;
    rd_cycle[ 3321] = 1'b1;  wr_cycle[ 3321] = 1'b0;  addr_rom[ 3321]='h00000df4;  wr_data_rom[ 3321]='h00000000;
    rd_cycle[ 3322] = 1'b0;  wr_cycle[ 3322] = 1'b1;  addr_rom[ 3322]='h00000628;  wr_data_rom[ 3322]='h0000021f;
    rd_cycle[ 3323] = 1'b1;  wr_cycle[ 3323] = 1'b0;  addr_rom[ 3323]='h00000bac;  wr_data_rom[ 3323]='h00000000;
    rd_cycle[ 3324] = 1'b1;  wr_cycle[ 3324] = 1'b0;  addr_rom[ 3324]='h00000580;  wr_data_rom[ 3324]='h00000000;
    rd_cycle[ 3325] = 1'b0;  wr_cycle[ 3325] = 1'b1;  addr_rom[ 3325]='h00000798;  wr_data_rom[ 3325]='h00000e7c;
    rd_cycle[ 3326] = 1'b1;  wr_cycle[ 3326] = 1'b0;  addr_rom[ 3326]='h0000095c;  wr_data_rom[ 3326]='h00000000;
    rd_cycle[ 3327] = 1'b1;  wr_cycle[ 3327] = 1'b0;  addr_rom[ 3327]='h0000086c;  wr_data_rom[ 3327]='h00000000;
    rd_cycle[ 3328] = 1'b0;  wr_cycle[ 3328] = 1'b1;  addr_rom[ 3328]='h0000076c;  wr_data_rom[ 3328]='h00000c25;
    rd_cycle[ 3329] = 1'b1;  wr_cycle[ 3329] = 1'b0;  addr_rom[ 3329]='h000006ec;  wr_data_rom[ 3329]='h00000000;
    rd_cycle[ 3330] = 1'b1;  wr_cycle[ 3330] = 1'b0;  addr_rom[ 3330]='h00000c54;  wr_data_rom[ 3330]='h00000000;
    rd_cycle[ 3331] = 1'b1;  wr_cycle[ 3331] = 1'b0;  addr_rom[ 3331]='h000004e0;  wr_data_rom[ 3331]='h00000000;
    rd_cycle[ 3332] = 1'b1;  wr_cycle[ 3332] = 1'b0;  addr_rom[ 3332]='h00000910;  wr_data_rom[ 3332]='h00000000;
    rd_cycle[ 3333] = 1'b0;  wr_cycle[ 3333] = 1'b1;  addr_rom[ 3333]='h00000c50;  wr_data_rom[ 3333]='h000004e5;
    rd_cycle[ 3334] = 1'b1;  wr_cycle[ 3334] = 1'b0;  addr_rom[ 3334]='h00000670;  wr_data_rom[ 3334]='h00000000;
    rd_cycle[ 3335] = 1'b1;  wr_cycle[ 3335] = 1'b0;  addr_rom[ 3335]='h00000a90;  wr_data_rom[ 3335]='h00000000;
    rd_cycle[ 3336] = 1'b0;  wr_cycle[ 3336] = 1'b1;  addr_rom[ 3336]='h00000930;  wr_data_rom[ 3336]='h00000250;
    rd_cycle[ 3337] = 1'b0;  wr_cycle[ 3337] = 1'b1;  addr_rom[ 3337]='h0000056c;  wr_data_rom[ 3337]='h000006a0;
    rd_cycle[ 3338] = 1'b1;  wr_cycle[ 3338] = 1'b0;  addr_rom[ 3338]='h00000744;  wr_data_rom[ 3338]='h00000000;
    rd_cycle[ 3339] = 1'b0;  wr_cycle[ 3339] = 1'b1;  addr_rom[ 3339]='h00000530;  wr_data_rom[ 3339]='h000002fa;
    rd_cycle[ 3340] = 1'b1;  wr_cycle[ 3340] = 1'b0;  addr_rom[ 3340]='h00000e28;  wr_data_rom[ 3340]='h00000000;
    rd_cycle[ 3341] = 1'b1;  wr_cycle[ 3341] = 1'b0;  addr_rom[ 3341]='h00000ee4;  wr_data_rom[ 3341]='h00000000;
    rd_cycle[ 3342] = 1'b0;  wr_cycle[ 3342] = 1'b1;  addr_rom[ 3342]='h00000c24;  wr_data_rom[ 3342]='h00000579;
    rd_cycle[ 3343] = 1'b1;  wr_cycle[ 3343] = 1'b0;  addr_rom[ 3343]='h00000990;  wr_data_rom[ 3343]='h00000000;
    rd_cycle[ 3344] = 1'b1;  wr_cycle[ 3344] = 1'b0;  addr_rom[ 3344]='h00000cc0;  wr_data_rom[ 3344]='h00000000;
    rd_cycle[ 3345] = 1'b0;  wr_cycle[ 3345] = 1'b1;  addr_rom[ 3345]='h0000060c;  wr_data_rom[ 3345]='h00000477;
    rd_cycle[ 3346] = 1'b1;  wr_cycle[ 3346] = 1'b0;  addr_rom[ 3346]='h000008a8;  wr_data_rom[ 3346]='h00000000;
    rd_cycle[ 3347] = 1'b0;  wr_cycle[ 3347] = 1'b1;  addr_rom[ 3347]='h0000057c;  wr_data_rom[ 3347]='h00000e1b;
    rd_cycle[ 3348] = 1'b0;  wr_cycle[ 3348] = 1'b1;  addr_rom[ 3348]='h000006fc;  wr_data_rom[ 3348]='h000000a1;
    rd_cycle[ 3349] = 1'b0;  wr_cycle[ 3349] = 1'b1;  addr_rom[ 3349]='h00000848;  wr_data_rom[ 3349]='h00000d3f;
    rd_cycle[ 3350] = 1'b0;  wr_cycle[ 3350] = 1'b1;  addr_rom[ 3350]='h0000022c;  wr_data_rom[ 3350]='h00000ef3;
    rd_cycle[ 3351] = 1'b1;  wr_cycle[ 3351] = 1'b0;  addr_rom[ 3351]='h00000c94;  wr_data_rom[ 3351]='h00000000;
    rd_cycle[ 3352] = 1'b0;  wr_cycle[ 3352] = 1'b1;  addr_rom[ 3352]='h0000058c;  wr_data_rom[ 3352]='h00000287;
    rd_cycle[ 3353] = 1'b1;  wr_cycle[ 3353] = 1'b0;  addr_rom[ 3353]='h00000954;  wr_data_rom[ 3353]='h00000000;
    rd_cycle[ 3354] = 1'b0;  wr_cycle[ 3354] = 1'b1;  addr_rom[ 3354]='h00000410;  wr_data_rom[ 3354]='h000000d9;
    rd_cycle[ 3355] = 1'b1;  wr_cycle[ 3355] = 1'b0;  addr_rom[ 3355]='h00000680;  wr_data_rom[ 3355]='h00000000;
    rd_cycle[ 3356] = 1'b1;  wr_cycle[ 3356] = 1'b0;  addr_rom[ 3356]='h000004ac;  wr_data_rom[ 3356]='h00000000;
    rd_cycle[ 3357] = 1'b0;  wr_cycle[ 3357] = 1'b1;  addr_rom[ 3357]='h000004dc;  wr_data_rom[ 3357]='h000002f0;
    rd_cycle[ 3358] = 1'b0;  wr_cycle[ 3358] = 1'b1;  addr_rom[ 3358]='h00000c90;  wr_data_rom[ 3358]='h00000eec;
    rd_cycle[ 3359] = 1'b0;  wr_cycle[ 3359] = 1'b1;  addr_rom[ 3359]='h000007f8;  wr_data_rom[ 3359]='h00000ad9;
    rd_cycle[ 3360] = 1'b1;  wr_cycle[ 3360] = 1'b0;  addr_rom[ 3360]='h00000b4c;  wr_data_rom[ 3360]='h00000000;
    rd_cycle[ 3361] = 1'b1;  wr_cycle[ 3361] = 1'b0;  addr_rom[ 3361]='h00000a08;  wr_data_rom[ 3361]='h00000000;
    rd_cycle[ 3362] = 1'b1;  wr_cycle[ 3362] = 1'b0;  addr_rom[ 3362]='h00000e04;  wr_data_rom[ 3362]='h00000000;
    rd_cycle[ 3363] = 1'b1;  wr_cycle[ 3363] = 1'b0;  addr_rom[ 3363]='h00000d64;  wr_data_rom[ 3363]='h00000000;
    rd_cycle[ 3364] = 1'b0;  wr_cycle[ 3364] = 1'b1;  addr_rom[ 3364]='h0000016c;  wr_data_rom[ 3364]='h00000c74;
    rd_cycle[ 3365] = 1'b0;  wr_cycle[ 3365] = 1'b1;  addr_rom[ 3365]='h00000be4;  wr_data_rom[ 3365]='h0000003e;
    rd_cycle[ 3366] = 1'b1;  wr_cycle[ 3366] = 1'b0;  addr_rom[ 3366]='h00000704;  wr_data_rom[ 3366]='h00000000;
    rd_cycle[ 3367] = 1'b1;  wr_cycle[ 3367] = 1'b0;  addr_rom[ 3367]='h00000ef0;  wr_data_rom[ 3367]='h00000000;
    rd_cycle[ 3368] = 1'b0;  wr_cycle[ 3368] = 1'b1;  addr_rom[ 3368]='h000009f4;  wr_data_rom[ 3368]='h0000038b;
    rd_cycle[ 3369] = 1'b0;  wr_cycle[ 3369] = 1'b1;  addr_rom[ 3369]='h00000678;  wr_data_rom[ 3369]='h00000bc2;
    rd_cycle[ 3370] = 1'b1;  wr_cycle[ 3370] = 1'b0;  addr_rom[ 3370]='h00000b88;  wr_data_rom[ 3370]='h00000000;
    rd_cycle[ 3371] = 1'b1;  wr_cycle[ 3371] = 1'b0;  addr_rom[ 3371]='h00000b30;  wr_data_rom[ 3371]='h00000000;
    rd_cycle[ 3372] = 1'b1;  wr_cycle[ 3372] = 1'b0;  addr_rom[ 3372]='h00000624;  wr_data_rom[ 3372]='h00000000;
    rd_cycle[ 3373] = 1'b1;  wr_cycle[ 3373] = 1'b0;  addr_rom[ 3373]='h00000b04;  wr_data_rom[ 3373]='h00000000;
    rd_cycle[ 3374] = 1'b1;  wr_cycle[ 3374] = 1'b0;  addr_rom[ 3374]='h00000cec;  wr_data_rom[ 3374]='h00000000;
    rd_cycle[ 3375] = 1'b0;  wr_cycle[ 3375] = 1'b1;  addr_rom[ 3375]='h00000ce8;  wr_data_rom[ 3375]='h00000926;
    rd_cycle[ 3376] = 1'b0;  wr_cycle[ 3376] = 1'b1;  addr_rom[ 3376]='h000002b8;  wr_data_rom[ 3376]='h00000bd3;
    rd_cycle[ 3377] = 1'b0;  wr_cycle[ 3377] = 1'b1;  addr_rom[ 3377]='h000001d8;  wr_data_rom[ 3377]='h0000028c;
    rd_cycle[ 3378] = 1'b0;  wr_cycle[ 3378] = 1'b1;  addr_rom[ 3378]='h00000a3c;  wr_data_rom[ 3378]='h00000b87;
    rd_cycle[ 3379] = 1'b1;  wr_cycle[ 3379] = 1'b0;  addr_rom[ 3379]='h00000ce4;  wr_data_rom[ 3379]='h00000000;
    rd_cycle[ 3380] = 1'b1;  wr_cycle[ 3380] = 1'b0;  addr_rom[ 3380]='h00000a1c;  wr_data_rom[ 3380]='h00000000;
    rd_cycle[ 3381] = 1'b1;  wr_cycle[ 3381] = 1'b0;  addr_rom[ 3381]='h00000a70;  wr_data_rom[ 3381]='h00000000;
    rd_cycle[ 3382] = 1'b0;  wr_cycle[ 3382] = 1'b1;  addr_rom[ 3382]='h00000704;  wr_data_rom[ 3382]='h00000197;
    rd_cycle[ 3383] = 1'b1;  wr_cycle[ 3383] = 1'b0;  addr_rom[ 3383]='h00000da4;  wr_data_rom[ 3383]='h00000000;
    rd_cycle[ 3384] = 1'b1;  wr_cycle[ 3384] = 1'b0;  addr_rom[ 3384]='h00000a60;  wr_data_rom[ 3384]='h00000000;
    rd_cycle[ 3385] = 1'b0;  wr_cycle[ 3385] = 1'b1;  addr_rom[ 3385]='h00000a68;  wr_data_rom[ 3385]='h0000071f;
    rd_cycle[ 3386] = 1'b1;  wr_cycle[ 3386] = 1'b0;  addr_rom[ 3386]='h0000093c;  wr_data_rom[ 3386]='h00000000;
    rd_cycle[ 3387] = 1'b1;  wr_cycle[ 3387] = 1'b0;  addr_rom[ 3387]='h00000cf8;  wr_data_rom[ 3387]='h00000000;
    rd_cycle[ 3388] = 1'b0;  wr_cycle[ 3388] = 1'b1;  addr_rom[ 3388]='h000000e8;  wr_data_rom[ 3388]='h000000de;
    rd_cycle[ 3389] = 1'b1;  wr_cycle[ 3389] = 1'b0;  addr_rom[ 3389]='h00000964;  wr_data_rom[ 3389]='h00000000;
    rd_cycle[ 3390] = 1'b1;  wr_cycle[ 3390] = 1'b0;  addr_rom[ 3390]='h00000dc4;  wr_data_rom[ 3390]='h00000000;
    rd_cycle[ 3391] = 1'b0;  wr_cycle[ 3391] = 1'b1;  addr_rom[ 3391]='h00000808;  wr_data_rom[ 3391]='h0000038d;
    rd_cycle[ 3392] = 1'b0;  wr_cycle[ 3392] = 1'b1;  addr_rom[ 3392]='h000000cc;  wr_data_rom[ 3392]='h00000ddf;
    rd_cycle[ 3393] = 1'b1;  wr_cycle[ 3393] = 1'b0;  addr_rom[ 3393]='h0000087c;  wr_data_rom[ 3393]='h00000000;
    rd_cycle[ 3394] = 1'b0;  wr_cycle[ 3394] = 1'b1;  addr_rom[ 3394]='h00000e74;  wr_data_rom[ 3394]='h00000212;
    rd_cycle[ 3395] = 1'b0;  wr_cycle[ 3395] = 1'b1;  addr_rom[ 3395]='h00000ccc;  wr_data_rom[ 3395]='h000007b2;
    rd_cycle[ 3396] = 1'b0;  wr_cycle[ 3396] = 1'b1;  addr_rom[ 3396]='h00000264;  wr_data_rom[ 3396]='h00000565;
    rd_cycle[ 3397] = 1'b1;  wr_cycle[ 3397] = 1'b0;  addr_rom[ 3397]='h00000e30;  wr_data_rom[ 3397]='h00000000;
    rd_cycle[ 3398] = 1'b0;  wr_cycle[ 3398] = 1'b1;  addr_rom[ 3398]='h000004ec;  wr_data_rom[ 3398]='h000004b8;
    rd_cycle[ 3399] = 1'b1;  wr_cycle[ 3399] = 1'b0;  addr_rom[ 3399]='h00000d48;  wr_data_rom[ 3399]='h00000000;
    rd_cycle[ 3400] = 1'b1;  wr_cycle[ 3400] = 1'b0;  addr_rom[ 3400]='h00000534;  wr_data_rom[ 3400]='h00000000;
    rd_cycle[ 3401] = 1'b0;  wr_cycle[ 3401] = 1'b1;  addr_rom[ 3401]='h00000bec;  wr_data_rom[ 3401]='h000009c9;
    rd_cycle[ 3402] = 1'b0;  wr_cycle[ 3402] = 1'b1;  addr_rom[ 3402]='h00000278;  wr_data_rom[ 3402]='h00000708;
    rd_cycle[ 3403] = 1'b0;  wr_cycle[ 3403] = 1'b1;  addr_rom[ 3403]='h00000b94;  wr_data_rom[ 3403]='h000000ba;
    rd_cycle[ 3404] = 1'b1;  wr_cycle[ 3404] = 1'b0;  addr_rom[ 3404]='h00000810;  wr_data_rom[ 3404]='h00000000;
    rd_cycle[ 3405] = 1'b0;  wr_cycle[ 3405] = 1'b1;  addr_rom[ 3405]='h000003ec;  wr_data_rom[ 3405]='h0000000e;
    rd_cycle[ 3406] = 1'b0;  wr_cycle[ 3406] = 1'b1;  addr_rom[ 3406]='h00000d40;  wr_data_rom[ 3406]='h00000448;
    rd_cycle[ 3407] = 1'b1;  wr_cycle[ 3407] = 1'b0;  addr_rom[ 3407]='h00000178;  wr_data_rom[ 3407]='h00000000;
    rd_cycle[ 3408] = 1'b1;  wr_cycle[ 3408] = 1'b0;  addr_rom[ 3408]='h00000720;  wr_data_rom[ 3408]='h00000000;
    rd_cycle[ 3409] = 1'b0;  wr_cycle[ 3409] = 1'b1;  addr_rom[ 3409]='h000008f0;  wr_data_rom[ 3409]='h00000334;
    rd_cycle[ 3410] = 1'b1;  wr_cycle[ 3410] = 1'b0;  addr_rom[ 3410]='h00000750;  wr_data_rom[ 3410]='h00000000;
    rd_cycle[ 3411] = 1'b1;  wr_cycle[ 3411] = 1'b0;  addr_rom[ 3411]='h00000ea4;  wr_data_rom[ 3411]='h00000000;
    rd_cycle[ 3412] = 1'b0;  wr_cycle[ 3412] = 1'b1;  addr_rom[ 3412]='h00000924;  wr_data_rom[ 3412]='h00000b03;
    rd_cycle[ 3413] = 1'b1;  wr_cycle[ 3413] = 1'b0;  addr_rom[ 3413]='h00000838;  wr_data_rom[ 3413]='h00000000;
    rd_cycle[ 3414] = 1'b1;  wr_cycle[ 3414] = 1'b0;  addr_rom[ 3414]='h00000f50;  wr_data_rom[ 3414]='h00000000;
    rd_cycle[ 3415] = 1'b0;  wr_cycle[ 3415] = 1'b1;  addr_rom[ 3415]='h000003e0;  wr_data_rom[ 3415]='h0000011c;
    rd_cycle[ 3416] = 1'b1;  wr_cycle[ 3416] = 1'b0;  addr_rom[ 3416]='h00000f74;  wr_data_rom[ 3416]='h00000000;
    rd_cycle[ 3417] = 1'b0;  wr_cycle[ 3417] = 1'b1;  addr_rom[ 3417]='h00000db8;  wr_data_rom[ 3417]='h00000f20;
    rd_cycle[ 3418] = 1'b1;  wr_cycle[ 3418] = 1'b0;  addr_rom[ 3418]='h00000d8c;  wr_data_rom[ 3418]='h00000000;
    rd_cycle[ 3419] = 1'b0;  wr_cycle[ 3419] = 1'b1;  addr_rom[ 3419]='h00000e50;  wr_data_rom[ 3419]='h00000269;
    rd_cycle[ 3420] = 1'b1;  wr_cycle[ 3420] = 1'b0;  addr_rom[ 3420]='h00000df4;  wr_data_rom[ 3420]='h00000000;
    rd_cycle[ 3421] = 1'b1;  wr_cycle[ 3421] = 1'b0;  addr_rom[ 3421]='h00000a6c;  wr_data_rom[ 3421]='h00000000;
    rd_cycle[ 3422] = 1'b1;  wr_cycle[ 3422] = 1'b0;  addr_rom[ 3422]='h00000774;  wr_data_rom[ 3422]='h00000000;
    rd_cycle[ 3423] = 1'b0;  wr_cycle[ 3423] = 1'b1;  addr_rom[ 3423]='h00000308;  wr_data_rom[ 3423]='h00000217;
    rd_cycle[ 3424] = 1'b0;  wr_cycle[ 3424] = 1'b1;  addr_rom[ 3424]='h00000e04;  wr_data_rom[ 3424]='h00000baa;
    rd_cycle[ 3425] = 1'b0;  wr_cycle[ 3425] = 1'b1;  addr_rom[ 3425]='h00000f2c;  wr_data_rom[ 3425]='h000008c3;
    rd_cycle[ 3426] = 1'b1;  wr_cycle[ 3426] = 1'b0;  addr_rom[ 3426]='h00000694;  wr_data_rom[ 3426]='h00000000;
    rd_cycle[ 3427] = 1'b0;  wr_cycle[ 3427] = 1'b1;  addr_rom[ 3427]='h00000aa4;  wr_data_rom[ 3427]='h0000008f;
    rd_cycle[ 3428] = 1'b1;  wr_cycle[ 3428] = 1'b0;  addr_rom[ 3428]='h00000634;  wr_data_rom[ 3428]='h00000000;
    rd_cycle[ 3429] = 1'b1;  wr_cycle[ 3429] = 1'b0;  addr_rom[ 3429]='h000002d8;  wr_data_rom[ 3429]='h00000000;
    rd_cycle[ 3430] = 1'b1;  wr_cycle[ 3430] = 1'b0;  addr_rom[ 3430]='h00000f84;  wr_data_rom[ 3430]='h00000000;
    rd_cycle[ 3431] = 1'b0;  wr_cycle[ 3431] = 1'b1;  addr_rom[ 3431]='h00000f0c;  wr_data_rom[ 3431]='h00000d6e;
    rd_cycle[ 3432] = 1'b0;  wr_cycle[ 3432] = 1'b1;  addr_rom[ 3432]='h00000818;  wr_data_rom[ 3432]='h0000091f;
    rd_cycle[ 3433] = 1'b1;  wr_cycle[ 3433] = 1'b0;  addr_rom[ 3433]='h00000494;  wr_data_rom[ 3433]='h00000000;
    rd_cycle[ 3434] = 1'b0;  wr_cycle[ 3434] = 1'b1;  addr_rom[ 3434]='h000008a8;  wr_data_rom[ 3434]='h00000699;
    rd_cycle[ 3435] = 1'b1;  wr_cycle[ 3435] = 1'b0;  addr_rom[ 3435]='h00000d14;  wr_data_rom[ 3435]='h00000000;
    rd_cycle[ 3436] = 1'b1;  wr_cycle[ 3436] = 1'b0;  addr_rom[ 3436]='h00000424;  wr_data_rom[ 3436]='h00000000;
    rd_cycle[ 3437] = 1'b0;  wr_cycle[ 3437] = 1'b1;  addr_rom[ 3437]='h00000838;  wr_data_rom[ 3437]='h00000b4b;
    rd_cycle[ 3438] = 1'b0;  wr_cycle[ 3438] = 1'b1;  addr_rom[ 3438]='h000005f4;  wr_data_rom[ 3438]='h00000f9b;
    rd_cycle[ 3439] = 1'b1;  wr_cycle[ 3439] = 1'b0;  addr_rom[ 3439]='h00000728;  wr_data_rom[ 3439]='h00000000;
    rd_cycle[ 3440] = 1'b0;  wr_cycle[ 3440] = 1'b1;  addr_rom[ 3440]='h00000554;  wr_data_rom[ 3440]='h000007ab;
    rd_cycle[ 3441] = 1'b0;  wr_cycle[ 3441] = 1'b1;  addr_rom[ 3441]='h00000c48;  wr_data_rom[ 3441]='h00000711;
    rd_cycle[ 3442] = 1'b0;  wr_cycle[ 3442] = 1'b1;  addr_rom[ 3442]='h00000830;  wr_data_rom[ 3442]='h00000c3c;
    rd_cycle[ 3443] = 1'b0;  wr_cycle[ 3443] = 1'b1;  addr_rom[ 3443]='h00000984;  wr_data_rom[ 3443]='h0000071a;
    rd_cycle[ 3444] = 1'b0;  wr_cycle[ 3444] = 1'b1;  addr_rom[ 3444]='h00000474;  wr_data_rom[ 3444]='h000000b6;
    rd_cycle[ 3445] = 1'b0;  wr_cycle[ 3445] = 1'b1;  addr_rom[ 3445]='h00000e80;  wr_data_rom[ 3445]='h00000884;
    rd_cycle[ 3446] = 1'b1;  wr_cycle[ 3446] = 1'b0;  addr_rom[ 3446]='h00000030;  wr_data_rom[ 3446]='h00000000;
    rd_cycle[ 3447] = 1'b0;  wr_cycle[ 3447] = 1'b1;  addr_rom[ 3447]='h00000064;  wr_data_rom[ 3447]='h00000885;
    rd_cycle[ 3448] = 1'b1;  wr_cycle[ 3448] = 1'b0;  addr_rom[ 3448]='h00000098;  wr_data_rom[ 3448]='h00000000;
    rd_cycle[ 3449] = 1'b0;  wr_cycle[ 3449] = 1'b1;  addr_rom[ 3449]='h00000424;  wr_data_rom[ 3449]='h000004a6;
    rd_cycle[ 3450] = 1'b0;  wr_cycle[ 3450] = 1'b1;  addr_rom[ 3450]='h00000870;  wr_data_rom[ 3450]='h000007a6;
    rd_cycle[ 3451] = 1'b0;  wr_cycle[ 3451] = 1'b1;  addr_rom[ 3451]='h000004dc;  wr_data_rom[ 3451]='h00000405;
    rd_cycle[ 3452] = 1'b1;  wr_cycle[ 3452] = 1'b0;  addr_rom[ 3452]='h00000c58;  wr_data_rom[ 3452]='h00000000;
    rd_cycle[ 3453] = 1'b0;  wr_cycle[ 3453] = 1'b1;  addr_rom[ 3453]='h000005dc;  wr_data_rom[ 3453]='h00000e1a;
    rd_cycle[ 3454] = 1'b1;  wr_cycle[ 3454] = 1'b0;  addr_rom[ 3454]='h000000cc;  wr_data_rom[ 3454]='h00000000;
    rd_cycle[ 3455] = 1'b0;  wr_cycle[ 3455] = 1'b1;  addr_rom[ 3455]='h000000f4;  wr_data_rom[ 3455]='h00000867;
    rd_cycle[ 3456] = 1'b1;  wr_cycle[ 3456] = 1'b0;  addr_rom[ 3456]='h00000bc0;  wr_data_rom[ 3456]='h00000000;
    rd_cycle[ 3457] = 1'b1;  wr_cycle[ 3457] = 1'b0;  addr_rom[ 3457]='h000008b4;  wr_data_rom[ 3457]='h00000000;
    rd_cycle[ 3458] = 1'b1;  wr_cycle[ 3458] = 1'b0;  addr_rom[ 3458]='h000002dc;  wr_data_rom[ 3458]='h00000000;
    rd_cycle[ 3459] = 1'b1;  wr_cycle[ 3459] = 1'b0;  addr_rom[ 3459]='h00000654;  wr_data_rom[ 3459]='h00000000;
    rd_cycle[ 3460] = 1'b1;  wr_cycle[ 3460] = 1'b0;  addr_rom[ 3460]='h000007c8;  wr_data_rom[ 3460]='h00000000;
    rd_cycle[ 3461] = 1'b0;  wr_cycle[ 3461] = 1'b1;  addr_rom[ 3461]='h000006c4;  wr_data_rom[ 3461]='h000003b7;
    rd_cycle[ 3462] = 1'b1;  wr_cycle[ 3462] = 1'b0;  addr_rom[ 3462]='h00000c54;  wr_data_rom[ 3462]='h00000000;
    rd_cycle[ 3463] = 1'b0;  wr_cycle[ 3463] = 1'b1;  addr_rom[ 3463]='h00000128;  wr_data_rom[ 3463]='h00000cd7;
    rd_cycle[ 3464] = 1'b0;  wr_cycle[ 3464] = 1'b1;  addr_rom[ 3464]='h00000b94;  wr_data_rom[ 3464]='h000007be;
    rd_cycle[ 3465] = 1'b0;  wr_cycle[ 3465] = 1'b1;  addr_rom[ 3465]='h000001f4;  wr_data_rom[ 3465]='h00000750;
    rd_cycle[ 3466] = 1'b1;  wr_cycle[ 3466] = 1'b0;  addr_rom[ 3466]='h000000a4;  wr_data_rom[ 3466]='h00000000;
    rd_cycle[ 3467] = 1'b1;  wr_cycle[ 3467] = 1'b0;  addr_rom[ 3467]='h00000d20;  wr_data_rom[ 3467]='h00000000;
    rd_cycle[ 3468] = 1'b0;  wr_cycle[ 3468] = 1'b1;  addr_rom[ 3468]='h00000ed4;  wr_data_rom[ 3468]='h00000dd9;
    rd_cycle[ 3469] = 1'b0;  wr_cycle[ 3469] = 1'b1;  addr_rom[ 3469]='h00000af8;  wr_data_rom[ 3469]='h00000d02;
    rd_cycle[ 3470] = 1'b1;  wr_cycle[ 3470] = 1'b0;  addr_rom[ 3470]='h00000818;  wr_data_rom[ 3470]='h00000000;
    rd_cycle[ 3471] = 1'b1;  wr_cycle[ 3471] = 1'b0;  addr_rom[ 3471]='h00000294;  wr_data_rom[ 3471]='h00000000;
    rd_cycle[ 3472] = 1'b1;  wr_cycle[ 3472] = 1'b0;  addr_rom[ 3472]='h00000314;  wr_data_rom[ 3472]='h00000000;
    rd_cycle[ 3473] = 1'b1;  wr_cycle[ 3473] = 1'b0;  addr_rom[ 3473]='h000001cc;  wr_data_rom[ 3473]='h00000000;
    rd_cycle[ 3474] = 1'b1;  wr_cycle[ 3474] = 1'b0;  addr_rom[ 3474]='h0000010c;  wr_data_rom[ 3474]='h00000000;
    rd_cycle[ 3475] = 1'b0;  wr_cycle[ 3475] = 1'b1;  addr_rom[ 3475]='h00000eac;  wr_data_rom[ 3475]='h000006a4;
    rd_cycle[ 3476] = 1'b1;  wr_cycle[ 3476] = 1'b0;  addr_rom[ 3476]='h000000f8;  wr_data_rom[ 3476]='h00000000;
    rd_cycle[ 3477] = 1'b0;  wr_cycle[ 3477] = 1'b1;  addr_rom[ 3477]='h00000a20;  wr_data_rom[ 3477]='h000003bd;
    rd_cycle[ 3478] = 1'b0;  wr_cycle[ 3478] = 1'b1;  addr_rom[ 3478]='h000007d0;  wr_data_rom[ 3478]='h00000559;
    rd_cycle[ 3479] = 1'b0;  wr_cycle[ 3479] = 1'b1;  addr_rom[ 3479]='h00000d7c;  wr_data_rom[ 3479]='h00000c73;
    rd_cycle[ 3480] = 1'b0;  wr_cycle[ 3480] = 1'b1;  addr_rom[ 3480]='h000009c0;  wr_data_rom[ 3480]='h000009bd;
    rd_cycle[ 3481] = 1'b0;  wr_cycle[ 3481] = 1'b1;  addr_rom[ 3481]='h000007bc;  wr_data_rom[ 3481]='h000006fb;
    rd_cycle[ 3482] = 1'b1;  wr_cycle[ 3482] = 1'b0;  addr_rom[ 3482]='h0000074c;  wr_data_rom[ 3482]='h00000000;
    rd_cycle[ 3483] = 1'b1;  wr_cycle[ 3483] = 1'b0;  addr_rom[ 3483]='h000007e8;  wr_data_rom[ 3483]='h00000000;
    rd_cycle[ 3484] = 1'b1;  wr_cycle[ 3484] = 1'b0;  addr_rom[ 3484]='h00000ce8;  wr_data_rom[ 3484]='h00000000;
    rd_cycle[ 3485] = 1'b0;  wr_cycle[ 3485] = 1'b1;  addr_rom[ 3485]='h00000654;  wr_data_rom[ 3485]='h0000007f;
    rd_cycle[ 3486] = 1'b1;  wr_cycle[ 3486] = 1'b0;  addr_rom[ 3486]='h00000760;  wr_data_rom[ 3486]='h00000000;
    rd_cycle[ 3487] = 1'b1;  wr_cycle[ 3487] = 1'b0;  addr_rom[ 3487]='h00000264;  wr_data_rom[ 3487]='h00000000;
    rd_cycle[ 3488] = 1'b0;  wr_cycle[ 3488] = 1'b1;  addr_rom[ 3488]='h0000037c;  wr_data_rom[ 3488]='h000003cc;
    rd_cycle[ 3489] = 1'b1;  wr_cycle[ 3489] = 1'b0;  addr_rom[ 3489]='h0000069c;  wr_data_rom[ 3489]='h00000000;
    rd_cycle[ 3490] = 1'b1;  wr_cycle[ 3490] = 1'b0;  addr_rom[ 3490]='h00000a04;  wr_data_rom[ 3490]='h00000000;
    rd_cycle[ 3491] = 1'b0;  wr_cycle[ 3491] = 1'b1;  addr_rom[ 3491]='h00000aec;  wr_data_rom[ 3491]='h00000883;
    rd_cycle[ 3492] = 1'b0;  wr_cycle[ 3492] = 1'b1;  addr_rom[ 3492]='h00000558;  wr_data_rom[ 3492]='h000000f6;
    rd_cycle[ 3493] = 1'b1;  wr_cycle[ 3493] = 1'b0;  addr_rom[ 3493]='h00000dbc;  wr_data_rom[ 3493]='h00000000;
    rd_cycle[ 3494] = 1'b0;  wr_cycle[ 3494] = 1'b1;  addr_rom[ 3494]='h0000043c;  wr_data_rom[ 3494]='h00000e34;
    rd_cycle[ 3495] = 1'b0;  wr_cycle[ 3495] = 1'b1;  addr_rom[ 3495]='h00000cc0;  wr_data_rom[ 3495]='h00000384;
    rd_cycle[ 3496] = 1'b0;  wr_cycle[ 3496] = 1'b1;  addr_rom[ 3496]='h00000528;  wr_data_rom[ 3496]='h00000405;
    rd_cycle[ 3497] = 1'b1;  wr_cycle[ 3497] = 1'b0;  addr_rom[ 3497]='h00000be4;  wr_data_rom[ 3497]='h00000000;
    rd_cycle[ 3498] = 1'b1;  wr_cycle[ 3498] = 1'b0;  addr_rom[ 3498]='h00000428;  wr_data_rom[ 3498]='h00000000;
    rd_cycle[ 3499] = 1'b0;  wr_cycle[ 3499] = 1'b1;  addr_rom[ 3499]='h00000f64;  wr_data_rom[ 3499]='h00000512;
    rd_cycle[ 3500] = 1'b1;  wr_cycle[ 3500] = 1'b0;  addr_rom[ 3500]='h000008e0;  wr_data_rom[ 3500]='h00000000;
    rd_cycle[ 3501] = 1'b0;  wr_cycle[ 3501] = 1'b1;  addr_rom[ 3501]='h0000042c;  wr_data_rom[ 3501]='h00000473;
    rd_cycle[ 3502] = 1'b1;  wr_cycle[ 3502] = 1'b0;  addr_rom[ 3502]='h00000248;  wr_data_rom[ 3502]='h00000000;
    rd_cycle[ 3503] = 1'b0;  wr_cycle[ 3503] = 1'b1;  addr_rom[ 3503]='h00000860;  wr_data_rom[ 3503]='h00000068;
    rd_cycle[ 3504] = 1'b1;  wr_cycle[ 3504] = 1'b0;  addr_rom[ 3504]='h000005c8;  wr_data_rom[ 3504]='h00000000;
    rd_cycle[ 3505] = 1'b1;  wr_cycle[ 3505] = 1'b0;  addr_rom[ 3505]='h00000b54;  wr_data_rom[ 3505]='h00000000;
    rd_cycle[ 3506] = 1'b1;  wr_cycle[ 3506] = 1'b0;  addr_rom[ 3506]='h0000092c;  wr_data_rom[ 3506]='h00000000;
    rd_cycle[ 3507] = 1'b0;  wr_cycle[ 3507] = 1'b1;  addr_rom[ 3507]='h00000a5c;  wr_data_rom[ 3507]='h0000028a;
    rd_cycle[ 3508] = 1'b1;  wr_cycle[ 3508] = 1'b0;  addr_rom[ 3508]='h00000250;  wr_data_rom[ 3508]='h00000000;
    rd_cycle[ 3509] = 1'b1;  wr_cycle[ 3509] = 1'b0;  addr_rom[ 3509]='h00000dd0;  wr_data_rom[ 3509]='h00000000;
    rd_cycle[ 3510] = 1'b0;  wr_cycle[ 3510] = 1'b1;  addr_rom[ 3510]='h00000544;  wr_data_rom[ 3510]='h00000a7f;
    rd_cycle[ 3511] = 1'b0;  wr_cycle[ 3511] = 1'b1;  addr_rom[ 3511]='h00000d30;  wr_data_rom[ 3511]='h000003f5;
    rd_cycle[ 3512] = 1'b0;  wr_cycle[ 3512] = 1'b1;  addr_rom[ 3512]='h00000b58;  wr_data_rom[ 3512]='h00000f36;
    rd_cycle[ 3513] = 1'b0;  wr_cycle[ 3513] = 1'b1;  addr_rom[ 3513]='h00000b80;  wr_data_rom[ 3513]='h00000030;
    rd_cycle[ 3514] = 1'b1;  wr_cycle[ 3514] = 1'b0;  addr_rom[ 3514]='h00000ac8;  wr_data_rom[ 3514]='h00000000;
    rd_cycle[ 3515] = 1'b1;  wr_cycle[ 3515] = 1'b0;  addr_rom[ 3515]='h000001b0;  wr_data_rom[ 3515]='h00000000;
    rd_cycle[ 3516] = 1'b0;  wr_cycle[ 3516] = 1'b1;  addr_rom[ 3516]='h00000818;  wr_data_rom[ 3516]='h0000004a;
    rd_cycle[ 3517] = 1'b1;  wr_cycle[ 3517] = 1'b0;  addr_rom[ 3517]='h00000074;  wr_data_rom[ 3517]='h00000000;
    rd_cycle[ 3518] = 1'b0;  wr_cycle[ 3518] = 1'b1;  addr_rom[ 3518]='h00000078;  wr_data_rom[ 3518]='h000008f1;
    rd_cycle[ 3519] = 1'b1;  wr_cycle[ 3519] = 1'b0;  addr_rom[ 3519]='h0000047c;  wr_data_rom[ 3519]='h00000000;
    rd_cycle[ 3520] = 1'b0;  wr_cycle[ 3520] = 1'b1;  addr_rom[ 3520]='h000008c0;  wr_data_rom[ 3520]='h0000011c;
    rd_cycle[ 3521] = 1'b1;  wr_cycle[ 3521] = 1'b0;  addr_rom[ 3521]='h000007a4;  wr_data_rom[ 3521]='h00000000;
    rd_cycle[ 3522] = 1'b1;  wr_cycle[ 3522] = 1'b0;  addr_rom[ 3522]='h00000b74;  wr_data_rom[ 3522]='h00000000;
    rd_cycle[ 3523] = 1'b0;  wr_cycle[ 3523] = 1'b1;  addr_rom[ 3523]='h00000094;  wr_data_rom[ 3523]='h0000073d;
    rd_cycle[ 3524] = 1'b0;  wr_cycle[ 3524] = 1'b1;  addr_rom[ 3524]='h00000220;  wr_data_rom[ 3524]='h000009db;
    rd_cycle[ 3525] = 1'b1;  wr_cycle[ 3525] = 1'b0;  addr_rom[ 3525]='h00000778;  wr_data_rom[ 3525]='h00000000;
    rd_cycle[ 3526] = 1'b0;  wr_cycle[ 3526] = 1'b1;  addr_rom[ 3526]='h00000358;  wr_data_rom[ 3526]='h00000317;
    rd_cycle[ 3527] = 1'b1;  wr_cycle[ 3527] = 1'b0;  addr_rom[ 3527]='h000006e4;  wr_data_rom[ 3527]='h00000000;
    rd_cycle[ 3528] = 1'b1;  wr_cycle[ 3528] = 1'b0;  addr_rom[ 3528]='h00000224;  wr_data_rom[ 3528]='h00000000;
    rd_cycle[ 3529] = 1'b1;  wr_cycle[ 3529] = 1'b0;  addr_rom[ 3529]='h0000075c;  wr_data_rom[ 3529]='h00000000;
    rd_cycle[ 3530] = 1'b0;  wr_cycle[ 3530] = 1'b1;  addr_rom[ 3530]='h00000a8c;  wr_data_rom[ 3530]='h00000edb;
    rd_cycle[ 3531] = 1'b0;  wr_cycle[ 3531] = 1'b1;  addr_rom[ 3531]='h000008f8;  wr_data_rom[ 3531]='h00000bec;
    rd_cycle[ 3532] = 1'b1;  wr_cycle[ 3532] = 1'b0;  addr_rom[ 3532]='h000002bc;  wr_data_rom[ 3532]='h00000000;
    rd_cycle[ 3533] = 1'b0;  wr_cycle[ 3533] = 1'b1;  addr_rom[ 3533]='h000005dc;  wr_data_rom[ 3533]='h00000659;
    rd_cycle[ 3534] = 1'b1;  wr_cycle[ 3534] = 1'b0;  addr_rom[ 3534]='h000003a8;  wr_data_rom[ 3534]='h00000000;
    rd_cycle[ 3535] = 1'b0;  wr_cycle[ 3535] = 1'b1;  addr_rom[ 3535]='h00000b64;  wr_data_rom[ 3535]='h000000af;
    rd_cycle[ 3536] = 1'b0;  wr_cycle[ 3536] = 1'b1;  addr_rom[ 3536]='h00000c44;  wr_data_rom[ 3536]='h00000253;
    rd_cycle[ 3537] = 1'b1;  wr_cycle[ 3537] = 1'b0;  addr_rom[ 3537]='h00000704;  wr_data_rom[ 3537]='h00000000;
    rd_cycle[ 3538] = 1'b0;  wr_cycle[ 3538] = 1'b1;  addr_rom[ 3538]='h00000e6c;  wr_data_rom[ 3538]='h000004b0;
    rd_cycle[ 3539] = 1'b0;  wr_cycle[ 3539] = 1'b1;  addr_rom[ 3539]='h00000a1c;  wr_data_rom[ 3539]='h00000d22;
    rd_cycle[ 3540] = 1'b1;  wr_cycle[ 3540] = 1'b0;  addr_rom[ 3540]='h00000a38;  wr_data_rom[ 3540]='h00000000;
    rd_cycle[ 3541] = 1'b0;  wr_cycle[ 3541] = 1'b1;  addr_rom[ 3541]='h00000dcc;  wr_data_rom[ 3541]='h00000a5d;
    rd_cycle[ 3542] = 1'b0;  wr_cycle[ 3542] = 1'b1;  addr_rom[ 3542]='h000007e8;  wr_data_rom[ 3542]='h00000086;
    rd_cycle[ 3543] = 1'b0;  wr_cycle[ 3543] = 1'b1;  addr_rom[ 3543]='h00000594;  wr_data_rom[ 3543]='h00000a9a;
    rd_cycle[ 3544] = 1'b0;  wr_cycle[ 3544] = 1'b1;  addr_rom[ 3544]='h00000518;  wr_data_rom[ 3544]='h000005de;
    rd_cycle[ 3545] = 1'b1;  wr_cycle[ 3545] = 1'b0;  addr_rom[ 3545]='h00000a4c;  wr_data_rom[ 3545]='h00000000;
    rd_cycle[ 3546] = 1'b1;  wr_cycle[ 3546] = 1'b0;  addr_rom[ 3546]='h00000c08;  wr_data_rom[ 3546]='h00000000;
    rd_cycle[ 3547] = 1'b0;  wr_cycle[ 3547] = 1'b1;  addr_rom[ 3547]='h000003cc;  wr_data_rom[ 3547]='h00000451;
    rd_cycle[ 3548] = 1'b0;  wr_cycle[ 3548] = 1'b1;  addr_rom[ 3548]='h00000898;  wr_data_rom[ 3548]='h00000748;
    rd_cycle[ 3549] = 1'b0;  wr_cycle[ 3549] = 1'b1;  addr_rom[ 3549]='h00000dcc;  wr_data_rom[ 3549]='h00000419;
    rd_cycle[ 3550] = 1'b1;  wr_cycle[ 3550] = 1'b0;  addr_rom[ 3550]='h00000cb4;  wr_data_rom[ 3550]='h00000000;
    rd_cycle[ 3551] = 1'b1;  wr_cycle[ 3551] = 1'b0;  addr_rom[ 3551]='h00000f2c;  wr_data_rom[ 3551]='h00000000;
    rd_cycle[ 3552] = 1'b1;  wr_cycle[ 3552] = 1'b0;  addr_rom[ 3552]='h000008b8;  wr_data_rom[ 3552]='h00000000;
    rd_cycle[ 3553] = 1'b0;  wr_cycle[ 3553] = 1'b1;  addr_rom[ 3553]='h00000ab4;  wr_data_rom[ 3553]='h0000018b;
    rd_cycle[ 3554] = 1'b1;  wr_cycle[ 3554] = 1'b0;  addr_rom[ 3554]='h00000188;  wr_data_rom[ 3554]='h00000000;
    rd_cycle[ 3555] = 1'b1;  wr_cycle[ 3555] = 1'b0;  addr_rom[ 3555]='h00000f78;  wr_data_rom[ 3555]='h00000000;
    rd_cycle[ 3556] = 1'b0;  wr_cycle[ 3556] = 1'b1;  addr_rom[ 3556]='h000006f8;  wr_data_rom[ 3556]='h00000c0a;
    rd_cycle[ 3557] = 1'b0;  wr_cycle[ 3557] = 1'b1;  addr_rom[ 3557]='h0000062c;  wr_data_rom[ 3557]='h00000a64;
    rd_cycle[ 3558] = 1'b0;  wr_cycle[ 3558] = 1'b1;  addr_rom[ 3558]='h000000c4;  wr_data_rom[ 3558]='h00000472;
    rd_cycle[ 3559] = 1'b0;  wr_cycle[ 3559] = 1'b1;  addr_rom[ 3559]='h0000052c;  wr_data_rom[ 3559]='h0000027f;
    rd_cycle[ 3560] = 1'b1;  wr_cycle[ 3560] = 1'b0;  addr_rom[ 3560]='h00000eb8;  wr_data_rom[ 3560]='h00000000;
    rd_cycle[ 3561] = 1'b0;  wr_cycle[ 3561] = 1'b1;  addr_rom[ 3561]='h0000095c;  wr_data_rom[ 3561]='h00000f41;
    rd_cycle[ 3562] = 1'b0;  wr_cycle[ 3562] = 1'b1;  addr_rom[ 3562]='h000001b4;  wr_data_rom[ 3562]='h0000036e;
    rd_cycle[ 3563] = 1'b1;  wr_cycle[ 3563] = 1'b0;  addr_rom[ 3563]='h000007d8;  wr_data_rom[ 3563]='h00000000;
    rd_cycle[ 3564] = 1'b0;  wr_cycle[ 3564] = 1'b1;  addr_rom[ 3564]='h00000478;  wr_data_rom[ 3564]='h00000017;
    rd_cycle[ 3565] = 1'b0;  wr_cycle[ 3565] = 1'b1;  addr_rom[ 3565]='h00000664;  wr_data_rom[ 3565]='h00000a36;
    rd_cycle[ 3566] = 1'b1;  wr_cycle[ 3566] = 1'b0;  addr_rom[ 3566]='h00000e58;  wr_data_rom[ 3566]='h00000000;
    rd_cycle[ 3567] = 1'b1;  wr_cycle[ 3567] = 1'b0;  addr_rom[ 3567]='h00000b00;  wr_data_rom[ 3567]='h00000000;
    rd_cycle[ 3568] = 1'b1;  wr_cycle[ 3568] = 1'b0;  addr_rom[ 3568]='h00000560;  wr_data_rom[ 3568]='h00000000;
    rd_cycle[ 3569] = 1'b0;  wr_cycle[ 3569] = 1'b1;  addr_rom[ 3569]='h000007c8;  wr_data_rom[ 3569]='h00000ea2;
    rd_cycle[ 3570] = 1'b0;  wr_cycle[ 3570] = 1'b1;  addr_rom[ 3570]='h000009d8;  wr_data_rom[ 3570]='h0000096b;
    rd_cycle[ 3571] = 1'b1;  wr_cycle[ 3571] = 1'b0;  addr_rom[ 3571]='h00000c78;  wr_data_rom[ 3571]='h00000000;
    rd_cycle[ 3572] = 1'b0;  wr_cycle[ 3572] = 1'b1;  addr_rom[ 3572]='h00000274;  wr_data_rom[ 3572]='h000004d9;
    rd_cycle[ 3573] = 1'b0;  wr_cycle[ 3573] = 1'b1;  addr_rom[ 3573]='h00000954;  wr_data_rom[ 3573]='h000004d0;
    rd_cycle[ 3574] = 1'b1;  wr_cycle[ 3574] = 1'b0;  addr_rom[ 3574]='h0000051c;  wr_data_rom[ 3574]='h00000000;
    rd_cycle[ 3575] = 1'b0;  wr_cycle[ 3575] = 1'b1;  addr_rom[ 3575]='h00000110;  wr_data_rom[ 3575]='h00000831;
    rd_cycle[ 3576] = 1'b0;  wr_cycle[ 3576] = 1'b1;  addr_rom[ 3576]='h00000848;  wr_data_rom[ 3576]='h00000d31;
    rd_cycle[ 3577] = 1'b1;  wr_cycle[ 3577] = 1'b0;  addr_rom[ 3577]='h00000c58;  wr_data_rom[ 3577]='h00000000;
    rd_cycle[ 3578] = 1'b1;  wr_cycle[ 3578] = 1'b0;  addr_rom[ 3578]='h000003e0;  wr_data_rom[ 3578]='h00000000;
    rd_cycle[ 3579] = 1'b0;  wr_cycle[ 3579] = 1'b1;  addr_rom[ 3579]='h000008a0;  wr_data_rom[ 3579]='h00000932;
    rd_cycle[ 3580] = 1'b1;  wr_cycle[ 3580] = 1'b0;  addr_rom[ 3580]='h00000100;  wr_data_rom[ 3580]='h00000000;
    rd_cycle[ 3581] = 1'b1;  wr_cycle[ 3581] = 1'b0;  addr_rom[ 3581]='h00000ef4;  wr_data_rom[ 3581]='h00000000;
    rd_cycle[ 3582] = 1'b1;  wr_cycle[ 3582] = 1'b0;  addr_rom[ 3582]='h00000f70;  wr_data_rom[ 3582]='h00000000;
    rd_cycle[ 3583] = 1'b1;  wr_cycle[ 3583] = 1'b0;  addr_rom[ 3583]='h000002f4;  wr_data_rom[ 3583]='h00000000;
    rd_cycle[ 3584] = 1'b1;  wr_cycle[ 3584] = 1'b0;  addr_rom[ 3584]='h0000047c;  wr_data_rom[ 3584]='h00000000;
    rd_cycle[ 3585] = 1'b1;  wr_cycle[ 3585] = 1'b0;  addr_rom[ 3585]='h000003fc;  wr_data_rom[ 3585]='h00000000;
    rd_cycle[ 3586] = 1'b0;  wr_cycle[ 3586] = 1'b1;  addr_rom[ 3586]='h00000e70;  wr_data_rom[ 3586]='h00000519;
    rd_cycle[ 3587] = 1'b0;  wr_cycle[ 3587] = 1'b1;  addr_rom[ 3587]='h00000104;  wr_data_rom[ 3587]='h00000276;
    rd_cycle[ 3588] = 1'b0;  wr_cycle[ 3588] = 1'b1;  addr_rom[ 3588]='h000003e8;  wr_data_rom[ 3588]='h00000b35;
    rd_cycle[ 3589] = 1'b1;  wr_cycle[ 3589] = 1'b0;  addr_rom[ 3589]='h0000026c;  wr_data_rom[ 3589]='h00000000;
    rd_cycle[ 3590] = 1'b0;  wr_cycle[ 3590] = 1'b1;  addr_rom[ 3590]='h00000a7c;  wr_data_rom[ 3590]='h0000096f;
    rd_cycle[ 3591] = 1'b1;  wr_cycle[ 3591] = 1'b0;  addr_rom[ 3591]='h00000ce8;  wr_data_rom[ 3591]='h00000000;
    rd_cycle[ 3592] = 1'b0;  wr_cycle[ 3592] = 1'b1;  addr_rom[ 3592]='h000009cc;  wr_data_rom[ 3592]='h00000e89;
    rd_cycle[ 3593] = 1'b0;  wr_cycle[ 3593] = 1'b1;  addr_rom[ 3593]='h00000a3c;  wr_data_rom[ 3593]='h00000201;
    rd_cycle[ 3594] = 1'b0;  wr_cycle[ 3594] = 1'b1;  addr_rom[ 3594]='h00000600;  wr_data_rom[ 3594]='h00000e07;
    rd_cycle[ 3595] = 1'b1;  wr_cycle[ 3595] = 1'b0;  addr_rom[ 3595]='h00000dac;  wr_data_rom[ 3595]='h00000000;
    rd_cycle[ 3596] = 1'b1;  wr_cycle[ 3596] = 1'b0;  addr_rom[ 3596]='h000003d0;  wr_data_rom[ 3596]='h00000000;
    rd_cycle[ 3597] = 1'b1;  wr_cycle[ 3597] = 1'b0;  addr_rom[ 3597]='h000008a0;  wr_data_rom[ 3597]='h00000000;
    rd_cycle[ 3598] = 1'b1;  wr_cycle[ 3598] = 1'b0;  addr_rom[ 3598]='h00000318;  wr_data_rom[ 3598]='h00000000;
    rd_cycle[ 3599] = 1'b1;  wr_cycle[ 3599] = 1'b0;  addr_rom[ 3599]='h00000e04;  wr_data_rom[ 3599]='h00000000;
    rd_cycle[ 3600] = 1'b1;  wr_cycle[ 3600] = 1'b0;  addr_rom[ 3600]='h000006b8;  wr_data_rom[ 3600]='h00000000;
    rd_cycle[ 3601] = 1'b1;  wr_cycle[ 3601] = 1'b0;  addr_rom[ 3601]='h00000828;  wr_data_rom[ 3601]='h00000000;
    rd_cycle[ 3602] = 1'b0;  wr_cycle[ 3602] = 1'b1;  addr_rom[ 3602]='h00000acc;  wr_data_rom[ 3602]='h00000b93;
    rd_cycle[ 3603] = 1'b1;  wr_cycle[ 3603] = 1'b0;  addr_rom[ 3603]='h00000b4c;  wr_data_rom[ 3603]='h00000000;
    rd_cycle[ 3604] = 1'b0;  wr_cycle[ 3604] = 1'b1;  addr_rom[ 3604]='h00000f00;  wr_data_rom[ 3604]='h0000039f;
    rd_cycle[ 3605] = 1'b1;  wr_cycle[ 3605] = 1'b0;  addr_rom[ 3605]='h00000848;  wr_data_rom[ 3605]='h00000000;
    rd_cycle[ 3606] = 1'b0;  wr_cycle[ 3606] = 1'b1;  addr_rom[ 3606]='h000002f4;  wr_data_rom[ 3606]='h00000038;
    rd_cycle[ 3607] = 1'b0;  wr_cycle[ 3607] = 1'b1;  addr_rom[ 3607]='h00000208;  wr_data_rom[ 3607]='h00000ad3;
    rd_cycle[ 3608] = 1'b0;  wr_cycle[ 3608] = 1'b1;  addr_rom[ 3608]='h00000160;  wr_data_rom[ 3608]='h00000c5e;
    rd_cycle[ 3609] = 1'b0;  wr_cycle[ 3609] = 1'b1;  addr_rom[ 3609]='h00000a80;  wr_data_rom[ 3609]='h00000194;
    rd_cycle[ 3610] = 1'b0;  wr_cycle[ 3610] = 1'b1;  addr_rom[ 3610]='h000006a0;  wr_data_rom[ 3610]='h0000069f;
    rd_cycle[ 3611] = 1'b0;  wr_cycle[ 3611] = 1'b1;  addr_rom[ 3611]='h00000724;  wr_data_rom[ 3611]='h00000c4d;
    rd_cycle[ 3612] = 1'b1;  wr_cycle[ 3612] = 1'b0;  addr_rom[ 3612]='h00000c4c;  wr_data_rom[ 3612]='h00000000;
    rd_cycle[ 3613] = 1'b0;  wr_cycle[ 3613] = 1'b1;  addr_rom[ 3613]='h00000c40;  wr_data_rom[ 3613]='h00000867;
    rd_cycle[ 3614] = 1'b1;  wr_cycle[ 3614] = 1'b0;  addr_rom[ 3614]='h00000be0;  wr_data_rom[ 3614]='h00000000;
    rd_cycle[ 3615] = 1'b0;  wr_cycle[ 3615] = 1'b1;  addr_rom[ 3615]='h000002a8;  wr_data_rom[ 3615]='h0000086f;
    rd_cycle[ 3616] = 1'b0;  wr_cycle[ 3616] = 1'b1;  addr_rom[ 3616]='h00000860;  wr_data_rom[ 3616]='h000004a0;
    rd_cycle[ 3617] = 1'b0;  wr_cycle[ 3617] = 1'b1;  addr_rom[ 3617]='h00000e4c;  wr_data_rom[ 3617]='h00000b91;
    rd_cycle[ 3618] = 1'b0;  wr_cycle[ 3618] = 1'b1;  addr_rom[ 3618]='h0000063c;  wr_data_rom[ 3618]='h00000f3d;
    rd_cycle[ 3619] = 1'b0;  wr_cycle[ 3619] = 1'b1;  addr_rom[ 3619]='h00000440;  wr_data_rom[ 3619]='h000006be;
    rd_cycle[ 3620] = 1'b1;  wr_cycle[ 3620] = 1'b0;  addr_rom[ 3620]='h0000014c;  wr_data_rom[ 3620]='h00000000;
    rd_cycle[ 3621] = 1'b1;  wr_cycle[ 3621] = 1'b0;  addr_rom[ 3621]='h00000308;  wr_data_rom[ 3621]='h00000000;
    rd_cycle[ 3622] = 1'b1;  wr_cycle[ 3622] = 1'b0;  addr_rom[ 3622]='h00000144;  wr_data_rom[ 3622]='h00000000;
    rd_cycle[ 3623] = 1'b1;  wr_cycle[ 3623] = 1'b0;  addr_rom[ 3623]='h00000c5c;  wr_data_rom[ 3623]='h00000000;
    rd_cycle[ 3624] = 1'b1;  wr_cycle[ 3624] = 1'b0;  addr_rom[ 3624]='h00000c20;  wr_data_rom[ 3624]='h00000000;
    rd_cycle[ 3625] = 1'b0;  wr_cycle[ 3625] = 1'b1;  addr_rom[ 3625]='h000001fc;  wr_data_rom[ 3625]='h000003fc;
    rd_cycle[ 3626] = 1'b0;  wr_cycle[ 3626] = 1'b1;  addr_rom[ 3626]='h000006e0;  wr_data_rom[ 3626]='h00000e81;
    rd_cycle[ 3627] = 1'b0;  wr_cycle[ 3627] = 1'b1;  addr_rom[ 3627]='h0000033c;  wr_data_rom[ 3627]='h00000351;
    rd_cycle[ 3628] = 1'b0;  wr_cycle[ 3628] = 1'b1;  addr_rom[ 3628]='h0000039c;  wr_data_rom[ 3628]='h00000b69;
    rd_cycle[ 3629] = 1'b0;  wr_cycle[ 3629] = 1'b1;  addr_rom[ 3629]='h000003a8;  wr_data_rom[ 3629]='h00000d12;
    rd_cycle[ 3630] = 1'b1;  wr_cycle[ 3630] = 1'b0;  addr_rom[ 3630]='h00000554;  wr_data_rom[ 3630]='h00000000;
    rd_cycle[ 3631] = 1'b0;  wr_cycle[ 3631] = 1'b1;  addr_rom[ 3631]='h00000b8c;  wr_data_rom[ 3631]='h00000862;
    rd_cycle[ 3632] = 1'b1;  wr_cycle[ 3632] = 1'b0;  addr_rom[ 3632]='h00000560;  wr_data_rom[ 3632]='h00000000;
    rd_cycle[ 3633] = 1'b0;  wr_cycle[ 3633] = 1'b1;  addr_rom[ 3633]='h000003d0;  wr_data_rom[ 3633]='h00000df5;
    rd_cycle[ 3634] = 1'b0;  wr_cycle[ 3634] = 1'b1;  addr_rom[ 3634]='h00000b58;  wr_data_rom[ 3634]='h0000036d;
    rd_cycle[ 3635] = 1'b1;  wr_cycle[ 3635] = 1'b0;  addr_rom[ 3635]='h000000fc;  wr_data_rom[ 3635]='h00000000;
    rd_cycle[ 3636] = 1'b0;  wr_cycle[ 3636] = 1'b1;  addr_rom[ 3636]='h00000e50;  wr_data_rom[ 3636]='h00000acc;
    rd_cycle[ 3637] = 1'b0;  wr_cycle[ 3637] = 1'b1;  addr_rom[ 3637]='h0000038c;  wr_data_rom[ 3637]='h00000b1f;
    rd_cycle[ 3638] = 1'b0;  wr_cycle[ 3638] = 1'b1;  addr_rom[ 3638]='h00000760;  wr_data_rom[ 3638]='h00000aa0;
    rd_cycle[ 3639] = 1'b0;  wr_cycle[ 3639] = 1'b1;  addr_rom[ 3639]='h00000f4c;  wr_data_rom[ 3639]='h00000133;
    rd_cycle[ 3640] = 1'b1;  wr_cycle[ 3640] = 1'b0;  addr_rom[ 3640]='h000004a4;  wr_data_rom[ 3640]='h00000000;
    rd_cycle[ 3641] = 1'b1;  wr_cycle[ 3641] = 1'b0;  addr_rom[ 3641]='h000001f0;  wr_data_rom[ 3641]='h00000000;
    rd_cycle[ 3642] = 1'b0;  wr_cycle[ 3642] = 1'b1;  addr_rom[ 3642]='h000001f0;  wr_data_rom[ 3642]='h00000ba3;
    rd_cycle[ 3643] = 1'b0;  wr_cycle[ 3643] = 1'b1;  addr_rom[ 3643]='h00000678;  wr_data_rom[ 3643]='h000006d7;
    rd_cycle[ 3644] = 1'b0;  wr_cycle[ 3644] = 1'b1;  addr_rom[ 3644]='h0000071c;  wr_data_rom[ 3644]='h00000b54;
    rd_cycle[ 3645] = 1'b1;  wr_cycle[ 3645] = 1'b0;  addr_rom[ 3645]='h00000800;  wr_data_rom[ 3645]='h00000000;
    rd_cycle[ 3646] = 1'b1;  wr_cycle[ 3646] = 1'b0;  addr_rom[ 3646]='h00000a40;  wr_data_rom[ 3646]='h00000000;
    rd_cycle[ 3647] = 1'b0;  wr_cycle[ 3647] = 1'b1;  addr_rom[ 3647]='h000003b8;  wr_data_rom[ 3647]='h00000289;
    rd_cycle[ 3648] = 1'b1;  wr_cycle[ 3648] = 1'b0;  addr_rom[ 3648]='h00000354;  wr_data_rom[ 3648]='h00000000;
    rd_cycle[ 3649] = 1'b0;  wr_cycle[ 3649] = 1'b1;  addr_rom[ 3649]='h00000b90;  wr_data_rom[ 3649]='h00000f10;
    rd_cycle[ 3650] = 1'b0;  wr_cycle[ 3650] = 1'b1;  addr_rom[ 3650]='h00000f40;  wr_data_rom[ 3650]='h00000bcd;
    rd_cycle[ 3651] = 1'b1;  wr_cycle[ 3651] = 1'b0;  addr_rom[ 3651]='h00000b68;  wr_data_rom[ 3651]='h00000000;
    rd_cycle[ 3652] = 1'b0;  wr_cycle[ 3652] = 1'b1;  addr_rom[ 3652]='h00000858;  wr_data_rom[ 3652]='h000001e7;
    rd_cycle[ 3653] = 1'b1;  wr_cycle[ 3653] = 1'b0;  addr_rom[ 3653]='h00000384;  wr_data_rom[ 3653]='h00000000;
    rd_cycle[ 3654] = 1'b1;  wr_cycle[ 3654] = 1'b0;  addr_rom[ 3654]='h0000069c;  wr_data_rom[ 3654]='h00000000;
    rd_cycle[ 3655] = 1'b1;  wr_cycle[ 3655] = 1'b0;  addr_rom[ 3655]='h00000994;  wr_data_rom[ 3655]='h00000000;
    rd_cycle[ 3656] = 1'b1;  wr_cycle[ 3656] = 1'b0;  addr_rom[ 3656]='h000000f4;  wr_data_rom[ 3656]='h00000000;
    rd_cycle[ 3657] = 1'b1;  wr_cycle[ 3657] = 1'b0;  addr_rom[ 3657]='h000004b8;  wr_data_rom[ 3657]='h00000000;
    rd_cycle[ 3658] = 1'b1;  wr_cycle[ 3658] = 1'b0;  addr_rom[ 3658]='h00000b00;  wr_data_rom[ 3658]='h00000000;
    rd_cycle[ 3659] = 1'b1;  wr_cycle[ 3659] = 1'b0;  addr_rom[ 3659]='h000001f4;  wr_data_rom[ 3659]='h00000000;
    rd_cycle[ 3660] = 1'b1;  wr_cycle[ 3660] = 1'b0;  addr_rom[ 3660]='h00000a50;  wr_data_rom[ 3660]='h00000000;
    rd_cycle[ 3661] = 1'b0;  wr_cycle[ 3661] = 1'b1;  addr_rom[ 3661]='h00000b4c;  wr_data_rom[ 3661]='h00000cea;
    rd_cycle[ 3662] = 1'b0;  wr_cycle[ 3662] = 1'b1;  addr_rom[ 3662]='h000000f8;  wr_data_rom[ 3662]='h0000086d;
    rd_cycle[ 3663] = 1'b1;  wr_cycle[ 3663] = 1'b0;  addr_rom[ 3663]='h00000924;  wr_data_rom[ 3663]='h00000000;
    rd_cycle[ 3664] = 1'b0;  wr_cycle[ 3664] = 1'b1;  addr_rom[ 3664]='h00000288;  wr_data_rom[ 3664]='h0000094c;
    rd_cycle[ 3665] = 1'b1;  wr_cycle[ 3665] = 1'b0;  addr_rom[ 3665]='h00000518;  wr_data_rom[ 3665]='h00000000;
    rd_cycle[ 3666] = 1'b0;  wr_cycle[ 3666] = 1'b1;  addr_rom[ 3666]='h000009ac;  wr_data_rom[ 3666]='h00000c15;
    rd_cycle[ 3667] = 1'b1;  wr_cycle[ 3667] = 1'b0;  addr_rom[ 3667]='h000008bc;  wr_data_rom[ 3667]='h00000000;
    rd_cycle[ 3668] = 1'b0;  wr_cycle[ 3668] = 1'b1;  addr_rom[ 3668]='h000008d0;  wr_data_rom[ 3668]='h0000027b;
    rd_cycle[ 3669] = 1'b1;  wr_cycle[ 3669] = 1'b0;  addr_rom[ 3669]='h00000d9c;  wr_data_rom[ 3669]='h00000000;
    rd_cycle[ 3670] = 1'b0;  wr_cycle[ 3670] = 1'b1;  addr_rom[ 3670]='h00000250;  wr_data_rom[ 3670]='h000007e0;
    rd_cycle[ 3671] = 1'b1;  wr_cycle[ 3671] = 1'b0;  addr_rom[ 3671]='h0000002c;  wr_data_rom[ 3671]='h00000000;
    rd_cycle[ 3672] = 1'b1;  wr_cycle[ 3672] = 1'b0;  addr_rom[ 3672]='h000002f4;  wr_data_rom[ 3672]='h00000000;
    rd_cycle[ 3673] = 1'b0;  wr_cycle[ 3673] = 1'b1;  addr_rom[ 3673]='h000003e8;  wr_data_rom[ 3673]='h00000660;
    rd_cycle[ 3674] = 1'b1;  wr_cycle[ 3674] = 1'b0;  addr_rom[ 3674]='h000001f8;  wr_data_rom[ 3674]='h00000000;
    rd_cycle[ 3675] = 1'b1;  wr_cycle[ 3675] = 1'b0;  addr_rom[ 3675]='h00000258;  wr_data_rom[ 3675]='h00000000;
    rd_cycle[ 3676] = 1'b1;  wr_cycle[ 3676] = 1'b0;  addr_rom[ 3676]='h0000078c;  wr_data_rom[ 3676]='h00000000;
    rd_cycle[ 3677] = 1'b1;  wr_cycle[ 3677] = 1'b0;  addr_rom[ 3677]='h000004a0;  wr_data_rom[ 3677]='h00000000;
    rd_cycle[ 3678] = 1'b1;  wr_cycle[ 3678] = 1'b0;  addr_rom[ 3678]='h00000d30;  wr_data_rom[ 3678]='h00000000;
    rd_cycle[ 3679] = 1'b0;  wr_cycle[ 3679] = 1'b1;  addr_rom[ 3679]='h00000180;  wr_data_rom[ 3679]='h000001c8;
    rd_cycle[ 3680] = 1'b1;  wr_cycle[ 3680] = 1'b0;  addr_rom[ 3680]='h00000914;  wr_data_rom[ 3680]='h00000000;
    rd_cycle[ 3681] = 1'b0;  wr_cycle[ 3681] = 1'b1;  addr_rom[ 3681]='h00000a3c;  wr_data_rom[ 3681]='h00000a79;
    rd_cycle[ 3682] = 1'b0;  wr_cycle[ 3682] = 1'b1;  addr_rom[ 3682]='h00000cf4;  wr_data_rom[ 3682]='h00000415;
    rd_cycle[ 3683] = 1'b1;  wr_cycle[ 3683] = 1'b0;  addr_rom[ 3683]='h00000008;  wr_data_rom[ 3683]='h00000000;
    rd_cycle[ 3684] = 1'b0;  wr_cycle[ 3684] = 1'b1;  addr_rom[ 3684]='h00000508;  wr_data_rom[ 3684]='h0000025f;
    rd_cycle[ 3685] = 1'b1;  wr_cycle[ 3685] = 1'b0;  addr_rom[ 3685]='h00000da4;  wr_data_rom[ 3685]='h00000000;
    rd_cycle[ 3686] = 1'b1;  wr_cycle[ 3686] = 1'b0;  addr_rom[ 3686]='h000007bc;  wr_data_rom[ 3686]='h00000000;
    rd_cycle[ 3687] = 1'b1;  wr_cycle[ 3687] = 1'b0;  addr_rom[ 3687]='h00000e74;  wr_data_rom[ 3687]='h00000000;
    rd_cycle[ 3688] = 1'b1;  wr_cycle[ 3688] = 1'b0;  addr_rom[ 3688]='h000002a4;  wr_data_rom[ 3688]='h00000000;
    rd_cycle[ 3689] = 1'b1;  wr_cycle[ 3689] = 1'b0;  addr_rom[ 3689]='h00000350;  wr_data_rom[ 3689]='h00000000;
    rd_cycle[ 3690] = 1'b0;  wr_cycle[ 3690] = 1'b1;  addr_rom[ 3690]='h00000f30;  wr_data_rom[ 3690]='h0000073e;
    rd_cycle[ 3691] = 1'b1;  wr_cycle[ 3691] = 1'b0;  addr_rom[ 3691]='h00000f48;  wr_data_rom[ 3691]='h00000000;
    rd_cycle[ 3692] = 1'b0;  wr_cycle[ 3692] = 1'b1;  addr_rom[ 3692]='h0000096c;  wr_data_rom[ 3692]='h0000032d;
    rd_cycle[ 3693] = 1'b1;  wr_cycle[ 3693] = 1'b0;  addr_rom[ 3693]='h0000050c;  wr_data_rom[ 3693]='h00000000;
    rd_cycle[ 3694] = 1'b0;  wr_cycle[ 3694] = 1'b1;  addr_rom[ 3694]='h0000008c;  wr_data_rom[ 3694]='h00000c68;
    rd_cycle[ 3695] = 1'b0;  wr_cycle[ 3695] = 1'b1;  addr_rom[ 3695]='h00000f00;  wr_data_rom[ 3695]='h000009a6;
    rd_cycle[ 3696] = 1'b0;  wr_cycle[ 3696] = 1'b1;  addr_rom[ 3696]='h0000067c;  wr_data_rom[ 3696]='h00000a3c;
    rd_cycle[ 3697] = 1'b1;  wr_cycle[ 3697] = 1'b0;  addr_rom[ 3697]='h0000044c;  wr_data_rom[ 3697]='h00000000;
    rd_cycle[ 3698] = 1'b0;  wr_cycle[ 3698] = 1'b1;  addr_rom[ 3698]='h0000011c;  wr_data_rom[ 3698]='h00000e4b;
    rd_cycle[ 3699] = 1'b0;  wr_cycle[ 3699] = 1'b1;  addr_rom[ 3699]='h00000ed4;  wr_data_rom[ 3699]='h000005a1;
    rd_cycle[ 3700] = 1'b0;  wr_cycle[ 3700] = 1'b1;  addr_rom[ 3700]='h00000aa8;  wr_data_rom[ 3700]='h00000383;
    rd_cycle[ 3701] = 1'b0;  wr_cycle[ 3701] = 1'b1;  addr_rom[ 3701]='h000003d8;  wr_data_rom[ 3701]='h00000e76;
    rd_cycle[ 3702] = 1'b1;  wr_cycle[ 3702] = 1'b0;  addr_rom[ 3702]='h00000ac4;  wr_data_rom[ 3702]='h00000000;
    rd_cycle[ 3703] = 1'b0;  wr_cycle[ 3703] = 1'b1;  addr_rom[ 3703]='h00000954;  wr_data_rom[ 3703]='h0000075c;
    rd_cycle[ 3704] = 1'b1;  wr_cycle[ 3704] = 1'b0;  addr_rom[ 3704]='h00000260;  wr_data_rom[ 3704]='h00000000;
    rd_cycle[ 3705] = 1'b0;  wr_cycle[ 3705] = 1'b1;  addr_rom[ 3705]='h00000aec;  wr_data_rom[ 3705]='h00000362;
    rd_cycle[ 3706] = 1'b0;  wr_cycle[ 3706] = 1'b1;  addr_rom[ 3706]='h00000e08;  wr_data_rom[ 3706]='h000002f5;
    rd_cycle[ 3707] = 1'b1;  wr_cycle[ 3707] = 1'b0;  addr_rom[ 3707]='h00000c5c;  wr_data_rom[ 3707]='h00000000;
    rd_cycle[ 3708] = 1'b1;  wr_cycle[ 3708] = 1'b0;  addr_rom[ 3708]='h00000e44;  wr_data_rom[ 3708]='h00000000;
    rd_cycle[ 3709] = 1'b1;  wr_cycle[ 3709] = 1'b0;  addr_rom[ 3709]='h000005d0;  wr_data_rom[ 3709]='h00000000;
    rd_cycle[ 3710] = 1'b0;  wr_cycle[ 3710] = 1'b1;  addr_rom[ 3710]='h00000ea4;  wr_data_rom[ 3710]='h00000ba0;
    rd_cycle[ 3711] = 1'b1;  wr_cycle[ 3711] = 1'b0;  addr_rom[ 3711]='h00000dfc;  wr_data_rom[ 3711]='h00000000;
    rd_cycle[ 3712] = 1'b1;  wr_cycle[ 3712] = 1'b0;  addr_rom[ 3712]='h00000464;  wr_data_rom[ 3712]='h00000000;
    rd_cycle[ 3713] = 1'b0;  wr_cycle[ 3713] = 1'b1;  addr_rom[ 3713]='h0000089c;  wr_data_rom[ 3713]='h000001e5;
    rd_cycle[ 3714] = 1'b1;  wr_cycle[ 3714] = 1'b0;  addr_rom[ 3714]='h00000e0c;  wr_data_rom[ 3714]='h00000000;
    rd_cycle[ 3715] = 1'b0;  wr_cycle[ 3715] = 1'b1;  addr_rom[ 3715]='h0000051c;  wr_data_rom[ 3715]='h00000663;
    rd_cycle[ 3716] = 1'b1;  wr_cycle[ 3716] = 1'b0;  addr_rom[ 3716]='h000003b0;  wr_data_rom[ 3716]='h00000000;
    rd_cycle[ 3717] = 1'b1;  wr_cycle[ 3717] = 1'b0;  addr_rom[ 3717]='h00000c48;  wr_data_rom[ 3717]='h00000000;
    rd_cycle[ 3718] = 1'b1;  wr_cycle[ 3718] = 1'b0;  addr_rom[ 3718]='h00000500;  wr_data_rom[ 3718]='h00000000;
    rd_cycle[ 3719] = 1'b1;  wr_cycle[ 3719] = 1'b0;  addr_rom[ 3719]='h000004c4;  wr_data_rom[ 3719]='h00000000;
    rd_cycle[ 3720] = 1'b0;  wr_cycle[ 3720] = 1'b1;  addr_rom[ 3720]='h00000578;  wr_data_rom[ 3720]='h00000bfb;
    rd_cycle[ 3721] = 1'b0;  wr_cycle[ 3721] = 1'b1;  addr_rom[ 3721]='h00000940;  wr_data_rom[ 3721]='h00000c28;
    rd_cycle[ 3722] = 1'b0;  wr_cycle[ 3722] = 1'b1;  addr_rom[ 3722]='h000009fc;  wr_data_rom[ 3722]='h00000751;
    rd_cycle[ 3723] = 1'b0;  wr_cycle[ 3723] = 1'b1;  addr_rom[ 3723]='h00000b80;  wr_data_rom[ 3723]='h00000ed1;
    rd_cycle[ 3724] = 1'b1;  wr_cycle[ 3724] = 1'b0;  addr_rom[ 3724]='h00000120;  wr_data_rom[ 3724]='h00000000;
    rd_cycle[ 3725] = 1'b1;  wr_cycle[ 3725] = 1'b0;  addr_rom[ 3725]='h000008f0;  wr_data_rom[ 3725]='h00000000;
    rd_cycle[ 3726] = 1'b0;  wr_cycle[ 3726] = 1'b1;  addr_rom[ 3726]='h00000f30;  wr_data_rom[ 3726]='h00000e92;
    rd_cycle[ 3727] = 1'b1;  wr_cycle[ 3727] = 1'b0;  addr_rom[ 3727]='h00000ce8;  wr_data_rom[ 3727]='h00000000;
    rd_cycle[ 3728] = 1'b0;  wr_cycle[ 3728] = 1'b1;  addr_rom[ 3728]='h00000310;  wr_data_rom[ 3728]='h00000b94;
    rd_cycle[ 3729] = 1'b0;  wr_cycle[ 3729] = 1'b1;  addr_rom[ 3729]='h000005a4;  wr_data_rom[ 3729]='h00000b1d;
    rd_cycle[ 3730] = 1'b0;  wr_cycle[ 3730] = 1'b1;  addr_rom[ 3730]='h00000c6c;  wr_data_rom[ 3730]='h00000cc9;
    rd_cycle[ 3731] = 1'b1;  wr_cycle[ 3731] = 1'b0;  addr_rom[ 3731]='h00000c7c;  wr_data_rom[ 3731]='h00000000;
    rd_cycle[ 3732] = 1'b1;  wr_cycle[ 3732] = 1'b0;  addr_rom[ 3732]='h000009a4;  wr_data_rom[ 3732]='h00000000;
    rd_cycle[ 3733] = 1'b1;  wr_cycle[ 3733] = 1'b0;  addr_rom[ 3733]='h0000024c;  wr_data_rom[ 3733]='h00000000;
    rd_cycle[ 3734] = 1'b1;  wr_cycle[ 3734] = 1'b0;  addr_rom[ 3734]='h00000620;  wr_data_rom[ 3734]='h00000000;
    rd_cycle[ 3735] = 1'b1;  wr_cycle[ 3735] = 1'b0;  addr_rom[ 3735]='h00000768;  wr_data_rom[ 3735]='h00000000;
    rd_cycle[ 3736] = 1'b1;  wr_cycle[ 3736] = 1'b0;  addr_rom[ 3736]='h00000b58;  wr_data_rom[ 3736]='h00000000;
    rd_cycle[ 3737] = 1'b0;  wr_cycle[ 3737] = 1'b1;  addr_rom[ 3737]='h00000f0c;  wr_data_rom[ 3737]='h00000ace;
    rd_cycle[ 3738] = 1'b0;  wr_cycle[ 3738] = 1'b1;  addr_rom[ 3738]='h00000398;  wr_data_rom[ 3738]='h00000236;
    rd_cycle[ 3739] = 1'b1;  wr_cycle[ 3739] = 1'b0;  addr_rom[ 3739]='h00000314;  wr_data_rom[ 3739]='h00000000;
    rd_cycle[ 3740] = 1'b0;  wr_cycle[ 3740] = 1'b1;  addr_rom[ 3740]='h00000244;  wr_data_rom[ 3740]='h0000085d;
    rd_cycle[ 3741] = 1'b0;  wr_cycle[ 3741] = 1'b1;  addr_rom[ 3741]='h00000264;  wr_data_rom[ 3741]='h00000e05;
    rd_cycle[ 3742] = 1'b0;  wr_cycle[ 3742] = 1'b1;  addr_rom[ 3742]='h00000918;  wr_data_rom[ 3742]='h00000dcb;
    rd_cycle[ 3743] = 1'b1;  wr_cycle[ 3743] = 1'b0;  addr_rom[ 3743]='h00000e80;  wr_data_rom[ 3743]='h00000000;
    rd_cycle[ 3744] = 1'b1;  wr_cycle[ 3744] = 1'b0;  addr_rom[ 3744]='h00000d18;  wr_data_rom[ 3744]='h00000000;
    rd_cycle[ 3745] = 1'b0;  wr_cycle[ 3745] = 1'b1;  addr_rom[ 3745]='h00000d18;  wr_data_rom[ 3745]='h00000f52;
    rd_cycle[ 3746] = 1'b0;  wr_cycle[ 3746] = 1'b1;  addr_rom[ 3746]='h00000b80;  wr_data_rom[ 3746]='h00000dc3;
    rd_cycle[ 3747] = 1'b1;  wr_cycle[ 3747] = 1'b0;  addr_rom[ 3747]='h00000e44;  wr_data_rom[ 3747]='h00000000;
    rd_cycle[ 3748] = 1'b0;  wr_cycle[ 3748] = 1'b1;  addr_rom[ 3748]='h00000ae4;  wr_data_rom[ 3748]='h00000074;
    rd_cycle[ 3749] = 1'b0;  wr_cycle[ 3749] = 1'b1;  addr_rom[ 3749]='h000005ac;  wr_data_rom[ 3749]='h00000677;
    rd_cycle[ 3750] = 1'b0;  wr_cycle[ 3750] = 1'b1;  addr_rom[ 3750]='h0000016c;  wr_data_rom[ 3750]='h00000358;
    rd_cycle[ 3751] = 1'b1;  wr_cycle[ 3751] = 1'b0;  addr_rom[ 3751]='h00000ad0;  wr_data_rom[ 3751]='h00000000;
    rd_cycle[ 3752] = 1'b0;  wr_cycle[ 3752] = 1'b1;  addr_rom[ 3752]='h000006d0;  wr_data_rom[ 3752]='h00000e0d;
    rd_cycle[ 3753] = 1'b0;  wr_cycle[ 3753] = 1'b1;  addr_rom[ 3753]='h00000454;  wr_data_rom[ 3753]='h000001e2;
    rd_cycle[ 3754] = 1'b1;  wr_cycle[ 3754] = 1'b0;  addr_rom[ 3754]='h00000ec0;  wr_data_rom[ 3754]='h00000000;
    rd_cycle[ 3755] = 1'b0;  wr_cycle[ 3755] = 1'b1;  addr_rom[ 3755]='h00000348;  wr_data_rom[ 3755]='h00000992;
    rd_cycle[ 3756] = 1'b0;  wr_cycle[ 3756] = 1'b1;  addr_rom[ 3756]='h00000470;  wr_data_rom[ 3756]='h000000c0;
    rd_cycle[ 3757] = 1'b1;  wr_cycle[ 3757] = 1'b0;  addr_rom[ 3757]='h000001c4;  wr_data_rom[ 3757]='h00000000;
    rd_cycle[ 3758] = 1'b0;  wr_cycle[ 3758] = 1'b1;  addr_rom[ 3758]='h00000a38;  wr_data_rom[ 3758]='h00000870;
    rd_cycle[ 3759] = 1'b0;  wr_cycle[ 3759] = 1'b1;  addr_rom[ 3759]='h000001a4;  wr_data_rom[ 3759]='h00000f3a;
    rd_cycle[ 3760] = 1'b1;  wr_cycle[ 3760] = 1'b0;  addr_rom[ 3760]='h000007a8;  wr_data_rom[ 3760]='h00000000;
    rd_cycle[ 3761] = 1'b1;  wr_cycle[ 3761] = 1'b0;  addr_rom[ 3761]='h0000017c;  wr_data_rom[ 3761]='h00000000;
    rd_cycle[ 3762] = 1'b0;  wr_cycle[ 3762] = 1'b1;  addr_rom[ 3762]='h0000051c;  wr_data_rom[ 3762]='h000000c9;
    rd_cycle[ 3763] = 1'b0;  wr_cycle[ 3763] = 1'b1;  addr_rom[ 3763]='h00000e08;  wr_data_rom[ 3763]='h000007f4;
    rd_cycle[ 3764] = 1'b0;  wr_cycle[ 3764] = 1'b1;  addr_rom[ 3764]='h00000904;  wr_data_rom[ 3764]='h00000461;
    rd_cycle[ 3765] = 1'b1;  wr_cycle[ 3765] = 1'b0;  addr_rom[ 3765]='h00000d08;  wr_data_rom[ 3765]='h00000000;
    rd_cycle[ 3766] = 1'b1;  wr_cycle[ 3766] = 1'b0;  addr_rom[ 3766]='h00000108;  wr_data_rom[ 3766]='h00000000;
    rd_cycle[ 3767] = 1'b1;  wr_cycle[ 3767] = 1'b0;  addr_rom[ 3767]='h00000e20;  wr_data_rom[ 3767]='h00000000;
    rd_cycle[ 3768] = 1'b1;  wr_cycle[ 3768] = 1'b0;  addr_rom[ 3768]='h00000c9c;  wr_data_rom[ 3768]='h00000000;
    rd_cycle[ 3769] = 1'b0;  wr_cycle[ 3769] = 1'b1;  addr_rom[ 3769]='h000006c0;  wr_data_rom[ 3769]='h0000070c;
    rd_cycle[ 3770] = 1'b0;  wr_cycle[ 3770] = 1'b1;  addr_rom[ 3770]='h00000ae8;  wr_data_rom[ 3770]='h00000cb4;
    rd_cycle[ 3771] = 1'b0;  wr_cycle[ 3771] = 1'b1;  addr_rom[ 3771]='h00000ec0;  wr_data_rom[ 3771]='h0000052e;
    rd_cycle[ 3772] = 1'b0;  wr_cycle[ 3772] = 1'b1;  addr_rom[ 3772]='h000007e0;  wr_data_rom[ 3772]='h000007c8;
    rd_cycle[ 3773] = 1'b1;  wr_cycle[ 3773] = 1'b0;  addr_rom[ 3773]='h00000a38;  wr_data_rom[ 3773]='h00000000;
    rd_cycle[ 3774] = 1'b0;  wr_cycle[ 3774] = 1'b1;  addr_rom[ 3774]='h00000420;  wr_data_rom[ 3774]='h0000031c;
    rd_cycle[ 3775] = 1'b0;  wr_cycle[ 3775] = 1'b1;  addr_rom[ 3775]='h00000670;  wr_data_rom[ 3775]='h00000cf8;
    rd_cycle[ 3776] = 1'b0;  wr_cycle[ 3776] = 1'b1;  addr_rom[ 3776]='h00000da0;  wr_data_rom[ 3776]='h000005a6;
    rd_cycle[ 3777] = 1'b1;  wr_cycle[ 3777] = 1'b0;  addr_rom[ 3777]='h00000d48;  wr_data_rom[ 3777]='h00000000;
    rd_cycle[ 3778] = 1'b1;  wr_cycle[ 3778] = 1'b0;  addr_rom[ 3778]='h000005c0;  wr_data_rom[ 3778]='h00000000;
    rd_cycle[ 3779] = 1'b1;  wr_cycle[ 3779] = 1'b0;  addr_rom[ 3779]='h00000440;  wr_data_rom[ 3779]='h00000000;
    rd_cycle[ 3780] = 1'b1;  wr_cycle[ 3780] = 1'b0;  addr_rom[ 3780]='h00000780;  wr_data_rom[ 3780]='h00000000;
    rd_cycle[ 3781] = 1'b0;  wr_cycle[ 3781] = 1'b1;  addr_rom[ 3781]='h00000690;  wr_data_rom[ 3781]='h0000083c;
    rd_cycle[ 3782] = 1'b0;  wr_cycle[ 3782] = 1'b1;  addr_rom[ 3782]='h00000b70;  wr_data_rom[ 3782]='h00000137;
    rd_cycle[ 3783] = 1'b1;  wr_cycle[ 3783] = 1'b0;  addr_rom[ 3783]='h000003bc;  wr_data_rom[ 3783]='h00000000;
    rd_cycle[ 3784] = 1'b1;  wr_cycle[ 3784] = 1'b0;  addr_rom[ 3784]='h00000d1c;  wr_data_rom[ 3784]='h00000000;
    rd_cycle[ 3785] = 1'b0;  wr_cycle[ 3785] = 1'b1;  addr_rom[ 3785]='h00000d14;  wr_data_rom[ 3785]='h0000072c;
    rd_cycle[ 3786] = 1'b1;  wr_cycle[ 3786] = 1'b0;  addr_rom[ 3786]='h00000768;  wr_data_rom[ 3786]='h00000000;
    rd_cycle[ 3787] = 1'b0;  wr_cycle[ 3787] = 1'b1;  addr_rom[ 3787]='h000003e4;  wr_data_rom[ 3787]='h00000d46;
    rd_cycle[ 3788] = 1'b1;  wr_cycle[ 3788] = 1'b0;  addr_rom[ 3788]='h00000234;  wr_data_rom[ 3788]='h00000000;
    rd_cycle[ 3789] = 1'b1;  wr_cycle[ 3789] = 1'b0;  addr_rom[ 3789]='h00000a2c;  wr_data_rom[ 3789]='h00000000;
    rd_cycle[ 3790] = 1'b0;  wr_cycle[ 3790] = 1'b1;  addr_rom[ 3790]='h00000ab4;  wr_data_rom[ 3790]='h0000077f;
    rd_cycle[ 3791] = 1'b0;  wr_cycle[ 3791] = 1'b1;  addr_rom[ 3791]='h00000608;  wr_data_rom[ 3791]='h000008e8;
    rd_cycle[ 3792] = 1'b0;  wr_cycle[ 3792] = 1'b1;  addr_rom[ 3792]='h00000964;  wr_data_rom[ 3792]='h0000057a;
    rd_cycle[ 3793] = 1'b0;  wr_cycle[ 3793] = 1'b1;  addr_rom[ 3793]='h0000075c;  wr_data_rom[ 3793]='h00000f1d;
    rd_cycle[ 3794] = 1'b0;  wr_cycle[ 3794] = 1'b1;  addr_rom[ 3794]='h000007b4;  wr_data_rom[ 3794]='h000001c2;
    rd_cycle[ 3795] = 1'b0;  wr_cycle[ 3795] = 1'b1;  addr_rom[ 3795]='h0000097c;  wr_data_rom[ 3795]='h00000bab;
    rd_cycle[ 3796] = 1'b1;  wr_cycle[ 3796] = 1'b0;  addr_rom[ 3796]='h00000c64;  wr_data_rom[ 3796]='h00000000;
    rd_cycle[ 3797] = 1'b1;  wr_cycle[ 3797] = 1'b0;  addr_rom[ 3797]='h00000adc;  wr_data_rom[ 3797]='h00000000;
    rd_cycle[ 3798] = 1'b0;  wr_cycle[ 3798] = 1'b1;  addr_rom[ 3798]='h00000e74;  wr_data_rom[ 3798]='h00000bb3;
    rd_cycle[ 3799] = 1'b0;  wr_cycle[ 3799] = 1'b1;  addr_rom[ 3799]='h0000035c;  wr_data_rom[ 3799]='h000003c4;
    rd_cycle[ 3800] = 1'b0;  wr_cycle[ 3800] = 1'b1;  addr_rom[ 3800]='h00000c10;  wr_data_rom[ 3800]='h00000f60;
    rd_cycle[ 3801] = 1'b0;  wr_cycle[ 3801] = 1'b1;  addr_rom[ 3801]='h000006bc;  wr_data_rom[ 3801]='h00000d81;
    rd_cycle[ 3802] = 1'b1;  wr_cycle[ 3802] = 1'b0;  addr_rom[ 3802]='h0000092c;  wr_data_rom[ 3802]='h00000000;
    rd_cycle[ 3803] = 1'b0;  wr_cycle[ 3803] = 1'b1;  addr_rom[ 3803]='h000003f4;  wr_data_rom[ 3803]='h0000006f;
    rd_cycle[ 3804] = 1'b0;  wr_cycle[ 3804] = 1'b1;  addr_rom[ 3804]='h00000ca8;  wr_data_rom[ 3804]='h00000dd1;
    rd_cycle[ 3805] = 1'b0;  wr_cycle[ 3805] = 1'b1;  addr_rom[ 3805]='h000005c0;  wr_data_rom[ 3805]='h00000cb8;
    rd_cycle[ 3806] = 1'b1;  wr_cycle[ 3806] = 1'b0;  addr_rom[ 3806]='h00000ca8;  wr_data_rom[ 3806]='h00000000;
    rd_cycle[ 3807] = 1'b1;  wr_cycle[ 3807] = 1'b0;  addr_rom[ 3807]='h0000017c;  wr_data_rom[ 3807]='h00000000;
    rd_cycle[ 3808] = 1'b0;  wr_cycle[ 3808] = 1'b1;  addr_rom[ 3808]='h0000093c;  wr_data_rom[ 3808]='h000007f5;
    rd_cycle[ 3809] = 1'b0;  wr_cycle[ 3809] = 1'b1;  addr_rom[ 3809]='h000003e4;  wr_data_rom[ 3809]='h00000097;
    rd_cycle[ 3810] = 1'b0;  wr_cycle[ 3810] = 1'b1;  addr_rom[ 3810]='h00000dd8;  wr_data_rom[ 3810]='h00000eef;
    rd_cycle[ 3811] = 1'b1;  wr_cycle[ 3811] = 1'b0;  addr_rom[ 3811]='h00000638;  wr_data_rom[ 3811]='h00000000;
    rd_cycle[ 3812] = 1'b0;  wr_cycle[ 3812] = 1'b1;  addr_rom[ 3812]='h0000046c;  wr_data_rom[ 3812]='h00000549;
    rd_cycle[ 3813] = 1'b1;  wr_cycle[ 3813] = 1'b0;  addr_rom[ 3813]='h00000b78;  wr_data_rom[ 3813]='h00000000;
    rd_cycle[ 3814] = 1'b1;  wr_cycle[ 3814] = 1'b0;  addr_rom[ 3814]='h00000c08;  wr_data_rom[ 3814]='h00000000;
    rd_cycle[ 3815] = 1'b1;  wr_cycle[ 3815] = 1'b0;  addr_rom[ 3815]='h00000564;  wr_data_rom[ 3815]='h00000000;
    rd_cycle[ 3816] = 1'b0;  wr_cycle[ 3816] = 1'b1;  addr_rom[ 3816]='h00000a4c;  wr_data_rom[ 3816]='h000001a5;
    rd_cycle[ 3817] = 1'b1;  wr_cycle[ 3817] = 1'b0;  addr_rom[ 3817]='h00000d24;  wr_data_rom[ 3817]='h00000000;
    rd_cycle[ 3818] = 1'b1;  wr_cycle[ 3818] = 1'b0;  addr_rom[ 3818]='h00000298;  wr_data_rom[ 3818]='h00000000;
    rd_cycle[ 3819] = 1'b0;  wr_cycle[ 3819] = 1'b1;  addr_rom[ 3819]='h00000b88;  wr_data_rom[ 3819]='h00000563;
    rd_cycle[ 3820] = 1'b1;  wr_cycle[ 3820] = 1'b0;  addr_rom[ 3820]='h000003a4;  wr_data_rom[ 3820]='h00000000;
    rd_cycle[ 3821] = 1'b0;  wr_cycle[ 3821] = 1'b1;  addr_rom[ 3821]='h000006fc;  wr_data_rom[ 3821]='h00000011;
    rd_cycle[ 3822] = 1'b0;  wr_cycle[ 3822] = 1'b1;  addr_rom[ 3822]='h00000a90;  wr_data_rom[ 3822]='h00000ee5;
    rd_cycle[ 3823] = 1'b1;  wr_cycle[ 3823] = 1'b0;  addr_rom[ 3823]='h000009d8;  wr_data_rom[ 3823]='h00000000;
    rd_cycle[ 3824] = 1'b1;  wr_cycle[ 3824] = 1'b0;  addr_rom[ 3824]='h00000d2c;  wr_data_rom[ 3824]='h00000000;
    rd_cycle[ 3825] = 1'b0;  wr_cycle[ 3825] = 1'b1;  addr_rom[ 3825]='h00000ac4;  wr_data_rom[ 3825]='h00000b04;
    rd_cycle[ 3826] = 1'b1;  wr_cycle[ 3826] = 1'b0;  addr_rom[ 3826]='h00000320;  wr_data_rom[ 3826]='h00000000;
    rd_cycle[ 3827] = 1'b0;  wr_cycle[ 3827] = 1'b1;  addr_rom[ 3827]='h00000640;  wr_data_rom[ 3827]='h000005d7;
    rd_cycle[ 3828] = 1'b1;  wr_cycle[ 3828] = 1'b0;  addr_rom[ 3828]='h00000ab8;  wr_data_rom[ 3828]='h00000000;
    rd_cycle[ 3829] = 1'b1;  wr_cycle[ 3829] = 1'b0;  addr_rom[ 3829]='h00000784;  wr_data_rom[ 3829]='h00000000;
    rd_cycle[ 3830] = 1'b1;  wr_cycle[ 3830] = 1'b0;  addr_rom[ 3830]='h00000564;  wr_data_rom[ 3830]='h00000000;
    rd_cycle[ 3831] = 1'b1;  wr_cycle[ 3831] = 1'b0;  addr_rom[ 3831]='h000004b8;  wr_data_rom[ 3831]='h00000000;
    rd_cycle[ 3832] = 1'b1;  wr_cycle[ 3832] = 1'b0;  addr_rom[ 3832]='h00000594;  wr_data_rom[ 3832]='h00000000;
    rd_cycle[ 3833] = 1'b0;  wr_cycle[ 3833] = 1'b1;  addr_rom[ 3833]='h00000920;  wr_data_rom[ 3833]='h0000052d;
    rd_cycle[ 3834] = 1'b0;  wr_cycle[ 3834] = 1'b1;  addr_rom[ 3834]='h000003a0;  wr_data_rom[ 3834]='h000001df;
    rd_cycle[ 3835] = 1'b0;  wr_cycle[ 3835] = 1'b1;  addr_rom[ 3835]='h00000624;  wr_data_rom[ 3835]='h00000d0c;
    rd_cycle[ 3836] = 1'b1;  wr_cycle[ 3836] = 1'b0;  addr_rom[ 3836]='h00000ad4;  wr_data_rom[ 3836]='h00000000;
    rd_cycle[ 3837] = 1'b1;  wr_cycle[ 3837] = 1'b0;  addr_rom[ 3837]='h00000038;  wr_data_rom[ 3837]='h00000000;
    rd_cycle[ 3838] = 1'b0;  wr_cycle[ 3838] = 1'b1;  addr_rom[ 3838]='h00000024;  wr_data_rom[ 3838]='h00000731;
    rd_cycle[ 3839] = 1'b1;  wr_cycle[ 3839] = 1'b0;  addr_rom[ 3839]='h00000dc0;  wr_data_rom[ 3839]='h00000000;
    rd_cycle[ 3840] = 1'b1;  wr_cycle[ 3840] = 1'b0;  addr_rom[ 3840]='h000008a4;  wr_data_rom[ 3840]='h00000000;
    rd_cycle[ 3841] = 1'b1;  wr_cycle[ 3841] = 1'b0;  addr_rom[ 3841]='h00000918;  wr_data_rom[ 3841]='h00000000;
    rd_cycle[ 3842] = 1'b0;  wr_cycle[ 3842] = 1'b1;  addr_rom[ 3842]='h000003f4;  wr_data_rom[ 3842]='h0000011d;
    rd_cycle[ 3843] = 1'b1;  wr_cycle[ 3843] = 1'b0;  addr_rom[ 3843]='h000005e4;  wr_data_rom[ 3843]='h00000000;
    rd_cycle[ 3844] = 1'b1;  wr_cycle[ 3844] = 1'b0;  addr_rom[ 3844]='h00000a88;  wr_data_rom[ 3844]='h00000000;
    rd_cycle[ 3845] = 1'b1;  wr_cycle[ 3845] = 1'b0;  addr_rom[ 3845]='h00000b74;  wr_data_rom[ 3845]='h00000000;
    rd_cycle[ 3846] = 1'b1;  wr_cycle[ 3846] = 1'b0;  addr_rom[ 3846]='h00000f54;  wr_data_rom[ 3846]='h00000000;
    rd_cycle[ 3847] = 1'b1;  wr_cycle[ 3847] = 1'b0;  addr_rom[ 3847]='h000002b0;  wr_data_rom[ 3847]='h00000000;
    rd_cycle[ 3848] = 1'b1;  wr_cycle[ 3848] = 1'b0;  addr_rom[ 3848]='h00000b38;  wr_data_rom[ 3848]='h00000000;
    rd_cycle[ 3849] = 1'b1;  wr_cycle[ 3849] = 1'b0;  addr_rom[ 3849]='h000005c0;  wr_data_rom[ 3849]='h00000000;
    rd_cycle[ 3850] = 1'b1;  wr_cycle[ 3850] = 1'b0;  addr_rom[ 3850]='h000009c0;  wr_data_rom[ 3850]='h00000000;
    rd_cycle[ 3851] = 1'b1;  wr_cycle[ 3851] = 1'b0;  addr_rom[ 3851]='h000001e4;  wr_data_rom[ 3851]='h00000000;
    rd_cycle[ 3852] = 1'b0;  wr_cycle[ 3852] = 1'b1;  addr_rom[ 3852]='h000007b8;  wr_data_rom[ 3852]='h00000a99;
    rd_cycle[ 3853] = 1'b1;  wr_cycle[ 3853] = 1'b0;  addr_rom[ 3853]='h00000be4;  wr_data_rom[ 3853]='h00000000;
    rd_cycle[ 3854] = 1'b0;  wr_cycle[ 3854] = 1'b1;  addr_rom[ 3854]='h0000040c;  wr_data_rom[ 3854]='h000006f8;
    rd_cycle[ 3855] = 1'b1;  wr_cycle[ 3855] = 1'b0;  addr_rom[ 3855]='h000009a4;  wr_data_rom[ 3855]='h00000000;
    rd_cycle[ 3856] = 1'b1;  wr_cycle[ 3856] = 1'b0;  addr_rom[ 3856]='h00000304;  wr_data_rom[ 3856]='h00000000;
    rd_cycle[ 3857] = 1'b0;  wr_cycle[ 3857] = 1'b1;  addr_rom[ 3857]='h00000f70;  wr_data_rom[ 3857]='h00000a23;
    rd_cycle[ 3858] = 1'b1;  wr_cycle[ 3858] = 1'b0;  addr_rom[ 3858]='h00000290;  wr_data_rom[ 3858]='h00000000;
    rd_cycle[ 3859] = 1'b1;  wr_cycle[ 3859] = 1'b0;  addr_rom[ 3859]='h00000f78;  wr_data_rom[ 3859]='h00000000;
    rd_cycle[ 3860] = 1'b0;  wr_cycle[ 3860] = 1'b1;  addr_rom[ 3860]='h00000044;  wr_data_rom[ 3860]='h00000251;
    rd_cycle[ 3861] = 1'b1;  wr_cycle[ 3861] = 1'b0;  addr_rom[ 3861]='h000001ac;  wr_data_rom[ 3861]='h00000000;
    rd_cycle[ 3862] = 1'b1;  wr_cycle[ 3862] = 1'b0;  addr_rom[ 3862]='h000004f8;  wr_data_rom[ 3862]='h00000000;
    rd_cycle[ 3863] = 1'b1;  wr_cycle[ 3863] = 1'b0;  addr_rom[ 3863]='h00000b0c;  wr_data_rom[ 3863]='h00000000;
    rd_cycle[ 3864] = 1'b0;  wr_cycle[ 3864] = 1'b1;  addr_rom[ 3864]='h00000610;  wr_data_rom[ 3864]='h00000897;
    rd_cycle[ 3865] = 1'b0;  wr_cycle[ 3865] = 1'b1;  addr_rom[ 3865]='h00000398;  wr_data_rom[ 3865]='h00000447;
    rd_cycle[ 3866] = 1'b0;  wr_cycle[ 3866] = 1'b1;  addr_rom[ 3866]='h000009d4;  wr_data_rom[ 3866]='h000008aa;
    rd_cycle[ 3867] = 1'b0;  wr_cycle[ 3867] = 1'b1;  addr_rom[ 3867]='h00000050;  wr_data_rom[ 3867]='h00000d8a;
    rd_cycle[ 3868] = 1'b1;  wr_cycle[ 3868] = 1'b0;  addr_rom[ 3868]='h000002a0;  wr_data_rom[ 3868]='h00000000;
    rd_cycle[ 3869] = 1'b0;  wr_cycle[ 3869] = 1'b1;  addr_rom[ 3869]='h000008cc;  wr_data_rom[ 3869]='h000001a9;
    rd_cycle[ 3870] = 1'b1;  wr_cycle[ 3870] = 1'b0;  addr_rom[ 3870]='h0000089c;  wr_data_rom[ 3870]='h00000000;
    rd_cycle[ 3871] = 1'b0;  wr_cycle[ 3871] = 1'b1;  addr_rom[ 3871]='h00000acc;  wr_data_rom[ 3871]='h00000f92;
    rd_cycle[ 3872] = 1'b1;  wr_cycle[ 3872] = 1'b0;  addr_rom[ 3872]='h00000cc8;  wr_data_rom[ 3872]='h00000000;
    rd_cycle[ 3873] = 1'b1;  wr_cycle[ 3873] = 1'b0;  addr_rom[ 3873]='h00000b8c;  wr_data_rom[ 3873]='h00000000;
    rd_cycle[ 3874] = 1'b0;  wr_cycle[ 3874] = 1'b1;  addr_rom[ 3874]='h00000eac;  wr_data_rom[ 3874]='h000000c1;
    rd_cycle[ 3875] = 1'b0;  wr_cycle[ 3875] = 1'b1;  addr_rom[ 3875]='h00000848;  wr_data_rom[ 3875]='h00000e8a;
    rd_cycle[ 3876] = 1'b1;  wr_cycle[ 3876] = 1'b0;  addr_rom[ 3876]='h00000d10;  wr_data_rom[ 3876]='h00000000;
    rd_cycle[ 3877] = 1'b1;  wr_cycle[ 3877] = 1'b0;  addr_rom[ 3877]='h00000468;  wr_data_rom[ 3877]='h00000000;
    rd_cycle[ 3878] = 1'b1;  wr_cycle[ 3878] = 1'b0;  addr_rom[ 3878]='h000002cc;  wr_data_rom[ 3878]='h00000000;
    rd_cycle[ 3879] = 1'b1;  wr_cycle[ 3879] = 1'b0;  addr_rom[ 3879]='h00000584;  wr_data_rom[ 3879]='h00000000;
    rd_cycle[ 3880] = 1'b1;  wr_cycle[ 3880] = 1'b0;  addr_rom[ 3880]='h00000a88;  wr_data_rom[ 3880]='h00000000;
    rd_cycle[ 3881] = 1'b0;  wr_cycle[ 3881] = 1'b1;  addr_rom[ 3881]='h000005ec;  wr_data_rom[ 3881]='h0000063e;
    rd_cycle[ 3882] = 1'b0;  wr_cycle[ 3882] = 1'b1;  addr_rom[ 3882]='h00000bf4;  wr_data_rom[ 3882]='h00000f78;
    rd_cycle[ 3883] = 1'b0;  wr_cycle[ 3883] = 1'b1;  addr_rom[ 3883]='h00000278;  wr_data_rom[ 3883]='h000003d4;
    rd_cycle[ 3884] = 1'b0;  wr_cycle[ 3884] = 1'b1;  addr_rom[ 3884]='h00000304;  wr_data_rom[ 3884]='h00000c6e;
    rd_cycle[ 3885] = 1'b0;  wr_cycle[ 3885] = 1'b1;  addr_rom[ 3885]='h00000428;  wr_data_rom[ 3885]='h00000766;
    rd_cycle[ 3886] = 1'b0;  wr_cycle[ 3886] = 1'b1;  addr_rom[ 3886]='h00000dbc;  wr_data_rom[ 3886]='h0000047c;
    rd_cycle[ 3887] = 1'b0;  wr_cycle[ 3887] = 1'b1;  addr_rom[ 3887]='h00000ac4;  wr_data_rom[ 3887]='h00000d3e;
    rd_cycle[ 3888] = 1'b0;  wr_cycle[ 3888] = 1'b1;  addr_rom[ 3888]='h00000318;  wr_data_rom[ 3888]='h00000359;
    rd_cycle[ 3889] = 1'b1;  wr_cycle[ 3889] = 1'b0;  addr_rom[ 3889]='h000000a8;  wr_data_rom[ 3889]='h00000000;
    rd_cycle[ 3890] = 1'b1;  wr_cycle[ 3890] = 1'b0;  addr_rom[ 3890]='h0000054c;  wr_data_rom[ 3890]='h00000000;
    rd_cycle[ 3891] = 1'b0;  wr_cycle[ 3891] = 1'b1;  addr_rom[ 3891]='h000004dc;  wr_data_rom[ 3891]='h00000919;
    rd_cycle[ 3892] = 1'b0;  wr_cycle[ 3892] = 1'b1;  addr_rom[ 3892]='h00000bf0;  wr_data_rom[ 3892]='h00000b7d;
    rd_cycle[ 3893] = 1'b1;  wr_cycle[ 3893] = 1'b0;  addr_rom[ 3893]='h000004a4;  wr_data_rom[ 3893]='h00000000;
    rd_cycle[ 3894] = 1'b0;  wr_cycle[ 3894] = 1'b1;  addr_rom[ 3894]='h00000534;  wr_data_rom[ 3894]='h00000bdc;
    rd_cycle[ 3895] = 1'b0;  wr_cycle[ 3895] = 1'b1;  addr_rom[ 3895]='h00000720;  wr_data_rom[ 3895]='h00000107;
    rd_cycle[ 3896] = 1'b1;  wr_cycle[ 3896] = 1'b0;  addr_rom[ 3896]='h000008d4;  wr_data_rom[ 3896]='h00000000;
    rd_cycle[ 3897] = 1'b0;  wr_cycle[ 3897] = 1'b1;  addr_rom[ 3897]='h00000ab8;  wr_data_rom[ 3897]='h00000c41;
    rd_cycle[ 3898] = 1'b0;  wr_cycle[ 3898] = 1'b1;  addr_rom[ 3898]='h000002a8;  wr_data_rom[ 3898]='h000009ce;
    rd_cycle[ 3899] = 1'b1;  wr_cycle[ 3899] = 1'b0;  addr_rom[ 3899]='h00000530;  wr_data_rom[ 3899]='h00000000;
    rd_cycle[ 3900] = 1'b0;  wr_cycle[ 3900] = 1'b1;  addr_rom[ 3900]='h00000b64;  wr_data_rom[ 3900]='h00000ce9;
    rd_cycle[ 3901] = 1'b0;  wr_cycle[ 3901] = 1'b1;  addr_rom[ 3901]='h00000698;  wr_data_rom[ 3901]='h0000098b;
    rd_cycle[ 3902] = 1'b1;  wr_cycle[ 3902] = 1'b0;  addr_rom[ 3902]='h00000bc4;  wr_data_rom[ 3902]='h00000000;
    rd_cycle[ 3903] = 1'b1;  wr_cycle[ 3903] = 1'b0;  addr_rom[ 3903]='h00000914;  wr_data_rom[ 3903]='h00000000;
    rd_cycle[ 3904] = 1'b1;  wr_cycle[ 3904] = 1'b0;  addr_rom[ 3904]='h00000854;  wr_data_rom[ 3904]='h00000000;
    rd_cycle[ 3905] = 1'b1;  wr_cycle[ 3905] = 1'b0;  addr_rom[ 3905]='h00000a9c;  wr_data_rom[ 3905]='h00000000;
    rd_cycle[ 3906] = 1'b0;  wr_cycle[ 3906] = 1'b1;  addr_rom[ 3906]='h000004e4;  wr_data_rom[ 3906]='h00000f65;
    rd_cycle[ 3907] = 1'b0;  wr_cycle[ 3907] = 1'b1;  addr_rom[ 3907]='h0000004c;  wr_data_rom[ 3907]='h00000c1e;
    rd_cycle[ 3908] = 1'b0;  wr_cycle[ 3908] = 1'b1;  addr_rom[ 3908]='h000008a0;  wr_data_rom[ 3908]='h00000970;
    rd_cycle[ 3909] = 1'b1;  wr_cycle[ 3909] = 1'b0;  addr_rom[ 3909]='h00000e74;  wr_data_rom[ 3909]='h00000000;
    rd_cycle[ 3910] = 1'b1;  wr_cycle[ 3910] = 1'b0;  addr_rom[ 3910]='h00000660;  wr_data_rom[ 3910]='h00000000;
    rd_cycle[ 3911] = 1'b1;  wr_cycle[ 3911] = 1'b0;  addr_rom[ 3911]='h000004d0;  wr_data_rom[ 3911]='h00000000;
    rd_cycle[ 3912] = 1'b0;  wr_cycle[ 3912] = 1'b1;  addr_rom[ 3912]='h00000798;  wr_data_rom[ 3912]='h00000e6b;
    rd_cycle[ 3913] = 1'b0;  wr_cycle[ 3913] = 1'b1;  addr_rom[ 3913]='h00000af4;  wr_data_rom[ 3913]='h00000c50;
    rd_cycle[ 3914] = 1'b1;  wr_cycle[ 3914] = 1'b0;  addr_rom[ 3914]='h00000494;  wr_data_rom[ 3914]='h00000000;
    rd_cycle[ 3915] = 1'b0;  wr_cycle[ 3915] = 1'b1;  addr_rom[ 3915]='h00000cd4;  wr_data_rom[ 3915]='h00000cef;
    rd_cycle[ 3916] = 1'b0;  wr_cycle[ 3916] = 1'b1;  addr_rom[ 3916]='h00000758;  wr_data_rom[ 3916]='h00000eaf;
    rd_cycle[ 3917] = 1'b0;  wr_cycle[ 3917] = 1'b1;  addr_rom[ 3917]='h00000bd4;  wr_data_rom[ 3917]='h00000f87;
    rd_cycle[ 3918] = 1'b0;  wr_cycle[ 3918] = 1'b1;  addr_rom[ 3918]='h00000d60;  wr_data_rom[ 3918]='h000008d0;
    rd_cycle[ 3919] = 1'b0;  wr_cycle[ 3919] = 1'b1;  addr_rom[ 3919]='h00000790;  wr_data_rom[ 3919]='h000003de;
    rd_cycle[ 3920] = 1'b1;  wr_cycle[ 3920] = 1'b0;  addr_rom[ 3920]='h00000dd4;  wr_data_rom[ 3920]='h00000000;
    rd_cycle[ 3921] = 1'b0;  wr_cycle[ 3921] = 1'b1;  addr_rom[ 3921]='h00000a4c;  wr_data_rom[ 3921]='h00000a23;
    rd_cycle[ 3922] = 1'b0;  wr_cycle[ 3922] = 1'b1;  addr_rom[ 3922]='h000000fc;  wr_data_rom[ 3922]='h000002c1;
    rd_cycle[ 3923] = 1'b0;  wr_cycle[ 3923] = 1'b1;  addr_rom[ 3923]='h000006cc;  wr_data_rom[ 3923]='h00000036;
    rd_cycle[ 3924] = 1'b0;  wr_cycle[ 3924] = 1'b1;  addr_rom[ 3924]='h00000d58;  wr_data_rom[ 3924]='h00000826;
    rd_cycle[ 3925] = 1'b0;  wr_cycle[ 3925] = 1'b1;  addr_rom[ 3925]='h00000064;  wr_data_rom[ 3925]='h00000f34;
    rd_cycle[ 3926] = 1'b0;  wr_cycle[ 3926] = 1'b1;  addr_rom[ 3926]='h00000300;  wr_data_rom[ 3926]='h000001d1;
    rd_cycle[ 3927] = 1'b0;  wr_cycle[ 3927] = 1'b1;  addr_rom[ 3927]='h000002c0;  wr_data_rom[ 3927]='h000009b7;
    rd_cycle[ 3928] = 1'b1;  wr_cycle[ 3928] = 1'b0;  addr_rom[ 3928]='h00000c64;  wr_data_rom[ 3928]='h00000000;
    rd_cycle[ 3929] = 1'b1;  wr_cycle[ 3929] = 1'b0;  addr_rom[ 3929]='h000006c4;  wr_data_rom[ 3929]='h00000000;
    rd_cycle[ 3930] = 1'b0;  wr_cycle[ 3930] = 1'b1;  addr_rom[ 3930]='h000009bc;  wr_data_rom[ 3930]='h00000ed3;
    rd_cycle[ 3931] = 1'b0;  wr_cycle[ 3931] = 1'b1;  addr_rom[ 3931]='h00000210;  wr_data_rom[ 3931]='h00000f81;
    rd_cycle[ 3932] = 1'b0;  wr_cycle[ 3932] = 1'b1;  addr_rom[ 3932]='h00000420;  wr_data_rom[ 3932]='h00000118;
    rd_cycle[ 3933] = 1'b0;  wr_cycle[ 3933] = 1'b1;  addr_rom[ 3933]='h000003c4;  wr_data_rom[ 3933]='h0000028d;
    rd_cycle[ 3934] = 1'b1;  wr_cycle[ 3934] = 1'b0;  addr_rom[ 3934]='h00000b40;  wr_data_rom[ 3934]='h00000000;
    rd_cycle[ 3935] = 1'b0;  wr_cycle[ 3935] = 1'b1;  addr_rom[ 3935]='h00000a18;  wr_data_rom[ 3935]='h000007db;
    rd_cycle[ 3936] = 1'b1;  wr_cycle[ 3936] = 1'b0;  addr_rom[ 3936]='h00000c8c;  wr_data_rom[ 3936]='h00000000;
    rd_cycle[ 3937] = 1'b0;  wr_cycle[ 3937] = 1'b1;  addr_rom[ 3937]='h00000008;  wr_data_rom[ 3937]='h00000221;
    rd_cycle[ 3938] = 1'b1;  wr_cycle[ 3938] = 1'b0;  addr_rom[ 3938]='h000006a8;  wr_data_rom[ 3938]='h00000000;
    rd_cycle[ 3939] = 1'b1;  wr_cycle[ 3939] = 1'b0;  addr_rom[ 3939]='h00000518;  wr_data_rom[ 3939]='h00000000;
    rd_cycle[ 3940] = 1'b0;  wr_cycle[ 3940] = 1'b1;  addr_rom[ 3940]='h00000134;  wr_data_rom[ 3940]='h000000e1;
    rd_cycle[ 3941] = 1'b0;  wr_cycle[ 3941] = 1'b1;  addr_rom[ 3941]='h0000010c;  wr_data_rom[ 3941]='h00000bbb;
    rd_cycle[ 3942] = 1'b0;  wr_cycle[ 3942] = 1'b1;  addr_rom[ 3942]='h00000724;  wr_data_rom[ 3942]='h00000598;
    rd_cycle[ 3943] = 1'b0;  wr_cycle[ 3943] = 1'b1;  addr_rom[ 3943]='h000007d4;  wr_data_rom[ 3943]='h00000264;
    rd_cycle[ 3944] = 1'b0;  wr_cycle[ 3944] = 1'b1;  addr_rom[ 3944]='h00000458;  wr_data_rom[ 3944]='h00000439;
    rd_cycle[ 3945] = 1'b1;  wr_cycle[ 3945] = 1'b0;  addr_rom[ 3945]='h00000a64;  wr_data_rom[ 3945]='h00000000;
    rd_cycle[ 3946] = 1'b1;  wr_cycle[ 3946] = 1'b0;  addr_rom[ 3946]='h00000a08;  wr_data_rom[ 3946]='h00000000;
    rd_cycle[ 3947] = 1'b1;  wr_cycle[ 3947] = 1'b0;  addr_rom[ 3947]='h00000978;  wr_data_rom[ 3947]='h00000000;
    rd_cycle[ 3948] = 1'b1;  wr_cycle[ 3948] = 1'b0;  addr_rom[ 3948]='h000004f4;  wr_data_rom[ 3948]='h00000000;
    rd_cycle[ 3949] = 1'b0;  wr_cycle[ 3949] = 1'b1;  addr_rom[ 3949]='h00000214;  wr_data_rom[ 3949]='h000000f3;
    rd_cycle[ 3950] = 1'b1;  wr_cycle[ 3950] = 1'b0;  addr_rom[ 3950]='h00000e7c;  wr_data_rom[ 3950]='h00000000;
    rd_cycle[ 3951] = 1'b0;  wr_cycle[ 3951] = 1'b1;  addr_rom[ 3951]='h00000b44;  wr_data_rom[ 3951]='h000000e4;
    rd_cycle[ 3952] = 1'b1;  wr_cycle[ 3952] = 1'b0;  addr_rom[ 3952]='h0000016c;  wr_data_rom[ 3952]='h00000000;
    rd_cycle[ 3953] = 1'b1;  wr_cycle[ 3953] = 1'b0;  addr_rom[ 3953]='h00000c50;  wr_data_rom[ 3953]='h00000000;
    rd_cycle[ 3954] = 1'b0;  wr_cycle[ 3954] = 1'b1;  addr_rom[ 3954]='h000001bc;  wr_data_rom[ 3954]='h0000028f;
    rd_cycle[ 3955] = 1'b1;  wr_cycle[ 3955] = 1'b0;  addr_rom[ 3955]='h00000bac;  wr_data_rom[ 3955]='h00000000;
    rd_cycle[ 3956] = 1'b0;  wr_cycle[ 3956] = 1'b1;  addr_rom[ 3956]='h0000048c;  wr_data_rom[ 3956]='h00000973;
    rd_cycle[ 3957] = 1'b0;  wr_cycle[ 3957] = 1'b1;  addr_rom[ 3957]='h00000f2c;  wr_data_rom[ 3957]='h0000062f;
    rd_cycle[ 3958] = 1'b1;  wr_cycle[ 3958] = 1'b0;  addr_rom[ 3958]='h00000604;  wr_data_rom[ 3958]='h00000000;
    rd_cycle[ 3959] = 1'b1;  wr_cycle[ 3959] = 1'b0;  addr_rom[ 3959]='h0000031c;  wr_data_rom[ 3959]='h00000000;
    rd_cycle[ 3960] = 1'b0;  wr_cycle[ 3960] = 1'b1;  addr_rom[ 3960]='h000007ac;  wr_data_rom[ 3960]='h00000ad1;
    rd_cycle[ 3961] = 1'b0;  wr_cycle[ 3961] = 1'b1;  addr_rom[ 3961]='h00000910;  wr_data_rom[ 3961]='h00000870;
    rd_cycle[ 3962] = 1'b1;  wr_cycle[ 3962] = 1'b0;  addr_rom[ 3962]='h00000018;  wr_data_rom[ 3962]='h00000000;
    rd_cycle[ 3963] = 1'b1;  wr_cycle[ 3963] = 1'b0;  addr_rom[ 3963]='h00000560;  wr_data_rom[ 3963]='h00000000;
    rd_cycle[ 3964] = 1'b0;  wr_cycle[ 3964] = 1'b1;  addr_rom[ 3964]='h00000b58;  wr_data_rom[ 3964]='h00000aba;
    rd_cycle[ 3965] = 1'b1;  wr_cycle[ 3965] = 1'b0;  addr_rom[ 3965]='h00000204;  wr_data_rom[ 3965]='h00000000;
    rd_cycle[ 3966] = 1'b0;  wr_cycle[ 3966] = 1'b1;  addr_rom[ 3966]='h00000ad0;  wr_data_rom[ 3966]='h000000c6;
    rd_cycle[ 3967] = 1'b0;  wr_cycle[ 3967] = 1'b1;  addr_rom[ 3967]='h00000340;  wr_data_rom[ 3967]='h000004a6;
    rd_cycle[ 3968] = 1'b0;  wr_cycle[ 3968] = 1'b1;  addr_rom[ 3968]='h00000934;  wr_data_rom[ 3968]='h00000153;
    rd_cycle[ 3969] = 1'b1;  wr_cycle[ 3969] = 1'b0;  addr_rom[ 3969]='h00000ccc;  wr_data_rom[ 3969]='h00000000;
    rd_cycle[ 3970] = 1'b0;  wr_cycle[ 3970] = 1'b1;  addr_rom[ 3970]='h000003cc;  wr_data_rom[ 3970]='h000009f2;
    rd_cycle[ 3971] = 1'b0;  wr_cycle[ 3971] = 1'b1;  addr_rom[ 3971]='h00000214;  wr_data_rom[ 3971]='h00000121;
    rd_cycle[ 3972] = 1'b1;  wr_cycle[ 3972] = 1'b0;  addr_rom[ 3972]='h00000938;  wr_data_rom[ 3972]='h00000000;
    rd_cycle[ 3973] = 1'b1;  wr_cycle[ 3973] = 1'b0;  addr_rom[ 3973]='h00000114;  wr_data_rom[ 3973]='h00000000;
    rd_cycle[ 3974] = 1'b1;  wr_cycle[ 3974] = 1'b0;  addr_rom[ 3974]='h00000668;  wr_data_rom[ 3974]='h00000000;
    rd_cycle[ 3975] = 1'b0;  wr_cycle[ 3975] = 1'b1;  addr_rom[ 3975]='h000008c4;  wr_data_rom[ 3975]='h00000708;
    rd_cycle[ 3976] = 1'b1;  wr_cycle[ 3976] = 1'b0;  addr_rom[ 3976]='h0000087c;  wr_data_rom[ 3976]='h00000000;
    rd_cycle[ 3977] = 1'b0;  wr_cycle[ 3977] = 1'b1;  addr_rom[ 3977]='h00000f74;  wr_data_rom[ 3977]='h0000099b;
    rd_cycle[ 3978] = 1'b1;  wr_cycle[ 3978] = 1'b0;  addr_rom[ 3978]='h00000dc8;  wr_data_rom[ 3978]='h00000000;
    rd_cycle[ 3979] = 1'b0;  wr_cycle[ 3979] = 1'b1;  addr_rom[ 3979]='h00000adc;  wr_data_rom[ 3979]='h00000ee7;
    rd_cycle[ 3980] = 1'b0;  wr_cycle[ 3980] = 1'b1;  addr_rom[ 3980]='h00000964;  wr_data_rom[ 3980]='h0000075c;
    rd_cycle[ 3981] = 1'b0;  wr_cycle[ 3981] = 1'b1;  addr_rom[ 3981]='h000008a8;  wr_data_rom[ 3981]='h00000dbd;
    rd_cycle[ 3982] = 1'b0;  wr_cycle[ 3982] = 1'b1;  addr_rom[ 3982]='h00000f34;  wr_data_rom[ 3982]='h00000623;
    rd_cycle[ 3983] = 1'b0;  wr_cycle[ 3983] = 1'b1;  addr_rom[ 3983]='h000007dc;  wr_data_rom[ 3983]='h00000495;
    rd_cycle[ 3984] = 1'b0;  wr_cycle[ 3984] = 1'b1;  addr_rom[ 3984]='h00000740;  wr_data_rom[ 3984]='h00000aad;
    rd_cycle[ 3985] = 1'b1;  wr_cycle[ 3985] = 1'b0;  addr_rom[ 3985]='h00000e1c;  wr_data_rom[ 3985]='h00000000;
    rd_cycle[ 3986] = 1'b1;  wr_cycle[ 3986] = 1'b0;  addr_rom[ 3986]='h00000404;  wr_data_rom[ 3986]='h00000000;
    rd_cycle[ 3987] = 1'b1;  wr_cycle[ 3987] = 1'b0;  addr_rom[ 3987]='h00000f24;  wr_data_rom[ 3987]='h00000000;
    rd_cycle[ 3988] = 1'b0;  wr_cycle[ 3988] = 1'b1;  addr_rom[ 3988]='h00000298;  wr_data_rom[ 3988]='h00000926;
    rd_cycle[ 3989] = 1'b1;  wr_cycle[ 3989] = 1'b0;  addr_rom[ 3989]='h00000298;  wr_data_rom[ 3989]='h00000000;
    rd_cycle[ 3990] = 1'b1;  wr_cycle[ 3990] = 1'b0;  addr_rom[ 3990]='h00000a58;  wr_data_rom[ 3990]='h00000000;
    rd_cycle[ 3991] = 1'b1;  wr_cycle[ 3991] = 1'b0;  addr_rom[ 3991]='h00000874;  wr_data_rom[ 3991]='h00000000;
    rd_cycle[ 3992] = 1'b0;  wr_cycle[ 3992] = 1'b1;  addr_rom[ 3992]='h000009ec;  wr_data_rom[ 3992]='h000008d3;
    rd_cycle[ 3993] = 1'b0;  wr_cycle[ 3993] = 1'b1;  addr_rom[ 3993]='h0000085c;  wr_data_rom[ 3993]='h0000045a;
    rd_cycle[ 3994] = 1'b0;  wr_cycle[ 3994] = 1'b1;  addr_rom[ 3994]='h00000e04;  wr_data_rom[ 3994]='h0000026d;
    rd_cycle[ 3995] = 1'b0;  wr_cycle[ 3995] = 1'b1;  addr_rom[ 3995]='h00000d58;  wr_data_rom[ 3995]='h00000d1e;
    rd_cycle[ 3996] = 1'b1;  wr_cycle[ 3996] = 1'b0;  addr_rom[ 3996]='h000007e0;  wr_data_rom[ 3996]='h00000000;
    rd_cycle[ 3997] = 1'b0;  wr_cycle[ 3997] = 1'b1;  addr_rom[ 3997]='h000009e4;  wr_data_rom[ 3997]='h00000047;
    rd_cycle[ 3998] = 1'b0;  wr_cycle[ 3998] = 1'b1;  addr_rom[ 3998]='h00000674;  wr_data_rom[ 3998]='h00000400;
    rd_cycle[ 3999] = 1'b0;  wr_cycle[ 3999] = 1'b1;  addr_rom[ 3999]='h000005a4;  wr_data_rom[ 3999]='h000008cd;
    // 1000 silence cycles
    rd_cycle[ 4000] = 1'b0;  wr_cycle[ 4000] = 1'b0;  addr_rom[ 4000]='h00000000;  wr_data_rom[ 4000]='h00000000;
    rd_cycle[ 4001] = 1'b0;  wr_cycle[ 4001] = 1'b0;  addr_rom[ 4001]='h00000000;  wr_data_rom[ 4001]='h00000000;
    rd_cycle[ 4002] = 1'b0;  wr_cycle[ 4002] = 1'b0;  addr_rom[ 4002]='h00000000;  wr_data_rom[ 4002]='h00000000;
    rd_cycle[ 4003] = 1'b0;  wr_cycle[ 4003] = 1'b0;  addr_rom[ 4003]='h00000000;  wr_data_rom[ 4003]='h00000000;
    rd_cycle[ 4004] = 1'b0;  wr_cycle[ 4004] = 1'b0;  addr_rom[ 4004]='h00000000;  wr_data_rom[ 4004]='h00000000;
    rd_cycle[ 4005] = 1'b0;  wr_cycle[ 4005] = 1'b0;  addr_rom[ 4005]='h00000000;  wr_data_rom[ 4005]='h00000000;
    rd_cycle[ 4006] = 1'b0;  wr_cycle[ 4006] = 1'b0;  addr_rom[ 4006]='h00000000;  wr_data_rom[ 4006]='h00000000;
    rd_cycle[ 4007] = 1'b0;  wr_cycle[ 4007] = 1'b0;  addr_rom[ 4007]='h00000000;  wr_data_rom[ 4007]='h00000000;
    rd_cycle[ 4008] = 1'b0;  wr_cycle[ 4008] = 1'b0;  addr_rom[ 4008]='h00000000;  wr_data_rom[ 4008]='h00000000;
    rd_cycle[ 4009] = 1'b0;  wr_cycle[ 4009] = 1'b0;  addr_rom[ 4009]='h00000000;  wr_data_rom[ 4009]='h00000000;
    rd_cycle[ 4010] = 1'b0;  wr_cycle[ 4010] = 1'b0;  addr_rom[ 4010]='h00000000;  wr_data_rom[ 4010]='h00000000;
    rd_cycle[ 4011] = 1'b0;  wr_cycle[ 4011] = 1'b0;  addr_rom[ 4011]='h00000000;  wr_data_rom[ 4011]='h00000000;
    rd_cycle[ 4012] = 1'b0;  wr_cycle[ 4012] = 1'b0;  addr_rom[ 4012]='h00000000;  wr_data_rom[ 4012]='h00000000;
    rd_cycle[ 4013] = 1'b0;  wr_cycle[ 4013] = 1'b0;  addr_rom[ 4013]='h00000000;  wr_data_rom[ 4013]='h00000000;
    rd_cycle[ 4014] = 1'b0;  wr_cycle[ 4014] = 1'b0;  addr_rom[ 4014]='h00000000;  wr_data_rom[ 4014]='h00000000;
    rd_cycle[ 4015] = 1'b0;  wr_cycle[ 4015] = 1'b0;  addr_rom[ 4015]='h00000000;  wr_data_rom[ 4015]='h00000000;
    rd_cycle[ 4016] = 1'b0;  wr_cycle[ 4016] = 1'b0;  addr_rom[ 4016]='h00000000;  wr_data_rom[ 4016]='h00000000;
    rd_cycle[ 4017] = 1'b0;  wr_cycle[ 4017] = 1'b0;  addr_rom[ 4017]='h00000000;  wr_data_rom[ 4017]='h00000000;
    rd_cycle[ 4018] = 1'b0;  wr_cycle[ 4018] = 1'b0;  addr_rom[ 4018]='h00000000;  wr_data_rom[ 4018]='h00000000;
    rd_cycle[ 4019] = 1'b0;  wr_cycle[ 4019] = 1'b0;  addr_rom[ 4019]='h00000000;  wr_data_rom[ 4019]='h00000000;
    rd_cycle[ 4020] = 1'b0;  wr_cycle[ 4020] = 1'b0;  addr_rom[ 4020]='h00000000;  wr_data_rom[ 4020]='h00000000;
    rd_cycle[ 4021] = 1'b0;  wr_cycle[ 4021] = 1'b0;  addr_rom[ 4021]='h00000000;  wr_data_rom[ 4021]='h00000000;
    rd_cycle[ 4022] = 1'b0;  wr_cycle[ 4022] = 1'b0;  addr_rom[ 4022]='h00000000;  wr_data_rom[ 4022]='h00000000;
    rd_cycle[ 4023] = 1'b0;  wr_cycle[ 4023] = 1'b0;  addr_rom[ 4023]='h00000000;  wr_data_rom[ 4023]='h00000000;
    rd_cycle[ 4024] = 1'b0;  wr_cycle[ 4024] = 1'b0;  addr_rom[ 4024]='h00000000;  wr_data_rom[ 4024]='h00000000;
    rd_cycle[ 4025] = 1'b0;  wr_cycle[ 4025] = 1'b0;  addr_rom[ 4025]='h00000000;  wr_data_rom[ 4025]='h00000000;
    rd_cycle[ 4026] = 1'b0;  wr_cycle[ 4026] = 1'b0;  addr_rom[ 4026]='h00000000;  wr_data_rom[ 4026]='h00000000;
    rd_cycle[ 4027] = 1'b0;  wr_cycle[ 4027] = 1'b0;  addr_rom[ 4027]='h00000000;  wr_data_rom[ 4027]='h00000000;
    rd_cycle[ 4028] = 1'b0;  wr_cycle[ 4028] = 1'b0;  addr_rom[ 4028]='h00000000;  wr_data_rom[ 4028]='h00000000;
    rd_cycle[ 4029] = 1'b0;  wr_cycle[ 4029] = 1'b0;  addr_rom[ 4029]='h00000000;  wr_data_rom[ 4029]='h00000000;
    rd_cycle[ 4030] = 1'b0;  wr_cycle[ 4030] = 1'b0;  addr_rom[ 4030]='h00000000;  wr_data_rom[ 4030]='h00000000;
    rd_cycle[ 4031] = 1'b0;  wr_cycle[ 4031] = 1'b0;  addr_rom[ 4031]='h00000000;  wr_data_rom[ 4031]='h00000000;
    rd_cycle[ 4032] = 1'b0;  wr_cycle[ 4032] = 1'b0;  addr_rom[ 4032]='h00000000;  wr_data_rom[ 4032]='h00000000;
    rd_cycle[ 4033] = 1'b0;  wr_cycle[ 4033] = 1'b0;  addr_rom[ 4033]='h00000000;  wr_data_rom[ 4033]='h00000000;
    rd_cycle[ 4034] = 1'b0;  wr_cycle[ 4034] = 1'b0;  addr_rom[ 4034]='h00000000;  wr_data_rom[ 4034]='h00000000;
    rd_cycle[ 4035] = 1'b0;  wr_cycle[ 4035] = 1'b0;  addr_rom[ 4035]='h00000000;  wr_data_rom[ 4035]='h00000000;
    rd_cycle[ 4036] = 1'b0;  wr_cycle[ 4036] = 1'b0;  addr_rom[ 4036]='h00000000;  wr_data_rom[ 4036]='h00000000;
    rd_cycle[ 4037] = 1'b0;  wr_cycle[ 4037] = 1'b0;  addr_rom[ 4037]='h00000000;  wr_data_rom[ 4037]='h00000000;
    rd_cycle[ 4038] = 1'b0;  wr_cycle[ 4038] = 1'b0;  addr_rom[ 4038]='h00000000;  wr_data_rom[ 4038]='h00000000;
    rd_cycle[ 4039] = 1'b0;  wr_cycle[ 4039] = 1'b0;  addr_rom[ 4039]='h00000000;  wr_data_rom[ 4039]='h00000000;
    rd_cycle[ 4040] = 1'b0;  wr_cycle[ 4040] = 1'b0;  addr_rom[ 4040]='h00000000;  wr_data_rom[ 4040]='h00000000;
    rd_cycle[ 4041] = 1'b0;  wr_cycle[ 4041] = 1'b0;  addr_rom[ 4041]='h00000000;  wr_data_rom[ 4041]='h00000000;
    rd_cycle[ 4042] = 1'b0;  wr_cycle[ 4042] = 1'b0;  addr_rom[ 4042]='h00000000;  wr_data_rom[ 4042]='h00000000;
    rd_cycle[ 4043] = 1'b0;  wr_cycle[ 4043] = 1'b0;  addr_rom[ 4043]='h00000000;  wr_data_rom[ 4043]='h00000000;
    rd_cycle[ 4044] = 1'b0;  wr_cycle[ 4044] = 1'b0;  addr_rom[ 4044]='h00000000;  wr_data_rom[ 4044]='h00000000;
    rd_cycle[ 4045] = 1'b0;  wr_cycle[ 4045] = 1'b0;  addr_rom[ 4045]='h00000000;  wr_data_rom[ 4045]='h00000000;
    rd_cycle[ 4046] = 1'b0;  wr_cycle[ 4046] = 1'b0;  addr_rom[ 4046]='h00000000;  wr_data_rom[ 4046]='h00000000;
    rd_cycle[ 4047] = 1'b0;  wr_cycle[ 4047] = 1'b0;  addr_rom[ 4047]='h00000000;  wr_data_rom[ 4047]='h00000000;
    rd_cycle[ 4048] = 1'b0;  wr_cycle[ 4048] = 1'b0;  addr_rom[ 4048]='h00000000;  wr_data_rom[ 4048]='h00000000;
    rd_cycle[ 4049] = 1'b0;  wr_cycle[ 4049] = 1'b0;  addr_rom[ 4049]='h00000000;  wr_data_rom[ 4049]='h00000000;
    rd_cycle[ 4050] = 1'b0;  wr_cycle[ 4050] = 1'b0;  addr_rom[ 4050]='h00000000;  wr_data_rom[ 4050]='h00000000;
    rd_cycle[ 4051] = 1'b0;  wr_cycle[ 4051] = 1'b0;  addr_rom[ 4051]='h00000000;  wr_data_rom[ 4051]='h00000000;
    rd_cycle[ 4052] = 1'b0;  wr_cycle[ 4052] = 1'b0;  addr_rom[ 4052]='h00000000;  wr_data_rom[ 4052]='h00000000;
    rd_cycle[ 4053] = 1'b0;  wr_cycle[ 4053] = 1'b0;  addr_rom[ 4053]='h00000000;  wr_data_rom[ 4053]='h00000000;
    rd_cycle[ 4054] = 1'b0;  wr_cycle[ 4054] = 1'b0;  addr_rom[ 4054]='h00000000;  wr_data_rom[ 4054]='h00000000;
    rd_cycle[ 4055] = 1'b0;  wr_cycle[ 4055] = 1'b0;  addr_rom[ 4055]='h00000000;  wr_data_rom[ 4055]='h00000000;
    rd_cycle[ 4056] = 1'b0;  wr_cycle[ 4056] = 1'b0;  addr_rom[ 4056]='h00000000;  wr_data_rom[ 4056]='h00000000;
    rd_cycle[ 4057] = 1'b0;  wr_cycle[ 4057] = 1'b0;  addr_rom[ 4057]='h00000000;  wr_data_rom[ 4057]='h00000000;
    rd_cycle[ 4058] = 1'b0;  wr_cycle[ 4058] = 1'b0;  addr_rom[ 4058]='h00000000;  wr_data_rom[ 4058]='h00000000;
    rd_cycle[ 4059] = 1'b0;  wr_cycle[ 4059] = 1'b0;  addr_rom[ 4059]='h00000000;  wr_data_rom[ 4059]='h00000000;
    rd_cycle[ 4060] = 1'b0;  wr_cycle[ 4060] = 1'b0;  addr_rom[ 4060]='h00000000;  wr_data_rom[ 4060]='h00000000;
    rd_cycle[ 4061] = 1'b0;  wr_cycle[ 4061] = 1'b0;  addr_rom[ 4061]='h00000000;  wr_data_rom[ 4061]='h00000000;
    rd_cycle[ 4062] = 1'b0;  wr_cycle[ 4062] = 1'b0;  addr_rom[ 4062]='h00000000;  wr_data_rom[ 4062]='h00000000;
    rd_cycle[ 4063] = 1'b0;  wr_cycle[ 4063] = 1'b0;  addr_rom[ 4063]='h00000000;  wr_data_rom[ 4063]='h00000000;
    rd_cycle[ 4064] = 1'b0;  wr_cycle[ 4064] = 1'b0;  addr_rom[ 4064]='h00000000;  wr_data_rom[ 4064]='h00000000;
    rd_cycle[ 4065] = 1'b0;  wr_cycle[ 4065] = 1'b0;  addr_rom[ 4065]='h00000000;  wr_data_rom[ 4065]='h00000000;
    rd_cycle[ 4066] = 1'b0;  wr_cycle[ 4066] = 1'b0;  addr_rom[ 4066]='h00000000;  wr_data_rom[ 4066]='h00000000;
    rd_cycle[ 4067] = 1'b0;  wr_cycle[ 4067] = 1'b0;  addr_rom[ 4067]='h00000000;  wr_data_rom[ 4067]='h00000000;
    rd_cycle[ 4068] = 1'b0;  wr_cycle[ 4068] = 1'b0;  addr_rom[ 4068]='h00000000;  wr_data_rom[ 4068]='h00000000;
    rd_cycle[ 4069] = 1'b0;  wr_cycle[ 4069] = 1'b0;  addr_rom[ 4069]='h00000000;  wr_data_rom[ 4069]='h00000000;
    rd_cycle[ 4070] = 1'b0;  wr_cycle[ 4070] = 1'b0;  addr_rom[ 4070]='h00000000;  wr_data_rom[ 4070]='h00000000;
    rd_cycle[ 4071] = 1'b0;  wr_cycle[ 4071] = 1'b0;  addr_rom[ 4071]='h00000000;  wr_data_rom[ 4071]='h00000000;
    rd_cycle[ 4072] = 1'b0;  wr_cycle[ 4072] = 1'b0;  addr_rom[ 4072]='h00000000;  wr_data_rom[ 4072]='h00000000;
    rd_cycle[ 4073] = 1'b0;  wr_cycle[ 4073] = 1'b0;  addr_rom[ 4073]='h00000000;  wr_data_rom[ 4073]='h00000000;
    rd_cycle[ 4074] = 1'b0;  wr_cycle[ 4074] = 1'b0;  addr_rom[ 4074]='h00000000;  wr_data_rom[ 4074]='h00000000;
    rd_cycle[ 4075] = 1'b0;  wr_cycle[ 4075] = 1'b0;  addr_rom[ 4075]='h00000000;  wr_data_rom[ 4075]='h00000000;
    rd_cycle[ 4076] = 1'b0;  wr_cycle[ 4076] = 1'b0;  addr_rom[ 4076]='h00000000;  wr_data_rom[ 4076]='h00000000;
    rd_cycle[ 4077] = 1'b0;  wr_cycle[ 4077] = 1'b0;  addr_rom[ 4077]='h00000000;  wr_data_rom[ 4077]='h00000000;
    rd_cycle[ 4078] = 1'b0;  wr_cycle[ 4078] = 1'b0;  addr_rom[ 4078]='h00000000;  wr_data_rom[ 4078]='h00000000;
    rd_cycle[ 4079] = 1'b0;  wr_cycle[ 4079] = 1'b0;  addr_rom[ 4079]='h00000000;  wr_data_rom[ 4079]='h00000000;
    rd_cycle[ 4080] = 1'b0;  wr_cycle[ 4080] = 1'b0;  addr_rom[ 4080]='h00000000;  wr_data_rom[ 4080]='h00000000;
    rd_cycle[ 4081] = 1'b0;  wr_cycle[ 4081] = 1'b0;  addr_rom[ 4081]='h00000000;  wr_data_rom[ 4081]='h00000000;
    rd_cycle[ 4082] = 1'b0;  wr_cycle[ 4082] = 1'b0;  addr_rom[ 4082]='h00000000;  wr_data_rom[ 4082]='h00000000;
    rd_cycle[ 4083] = 1'b0;  wr_cycle[ 4083] = 1'b0;  addr_rom[ 4083]='h00000000;  wr_data_rom[ 4083]='h00000000;
    rd_cycle[ 4084] = 1'b0;  wr_cycle[ 4084] = 1'b0;  addr_rom[ 4084]='h00000000;  wr_data_rom[ 4084]='h00000000;
    rd_cycle[ 4085] = 1'b0;  wr_cycle[ 4085] = 1'b0;  addr_rom[ 4085]='h00000000;  wr_data_rom[ 4085]='h00000000;
    rd_cycle[ 4086] = 1'b0;  wr_cycle[ 4086] = 1'b0;  addr_rom[ 4086]='h00000000;  wr_data_rom[ 4086]='h00000000;
    rd_cycle[ 4087] = 1'b0;  wr_cycle[ 4087] = 1'b0;  addr_rom[ 4087]='h00000000;  wr_data_rom[ 4087]='h00000000;
    rd_cycle[ 4088] = 1'b0;  wr_cycle[ 4088] = 1'b0;  addr_rom[ 4088]='h00000000;  wr_data_rom[ 4088]='h00000000;
    rd_cycle[ 4089] = 1'b0;  wr_cycle[ 4089] = 1'b0;  addr_rom[ 4089]='h00000000;  wr_data_rom[ 4089]='h00000000;
    rd_cycle[ 4090] = 1'b0;  wr_cycle[ 4090] = 1'b0;  addr_rom[ 4090]='h00000000;  wr_data_rom[ 4090]='h00000000;
    rd_cycle[ 4091] = 1'b0;  wr_cycle[ 4091] = 1'b0;  addr_rom[ 4091]='h00000000;  wr_data_rom[ 4091]='h00000000;
    rd_cycle[ 4092] = 1'b0;  wr_cycle[ 4092] = 1'b0;  addr_rom[ 4092]='h00000000;  wr_data_rom[ 4092]='h00000000;
    rd_cycle[ 4093] = 1'b0;  wr_cycle[ 4093] = 1'b0;  addr_rom[ 4093]='h00000000;  wr_data_rom[ 4093]='h00000000;
    rd_cycle[ 4094] = 1'b0;  wr_cycle[ 4094] = 1'b0;  addr_rom[ 4094]='h00000000;  wr_data_rom[ 4094]='h00000000;
    rd_cycle[ 4095] = 1'b0;  wr_cycle[ 4095] = 1'b0;  addr_rom[ 4095]='h00000000;  wr_data_rom[ 4095]='h00000000;
    rd_cycle[ 4096] = 1'b0;  wr_cycle[ 4096] = 1'b0;  addr_rom[ 4096]='h00000000;  wr_data_rom[ 4096]='h00000000;
    rd_cycle[ 4097] = 1'b0;  wr_cycle[ 4097] = 1'b0;  addr_rom[ 4097]='h00000000;  wr_data_rom[ 4097]='h00000000;
    rd_cycle[ 4098] = 1'b0;  wr_cycle[ 4098] = 1'b0;  addr_rom[ 4098]='h00000000;  wr_data_rom[ 4098]='h00000000;
    rd_cycle[ 4099] = 1'b0;  wr_cycle[ 4099] = 1'b0;  addr_rom[ 4099]='h00000000;  wr_data_rom[ 4099]='h00000000;
    rd_cycle[ 4100] = 1'b0;  wr_cycle[ 4100] = 1'b0;  addr_rom[ 4100]='h00000000;  wr_data_rom[ 4100]='h00000000;
    rd_cycle[ 4101] = 1'b0;  wr_cycle[ 4101] = 1'b0;  addr_rom[ 4101]='h00000000;  wr_data_rom[ 4101]='h00000000;
    rd_cycle[ 4102] = 1'b0;  wr_cycle[ 4102] = 1'b0;  addr_rom[ 4102]='h00000000;  wr_data_rom[ 4102]='h00000000;
    rd_cycle[ 4103] = 1'b0;  wr_cycle[ 4103] = 1'b0;  addr_rom[ 4103]='h00000000;  wr_data_rom[ 4103]='h00000000;
    rd_cycle[ 4104] = 1'b0;  wr_cycle[ 4104] = 1'b0;  addr_rom[ 4104]='h00000000;  wr_data_rom[ 4104]='h00000000;
    rd_cycle[ 4105] = 1'b0;  wr_cycle[ 4105] = 1'b0;  addr_rom[ 4105]='h00000000;  wr_data_rom[ 4105]='h00000000;
    rd_cycle[ 4106] = 1'b0;  wr_cycle[ 4106] = 1'b0;  addr_rom[ 4106]='h00000000;  wr_data_rom[ 4106]='h00000000;
    rd_cycle[ 4107] = 1'b0;  wr_cycle[ 4107] = 1'b0;  addr_rom[ 4107]='h00000000;  wr_data_rom[ 4107]='h00000000;
    rd_cycle[ 4108] = 1'b0;  wr_cycle[ 4108] = 1'b0;  addr_rom[ 4108]='h00000000;  wr_data_rom[ 4108]='h00000000;
    rd_cycle[ 4109] = 1'b0;  wr_cycle[ 4109] = 1'b0;  addr_rom[ 4109]='h00000000;  wr_data_rom[ 4109]='h00000000;
    rd_cycle[ 4110] = 1'b0;  wr_cycle[ 4110] = 1'b0;  addr_rom[ 4110]='h00000000;  wr_data_rom[ 4110]='h00000000;
    rd_cycle[ 4111] = 1'b0;  wr_cycle[ 4111] = 1'b0;  addr_rom[ 4111]='h00000000;  wr_data_rom[ 4111]='h00000000;
    rd_cycle[ 4112] = 1'b0;  wr_cycle[ 4112] = 1'b0;  addr_rom[ 4112]='h00000000;  wr_data_rom[ 4112]='h00000000;
    rd_cycle[ 4113] = 1'b0;  wr_cycle[ 4113] = 1'b0;  addr_rom[ 4113]='h00000000;  wr_data_rom[ 4113]='h00000000;
    rd_cycle[ 4114] = 1'b0;  wr_cycle[ 4114] = 1'b0;  addr_rom[ 4114]='h00000000;  wr_data_rom[ 4114]='h00000000;
    rd_cycle[ 4115] = 1'b0;  wr_cycle[ 4115] = 1'b0;  addr_rom[ 4115]='h00000000;  wr_data_rom[ 4115]='h00000000;
    rd_cycle[ 4116] = 1'b0;  wr_cycle[ 4116] = 1'b0;  addr_rom[ 4116]='h00000000;  wr_data_rom[ 4116]='h00000000;
    rd_cycle[ 4117] = 1'b0;  wr_cycle[ 4117] = 1'b0;  addr_rom[ 4117]='h00000000;  wr_data_rom[ 4117]='h00000000;
    rd_cycle[ 4118] = 1'b0;  wr_cycle[ 4118] = 1'b0;  addr_rom[ 4118]='h00000000;  wr_data_rom[ 4118]='h00000000;
    rd_cycle[ 4119] = 1'b0;  wr_cycle[ 4119] = 1'b0;  addr_rom[ 4119]='h00000000;  wr_data_rom[ 4119]='h00000000;
    rd_cycle[ 4120] = 1'b0;  wr_cycle[ 4120] = 1'b0;  addr_rom[ 4120]='h00000000;  wr_data_rom[ 4120]='h00000000;
    rd_cycle[ 4121] = 1'b0;  wr_cycle[ 4121] = 1'b0;  addr_rom[ 4121]='h00000000;  wr_data_rom[ 4121]='h00000000;
    rd_cycle[ 4122] = 1'b0;  wr_cycle[ 4122] = 1'b0;  addr_rom[ 4122]='h00000000;  wr_data_rom[ 4122]='h00000000;
    rd_cycle[ 4123] = 1'b0;  wr_cycle[ 4123] = 1'b0;  addr_rom[ 4123]='h00000000;  wr_data_rom[ 4123]='h00000000;
    rd_cycle[ 4124] = 1'b0;  wr_cycle[ 4124] = 1'b0;  addr_rom[ 4124]='h00000000;  wr_data_rom[ 4124]='h00000000;
    rd_cycle[ 4125] = 1'b0;  wr_cycle[ 4125] = 1'b0;  addr_rom[ 4125]='h00000000;  wr_data_rom[ 4125]='h00000000;
    rd_cycle[ 4126] = 1'b0;  wr_cycle[ 4126] = 1'b0;  addr_rom[ 4126]='h00000000;  wr_data_rom[ 4126]='h00000000;
    rd_cycle[ 4127] = 1'b0;  wr_cycle[ 4127] = 1'b0;  addr_rom[ 4127]='h00000000;  wr_data_rom[ 4127]='h00000000;
    rd_cycle[ 4128] = 1'b0;  wr_cycle[ 4128] = 1'b0;  addr_rom[ 4128]='h00000000;  wr_data_rom[ 4128]='h00000000;
    rd_cycle[ 4129] = 1'b0;  wr_cycle[ 4129] = 1'b0;  addr_rom[ 4129]='h00000000;  wr_data_rom[ 4129]='h00000000;
    rd_cycle[ 4130] = 1'b0;  wr_cycle[ 4130] = 1'b0;  addr_rom[ 4130]='h00000000;  wr_data_rom[ 4130]='h00000000;
    rd_cycle[ 4131] = 1'b0;  wr_cycle[ 4131] = 1'b0;  addr_rom[ 4131]='h00000000;  wr_data_rom[ 4131]='h00000000;
    rd_cycle[ 4132] = 1'b0;  wr_cycle[ 4132] = 1'b0;  addr_rom[ 4132]='h00000000;  wr_data_rom[ 4132]='h00000000;
    rd_cycle[ 4133] = 1'b0;  wr_cycle[ 4133] = 1'b0;  addr_rom[ 4133]='h00000000;  wr_data_rom[ 4133]='h00000000;
    rd_cycle[ 4134] = 1'b0;  wr_cycle[ 4134] = 1'b0;  addr_rom[ 4134]='h00000000;  wr_data_rom[ 4134]='h00000000;
    rd_cycle[ 4135] = 1'b0;  wr_cycle[ 4135] = 1'b0;  addr_rom[ 4135]='h00000000;  wr_data_rom[ 4135]='h00000000;
    rd_cycle[ 4136] = 1'b0;  wr_cycle[ 4136] = 1'b0;  addr_rom[ 4136]='h00000000;  wr_data_rom[ 4136]='h00000000;
    rd_cycle[ 4137] = 1'b0;  wr_cycle[ 4137] = 1'b0;  addr_rom[ 4137]='h00000000;  wr_data_rom[ 4137]='h00000000;
    rd_cycle[ 4138] = 1'b0;  wr_cycle[ 4138] = 1'b0;  addr_rom[ 4138]='h00000000;  wr_data_rom[ 4138]='h00000000;
    rd_cycle[ 4139] = 1'b0;  wr_cycle[ 4139] = 1'b0;  addr_rom[ 4139]='h00000000;  wr_data_rom[ 4139]='h00000000;
    rd_cycle[ 4140] = 1'b0;  wr_cycle[ 4140] = 1'b0;  addr_rom[ 4140]='h00000000;  wr_data_rom[ 4140]='h00000000;
    rd_cycle[ 4141] = 1'b0;  wr_cycle[ 4141] = 1'b0;  addr_rom[ 4141]='h00000000;  wr_data_rom[ 4141]='h00000000;
    rd_cycle[ 4142] = 1'b0;  wr_cycle[ 4142] = 1'b0;  addr_rom[ 4142]='h00000000;  wr_data_rom[ 4142]='h00000000;
    rd_cycle[ 4143] = 1'b0;  wr_cycle[ 4143] = 1'b0;  addr_rom[ 4143]='h00000000;  wr_data_rom[ 4143]='h00000000;
    rd_cycle[ 4144] = 1'b0;  wr_cycle[ 4144] = 1'b0;  addr_rom[ 4144]='h00000000;  wr_data_rom[ 4144]='h00000000;
    rd_cycle[ 4145] = 1'b0;  wr_cycle[ 4145] = 1'b0;  addr_rom[ 4145]='h00000000;  wr_data_rom[ 4145]='h00000000;
    rd_cycle[ 4146] = 1'b0;  wr_cycle[ 4146] = 1'b0;  addr_rom[ 4146]='h00000000;  wr_data_rom[ 4146]='h00000000;
    rd_cycle[ 4147] = 1'b0;  wr_cycle[ 4147] = 1'b0;  addr_rom[ 4147]='h00000000;  wr_data_rom[ 4147]='h00000000;
    rd_cycle[ 4148] = 1'b0;  wr_cycle[ 4148] = 1'b0;  addr_rom[ 4148]='h00000000;  wr_data_rom[ 4148]='h00000000;
    rd_cycle[ 4149] = 1'b0;  wr_cycle[ 4149] = 1'b0;  addr_rom[ 4149]='h00000000;  wr_data_rom[ 4149]='h00000000;
    rd_cycle[ 4150] = 1'b0;  wr_cycle[ 4150] = 1'b0;  addr_rom[ 4150]='h00000000;  wr_data_rom[ 4150]='h00000000;
    rd_cycle[ 4151] = 1'b0;  wr_cycle[ 4151] = 1'b0;  addr_rom[ 4151]='h00000000;  wr_data_rom[ 4151]='h00000000;
    rd_cycle[ 4152] = 1'b0;  wr_cycle[ 4152] = 1'b0;  addr_rom[ 4152]='h00000000;  wr_data_rom[ 4152]='h00000000;
    rd_cycle[ 4153] = 1'b0;  wr_cycle[ 4153] = 1'b0;  addr_rom[ 4153]='h00000000;  wr_data_rom[ 4153]='h00000000;
    rd_cycle[ 4154] = 1'b0;  wr_cycle[ 4154] = 1'b0;  addr_rom[ 4154]='h00000000;  wr_data_rom[ 4154]='h00000000;
    rd_cycle[ 4155] = 1'b0;  wr_cycle[ 4155] = 1'b0;  addr_rom[ 4155]='h00000000;  wr_data_rom[ 4155]='h00000000;
    rd_cycle[ 4156] = 1'b0;  wr_cycle[ 4156] = 1'b0;  addr_rom[ 4156]='h00000000;  wr_data_rom[ 4156]='h00000000;
    rd_cycle[ 4157] = 1'b0;  wr_cycle[ 4157] = 1'b0;  addr_rom[ 4157]='h00000000;  wr_data_rom[ 4157]='h00000000;
    rd_cycle[ 4158] = 1'b0;  wr_cycle[ 4158] = 1'b0;  addr_rom[ 4158]='h00000000;  wr_data_rom[ 4158]='h00000000;
    rd_cycle[ 4159] = 1'b0;  wr_cycle[ 4159] = 1'b0;  addr_rom[ 4159]='h00000000;  wr_data_rom[ 4159]='h00000000;
    rd_cycle[ 4160] = 1'b0;  wr_cycle[ 4160] = 1'b0;  addr_rom[ 4160]='h00000000;  wr_data_rom[ 4160]='h00000000;
    rd_cycle[ 4161] = 1'b0;  wr_cycle[ 4161] = 1'b0;  addr_rom[ 4161]='h00000000;  wr_data_rom[ 4161]='h00000000;
    rd_cycle[ 4162] = 1'b0;  wr_cycle[ 4162] = 1'b0;  addr_rom[ 4162]='h00000000;  wr_data_rom[ 4162]='h00000000;
    rd_cycle[ 4163] = 1'b0;  wr_cycle[ 4163] = 1'b0;  addr_rom[ 4163]='h00000000;  wr_data_rom[ 4163]='h00000000;
    rd_cycle[ 4164] = 1'b0;  wr_cycle[ 4164] = 1'b0;  addr_rom[ 4164]='h00000000;  wr_data_rom[ 4164]='h00000000;
    rd_cycle[ 4165] = 1'b0;  wr_cycle[ 4165] = 1'b0;  addr_rom[ 4165]='h00000000;  wr_data_rom[ 4165]='h00000000;
    rd_cycle[ 4166] = 1'b0;  wr_cycle[ 4166] = 1'b0;  addr_rom[ 4166]='h00000000;  wr_data_rom[ 4166]='h00000000;
    rd_cycle[ 4167] = 1'b0;  wr_cycle[ 4167] = 1'b0;  addr_rom[ 4167]='h00000000;  wr_data_rom[ 4167]='h00000000;
    rd_cycle[ 4168] = 1'b0;  wr_cycle[ 4168] = 1'b0;  addr_rom[ 4168]='h00000000;  wr_data_rom[ 4168]='h00000000;
    rd_cycle[ 4169] = 1'b0;  wr_cycle[ 4169] = 1'b0;  addr_rom[ 4169]='h00000000;  wr_data_rom[ 4169]='h00000000;
    rd_cycle[ 4170] = 1'b0;  wr_cycle[ 4170] = 1'b0;  addr_rom[ 4170]='h00000000;  wr_data_rom[ 4170]='h00000000;
    rd_cycle[ 4171] = 1'b0;  wr_cycle[ 4171] = 1'b0;  addr_rom[ 4171]='h00000000;  wr_data_rom[ 4171]='h00000000;
    rd_cycle[ 4172] = 1'b0;  wr_cycle[ 4172] = 1'b0;  addr_rom[ 4172]='h00000000;  wr_data_rom[ 4172]='h00000000;
    rd_cycle[ 4173] = 1'b0;  wr_cycle[ 4173] = 1'b0;  addr_rom[ 4173]='h00000000;  wr_data_rom[ 4173]='h00000000;
    rd_cycle[ 4174] = 1'b0;  wr_cycle[ 4174] = 1'b0;  addr_rom[ 4174]='h00000000;  wr_data_rom[ 4174]='h00000000;
    rd_cycle[ 4175] = 1'b0;  wr_cycle[ 4175] = 1'b0;  addr_rom[ 4175]='h00000000;  wr_data_rom[ 4175]='h00000000;
    rd_cycle[ 4176] = 1'b0;  wr_cycle[ 4176] = 1'b0;  addr_rom[ 4176]='h00000000;  wr_data_rom[ 4176]='h00000000;
    rd_cycle[ 4177] = 1'b0;  wr_cycle[ 4177] = 1'b0;  addr_rom[ 4177]='h00000000;  wr_data_rom[ 4177]='h00000000;
    rd_cycle[ 4178] = 1'b0;  wr_cycle[ 4178] = 1'b0;  addr_rom[ 4178]='h00000000;  wr_data_rom[ 4178]='h00000000;
    rd_cycle[ 4179] = 1'b0;  wr_cycle[ 4179] = 1'b0;  addr_rom[ 4179]='h00000000;  wr_data_rom[ 4179]='h00000000;
    rd_cycle[ 4180] = 1'b0;  wr_cycle[ 4180] = 1'b0;  addr_rom[ 4180]='h00000000;  wr_data_rom[ 4180]='h00000000;
    rd_cycle[ 4181] = 1'b0;  wr_cycle[ 4181] = 1'b0;  addr_rom[ 4181]='h00000000;  wr_data_rom[ 4181]='h00000000;
    rd_cycle[ 4182] = 1'b0;  wr_cycle[ 4182] = 1'b0;  addr_rom[ 4182]='h00000000;  wr_data_rom[ 4182]='h00000000;
    rd_cycle[ 4183] = 1'b0;  wr_cycle[ 4183] = 1'b0;  addr_rom[ 4183]='h00000000;  wr_data_rom[ 4183]='h00000000;
    rd_cycle[ 4184] = 1'b0;  wr_cycle[ 4184] = 1'b0;  addr_rom[ 4184]='h00000000;  wr_data_rom[ 4184]='h00000000;
    rd_cycle[ 4185] = 1'b0;  wr_cycle[ 4185] = 1'b0;  addr_rom[ 4185]='h00000000;  wr_data_rom[ 4185]='h00000000;
    rd_cycle[ 4186] = 1'b0;  wr_cycle[ 4186] = 1'b0;  addr_rom[ 4186]='h00000000;  wr_data_rom[ 4186]='h00000000;
    rd_cycle[ 4187] = 1'b0;  wr_cycle[ 4187] = 1'b0;  addr_rom[ 4187]='h00000000;  wr_data_rom[ 4187]='h00000000;
    rd_cycle[ 4188] = 1'b0;  wr_cycle[ 4188] = 1'b0;  addr_rom[ 4188]='h00000000;  wr_data_rom[ 4188]='h00000000;
    rd_cycle[ 4189] = 1'b0;  wr_cycle[ 4189] = 1'b0;  addr_rom[ 4189]='h00000000;  wr_data_rom[ 4189]='h00000000;
    rd_cycle[ 4190] = 1'b0;  wr_cycle[ 4190] = 1'b0;  addr_rom[ 4190]='h00000000;  wr_data_rom[ 4190]='h00000000;
    rd_cycle[ 4191] = 1'b0;  wr_cycle[ 4191] = 1'b0;  addr_rom[ 4191]='h00000000;  wr_data_rom[ 4191]='h00000000;
    rd_cycle[ 4192] = 1'b0;  wr_cycle[ 4192] = 1'b0;  addr_rom[ 4192]='h00000000;  wr_data_rom[ 4192]='h00000000;
    rd_cycle[ 4193] = 1'b0;  wr_cycle[ 4193] = 1'b0;  addr_rom[ 4193]='h00000000;  wr_data_rom[ 4193]='h00000000;
    rd_cycle[ 4194] = 1'b0;  wr_cycle[ 4194] = 1'b0;  addr_rom[ 4194]='h00000000;  wr_data_rom[ 4194]='h00000000;
    rd_cycle[ 4195] = 1'b0;  wr_cycle[ 4195] = 1'b0;  addr_rom[ 4195]='h00000000;  wr_data_rom[ 4195]='h00000000;
    rd_cycle[ 4196] = 1'b0;  wr_cycle[ 4196] = 1'b0;  addr_rom[ 4196]='h00000000;  wr_data_rom[ 4196]='h00000000;
    rd_cycle[ 4197] = 1'b0;  wr_cycle[ 4197] = 1'b0;  addr_rom[ 4197]='h00000000;  wr_data_rom[ 4197]='h00000000;
    rd_cycle[ 4198] = 1'b0;  wr_cycle[ 4198] = 1'b0;  addr_rom[ 4198]='h00000000;  wr_data_rom[ 4198]='h00000000;
    rd_cycle[ 4199] = 1'b0;  wr_cycle[ 4199] = 1'b0;  addr_rom[ 4199]='h00000000;  wr_data_rom[ 4199]='h00000000;
    rd_cycle[ 4200] = 1'b0;  wr_cycle[ 4200] = 1'b0;  addr_rom[ 4200]='h00000000;  wr_data_rom[ 4200]='h00000000;
    rd_cycle[ 4201] = 1'b0;  wr_cycle[ 4201] = 1'b0;  addr_rom[ 4201]='h00000000;  wr_data_rom[ 4201]='h00000000;
    rd_cycle[ 4202] = 1'b0;  wr_cycle[ 4202] = 1'b0;  addr_rom[ 4202]='h00000000;  wr_data_rom[ 4202]='h00000000;
    rd_cycle[ 4203] = 1'b0;  wr_cycle[ 4203] = 1'b0;  addr_rom[ 4203]='h00000000;  wr_data_rom[ 4203]='h00000000;
    rd_cycle[ 4204] = 1'b0;  wr_cycle[ 4204] = 1'b0;  addr_rom[ 4204]='h00000000;  wr_data_rom[ 4204]='h00000000;
    rd_cycle[ 4205] = 1'b0;  wr_cycle[ 4205] = 1'b0;  addr_rom[ 4205]='h00000000;  wr_data_rom[ 4205]='h00000000;
    rd_cycle[ 4206] = 1'b0;  wr_cycle[ 4206] = 1'b0;  addr_rom[ 4206]='h00000000;  wr_data_rom[ 4206]='h00000000;
    rd_cycle[ 4207] = 1'b0;  wr_cycle[ 4207] = 1'b0;  addr_rom[ 4207]='h00000000;  wr_data_rom[ 4207]='h00000000;
    rd_cycle[ 4208] = 1'b0;  wr_cycle[ 4208] = 1'b0;  addr_rom[ 4208]='h00000000;  wr_data_rom[ 4208]='h00000000;
    rd_cycle[ 4209] = 1'b0;  wr_cycle[ 4209] = 1'b0;  addr_rom[ 4209]='h00000000;  wr_data_rom[ 4209]='h00000000;
    rd_cycle[ 4210] = 1'b0;  wr_cycle[ 4210] = 1'b0;  addr_rom[ 4210]='h00000000;  wr_data_rom[ 4210]='h00000000;
    rd_cycle[ 4211] = 1'b0;  wr_cycle[ 4211] = 1'b0;  addr_rom[ 4211]='h00000000;  wr_data_rom[ 4211]='h00000000;
    rd_cycle[ 4212] = 1'b0;  wr_cycle[ 4212] = 1'b0;  addr_rom[ 4212]='h00000000;  wr_data_rom[ 4212]='h00000000;
    rd_cycle[ 4213] = 1'b0;  wr_cycle[ 4213] = 1'b0;  addr_rom[ 4213]='h00000000;  wr_data_rom[ 4213]='h00000000;
    rd_cycle[ 4214] = 1'b0;  wr_cycle[ 4214] = 1'b0;  addr_rom[ 4214]='h00000000;  wr_data_rom[ 4214]='h00000000;
    rd_cycle[ 4215] = 1'b0;  wr_cycle[ 4215] = 1'b0;  addr_rom[ 4215]='h00000000;  wr_data_rom[ 4215]='h00000000;
    rd_cycle[ 4216] = 1'b0;  wr_cycle[ 4216] = 1'b0;  addr_rom[ 4216]='h00000000;  wr_data_rom[ 4216]='h00000000;
    rd_cycle[ 4217] = 1'b0;  wr_cycle[ 4217] = 1'b0;  addr_rom[ 4217]='h00000000;  wr_data_rom[ 4217]='h00000000;
    rd_cycle[ 4218] = 1'b0;  wr_cycle[ 4218] = 1'b0;  addr_rom[ 4218]='h00000000;  wr_data_rom[ 4218]='h00000000;
    rd_cycle[ 4219] = 1'b0;  wr_cycle[ 4219] = 1'b0;  addr_rom[ 4219]='h00000000;  wr_data_rom[ 4219]='h00000000;
    rd_cycle[ 4220] = 1'b0;  wr_cycle[ 4220] = 1'b0;  addr_rom[ 4220]='h00000000;  wr_data_rom[ 4220]='h00000000;
    rd_cycle[ 4221] = 1'b0;  wr_cycle[ 4221] = 1'b0;  addr_rom[ 4221]='h00000000;  wr_data_rom[ 4221]='h00000000;
    rd_cycle[ 4222] = 1'b0;  wr_cycle[ 4222] = 1'b0;  addr_rom[ 4222]='h00000000;  wr_data_rom[ 4222]='h00000000;
    rd_cycle[ 4223] = 1'b0;  wr_cycle[ 4223] = 1'b0;  addr_rom[ 4223]='h00000000;  wr_data_rom[ 4223]='h00000000;
    rd_cycle[ 4224] = 1'b0;  wr_cycle[ 4224] = 1'b0;  addr_rom[ 4224]='h00000000;  wr_data_rom[ 4224]='h00000000;
    rd_cycle[ 4225] = 1'b0;  wr_cycle[ 4225] = 1'b0;  addr_rom[ 4225]='h00000000;  wr_data_rom[ 4225]='h00000000;
    rd_cycle[ 4226] = 1'b0;  wr_cycle[ 4226] = 1'b0;  addr_rom[ 4226]='h00000000;  wr_data_rom[ 4226]='h00000000;
    rd_cycle[ 4227] = 1'b0;  wr_cycle[ 4227] = 1'b0;  addr_rom[ 4227]='h00000000;  wr_data_rom[ 4227]='h00000000;
    rd_cycle[ 4228] = 1'b0;  wr_cycle[ 4228] = 1'b0;  addr_rom[ 4228]='h00000000;  wr_data_rom[ 4228]='h00000000;
    rd_cycle[ 4229] = 1'b0;  wr_cycle[ 4229] = 1'b0;  addr_rom[ 4229]='h00000000;  wr_data_rom[ 4229]='h00000000;
    rd_cycle[ 4230] = 1'b0;  wr_cycle[ 4230] = 1'b0;  addr_rom[ 4230]='h00000000;  wr_data_rom[ 4230]='h00000000;
    rd_cycle[ 4231] = 1'b0;  wr_cycle[ 4231] = 1'b0;  addr_rom[ 4231]='h00000000;  wr_data_rom[ 4231]='h00000000;
    rd_cycle[ 4232] = 1'b0;  wr_cycle[ 4232] = 1'b0;  addr_rom[ 4232]='h00000000;  wr_data_rom[ 4232]='h00000000;
    rd_cycle[ 4233] = 1'b0;  wr_cycle[ 4233] = 1'b0;  addr_rom[ 4233]='h00000000;  wr_data_rom[ 4233]='h00000000;
    rd_cycle[ 4234] = 1'b0;  wr_cycle[ 4234] = 1'b0;  addr_rom[ 4234]='h00000000;  wr_data_rom[ 4234]='h00000000;
    rd_cycle[ 4235] = 1'b0;  wr_cycle[ 4235] = 1'b0;  addr_rom[ 4235]='h00000000;  wr_data_rom[ 4235]='h00000000;
    rd_cycle[ 4236] = 1'b0;  wr_cycle[ 4236] = 1'b0;  addr_rom[ 4236]='h00000000;  wr_data_rom[ 4236]='h00000000;
    rd_cycle[ 4237] = 1'b0;  wr_cycle[ 4237] = 1'b0;  addr_rom[ 4237]='h00000000;  wr_data_rom[ 4237]='h00000000;
    rd_cycle[ 4238] = 1'b0;  wr_cycle[ 4238] = 1'b0;  addr_rom[ 4238]='h00000000;  wr_data_rom[ 4238]='h00000000;
    rd_cycle[ 4239] = 1'b0;  wr_cycle[ 4239] = 1'b0;  addr_rom[ 4239]='h00000000;  wr_data_rom[ 4239]='h00000000;
    rd_cycle[ 4240] = 1'b0;  wr_cycle[ 4240] = 1'b0;  addr_rom[ 4240]='h00000000;  wr_data_rom[ 4240]='h00000000;
    rd_cycle[ 4241] = 1'b0;  wr_cycle[ 4241] = 1'b0;  addr_rom[ 4241]='h00000000;  wr_data_rom[ 4241]='h00000000;
    rd_cycle[ 4242] = 1'b0;  wr_cycle[ 4242] = 1'b0;  addr_rom[ 4242]='h00000000;  wr_data_rom[ 4242]='h00000000;
    rd_cycle[ 4243] = 1'b0;  wr_cycle[ 4243] = 1'b0;  addr_rom[ 4243]='h00000000;  wr_data_rom[ 4243]='h00000000;
    rd_cycle[ 4244] = 1'b0;  wr_cycle[ 4244] = 1'b0;  addr_rom[ 4244]='h00000000;  wr_data_rom[ 4244]='h00000000;
    rd_cycle[ 4245] = 1'b0;  wr_cycle[ 4245] = 1'b0;  addr_rom[ 4245]='h00000000;  wr_data_rom[ 4245]='h00000000;
    rd_cycle[ 4246] = 1'b0;  wr_cycle[ 4246] = 1'b0;  addr_rom[ 4246]='h00000000;  wr_data_rom[ 4246]='h00000000;
    rd_cycle[ 4247] = 1'b0;  wr_cycle[ 4247] = 1'b0;  addr_rom[ 4247]='h00000000;  wr_data_rom[ 4247]='h00000000;
    rd_cycle[ 4248] = 1'b0;  wr_cycle[ 4248] = 1'b0;  addr_rom[ 4248]='h00000000;  wr_data_rom[ 4248]='h00000000;
    rd_cycle[ 4249] = 1'b0;  wr_cycle[ 4249] = 1'b0;  addr_rom[ 4249]='h00000000;  wr_data_rom[ 4249]='h00000000;
    rd_cycle[ 4250] = 1'b0;  wr_cycle[ 4250] = 1'b0;  addr_rom[ 4250]='h00000000;  wr_data_rom[ 4250]='h00000000;
    rd_cycle[ 4251] = 1'b0;  wr_cycle[ 4251] = 1'b0;  addr_rom[ 4251]='h00000000;  wr_data_rom[ 4251]='h00000000;
    rd_cycle[ 4252] = 1'b0;  wr_cycle[ 4252] = 1'b0;  addr_rom[ 4252]='h00000000;  wr_data_rom[ 4252]='h00000000;
    rd_cycle[ 4253] = 1'b0;  wr_cycle[ 4253] = 1'b0;  addr_rom[ 4253]='h00000000;  wr_data_rom[ 4253]='h00000000;
    rd_cycle[ 4254] = 1'b0;  wr_cycle[ 4254] = 1'b0;  addr_rom[ 4254]='h00000000;  wr_data_rom[ 4254]='h00000000;
    rd_cycle[ 4255] = 1'b0;  wr_cycle[ 4255] = 1'b0;  addr_rom[ 4255]='h00000000;  wr_data_rom[ 4255]='h00000000;
    rd_cycle[ 4256] = 1'b0;  wr_cycle[ 4256] = 1'b0;  addr_rom[ 4256]='h00000000;  wr_data_rom[ 4256]='h00000000;
    rd_cycle[ 4257] = 1'b0;  wr_cycle[ 4257] = 1'b0;  addr_rom[ 4257]='h00000000;  wr_data_rom[ 4257]='h00000000;
    rd_cycle[ 4258] = 1'b0;  wr_cycle[ 4258] = 1'b0;  addr_rom[ 4258]='h00000000;  wr_data_rom[ 4258]='h00000000;
    rd_cycle[ 4259] = 1'b0;  wr_cycle[ 4259] = 1'b0;  addr_rom[ 4259]='h00000000;  wr_data_rom[ 4259]='h00000000;
    rd_cycle[ 4260] = 1'b0;  wr_cycle[ 4260] = 1'b0;  addr_rom[ 4260]='h00000000;  wr_data_rom[ 4260]='h00000000;
    rd_cycle[ 4261] = 1'b0;  wr_cycle[ 4261] = 1'b0;  addr_rom[ 4261]='h00000000;  wr_data_rom[ 4261]='h00000000;
    rd_cycle[ 4262] = 1'b0;  wr_cycle[ 4262] = 1'b0;  addr_rom[ 4262]='h00000000;  wr_data_rom[ 4262]='h00000000;
    rd_cycle[ 4263] = 1'b0;  wr_cycle[ 4263] = 1'b0;  addr_rom[ 4263]='h00000000;  wr_data_rom[ 4263]='h00000000;
    rd_cycle[ 4264] = 1'b0;  wr_cycle[ 4264] = 1'b0;  addr_rom[ 4264]='h00000000;  wr_data_rom[ 4264]='h00000000;
    rd_cycle[ 4265] = 1'b0;  wr_cycle[ 4265] = 1'b0;  addr_rom[ 4265]='h00000000;  wr_data_rom[ 4265]='h00000000;
    rd_cycle[ 4266] = 1'b0;  wr_cycle[ 4266] = 1'b0;  addr_rom[ 4266]='h00000000;  wr_data_rom[ 4266]='h00000000;
    rd_cycle[ 4267] = 1'b0;  wr_cycle[ 4267] = 1'b0;  addr_rom[ 4267]='h00000000;  wr_data_rom[ 4267]='h00000000;
    rd_cycle[ 4268] = 1'b0;  wr_cycle[ 4268] = 1'b0;  addr_rom[ 4268]='h00000000;  wr_data_rom[ 4268]='h00000000;
    rd_cycle[ 4269] = 1'b0;  wr_cycle[ 4269] = 1'b0;  addr_rom[ 4269]='h00000000;  wr_data_rom[ 4269]='h00000000;
    rd_cycle[ 4270] = 1'b0;  wr_cycle[ 4270] = 1'b0;  addr_rom[ 4270]='h00000000;  wr_data_rom[ 4270]='h00000000;
    rd_cycle[ 4271] = 1'b0;  wr_cycle[ 4271] = 1'b0;  addr_rom[ 4271]='h00000000;  wr_data_rom[ 4271]='h00000000;
    rd_cycle[ 4272] = 1'b0;  wr_cycle[ 4272] = 1'b0;  addr_rom[ 4272]='h00000000;  wr_data_rom[ 4272]='h00000000;
    rd_cycle[ 4273] = 1'b0;  wr_cycle[ 4273] = 1'b0;  addr_rom[ 4273]='h00000000;  wr_data_rom[ 4273]='h00000000;
    rd_cycle[ 4274] = 1'b0;  wr_cycle[ 4274] = 1'b0;  addr_rom[ 4274]='h00000000;  wr_data_rom[ 4274]='h00000000;
    rd_cycle[ 4275] = 1'b0;  wr_cycle[ 4275] = 1'b0;  addr_rom[ 4275]='h00000000;  wr_data_rom[ 4275]='h00000000;
    rd_cycle[ 4276] = 1'b0;  wr_cycle[ 4276] = 1'b0;  addr_rom[ 4276]='h00000000;  wr_data_rom[ 4276]='h00000000;
    rd_cycle[ 4277] = 1'b0;  wr_cycle[ 4277] = 1'b0;  addr_rom[ 4277]='h00000000;  wr_data_rom[ 4277]='h00000000;
    rd_cycle[ 4278] = 1'b0;  wr_cycle[ 4278] = 1'b0;  addr_rom[ 4278]='h00000000;  wr_data_rom[ 4278]='h00000000;
    rd_cycle[ 4279] = 1'b0;  wr_cycle[ 4279] = 1'b0;  addr_rom[ 4279]='h00000000;  wr_data_rom[ 4279]='h00000000;
    rd_cycle[ 4280] = 1'b0;  wr_cycle[ 4280] = 1'b0;  addr_rom[ 4280]='h00000000;  wr_data_rom[ 4280]='h00000000;
    rd_cycle[ 4281] = 1'b0;  wr_cycle[ 4281] = 1'b0;  addr_rom[ 4281]='h00000000;  wr_data_rom[ 4281]='h00000000;
    rd_cycle[ 4282] = 1'b0;  wr_cycle[ 4282] = 1'b0;  addr_rom[ 4282]='h00000000;  wr_data_rom[ 4282]='h00000000;
    rd_cycle[ 4283] = 1'b0;  wr_cycle[ 4283] = 1'b0;  addr_rom[ 4283]='h00000000;  wr_data_rom[ 4283]='h00000000;
    rd_cycle[ 4284] = 1'b0;  wr_cycle[ 4284] = 1'b0;  addr_rom[ 4284]='h00000000;  wr_data_rom[ 4284]='h00000000;
    rd_cycle[ 4285] = 1'b0;  wr_cycle[ 4285] = 1'b0;  addr_rom[ 4285]='h00000000;  wr_data_rom[ 4285]='h00000000;
    rd_cycle[ 4286] = 1'b0;  wr_cycle[ 4286] = 1'b0;  addr_rom[ 4286]='h00000000;  wr_data_rom[ 4286]='h00000000;
    rd_cycle[ 4287] = 1'b0;  wr_cycle[ 4287] = 1'b0;  addr_rom[ 4287]='h00000000;  wr_data_rom[ 4287]='h00000000;
    rd_cycle[ 4288] = 1'b0;  wr_cycle[ 4288] = 1'b0;  addr_rom[ 4288]='h00000000;  wr_data_rom[ 4288]='h00000000;
    rd_cycle[ 4289] = 1'b0;  wr_cycle[ 4289] = 1'b0;  addr_rom[ 4289]='h00000000;  wr_data_rom[ 4289]='h00000000;
    rd_cycle[ 4290] = 1'b0;  wr_cycle[ 4290] = 1'b0;  addr_rom[ 4290]='h00000000;  wr_data_rom[ 4290]='h00000000;
    rd_cycle[ 4291] = 1'b0;  wr_cycle[ 4291] = 1'b0;  addr_rom[ 4291]='h00000000;  wr_data_rom[ 4291]='h00000000;
    rd_cycle[ 4292] = 1'b0;  wr_cycle[ 4292] = 1'b0;  addr_rom[ 4292]='h00000000;  wr_data_rom[ 4292]='h00000000;
    rd_cycle[ 4293] = 1'b0;  wr_cycle[ 4293] = 1'b0;  addr_rom[ 4293]='h00000000;  wr_data_rom[ 4293]='h00000000;
    rd_cycle[ 4294] = 1'b0;  wr_cycle[ 4294] = 1'b0;  addr_rom[ 4294]='h00000000;  wr_data_rom[ 4294]='h00000000;
    rd_cycle[ 4295] = 1'b0;  wr_cycle[ 4295] = 1'b0;  addr_rom[ 4295]='h00000000;  wr_data_rom[ 4295]='h00000000;
    rd_cycle[ 4296] = 1'b0;  wr_cycle[ 4296] = 1'b0;  addr_rom[ 4296]='h00000000;  wr_data_rom[ 4296]='h00000000;
    rd_cycle[ 4297] = 1'b0;  wr_cycle[ 4297] = 1'b0;  addr_rom[ 4297]='h00000000;  wr_data_rom[ 4297]='h00000000;
    rd_cycle[ 4298] = 1'b0;  wr_cycle[ 4298] = 1'b0;  addr_rom[ 4298]='h00000000;  wr_data_rom[ 4298]='h00000000;
    rd_cycle[ 4299] = 1'b0;  wr_cycle[ 4299] = 1'b0;  addr_rom[ 4299]='h00000000;  wr_data_rom[ 4299]='h00000000;
    rd_cycle[ 4300] = 1'b0;  wr_cycle[ 4300] = 1'b0;  addr_rom[ 4300]='h00000000;  wr_data_rom[ 4300]='h00000000;
    rd_cycle[ 4301] = 1'b0;  wr_cycle[ 4301] = 1'b0;  addr_rom[ 4301]='h00000000;  wr_data_rom[ 4301]='h00000000;
    rd_cycle[ 4302] = 1'b0;  wr_cycle[ 4302] = 1'b0;  addr_rom[ 4302]='h00000000;  wr_data_rom[ 4302]='h00000000;
    rd_cycle[ 4303] = 1'b0;  wr_cycle[ 4303] = 1'b0;  addr_rom[ 4303]='h00000000;  wr_data_rom[ 4303]='h00000000;
    rd_cycle[ 4304] = 1'b0;  wr_cycle[ 4304] = 1'b0;  addr_rom[ 4304]='h00000000;  wr_data_rom[ 4304]='h00000000;
    rd_cycle[ 4305] = 1'b0;  wr_cycle[ 4305] = 1'b0;  addr_rom[ 4305]='h00000000;  wr_data_rom[ 4305]='h00000000;
    rd_cycle[ 4306] = 1'b0;  wr_cycle[ 4306] = 1'b0;  addr_rom[ 4306]='h00000000;  wr_data_rom[ 4306]='h00000000;
    rd_cycle[ 4307] = 1'b0;  wr_cycle[ 4307] = 1'b0;  addr_rom[ 4307]='h00000000;  wr_data_rom[ 4307]='h00000000;
    rd_cycle[ 4308] = 1'b0;  wr_cycle[ 4308] = 1'b0;  addr_rom[ 4308]='h00000000;  wr_data_rom[ 4308]='h00000000;
    rd_cycle[ 4309] = 1'b0;  wr_cycle[ 4309] = 1'b0;  addr_rom[ 4309]='h00000000;  wr_data_rom[ 4309]='h00000000;
    rd_cycle[ 4310] = 1'b0;  wr_cycle[ 4310] = 1'b0;  addr_rom[ 4310]='h00000000;  wr_data_rom[ 4310]='h00000000;
    rd_cycle[ 4311] = 1'b0;  wr_cycle[ 4311] = 1'b0;  addr_rom[ 4311]='h00000000;  wr_data_rom[ 4311]='h00000000;
    rd_cycle[ 4312] = 1'b0;  wr_cycle[ 4312] = 1'b0;  addr_rom[ 4312]='h00000000;  wr_data_rom[ 4312]='h00000000;
    rd_cycle[ 4313] = 1'b0;  wr_cycle[ 4313] = 1'b0;  addr_rom[ 4313]='h00000000;  wr_data_rom[ 4313]='h00000000;
    rd_cycle[ 4314] = 1'b0;  wr_cycle[ 4314] = 1'b0;  addr_rom[ 4314]='h00000000;  wr_data_rom[ 4314]='h00000000;
    rd_cycle[ 4315] = 1'b0;  wr_cycle[ 4315] = 1'b0;  addr_rom[ 4315]='h00000000;  wr_data_rom[ 4315]='h00000000;
    rd_cycle[ 4316] = 1'b0;  wr_cycle[ 4316] = 1'b0;  addr_rom[ 4316]='h00000000;  wr_data_rom[ 4316]='h00000000;
    rd_cycle[ 4317] = 1'b0;  wr_cycle[ 4317] = 1'b0;  addr_rom[ 4317]='h00000000;  wr_data_rom[ 4317]='h00000000;
    rd_cycle[ 4318] = 1'b0;  wr_cycle[ 4318] = 1'b0;  addr_rom[ 4318]='h00000000;  wr_data_rom[ 4318]='h00000000;
    rd_cycle[ 4319] = 1'b0;  wr_cycle[ 4319] = 1'b0;  addr_rom[ 4319]='h00000000;  wr_data_rom[ 4319]='h00000000;
    rd_cycle[ 4320] = 1'b0;  wr_cycle[ 4320] = 1'b0;  addr_rom[ 4320]='h00000000;  wr_data_rom[ 4320]='h00000000;
    rd_cycle[ 4321] = 1'b0;  wr_cycle[ 4321] = 1'b0;  addr_rom[ 4321]='h00000000;  wr_data_rom[ 4321]='h00000000;
    rd_cycle[ 4322] = 1'b0;  wr_cycle[ 4322] = 1'b0;  addr_rom[ 4322]='h00000000;  wr_data_rom[ 4322]='h00000000;
    rd_cycle[ 4323] = 1'b0;  wr_cycle[ 4323] = 1'b0;  addr_rom[ 4323]='h00000000;  wr_data_rom[ 4323]='h00000000;
    rd_cycle[ 4324] = 1'b0;  wr_cycle[ 4324] = 1'b0;  addr_rom[ 4324]='h00000000;  wr_data_rom[ 4324]='h00000000;
    rd_cycle[ 4325] = 1'b0;  wr_cycle[ 4325] = 1'b0;  addr_rom[ 4325]='h00000000;  wr_data_rom[ 4325]='h00000000;
    rd_cycle[ 4326] = 1'b0;  wr_cycle[ 4326] = 1'b0;  addr_rom[ 4326]='h00000000;  wr_data_rom[ 4326]='h00000000;
    rd_cycle[ 4327] = 1'b0;  wr_cycle[ 4327] = 1'b0;  addr_rom[ 4327]='h00000000;  wr_data_rom[ 4327]='h00000000;
    rd_cycle[ 4328] = 1'b0;  wr_cycle[ 4328] = 1'b0;  addr_rom[ 4328]='h00000000;  wr_data_rom[ 4328]='h00000000;
    rd_cycle[ 4329] = 1'b0;  wr_cycle[ 4329] = 1'b0;  addr_rom[ 4329]='h00000000;  wr_data_rom[ 4329]='h00000000;
    rd_cycle[ 4330] = 1'b0;  wr_cycle[ 4330] = 1'b0;  addr_rom[ 4330]='h00000000;  wr_data_rom[ 4330]='h00000000;
    rd_cycle[ 4331] = 1'b0;  wr_cycle[ 4331] = 1'b0;  addr_rom[ 4331]='h00000000;  wr_data_rom[ 4331]='h00000000;
    rd_cycle[ 4332] = 1'b0;  wr_cycle[ 4332] = 1'b0;  addr_rom[ 4332]='h00000000;  wr_data_rom[ 4332]='h00000000;
    rd_cycle[ 4333] = 1'b0;  wr_cycle[ 4333] = 1'b0;  addr_rom[ 4333]='h00000000;  wr_data_rom[ 4333]='h00000000;
    rd_cycle[ 4334] = 1'b0;  wr_cycle[ 4334] = 1'b0;  addr_rom[ 4334]='h00000000;  wr_data_rom[ 4334]='h00000000;
    rd_cycle[ 4335] = 1'b0;  wr_cycle[ 4335] = 1'b0;  addr_rom[ 4335]='h00000000;  wr_data_rom[ 4335]='h00000000;
    rd_cycle[ 4336] = 1'b0;  wr_cycle[ 4336] = 1'b0;  addr_rom[ 4336]='h00000000;  wr_data_rom[ 4336]='h00000000;
    rd_cycle[ 4337] = 1'b0;  wr_cycle[ 4337] = 1'b0;  addr_rom[ 4337]='h00000000;  wr_data_rom[ 4337]='h00000000;
    rd_cycle[ 4338] = 1'b0;  wr_cycle[ 4338] = 1'b0;  addr_rom[ 4338]='h00000000;  wr_data_rom[ 4338]='h00000000;
    rd_cycle[ 4339] = 1'b0;  wr_cycle[ 4339] = 1'b0;  addr_rom[ 4339]='h00000000;  wr_data_rom[ 4339]='h00000000;
    rd_cycle[ 4340] = 1'b0;  wr_cycle[ 4340] = 1'b0;  addr_rom[ 4340]='h00000000;  wr_data_rom[ 4340]='h00000000;
    rd_cycle[ 4341] = 1'b0;  wr_cycle[ 4341] = 1'b0;  addr_rom[ 4341]='h00000000;  wr_data_rom[ 4341]='h00000000;
    rd_cycle[ 4342] = 1'b0;  wr_cycle[ 4342] = 1'b0;  addr_rom[ 4342]='h00000000;  wr_data_rom[ 4342]='h00000000;
    rd_cycle[ 4343] = 1'b0;  wr_cycle[ 4343] = 1'b0;  addr_rom[ 4343]='h00000000;  wr_data_rom[ 4343]='h00000000;
    rd_cycle[ 4344] = 1'b0;  wr_cycle[ 4344] = 1'b0;  addr_rom[ 4344]='h00000000;  wr_data_rom[ 4344]='h00000000;
    rd_cycle[ 4345] = 1'b0;  wr_cycle[ 4345] = 1'b0;  addr_rom[ 4345]='h00000000;  wr_data_rom[ 4345]='h00000000;
    rd_cycle[ 4346] = 1'b0;  wr_cycle[ 4346] = 1'b0;  addr_rom[ 4346]='h00000000;  wr_data_rom[ 4346]='h00000000;
    rd_cycle[ 4347] = 1'b0;  wr_cycle[ 4347] = 1'b0;  addr_rom[ 4347]='h00000000;  wr_data_rom[ 4347]='h00000000;
    rd_cycle[ 4348] = 1'b0;  wr_cycle[ 4348] = 1'b0;  addr_rom[ 4348]='h00000000;  wr_data_rom[ 4348]='h00000000;
    rd_cycle[ 4349] = 1'b0;  wr_cycle[ 4349] = 1'b0;  addr_rom[ 4349]='h00000000;  wr_data_rom[ 4349]='h00000000;
    rd_cycle[ 4350] = 1'b0;  wr_cycle[ 4350] = 1'b0;  addr_rom[ 4350]='h00000000;  wr_data_rom[ 4350]='h00000000;
    rd_cycle[ 4351] = 1'b0;  wr_cycle[ 4351] = 1'b0;  addr_rom[ 4351]='h00000000;  wr_data_rom[ 4351]='h00000000;
    rd_cycle[ 4352] = 1'b0;  wr_cycle[ 4352] = 1'b0;  addr_rom[ 4352]='h00000000;  wr_data_rom[ 4352]='h00000000;
    rd_cycle[ 4353] = 1'b0;  wr_cycle[ 4353] = 1'b0;  addr_rom[ 4353]='h00000000;  wr_data_rom[ 4353]='h00000000;
    rd_cycle[ 4354] = 1'b0;  wr_cycle[ 4354] = 1'b0;  addr_rom[ 4354]='h00000000;  wr_data_rom[ 4354]='h00000000;
    rd_cycle[ 4355] = 1'b0;  wr_cycle[ 4355] = 1'b0;  addr_rom[ 4355]='h00000000;  wr_data_rom[ 4355]='h00000000;
    rd_cycle[ 4356] = 1'b0;  wr_cycle[ 4356] = 1'b0;  addr_rom[ 4356]='h00000000;  wr_data_rom[ 4356]='h00000000;
    rd_cycle[ 4357] = 1'b0;  wr_cycle[ 4357] = 1'b0;  addr_rom[ 4357]='h00000000;  wr_data_rom[ 4357]='h00000000;
    rd_cycle[ 4358] = 1'b0;  wr_cycle[ 4358] = 1'b0;  addr_rom[ 4358]='h00000000;  wr_data_rom[ 4358]='h00000000;
    rd_cycle[ 4359] = 1'b0;  wr_cycle[ 4359] = 1'b0;  addr_rom[ 4359]='h00000000;  wr_data_rom[ 4359]='h00000000;
    rd_cycle[ 4360] = 1'b0;  wr_cycle[ 4360] = 1'b0;  addr_rom[ 4360]='h00000000;  wr_data_rom[ 4360]='h00000000;
    rd_cycle[ 4361] = 1'b0;  wr_cycle[ 4361] = 1'b0;  addr_rom[ 4361]='h00000000;  wr_data_rom[ 4361]='h00000000;
    rd_cycle[ 4362] = 1'b0;  wr_cycle[ 4362] = 1'b0;  addr_rom[ 4362]='h00000000;  wr_data_rom[ 4362]='h00000000;
    rd_cycle[ 4363] = 1'b0;  wr_cycle[ 4363] = 1'b0;  addr_rom[ 4363]='h00000000;  wr_data_rom[ 4363]='h00000000;
    rd_cycle[ 4364] = 1'b0;  wr_cycle[ 4364] = 1'b0;  addr_rom[ 4364]='h00000000;  wr_data_rom[ 4364]='h00000000;
    rd_cycle[ 4365] = 1'b0;  wr_cycle[ 4365] = 1'b0;  addr_rom[ 4365]='h00000000;  wr_data_rom[ 4365]='h00000000;
    rd_cycle[ 4366] = 1'b0;  wr_cycle[ 4366] = 1'b0;  addr_rom[ 4366]='h00000000;  wr_data_rom[ 4366]='h00000000;
    rd_cycle[ 4367] = 1'b0;  wr_cycle[ 4367] = 1'b0;  addr_rom[ 4367]='h00000000;  wr_data_rom[ 4367]='h00000000;
    rd_cycle[ 4368] = 1'b0;  wr_cycle[ 4368] = 1'b0;  addr_rom[ 4368]='h00000000;  wr_data_rom[ 4368]='h00000000;
    rd_cycle[ 4369] = 1'b0;  wr_cycle[ 4369] = 1'b0;  addr_rom[ 4369]='h00000000;  wr_data_rom[ 4369]='h00000000;
    rd_cycle[ 4370] = 1'b0;  wr_cycle[ 4370] = 1'b0;  addr_rom[ 4370]='h00000000;  wr_data_rom[ 4370]='h00000000;
    rd_cycle[ 4371] = 1'b0;  wr_cycle[ 4371] = 1'b0;  addr_rom[ 4371]='h00000000;  wr_data_rom[ 4371]='h00000000;
    rd_cycle[ 4372] = 1'b0;  wr_cycle[ 4372] = 1'b0;  addr_rom[ 4372]='h00000000;  wr_data_rom[ 4372]='h00000000;
    rd_cycle[ 4373] = 1'b0;  wr_cycle[ 4373] = 1'b0;  addr_rom[ 4373]='h00000000;  wr_data_rom[ 4373]='h00000000;
    rd_cycle[ 4374] = 1'b0;  wr_cycle[ 4374] = 1'b0;  addr_rom[ 4374]='h00000000;  wr_data_rom[ 4374]='h00000000;
    rd_cycle[ 4375] = 1'b0;  wr_cycle[ 4375] = 1'b0;  addr_rom[ 4375]='h00000000;  wr_data_rom[ 4375]='h00000000;
    rd_cycle[ 4376] = 1'b0;  wr_cycle[ 4376] = 1'b0;  addr_rom[ 4376]='h00000000;  wr_data_rom[ 4376]='h00000000;
    rd_cycle[ 4377] = 1'b0;  wr_cycle[ 4377] = 1'b0;  addr_rom[ 4377]='h00000000;  wr_data_rom[ 4377]='h00000000;
    rd_cycle[ 4378] = 1'b0;  wr_cycle[ 4378] = 1'b0;  addr_rom[ 4378]='h00000000;  wr_data_rom[ 4378]='h00000000;
    rd_cycle[ 4379] = 1'b0;  wr_cycle[ 4379] = 1'b0;  addr_rom[ 4379]='h00000000;  wr_data_rom[ 4379]='h00000000;
    rd_cycle[ 4380] = 1'b0;  wr_cycle[ 4380] = 1'b0;  addr_rom[ 4380]='h00000000;  wr_data_rom[ 4380]='h00000000;
    rd_cycle[ 4381] = 1'b0;  wr_cycle[ 4381] = 1'b0;  addr_rom[ 4381]='h00000000;  wr_data_rom[ 4381]='h00000000;
    rd_cycle[ 4382] = 1'b0;  wr_cycle[ 4382] = 1'b0;  addr_rom[ 4382]='h00000000;  wr_data_rom[ 4382]='h00000000;
    rd_cycle[ 4383] = 1'b0;  wr_cycle[ 4383] = 1'b0;  addr_rom[ 4383]='h00000000;  wr_data_rom[ 4383]='h00000000;
    rd_cycle[ 4384] = 1'b0;  wr_cycle[ 4384] = 1'b0;  addr_rom[ 4384]='h00000000;  wr_data_rom[ 4384]='h00000000;
    rd_cycle[ 4385] = 1'b0;  wr_cycle[ 4385] = 1'b0;  addr_rom[ 4385]='h00000000;  wr_data_rom[ 4385]='h00000000;
    rd_cycle[ 4386] = 1'b0;  wr_cycle[ 4386] = 1'b0;  addr_rom[ 4386]='h00000000;  wr_data_rom[ 4386]='h00000000;
    rd_cycle[ 4387] = 1'b0;  wr_cycle[ 4387] = 1'b0;  addr_rom[ 4387]='h00000000;  wr_data_rom[ 4387]='h00000000;
    rd_cycle[ 4388] = 1'b0;  wr_cycle[ 4388] = 1'b0;  addr_rom[ 4388]='h00000000;  wr_data_rom[ 4388]='h00000000;
    rd_cycle[ 4389] = 1'b0;  wr_cycle[ 4389] = 1'b0;  addr_rom[ 4389]='h00000000;  wr_data_rom[ 4389]='h00000000;
    rd_cycle[ 4390] = 1'b0;  wr_cycle[ 4390] = 1'b0;  addr_rom[ 4390]='h00000000;  wr_data_rom[ 4390]='h00000000;
    rd_cycle[ 4391] = 1'b0;  wr_cycle[ 4391] = 1'b0;  addr_rom[ 4391]='h00000000;  wr_data_rom[ 4391]='h00000000;
    rd_cycle[ 4392] = 1'b0;  wr_cycle[ 4392] = 1'b0;  addr_rom[ 4392]='h00000000;  wr_data_rom[ 4392]='h00000000;
    rd_cycle[ 4393] = 1'b0;  wr_cycle[ 4393] = 1'b0;  addr_rom[ 4393]='h00000000;  wr_data_rom[ 4393]='h00000000;
    rd_cycle[ 4394] = 1'b0;  wr_cycle[ 4394] = 1'b0;  addr_rom[ 4394]='h00000000;  wr_data_rom[ 4394]='h00000000;
    rd_cycle[ 4395] = 1'b0;  wr_cycle[ 4395] = 1'b0;  addr_rom[ 4395]='h00000000;  wr_data_rom[ 4395]='h00000000;
    rd_cycle[ 4396] = 1'b0;  wr_cycle[ 4396] = 1'b0;  addr_rom[ 4396]='h00000000;  wr_data_rom[ 4396]='h00000000;
    rd_cycle[ 4397] = 1'b0;  wr_cycle[ 4397] = 1'b0;  addr_rom[ 4397]='h00000000;  wr_data_rom[ 4397]='h00000000;
    rd_cycle[ 4398] = 1'b0;  wr_cycle[ 4398] = 1'b0;  addr_rom[ 4398]='h00000000;  wr_data_rom[ 4398]='h00000000;
    rd_cycle[ 4399] = 1'b0;  wr_cycle[ 4399] = 1'b0;  addr_rom[ 4399]='h00000000;  wr_data_rom[ 4399]='h00000000;
    rd_cycle[ 4400] = 1'b0;  wr_cycle[ 4400] = 1'b0;  addr_rom[ 4400]='h00000000;  wr_data_rom[ 4400]='h00000000;
    rd_cycle[ 4401] = 1'b0;  wr_cycle[ 4401] = 1'b0;  addr_rom[ 4401]='h00000000;  wr_data_rom[ 4401]='h00000000;
    rd_cycle[ 4402] = 1'b0;  wr_cycle[ 4402] = 1'b0;  addr_rom[ 4402]='h00000000;  wr_data_rom[ 4402]='h00000000;
    rd_cycle[ 4403] = 1'b0;  wr_cycle[ 4403] = 1'b0;  addr_rom[ 4403]='h00000000;  wr_data_rom[ 4403]='h00000000;
    rd_cycle[ 4404] = 1'b0;  wr_cycle[ 4404] = 1'b0;  addr_rom[ 4404]='h00000000;  wr_data_rom[ 4404]='h00000000;
    rd_cycle[ 4405] = 1'b0;  wr_cycle[ 4405] = 1'b0;  addr_rom[ 4405]='h00000000;  wr_data_rom[ 4405]='h00000000;
    rd_cycle[ 4406] = 1'b0;  wr_cycle[ 4406] = 1'b0;  addr_rom[ 4406]='h00000000;  wr_data_rom[ 4406]='h00000000;
    rd_cycle[ 4407] = 1'b0;  wr_cycle[ 4407] = 1'b0;  addr_rom[ 4407]='h00000000;  wr_data_rom[ 4407]='h00000000;
    rd_cycle[ 4408] = 1'b0;  wr_cycle[ 4408] = 1'b0;  addr_rom[ 4408]='h00000000;  wr_data_rom[ 4408]='h00000000;
    rd_cycle[ 4409] = 1'b0;  wr_cycle[ 4409] = 1'b0;  addr_rom[ 4409]='h00000000;  wr_data_rom[ 4409]='h00000000;
    rd_cycle[ 4410] = 1'b0;  wr_cycle[ 4410] = 1'b0;  addr_rom[ 4410]='h00000000;  wr_data_rom[ 4410]='h00000000;
    rd_cycle[ 4411] = 1'b0;  wr_cycle[ 4411] = 1'b0;  addr_rom[ 4411]='h00000000;  wr_data_rom[ 4411]='h00000000;
    rd_cycle[ 4412] = 1'b0;  wr_cycle[ 4412] = 1'b0;  addr_rom[ 4412]='h00000000;  wr_data_rom[ 4412]='h00000000;
    rd_cycle[ 4413] = 1'b0;  wr_cycle[ 4413] = 1'b0;  addr_rom[ 4413]='h00000000;  wr_data_rom[ 4413]='h00000000;
    rd_cycle[ 4414] = 1'b0;  wr_cycle[ 4414] = 1'b0;  addr_rom[ 4414]='h00000000;  wr_data_rom[ 4414]='h00000000;
    rd_cycle[ 4415] = 1'b0;  wr_cycle[ 4415] = 1'b0;  addr_rom[ 4415]='h00000000;  wr_data_rom[ 4415]='h00000000;
    rd_cycle[ 4416] = 1'b0;  wr_cycle[ 4416] = 1'b0;  addr_rom[ 4416]='h00000000;  wr_data_rom[ 4416]='h00000000;
    rd_cycle[ 4417] = 1'b0;  wr_cycle[ 4417] = 1'b0;  addr_rom[ 4417]='h00000000;  wr_data_rom[ 4417]='h00000000;
    rd_cycle[ 4418] = 1'b0;  wr_cycle[ 4418] = 1'b0;  addr_rom[ 4418]='h00000000;  wr_data_rom[ 4418]='h00000000;
    rd_cycle[ 4419] = 1'b0;  wr_cycle[ 4419] = 1'b0;  addr_rom[ 4419]='h00000000;  wr_data_rom[ 4419]='h00000000;
    rd_cycle[ 4420] = 1'b0;  wr_cycle[ 4420] = 1'b0;  addr_rom[ 4420]='h00000000;  wr_data_rom[ 4420]='h00000000;
    rd_cycle[ 4421] = 1'b0;  wr_cycle[ 4421] = 1'b0;  addr_rom[ 4421]='h00000000;  wr_data_rom[ 4421]='h00000000;
    rd_cycle[ 4422] = 1'b0;  wr_cycle[ 4422] = 1'b0;  addr_rom[ 4422]='h00000000;  wr_data_rom[ 4422]='h00000000;
    rd_cycle[ 4423] = 1'b0;  wr_cycle[ 4423] = 1'b0;  addr_rom[ 4423]='h00000000;  wr_data_rom[ 4423]='h00000000;
    rd_cycle[ 4424] = 1'b0;  wr_cycle[ 4424] = 1'b0;  addr_rom[ 4424]='h00000000;  wr_data_rom[ 4424]='h00000000;
    rd_cycle[ 4425] = 1'b0;  wr_cycle[ 4425] = 1'b0;  addr_rom[ 4425]='h00000000;  wr_data_rom[ 4425]='h00000000;
    rd_cycle[ 4426] = 1'b0;  wr_cycle[ 4426] = 1'b0;  addr_rom[ 4426]='h00000000;  wr_data_rom[ 4426]='h00000000;
    rd_cycle[ 4427] = 1'b0;  wr_cycle[ 4427] = 1'b0;  addr_rom[ 4427]='h00000000;  wr_data_rom[ 4427]='h00000000;
    rd_cycle[ 4428] = 1'b0;  wr_cycle[ 4428] = 1'b0;  addr_rom[ 4428]='h00000000;  wr_data_rom[ 4428]='h00000000;
    rd_cycle[ 4429] = 1'b0;  wr_cycle[ 4429] = 1'b0;  addr_rom[ 4429]='h00000000;  wr_data_rom[ 4429]='h00000000;
    rd_cycle[ 4430] = 1'b0;  wr_cycle[ 4430] = 1'b0;  addr_rom[ 4430]='h00000000;  wr_data_rom[ 4430]='h00000000;
    rd_cycle[ 4431] = 1'b0;  wr_cycle[ 4431] = 1'b0;  addr_rom[ 4431]='h00000000;  wr_data_rom[ 4431]='h00000000;
    rd_cycle[ 4432] = 1'b0;  wr_cycle[ 4432] = 1'b0;  addr_rom[ 4432]='h00000000;  wr_data_rom[ 4432]='h00000000;
    rd_cycle[ 4433] = 1'b0;  wr_cycle[ 4433] = 1'b0;  addr_rom[ 4433]='h00000000;  wr_data_rom[ 4433]='h00000000;
    rd_cycle[ 4434] = 1'b0;  wr_cycle[ 4434] = 1'b0;  addr_rom[ 4434]='h00000000;  wr_data_rom[ 4434]='h00000000;
    rd_cycle[ 4435] = 1'b0;  wr_cycle[ 4435] = 1'b0;  addr_rom[ 4435]='h00000000;  wr_data_rom[ 4435]='h00000000;
    rd_cycle[ 4436] = 1'b0;  wr_cycle[ 4436] = 1'b0;  addr_rom[ 4436]='h00000000;  wr_data_rom[ 4436]='h00000000;
    rd_cycle[ 4437] = 1'b0;  wr_cycle[ 4437] = 1'b0;  addr_rom[ 4437]='h00000000;  wr_data_rom[ 4437]='h00000000;
    rd_cycle[ 4438] = 1'b0;  wr_cycle[ 4438] = 1'b0;  addr_rom[ 4438]='h00000000;  wr_data_rom[ 4438]='h00000000;
    rd_cycle[ 4439] = 1'b0;  wr_cycle[ 4439] = 1'b0;  addr_rom[ 4439]='h00000000;  wr_data_rom[ 4439]='h00000000;
    rd_cycle[ 4440] = 1'b0;  wr_cycle[ 4440] = 1'b0;  addr_rom[ 4440]='h00000000;  wr_data_rom[ 4440]='h00000000;
    rd_cycle[ 4441] = 1'b0;  wr_cycle[ 4441] = 1'b0;  addr_rom[ 4441]='h00000000;  wr_data_rom[ 4441]='h00000000;
    rd_cycle[ 4442] = 1'b0;  wr_cycle[ 4442] = 1'b0;  addr_rom[ 4442]='h00000000;  wr_data_rom[ 4442]='h00000000;
    rd_cycle[ 4443] = 1'b0;  wr_cycle[ 4443] = 1'b0;  addr_rom[ 4443]='h00000000;  wr_data_rom[ 4443]='h00000000;
    rd_cycle[ 4444] = 1'b0;  wr_cycle[ 4444] = 1'b0;  addr_rom[ 4444]='h00000000;  wr_data_rom[ 4444]='h00000000;
    rd_cycle[ 4445] = 1'b0;  wr_cycle[ 4445] = 1'b0;  addr_rom[ 4445]='h00000000;  wr_data_rom[ 4445]='h00000000;
    rd_cycle[ 4446] = 1'b0;  wr_cycle[ 4446] = 1'b0;  addr_rom[ 4446]='h00000000;  wr_data_rom[ 4446]='h00000000;
    rd_cycle[ 4447] = 1'b0;  wr_cycle[ 4447] = 1'b0;  addr_rom[ 4447]='h00000000;  wr_data_rom[ 4447]='h00000000;
    rd_cycle[ 4448] = 1'b0;  wr_cycle[ 4448] = 1'b0;  addr_rom[ 4448]='h00000000;  wr_data_rom[ 4448]='h00000000;
    rd_cycle[ 4449] = 1'b0;  wr_cycle[ 4449] = 1'b0;  addr_rom[ 4449]='h00000000;  wr_data_rom[ 4449]='h00000000;
    rd_cycle[ 4450] = 1'b0;  wr_cycle[ 4450] = 1'b0;  addr_rom[ 4450]='h00000000;  wr_data_rom[ 4450]='h00000000;
    rd_cycle[ 4451] = 1'b0;  wr_cycle[ 4451] = 1'b0;  addr_rom[ 4451]='h00000000;  wr_data_rom[ 4451]='h00000000;
    rd_cycle[ 4452] = 1'b0;  wr_cycle[ 4452] = 1'b0;  addr_rom[ 4452]='h00000000;  wr_data_rom[ 4452]='h00000000;
    rd_cycle[ 4453] = 1'b0;  wr_cycle[ 4453] = 1'b0;  addr_rom[ 4453]='h00000000;  wr_data_rom[ 4453]='h00000000;
    rd_cycle[ 4454] = 1'b0;  wr_cycle[ 4454] = 1'b0;  addr_rom[ 4454]='h00000000;  wr_data_rom[ 4454]='h00000000;
    rd_cycle[ 4455] = 1'b0;  wr_cycle[ 4455] = 1'b0;  addr_rom[ 4455]='h00000000;  wr_data_rom[ 4455]='h00000000;
    rd_cycle[ 4456] = 1'b0;  wr_cycle[ 4456] = 1'b0;  addr_rom[ 4456]='h00000000;  wr_data_rom[ 4456]='h00000000;
    rd_cycle[ 4457] = 1'b0;  wr_cycle[ 4457] = 1'b0;  addr_rom[ 4457]='h00000000;  wr_data_rom[ 4457]='h00000000;
    rd_cycle[ 4458] = 1'b0;  wr_cycle[ 4458] = 1'b0;  addr_rom[ 4458]='h00000000;  wr_data_rom[ 4458]='h00000000;
    rd_cycle[ 4459] = 1'b0;  wr_cycle[ 4459] = 1'b0;  addr_rom[ 4459]='h00000000;  wr_data_rom[ 4459]='h00000000;
    rd_cycle[ 4460] = 1'b0;  wr_cycle[ 4460] = 1'b0;  addr_rom[ 4460]='h00000000;  wr_data_rom[ 4460]='h00000000;
    rd_cycle[ 4461] = 1'b0;  wr_cycle[ 4461] = 1'b0;  addr_rom[ 4461]='h00000000;  wr_data_rom[ 4461]='h00000000;
    rd_cycle[ 4462] = 1'b0;  wr_cycle[ 4462] = 1'b0;  addr_rom[ 4462]='h00000000;  wr_data_rom[ 4462]='h00000000;
    rd_cycle[ 4463] = 1'b0;  wr_cycle[ 4463] = 1'b0;  addr_rom[ 4463]='h00000000;  wr_data_rom[ 4463]='h00000000;
    rd_cycle[ 4464] = 1'b0;  wr_cycle[ 4464] = 1'b0;  addr_rom[ 4464]='h00000000;  wr_data_rom[ 4464]='h00000000;
    rd_cycle[ 4465] = 1'b0;  wr_cycle[ 4465] = 1'b0;  addr_rom[ 4465]='h00000000;  wr_data_rom[ 4465]='h00000000;
    rd_cycle[ 4466] = 1'b0;  wr_cycle[ 4466] = 1'b0;  addr_rom[ 4466]='h00000000;  wr_data_rom[ 4466]='h00000000;
    rd_cycle[ 4467] = 1'b0;  wr_cycle[ 4467] = 1'b0;  addr_rom[ 4467]='h00000000;  wr_data_rom[ 4467]='h00000000;
    rd_cycle[ 4468] = 1'b0;  wr_cycle[ 4468] = 1'b0;  addr_rom[ 4468]='h00000000;  wr_data_rom[ 4468]='h00000000;
    rd_cycle[ 4469] = 1'b0;  wr_cycle[ 4469] = 1'b0;  addr_rom[ 4469]='h00000000;  wr_data_rom[ 4469]='h00000000;
    rd_cycle[ 4470] = 1'b0;  wr_cycle[ 4470] = 1'b0;  addr_rom[ 4470]='h00000000;  wr_data_rom[ 4470]='h00000000;
    rd_cycle[ 4471] = 1'b0;  wr_cycle[ 4471] = 1'b0;  addr_rom[ 4471]='h00000000;  wr_data_rom[ 4471]='h00000000;
    rd_cycle[ 4472] = 1'b0;  wr_cycle[ 4472] = 1'b0;  addr_rom[ 4472]='h00000000;  wr_data_rom[ 4472]='h00000000;
    rd_cycle[ 4473] = 1'b0;  wr_cycle[ 4473] = 1'b0;  addr_rom[ 4473]='h00000000;  wr_data_rom[ 4473]='h00000000;
    rd_cycle[ 4474] = 1'b0;  wr_cycle[ 4474] = 1'b0;  addr_rom[ 4474]='h00000000;  wr_data_rom[ 4474]='h00000000;
    rd_cycle[ 4475] = 1'b0;  wr_cycle[ 4475] = 1'b0;  addr_rom[ 4475]='h00000000;  wr_data_rom[ 4475]='h00000000;
    rd_cycle[ 4476] = 1'b0;  wr_cycle[ 4476] = 1'b0;  addr_rom[ 4476]='h00000000;  wr_data_rom[ 4476]='h00000000;
    rd_cycle[ 4477] = 1'b0;  wr_cycle[ 4477] = 1'b0;  addr_rom[ 4477]='h00000000;  wr_data_rom[ 4477]='h00000000;
    rd_cycle[ 4478] = 1'b0;  wr_cycle[ 4478] = 1'b0;  addr_rom[ 4478]='h00000000;  wr_data_rom[ 4478]='h00000000;
    rd_cycle[ 4479] = 1'b0;  wr_cycle[ 4479] = 1'b0;  addr_rom[ 4479]='h00000000;  wr_data_rom[ 4479]='h00000000;
    rd_cycle[ 4480] = 1'b0;  wr_cycle[ 4480] = 1'b0;  addr_rom[ 4480]='h00000000;  wr_data_rom[ 4480]='h00000000;
    rd_cycle[ 4481] = 1'b0;  wr_cycle[ 4481] = 1'b0;  addr_rom[ 4481]='h00000000;  wr_data_rom[ 4481]='h00000000;
    rd_cycle[ 4482] = 1'b0;  wr_cycle[ 4482] = 1'b0;  addr_rom[ 4482]='h00000000;  wr_data_rom[ 4482]='h00000000;
    rd_cycle[ 4483] = 1'b0;  wr_cycle[ 4483] = 1'b0;  addr_rom[ 4483]='h00000000;  wr_data_rom[ 4483]='h00000000;
    rd_cycle[ 4484] = 1'b0;  wr_cycle[ 4484] = 1'b0;  addr_rom[ 4484]='h00000000;  wr_data_rom[ 4484]='h00000000;
    rd_cycle[ 4485] = 1'b0;  wr_cycle[ 4485] = 1'b0;  addr_rom[ 4485]='h00000000;  wr_data_rom[ 4485]='h00000000;
    rd_cycle[ 4486] = 1'b0;  wr_cycle[ 4486] = 1'b0;  addr_rom[ 4486]='h00000000;  wr_data_rom[ 4486]='h00000000;
    rd_cycle[ 4487] = 1'b0;  wr_cycle[ 4487] = 1'b0;  addr_rom[ 4487]='h00000000;  wr_data_rom[ 4487]='h00000000;
    rd_cycle[ 4488] = 1'b0;  wr_cycle[ 4488] = 1'b0;  addr_rom[ 4488]='h00000000;  wr_data_rom[ 4488]='h00000000;
    rd_cycle[ 4489] = 1'b0;  wr_cycle[ 4489] = 1'b0;  addr_rom[ 4489]='h00000000;  wr_data_rom[ 4489]='h00000000;
    rd_cycle[ 4490] = 1'b0;  wr_cycle[ 4490] = 1'b0;  addr_rom[ 4490]='h00000000;  wr_data_rom[ 4490]='h00000000;
    rd_cycle[ 4491] = 1'b0;  wr_cycle[ 4491] = 1'b0;  addr_rom[ 4491]='h00000000;  wr_data_rom[ 4491]='h00000000;
    rd_cycle[ 4492] = 1'b0;  wr_cycle[ 4492] = 1'b0;  addr_rom[ 4492]='h00000000;  wr_data_rom[ 4492]='h00000000;
    rd_cycle[ 4493] = 1'b0;  wr_cycle[ 4493] = 1'b0;  addr_rom[ 4493]='h00000000;  wr_data_rom[ 4493]='h00000000;
    rd_cycle[ 4494] = 1'b0;  wr_cycle[ 4494] = 1'b0;  addr_rom[ 4494]='h00000000;  wr_data_rom[ 4494]='h00000000;
    rd_cycle[ 4495] = 1'b0;  wr_cycle[ 4495] = 1'b0;  addr_rom[ 4495]='h00000000;  wr_data_rom[ 4495]='h00000000;
    rd_cycle[ 4496] = 1'b0;  wr_cycle[ 4496] = 1'b0;  addr_rom[ 4496]='h00000000;  wr_data_rom[ 4496]='h00000000;
    rd_cycle[ 4497] = 1'b0;  wr_cycle[ 4497] = 1'b0;  addr_rom[ 4497]='h00000000;  wr_data_rom[ 4497]='h00000000;
    rd_cycle[ 4498] = 1'b0;  wr_cycle[ 4498] = 1'b0;  addr_rom[ 4498]='h00000000;  wr_data_rom[ 4498]='h00000000;
    rd_cycle[ 4499] = 1'b0;  wr_cycle[ 4499] = 1'b0;  addr_rom[ 4499]='h00000000;  wr_data_rom[ 4499]='h00000000;
    rd_cycle[ 4500] = 1'b0;  wr_cycle[ 4500] = 1'b0;  addr_rom[ 4500]='h00000000;  wr_data_rom[ 4500]='h00000000;
    rd_cycle[ 4501] = 1'b0;  wr_cycle[ 4501] = 1'b0;  addr_rom[ 4501]='h00000000;  wr_data_rom[ 4501]='h00000000;
    rd_cycle[ 4502] = 1'b0;  wr_cycle[ 4502] = 1'b0;  addr_rom[ 4502]='h00000000;  wr_data_rom[ 4502]='h00000000;
    rd_cycle[ 4503] = 1'b0;  wr_cycle[ 4503] = 1'b0;  addr_rom[ 4503]='h00000000;  wr_data_rom[ 4503]='h00000000;
    rd_cycle[ 4504] = 1'b0;  wr_cycle[ 4504] = 1'b0;  addr_rom[ 4504]='h00000000;  wr_data_rom[ 4504]='h00000000;
    rd_cycle[ 4505] = 1'b0;  wr_cycle[ 4505] = 1'b0;  addr_rom[ 4505]='h00000000;  wr_data_rom[ 4505]='h00000000;
    rd_cycle[ 4506] = 1'b0;  wr_cycle[ 4506] = 1'b0;  addr_rom[ 4506]='h00000000;  wr_data_rom[ 4506]='h00000000;
    rd_cycle[ 4507] = 1'b0;  wr_cycle[ 4507] = 1'b0;  addr_rom[ 4507]='h00000000;  wr_data_rom[ 4507]='h00000000;
    rd_cycle[ 4508] = 1'b0;  wr_cycle[ 4508] = 1'b0;  addr_rom[ 4508]='h00000000;  wr_data_rom[ 4508]='h00000000;
    rd_cycle[ 4509] = 1'b0;  wr_cycle[ 4509] = 1'b0;  addr_rom[ 4509]='h00000000;  wr_data_rom[ 4509]='h00000000;
    rd_cycle[ 4510] = 1'b0;  wr_cycle[ 4510] = 1'b0;  addr_rom[ 4510]='h00000000;  wr_data_rom[ 4510]='h00000000;
    rd_cycle[ 4511] = 1'b0;  wr_cycle[ 4511] = 1'b0;  addr_rom[ 4511]='h00000000;  wr_data_rom[ 4511]='h00000000;
    rd_cycle[ 4512] = 1'b0;  wr_cycle[ 4512] = 1'b0;  addr_rom[ 4512]='h00000000;  wr_data_rom[ 4512]='h00000000;
    rd_cycle[ 4513] = 1'b0;  wr_cycle[ 4513] = 1'b0;  addr_rom[ 4513]='h00000000;  wr_data_rom[ 4513]='h00000000;
    rd_cycle[ 4514] = 1'b0;  wr_cycle[ 4514] = 1'b0;  addr_rom[ 4514]='h00000000;  wr_data_rom[ 4514]='h00000000;
    rd_cycle[ 4515] = 1'b0;  wr_cycle[ 4515] = 1'b0;  addr_rom[ 4515]='h00000000;  wr_data_rom[ 4515]='h00000000;
    rd_cycle[ 4516] = 1'b0;  wr_cycle[ 4516] = 1'b0;  addr_rom[ 4516]='h00000000;  wr_data_rom[ 4516]='h00000000;
    rd_cycle[ 4517] = 1'b0;  wr_cycle[ 4517] = 1'b0;  addr_rom[ 4517]='h00000000;  wr_data_rom[ 4517]='h00000000;
    rd_cycle[ 4518] = 1'b0;  wr_cycle[ 4518] = 1'b0;  addr_rom[ 4518]='h00000000;  wr_data_rom[ 4518]='h00000000;
    rd_cycle[ 4519] = 1'b0;  wr_cycle[ 4519] = 1'b0;  addr_rom[ 4519]='h00000000;  wr_data_rom[ 4519]='h00000000;
    rd_cycle[ 4520] = 1'b0;  wr_cycle[ 4520] = 1'b0;  addr_rom[ 4520]='h00000000;  wr_data_rom[ 4520]='h00000000;
    rd_cycle[ 4521] = 1'b0;  wr_cycle[ 4521] = 1'b0;  addr_rom[ 4521]='h00000000;  wr_data_rom[ 4521]='h00000000;
    rd_cycle[ 4522] = 1'b0;  wr_cycle[ 4522] = 1'b0;  addr_rom[ 4522]='h00000000;  wr_data_rom[ 4522]='h00000000;
    rd_cycle[ 4523] = 1'b0;  wr_cycle[ 4523] = 1'b0;  addr_rom[ 4523]='h00000000;  wr_data_rom[ 4523]='h00000000;
    rd_cycle[ 4524] = 1'b0;  wr_cycle[ 4524] = 1'b0;  addr_rom[ 4524]='h00000000;  wr_data_rom[ 4524]='h00000000;
    rd_cycle[ 4525] = 1'b0;  wr_cycle[ 4525] = 1'b0;  addr_rom[ 4525]='h00000000;  wr_data_rom[ 4525]='h00000000;
    rd_cycle[ 4526] = 1'b0;  wr_cycle[ 4526] = 1'b0;  addr_rom[ 4526]='h00000000;  wr_data_rom[ 4526]='h00000000;
    rd_cycle[ 4527] = 1'b0;  wr_cycle[ 4527] = 1'b0;  addr_rom[ 4527]='h00000000;  wr_data_rom[ 4527]='h00000000;
    rd_cycle[ 4528] = 1'b0;  wr_cycle[ 4528] = 1'b0;  addr_rom[ 4528]='h00000000;  wr_data_rom[ 4528]='h00000000;
    rd_cycle[ 4529] = 1'b0;  wr_cycle[ 4529] = 1'b0;  addr_rom[ 4529]='h00000000;  wr_data_rom[ 4529]='h00000000;
    rd_cycle[ 4530] = 1'b0;  wr_cycle[ 4530] = 1'b0;  addr_rom[ 4530]='h00000000;  wr_data_rom[ 4530]='h00000000;
    rd_cycle[ 4531] = 1'b0;  wr_cycle[ 4531] = 1'b0;  addr_rom[ 4531]='h00000000;  wr_data_rom[ 4531]='h00000000;
    rd_cycle[ 4532] = 1'b0;  wr_cycle[ 4532] = 1'b0;  addr_rom[ 4532]='h00000000;  wr_data_rom[ 4532]='h00000000;
    rd_cycle[ 4533] = 1'b0;  wr_cycle[ 4533] = 1'b0;  addr_rom[ 4533]='h00000000;  wr_data_rom[ 4533]='h00000000;
    rd_cycle[ 4534] = 1'b0;  wr_cycle[ 4534] = 1'b0;  addr_rom[ 4534]='h00000000;  wr_data_rom[ 4534]='h00000000;
    rd_cycle[ 4535] = 1'b0;  wr_cycle[ 4535] = 1'b0;  addr_rom[ 4535]='h00000000;  wr_data_rom[ 4535]='h00000000;
    rd_cycle[ 4536] = 1'b0;  wr_cycle[ 4536] = 1'b0;  addr_rom[ 4536]='h00000000;  wr_data_rom[ 4536]='h00000000;
    rd_cycle[ 4537] = 1'b0;  wr_cycle[ 4537] = 1'b0;  addr_rom[ 4537]='h00000000;  wr_data_rom[ 4537]='h00000000;
    rd_cycle[ 4538] = 1'b0;  wr_cycle[ 4538] = 1'b0;  addr_rom[ 4538]='h00000000;  wr_data_rom[ 4538]='h00000000;
    rd_cycle[ 4539] = 1'b0;  wr_cycle[ 4539] = 1'b0;  addr_rom[ 4539]='h00000000;  wr_data_rom[ 4539]='h00000000;
    rd_cycle[ 4540] = 1'b0;  wr_cycle[ 4540] = 1'b0;  addr_rom[ 4540]='h00000000;  wr_data_rom[ 4540]='h00000000;
    rd_cycle[ 4541] = 1'b0;  wr_cycle[ 4541] = 1'b0;  addr_rom[ 4541]='h00000000;  wr_data_rom[ 4541]='h00000000;
    rd_cycle[ 4542] = 1'b0;  wr_cycle[ 4542] = 1'b0;  addr_rom[ 4542]='h00000000;  wr_data_rom[ 4542]='h00000000;
    rd_cycle[ 4543] = 1'b0;  wr_cycle[ 4543] = 1'b0;  addr_rom[ 4543]='h00000000;  wr_data_rom[ 4543]='h00000000;
    rd_cycle[ 4544] = 1'b0;  wr_cycle[ 4544] = 1'b0;  addr_rom[ 4544]='h00000000;  wr_data_rom[ 4544]='h00000000;
    rd_cycle[ 4545] = 1'b0;  wr_cycle[ 4545] = 1'b0;  addr_rom[ 4545]='h00000000;  wr_data_rom[ 4545]='h00000000;
    rd_cycle[ 4546] = 1'b0;  wr_cycle[ 4546] = 1'b0;  addr_rom[ 4546]='h00000000;  wr_data_rom[ 4546]='h00000000;
    rd_cycle[ 4547] = 1'b0;  wr_cycle[ 4547] = 1'b0;  addr_rom[ 4547]='h00000000;  wr_data_rom[ 4547]='h00000000;
    rd_cycle[ 4548] = 1'b0;  wr_cycle[ 4548] = 1'b0;  addr_rom[ 4548]='h00000000;  wr_data_rom[ 4548]='h00000000;
    rd_cycle[ 4549] = 1'b0;  wr_cycle[ 4549] = 1'b0;  addr_rom[ 4549]='h00000000;  wr_data_rom[ 4549]='h00000000;
    rd_cycle[ 4550] = 1'b0;  wr_cycle[ 4550] = 1'b0;  addr_rom[ 4550]='h00000000;  wr_data_rom[ 4550]='h00000000;
    rd_cycle[ 4551] = 1'b0;  wr_cycle[ 4551] = 1'b0;  addr_rom[ 4551]='h00000000;  wr_data_rom[ 4551]='h00000000;
    rd_cycle[ 4552] = 1'b0;  wr_cycle[ 4552] = 1'b0;  addr_rom[ 4552]='h00000000;  wr_data_rom[ 4552]='h00000000;
    rd_cycle[ 4553] = 1'b0;  wr_cycle[ 4553] = 1'b0;  addr_rom[ 4553]='h00000000;  wr_data_rom[ 4553]='h00000000;
    rd_cycle[ 4554] = 1'b0;  wr_cycle[ 4554] = 1'b0;  addr_rom[ 4554]='h00000000;  wr_data_rom[ 4554]='h00000000;
    rd_cycle[ 4555] = 1'b0;  wr_cycle[ 4555] = 1'b0;  addr_rom[ 4555]='h00000000;  wr_data_rom[ 4555]='h00000000;
    rd_cycle[ 4556] = 1'b0;  wr_cycle[ 4556] = 1'b0;  addr_rom[ 4556]='h00000000;  wr_data_rom[ 4556]='h00000000;
    rd_cycle[ 4557] = 1'b0;  wr_cycle[ 4557] = 1'b0;  addr_rom[ 4557]='h00000000;  wr_data_rom[ 4557]='h00000000;
    rd_cycle[ 4558] = 1'b0;  wr_cycle[ 4558] = 1'b0;  addr_rom[ 4558]='h00000000;  wr_data_rom[ 4558]='h00000000;
    rd_cycle[ 4559] = 1'b0;  wr_cycle[ 4559] = 1'b0;  addr_rom[ 4559]='h00000000;  wr_data_rom[ 4559]='h00000000;
    rd_cycle[ 4560] = 1'b0;  wr_cycle[ 4560] = 1'b0;  addr_rom[ 4560]='h00000000;  wr_data_rom[ 4560]='h00000000;
    rd_cycle[ 4561] = 1'b0;  wr_cycle[ 4561] = 1'b0;  addr_rom[ 4561]='h00000000;  wr_data_rom[ 4561]='h00000000;
    rd_cycle[ 4562] = 1'b0;  wr_cycle[ 4562] = 1'b0;  addr_rom[ 4562]='h00000000;  wr_data_rom[ 4562]='h00000000;
    rd_cycle[ 4563] = 1'b0;  wr_cycle[ 4563] = 1'b0;  addr_rom[ 4563]='h00000000;  wr_data_rom[ 4563]='h00000000;
    rd_cycle[ 4564] = 1'b0;  wr_cycle[ 4564] = 1'b0;  addr_rom[ 4564]='h00000000;  wr_data_rom[ 4564]='h00000000;
    rd_cycle[ 4565] = 1'b0;  wr_cycle[ 4565] = 1'b0;  addr_rom[ 4565]='h00000000;  wr_data_rom[ 4565]='h00000000;
    rd_cycle[ 4566] = 1'b0;  wr_cycle[ 4566] = 1'b0;  addr_rom[ 4566]='h00000000;  wr_data_rom[ 4566]='h00000000;
    rd_cycle[ 4567] = 1'b0;  wr_cycle[ 4567] = 1'b0;  addr_rom[ 4567]='h00000000;  wr_data_rom[ 4567]='h00000000;
    rd_cycle[ 4568] = 1'b0;  wr_cycle[ 4568] = 1'b0;  addr_rom[ 4568]='h00000000;  wr_data_rom[ 4568]='h00000000;
    rd_cycle[ 4569] = 1'b0;  wr_cycle[ 4569] = 1'b0;  addr_rom[ 4569]='h00000000;  wr_data_rom[ 4569]='h00000000;
    rd_cycle[ 4570] = 1'b0;  wr_cycle[ 4570] = 1'b0;  addr_rom[ 4570]='h00000000;  wr_data_rom[ 4570]='h00000000;
    rd_cycle[ 4571] = 1'b0;  wr_cycle[ 4571] = 1'b0;  addr_rom[ 4571]='h00000000;  wr_data_rom[ 4571]='h00000000;
    rd_cycle[ 4572] = 1'b0;  wr_cycle[ 4572] = 1'b0;  addr_rom[ 4572]='h00000000;  wr_data_rom[ 4572]='h00000000;
    rd_cycle[ 4573] = 1'b0;  wr_cycle[ 4573] = 1'b0;  addr_rom[ 4573]='h00000000;  wr_data_rom[ 4573]='h00000000;
    rd_cycle[ 4574] = 1'b0;  wr_cycle[ 4574] = 1'b0;  addr_rom[ 4574]='h00000000;  wr_data_rom[ 4574]='h00000000;
    rd_cycle[ 4575] = 1'b0;  wr_cycle[ 4575] = 1'b0;  addr_rom[ 4575]='h00000000;  wr_data_rom[ 4575]='h00000000;
    rd_cycle[ 4576] = 1'b0;  wr_cycle[ 4576] = 1'b0;  addr_rom[ 4576]='h00000000;  wr_data_rom[ 4576]='h00000000;
    rd_cycle[ 4577] = 1'b0;  wr_cycle[ 4577] = 1'b0;  addr_rom[ 4577]='h00000000;  wr_data_rom[ 4577]='h00000000;
    rd_cycle[ 4578] = 1'b0;  wr_cycle[ 4578] = 1'b0;  addr_rom[ 4578]='h00000000;  wr_data_rom[ 4578]='h00000000;
    rd_cycle[ 4579] = 1'b0;  wr_cycle[ 4579] = 1'b0;  addr_rom[ 4579]='h00000000;  wr_data_rom[ 4579]='h00000000;
    rd_cycle[ 4580] = 1'b0;  wr_cycle[ 4580] = 1'b0;  addr_rom[ 4580]='h00000000;  wr_data_rom[ 4580]='h00000000;
    rd_cycle[ 4581] = 1'b0;  wr_cycle[ 4581] = 1'b0;  addr_rom[ 4581]='h00000000;  wr_data_rom[ 4581]='h00000000;
    rd_cycle[ 4582] = 1'b0;  wr_cycle[ 4582] = 1'b0;  addr_rom[ 4582]='h00000000;  wr_data_rom[ 4582]='h00000000;
    rd_cycle[ 4583] = 1'b0;  wr_cycle[ 4583] = 1'b0;  addr_rom[ 4583]='h00000000;  wr_data_rom[ 4583]='h00000000;
    rd_cycle[ 4584] = 1'b0;  wr_cycle[ 4584] = 1'b0;  addr_rom[ 4584]='h00000000;  wr_data_rom[ 4584]='h00000000;
    rd_cycle[ 4585] = 1'b0;  wr_cycle[ 4585] = 1'b0;  addr_rom[ 4585]='h00000000;  wr_data_rom[ 4585]='h00000000;
    rd_cycle[ 4586] = 1'b0;  wr_cycle[ 4586] = 1'b0;  addr_rom[ 4586]='h00000000;  wr_data_rom[ 4586]='h00000000;
    rd_cycle[ 4587] = 1'b0;  wr_cycle[ 4587] = 1'b0;  addr_rom[ 4587]='h00000000;  wr_data_rom[ 4587]='h00000000;
    rd_cycle[ 4588] = 1'b0;  wr_cycle[ 4588] = 1'b0;  addr_rom[ 4588]='h00000000;  wr_data_rom[ 4588]='h00000000;
    rd_cycle[ 4589] = 1'b0;  wr_cycle[ 4589] = 1'b0;  addr_rom[ 4589]='h00000000;  wr_data_rom[ 4589]='h00000000;
    rd_cycle[ 4590] = 1'b0;  wr_cycle[ 4590] = 1'b0;  addr_rom[ 4590]='h00000000;  wr_data_rom[ 4590]='h00000000;
    rd_cycle[ 4591] = 1'b0;  wr_cycle[ 4591] = 1'b0;  addr_rom[ 4591]='h00000000;  wr_data_rom[ 4591]='h00000000;
    rd_cycle[ 4592] = 1'b0;  wr_cycle[ 4592] = 1'b0;  addr_rom[ 4592]='h00000000;  wr_data_rom[ 4592]='h00000000;
    rd_cycle[ 4593] = 1'b0;  wr_cycle[ 4593] = 1'b0;  addr_rom[ 4593]='h00000000;  wr_data_rom[ 4593]='h00000000;
    rd_cycle[ 4594] = 1'b0;  wr_cycle[ 4594] = 1'b0;  addr_rom[ 4594]='h00000000;  wr_data_rom[ 4594]='h00000000;
    rd_cycle[ 4595] = 1'b0;  wr_cycle[ 4595] = 1'b0;  addr_rom[ 4595]='h00000000;  wr_data_rom[ 4595]='h00000000;
    rd_cycle[ 4596] = 1'b0;  wr_cycle[ 4596] = 1'b0;  addr_rom[ 4596]='h00000000;  wr_data_rom[ 4596]='h00000000;
    rd_cycle[ 4597] = 1'b0;  wr_cycle[ 4597] = 1'b0;  addr_rom[ 4597]='h00000000;  wr_data_rom[ 4597]='h00000000;
    rd_cycle[ 4598] = 1'b0;  wr_cycle[ 4598] = 1'b0;  addr_rom[ 4598]='h00000000;  wr_data_rom[ 4598]='h00000000;
    rd_cycle[ 4599] = 1'b0;  wr_cycle[ 4599] = 1'b0;  addr_rom[ 4599]='h00000000;  wr_data_rom[ 4599]='h00000000;
    rd_cycle[ 4600] = 1'b0;  wr_cycle[ 4600] = 1'b0;  addr_rom[ 4600]='h00000000;  wr_data_rom[ 4600]='h00000000;
    rd_cycle[ 4601] = 1'b0;  wr_cycle[ 4601] = 1'b0;  addr_rom[ 4601]='h00000000;  wr_data_rom[ 4601]='h00000000;
    rd_cycle[ 4602] = 1'b0;  wr_cycle[ 4602] = 1'b0;  addr_rom[ 4602]='h00000000;  wr_data_rom[ 4602]='h00000000;
    rd_cycle[ 4603] = 1'b0;  wr_cycle[ 4603] = 1'b0;  addr_rom[ 4603]='h00000000;  wr_data_rom[ 4603]='h00000000;
    rd_cycle[ 4604] = 1'b0;  wr_cycle[ 4604] = 1'b0;  addr_rom[ 4604]='h00000000;  wr_data_rom[ 4604]='h00000000;
    rd_cycle[ 4605] = 1'b0;  wr_cycle[ 4605] = 1'b0;  addr_rom[ 4605]='h00000000;  wr_data_rom[ 4605]='h00000000;
    rd_cycle[ 4606] = 1'b0;  wr_cycle[ 4606] = 1'b0;  addr_rom[ 4606]='h00000000;  wr_data_rom[ 4606]='h00000000;
    rd_cycle[ 4607] = 1'b0;  wr_cycle[ 4607] = 1'b0;  addr_rom[ 4607]='h00000000;  wr_data_rom[ 4607]='h00000000;
    rd_cycle[ 4608] = 1'b0;  wr_cycle[ 4608] = 1'b0;  addr_rom[ 4608]='h00000000;  wr_data_rom[ 4608]='h00000000;
    rd_cycle[ 4609] = 1'b0;  wr_cycle[ 4609] = 1'b0;  addr_rom[ 4609]='h00000000;  wr_data_rom[ 4609]='h00000000;
    rd_cycle[ 4610] = 1'b0;  wr_cycle[ 4610] = 1'b0;  addr_rom[ 4610]='h00000000;  wr_data_rom[ 4610]='h00000000;
    rd_cycle[ 4611] = 1'b0;  wr_cycle[ 4611] = 1'b0;  addr_rom[ 4611]='h00000000;  wr_data_rom[ 4611]='h00000000;
    rd_cycle[ 4612] = 1'b0;  wr_cycle[ 4612] = 1'b0;  addr_rom[ 4612]='h00000000;  wr_data_rom[ 4612]='h00000000;
    rd_cycle[ 4613] = 1'b0;  wr_cycle[ 4613] = 1'b0;  addr_rom[ 4613]='h00000000;  wr_data_rom[ 4613]='h00000000;
    rd_cycle[ 4614] = 1'b0;  wr_cycle[ 4614] = 1'b0;  addr_rom[ 4614]='h00000000;  wr_data_rom[ 4614]='h00000000;
    rd_cycle[ 4615] = 1'b0;  wr_cycle[ 4615] = 1'b0;  addr_rom[ 4615]='h00000000;  wr_data_rom[ 4615]='h00000000;
    rd_cycle[ 4616] = 1'b0;  wr_cycle[ 4616] = 1'b0;  addr_rom[ 4616]='h00000000;  wr_data_rom[ 4616]='h00000000;
    rd_cycle[ 4617] = 1'b0;  wr_cycle[ 4617] = 1'b0;  addr_rom[ 4617]='h00000000;  wr_data_rom[ 4617]='h00000000;
    rd_cycle[ 4618] = 1'b0;  wr_cycle[ 4618] = 1'b0;  addr_rom[ 4618]='h00000000;  wr_data_rom[ 4618]='h00000000;
    rd_cycle[ 4619] = 1'b0;  wr_cycle[ 4619] = 1'b0;  addr_rom[ 4619]='h00000000;  wr_data_rom[ 4619]='h00000000;
    rd_cycle[ 4620] = 1'b0;  wr_cycle[ 4620] = 1'b0;  addr_rom[ 4620]='h00000000;  wr_data_rom[ 4620]='h00000000;
    rd_cycle[ 4621] = 1'b0;  wr_cycle[ 4621] = 1'b0;  addr_rom[ 4621]='h00000000;  wr_data_rom[ 4621]='h00000000;
    rd_cycle[ 4622] = 1'b0;  wr_cycle[ 4622] = 1'b0;  addr_rom[ 4622]='h00000000;  wr_data_rom[ 4622]='h00000000;
    rd_cycle[ 4623] = 1'b0;  wr_cycle[ 4623] = 1'b0;  addr_rom[ 4623]='h00000000;  wr_data_rom[ 4623]='h00000000;
    rd_cycle[ 4624] = 1'b0;  wr_cycle[ 4624] = 1'b0;  addr_rom[ 4624]='h00000000;  wr_data_rom[ 4624]='h00000000;
    rd_cycle[ 4625] = 1'b0;  wr_cycle[ 4625] = 1'b0;  addr_rom[ 4625]='h00000000;  wr_data_rom[ 4625]='h00000000;
    rd_cycle[ 4626] = 1'b0;  wr_cycle[ 4626] = 1'b0;  addr_rom[ 4626]='h00000000;  wr_data_rom[ 4626]='h00000000;
    rd_cycle[ 4627] = 1'b0;  wr_cycle[ 4627] = 1'b0;  addr_rom[ 4627]='h00000000;  wr_data_rom[ 4627]='h00000000;
    rd_cycle[ 4628] = 1'b0;  wr_cycle[ 4628] = 1'b0;  addr_rom[ 4628]='h00000000;  wr_data_rom[ 4628]='h00000000;
    rd_cycle[ 4629] = 1'b0;  wr_cycle[ 4629] = 1'b0;  addr_rom[ 4629]='h00000000;  wr_data_rom[ 4629]='h00000000;
    rd_cycle[ 4630] = 1'b0;  wr_cycle[ 4630] = 1'b0;  addr_rom[ 4630]='h00000000;  wr_data_rom[ 4630]='h00000000;
    rd_cycle[ 4631] = 1'b0;  wr_cycle[ 4631] = 1'b0;  addr_rom[ 4631]='h00000000;  wr_data_rom[ 4631]='h00000000;
    rd_cycle[ 4632] = 1'b0;  wr_cycle[ 4632] = 1'b0;  addr_rom[ 4632]='h00000000;  wr_data_rom[ 4632]='h00000000;
    rd_cycle[ 4633] = 1'b0;  wr_cycle[ 4633] = 1'b0;  addr_rom[ 4633]='h00000000;  wr_data_rom[ 4633]='h00000000;
    rd_cycle[ 4634] = 1'b0;  wr_cycle[ 4634] = 1'b0;  addr_rom[ 4634]='h00000000;  wr_data_rom[ 4634]='h00000000;
    rd_cycle[ 4635] = 1'b0;  wr_cycle[ 4635] = 1'b0;  addr_rom[ 4635]='h00000000;  wr_data_rom[ 4635]='h00000000;
    rd_cycle[ 4636] = 1'b0;  wr_cycle[ 4636] = 1'b0;  addr_rom[ 4636]='h00000000;  wr_data_rom[ 4636]='h00000000;
    rd_cycle[ 4637] = 1'b0;  wr_cycle[ 4637] = 1'b0;  addr_rom[ 4637]='h00000000;  wr_data_rom[ 4637]='h00000000;
    rd_cycle[ 4638] = 1'b0;  wr_cycle[ 4638] = 1'b0;  addr_rom[ 4638]='h00000000;  wr_data_rom[ 4638]='h00000000;
    rd_cycle[ 4639] = 1'b0;  wr_cycle[ 4639] = 1'b0;  addr_rom[ 4639]='h00000000;  wr_data_rom[ 4639]='h00000000;
    rd_cycle[ 4640] = 1'b0;  wr_cycle[ 4640] = 1'b0;  addr_rom[ 4640]='h00000000;  wr_data_rom[ 4640]='h00000000;
    rd_cycle[ 4641] = 1'b0;  wr_cycle[ 4641] = 1'b0;  addr_rom[ 4641]='h00000000;  wr_data_rom[ 4641]='h00000000;
    rd_cycle[ 4642] = 1'b0;  wr_cycle[ 4642] = 1'b0;  addr_rom[ 4642]='h00000000;  wr_data_rom[ 4642]='h00000000;
    rd_cycle[ 4643] = 1'b0;  wr_cycle[ 4643] = 1'b0;  addr_rom[ 4643]='h00000000;  wr_data_rom[ 4643]='h00000000;
    rd_cycle[ 4644] = 1'b0;  wr_cycle[ 4644] = 1'b0;  addr_rom[ 4644]='h00000000;  wr_data_rom[ 4644]='h00000000;
    rd_cycle[ 4645] = 1'b0;  wr_cycle[ 4645] = 1'b0;  addr_rom[ 4645]='h00000000;  wr_data_rom[ 4645]='h00000000;
    rd_cycle[ 4646] = 1'b0;  wr_cycle[ 4646] = 1'b0;  addr_rom[ 4646]='h00000000;  wr_data_rom[ 4646]='h00000000;
    rd_cycle[ 4647] = 1'b0;  wr_cycle[ 4647] = 1'b0;  addr_rom[ 4647]='h00000000;  wr_data_rom[ 4647]='h00000000;
    rd_cycle[ 4648] = 1'b0;  wr_cycle[ 4648] = 1'b0;  addr_rom[ 4648]='h00000000;  wr_data_rom[ 4648]='h00000000;
    rd_cycle[ 4649] = 1'b0;  wr_cycle[ 4649] = 1'b0;  addr_rom[ 4649]='h00000000;  wr_data_rom[ 4649]='h00000000;
    rd_cycle[ 4650] = 1'b0;  wr_cycle[ 4650] = 1'b0;  addr_rom[ 4650]='h00000000;  wr_data_rom[ 4650]='h00000000;
    rd_cycle[ 4651] = 1'b0;  wr_cycle[ 4651] = 1'b0;  addr_rom[ 4651]='h00000000;  wr_data_rom[ 4651]='h00000000;
    rd_cycle[ 4652] = 1'b0;  wr_cycle[ 4652] = 1'b0;  addr_rom[ 4652]='h00000000;  wr_data_rom[ 4652]='h00000000;
    rd_cycle[ 4653] = 1'b0;  wr_cycle[ 4653] = 1'b0;  addr_rom[ 4653]='h00000000;  wr_data_rom[ 4653]='h00000000;
    rd_cycle[ 4654] = 1'b0;  wr_cycle[ 4654] = 1'b0;  addr_rom[ 4654]='h00000000;  wr_data_rom[ 4654]='h00000000;
    rd_cycle[ 4655] = 1'b0;  wr_cycle[ 4655] = 1'b0;  addr_rom[ 4655]='h00000000;  wr_data_rom[ 4655]='h00000000;
    rd_cycle[ 4656] = 1'b0;  wr_cycle[ 4656] = 1'b0;  addr_rom[ 4656]='h00000000;  wr_data_rom[ 4656]='h00000000;
    rd_cycle[ 4657] = 1'b0;  wr_cycle[ 4657] = 1'b0;  addr_rom[ 4657]='h00000000;  wr_data_rom[ 4657]='h00000000;
    rd_cycle[ 4658] = 1'b0;  wr_cycle[ 4658] = 1'b0;  addr_rom[ 4658]='h00000000;  wr_data_rom[ 4658]='h00000000;
    rd_cycle[ 4659] = 1'b0;  wr_cycle[ 4659] = 1'b0;  addr_rom[ 4659]='h00000000;  wr_data_rom[ 4659]='h00000000;
    rd_cycle[ 4660] = 1'b0;  wr_cycle[ 4660] = 1'b0;  addr_rom[ 4660]='h00000000;  wr_data_rom[ 4660]='h00000000;
    rd_cycle[ 4661] = 1'b0;  wr_cycle[ 4661] = 1'b0;  addr_rom[ 4661]='h00000000;  wr_data_rom[ 4661]='h00000000;
    rd_cycle[ 4662] = 1'b0;  wr_cycle[ 4662] = 1'b0;  addr_rom[ 4662]='h00000000;  wr_data_rom[ 4662]='h00000000;
    rd_cycle[ 4663] = 1'b0;  wr_cycle[ 4663] = 1'b0;  addr_rom[ 4663]='h00000000;  wr_data_rom[ 4663]='h00000000;
    rd_cycle[ 4664] = 1'b0;  wr_cycle[ 4664] = 1'b0;  addr_rom[ 4664]='h00000000;  wr_data_rom[ 4664]='h00000000;
    rd_cycle[ 4665] = 1'b0;  wr_cycle[ 4665] = 1'b0;  addr_rom[ 4665]='h00000000;  wr_data_rom[ 4665]='h00000000;
    rd_cycle[ 4666] = 1'b0;  wr_cycle[ 4666] = 1'b0;  addr_rom[ 4666]='h00000000;  wr_data_rom[ 4666]='h00000000;
    rd_cycle[ 4667] = 1'b0;  wr_cycle[ 4667] = 1'b0;  addr_rom[ 4667]='h00000000;  wr_data_rom[ 4667]='h00000000;
    rd_cycle[ 4668] = 1'b0;  wr_cycle[ 4668] = 1'b0;  addr_rom[ 4668]='h00000000;  wr_data_rom[ 4668]='h00000000;
    rd_cycle[ 4669] = 1'b0;  wr_cycle[ 4669] = 1'b0;  addr_rom[ 4669]='h00000000;  wr_data_rom[ 4669]='h00000000;
    rd_cycle[ 4670] = 1'b0;  wr_cycle[ 4670] = 1'b0;  addr_rom[ 4670]='h00000000;  wr_data_rom[ 4670]='h00000000;
    rd_cycle[ 4671] = 1'b0;  wr_cycle[ 4671] = 1'b0;  addr_rom[ 4671]='h00000000;  wr_data_rom[ 4671]='h00000000;
    rd_cycle[ 4672] = 1'b0;  wr_cycle[ 4672] = 1'b0;  addr_rom[ 4672]='h00000000;  wr_data_rom[ 4672]='h00000000;
    rd_cycle[ 4673] = 1'b0;  wr_cycle[ 4673] = 1'b0;  addr_rom[ 4673]='h00000000;  wr_data_rom[ 4673]='h00000000;
    rd_cycle[ 4674] = 1'b0;  wr_cycle[ 4674] = 1'b0;  addr_rom[ 4674]='h00000000;  wr_data_rom[ 4674]='h00000000;
    rd_cycle[ 4675] = 1'b0;  wr_cycle[ 4675] = 1'b0;  addr_rom[ 4675]='h00000000;  wr_data_rom[ 4675]='h00000000;
    rd_cycle[ 4676] = 1'b0;  wr_cycle[ 4676] = 1'b0;  addr_rom[ 4676]='h00000000;  wr_data_rom[ 4676]='h00000000;
    rd_cycle[ 4677] = 1'b0;  wr_cycle[ 4677] = 1'b0;  addr_rom[ 4677]='h00000000;  wr_data_rom[ 4677]='h00000000;
    rd_cycle[ 4678] = 1'b0;  wr_cycle[ 4678] = 1'b0;  addr_rom[ 4678]='h00000000;  wr_data_rom[ 4678]='h00000000;
    rd_cycle[ 4679] = 1'b0;  wr_cycle[ 4679] = 1'b0;  addr_rom[ 4679]='h00000000;  wr_data_rom[ 4679]='h00000000;
    rd_cycle[ 4680] = 1'b0;  wr_cycle[ 4680] = 1'b0;  addr_rom[ 4680]='h00000000;  wr_data_rom[ 4680]='h00000000;
    rd_cycle[ 4681] = 1'b0;  wr_cycle[ 4681] = 1'b0;  addr_rom[ 4681]='h00000000;  wr_data_rom[ 4681]='h00000000;
    rd_cycle[ 4682] = 1'b0;  wr_cycle[ 4682] = 1'b0;  addr_rom[ 4682]='h00000000;  wr_data_rom[ 4682]='h00000000;
    rd_cycle[ 4683] = 1'b0;  wr_cycle[ 4683] = 1'b0;  addr_rom[ 4683]='h00000000;  wr_data_rom[ 4683]='h00000000;
    rd_cycle[ 4684] = 1'b0;  wr_cycle[ 4684] = 1'b0;  addr_rom[ 4684]='h00000000;  wr_data_rom[ 4684]='h00000000;
    rd_cycle[ 4685] = 1'b0;  wr_cycle[ 4685] = 1'b0;  addr_rom[ 4685]='h00000000;  wr_data_rom[ 4685]='h00000000;
    rd_cycle[ 4686] = 1'b0;  wr_cycle[ 4686] = 1'b0;  addr_rom[ 4686]='h00000000;  wr_data_rom[ 4686]='h00000000;
    rd_cycle[ 4687] = 1'b0;  wr_cycle[ 4687] = 1'b0;  addr_rom[ 4687]='h00000000;  wr_data_rom[ 4687]='h00000000;
    rd_cycle[ 4688] = 1'b0;  wr_cycle[ 4688] = 1'b0;  addr_rom[ 4688]='h00000000;  wr_data_rom[ 4688]='h00000000;
    rd_cycle[ 4689] = 1'b0;  wr_cycle[ 4689] = 1'b0;  addr_rom[ 4689]='h00000000;  wr_data_rom[ 4689]='h00000000;
    rd_cycle[ 4690] = 1'b0;  wr_cycle[ 4690] = 1'b0;  addr_rom[ 4690]='h00000000;  wr_data_rom[ 4690]='h00000000;
    rd_cycle[ 4691] = 1'b0;  wr_cycle[ 4691] = 1'b0;  addr_rom[ 4691]='h00000000;  wr_data_rom[ 4691]='h00000000;
    rd_cycle[ 4692] = 1'b0;  wr_cycle[ 4692] = 1'b0;  addr_rom[ 4692]='h00000000;  wr_data_rom[ 4692]='h00000000;
    rd_cycle[ 4693] = 1'b0;  wr_cycle[ 4693] = 1'b0;  addr_rom[ 4693]='h00000000;  wr_data_rom[ 4693]='h00000000;
    rd_cycle[ 4694] = 1'b0;  wr_cycle[ 4694] = 1'b0;  addr_rom[ 4694]='h00000000;  wr_data_rom[ 4694]='h00000000;
    rd_cycle[ 4695] = 1'b0;  wr_cycle[ 4695] = 1'b0;  addr_rom[ 4695]='h00000000;  wr_data_rom[ 4695]='h00000000;
    rd_cycle[ 4696] = 1'b0;  wr_cycle[ 4696] = 1'b0;  addr_rom[ 4696]='h00000000;  wr_data_rom[ 4696]='h00000000;
    rd_cycle[ 4697] = 1'b0;  wr_cycle[ 4697] = 1'b0;  addr_rom[ 4697]='h00000000;  wr_data_rom[ 4697]='h00000000;
    rd_cycle[ 4698] = 1'b0;  wr_cycle[ 4698] = 1'b0;  addr_rom[ 4698]='h00000000;  wr_data_rom[ 4698]='h00000000;
    rd_cycle[ 4699] = 1'b0;  wr_cycle[ 4699] = 1'b0;  addr_rom[ 4699]='h00000000;  wr_data_rom[ 4699]='h00000000;
    rd_cycle[ 4700] = 1'b0;  wr_cycle[ 4700] = 1'b0;  addr_rom[ 4700]='h00000000;  wr_data_rom[ 4700]='h00000000;
    rd_cycle[ 4701] = 1'b0;  wr_cycle[ 4701] = 1'b0;  addr_rom[ 4701]='h00000000;  wr_data_rom[ 4701]='h00000000;
    rd_cycle[ 4702] = 1'b0;  wr_cycle[ 4702] = 1'b0;  addr_rom[ 4702]='h00000000;  wr_data_rom[ 4702]='h00000000;
    rd_cycle[ 4703] = 1'b0;  wr_cycle[ 4703] = 1'b0;  addr_rom[ 4703]='h00000000;  wr_data_rom[ 4703]='h00000000;
    rd_cycle[ 4704] = 1'b0;  wr_cycle[ 4704] = 1'b0;  addr_rom[ 4704]='h00000000;  wr_data_rom[ 4704]='h00000000;
    rd_cycle[ 4705] = 1'b0;  wr_cycle[ 4705] = 1'b0;  addr_rom[ 4705]='h00000000;  wr_data_rom[ 4705]='h00000000;
    rd_cycle[ 4706] = 1'b0;  wr_cycle[ 4706] = 1'b0;  addr_rom[ 4706]='h00000000;  wr_data_rom[ 4706]='h00000000;
    rd_cycle[ 4707] = 1'b0;  wr_cycle[ 4707] = 1'b0;  addr_rom[ 4707]='h00000000;  wr_data_rom[ 4707]='h00000000;
    rd_cycle[ 4708] = 1'b0;  wr_cycle[ 4708] = 1'b0;  addr_rom[ 4708]='h00000000;  wr_data_rom[ 4708]='h00000000;
    rd_cycle[ 4709] = 1'b0;  wr_cycle[ 4709] = 1'b0;  addr_rom[ 4709]='h00000000;  wr_data_rom[ 4709]='h00000000;
    rd_cycle[ 4710] = 1'b0;  wr_cycle[ 4710] = 1'b0;  addr_rom[ 4710]='h00000000;  wr_data_rom[ 4710]='h00000000;
    rd_cycle[ 4711] = 1'b0;  wr_cycle[ 4711] = 1'b0;  addr_rom[ 4711]='h00000000;  wr_data_rom[ 4711]='h00000000;
    rd_cycle[ 4712] = 1'b0;  wr_cycle[ 4712] = 1'b0;  addr_rom[ 4712]='h00000000;  wr_data_rom[ 4712]='h00000000;
    rd_cycle[ 4713] = 1'b0;  wr_cycle[ 4713] = 1'b0;  addr_rom[ 4713]='h00000000;  wr_data_rom[ 4713]='h00000000;
    rd_cycle[ 4714] = 1'b0;  wr_cycle[ 4714] = 1'b0;  addr_rom[ 4714]='h00000000;  wr_data_rom[ 4714]='h00000000;
    rd_cycle[ 4715] = 1'b0;  wr_cycle[ 4715] = 1'b0;  addr_rom[ 4715]='h00000000;  wr_data_rom[ 4715]='h00000000;
    rd_cycle[ 4716] = 1'b0;  wr_cycle[ 4716] = 1'b0;  addr_rom[ 4716]='h00000000;  wr_data_rom[ 4716]='h00000000;
    rd_cycle[ 4717] = 1'b0;  wr_cycle[ 4717] = 1'b0;  addr_rom[ 4717]='h00000000;  wr_data_rom[ 4717]='h00000000;
    rd_cycle[ 4718] = 1'b0;  wr_cycle[ 4718] = 1'b0;  addr_rom[ 4718]='h00000000;  wr_data_rom[ 4718]='h00000000;
    rd_cycle[ 4719] = 1'b0;  wr_cycle[ 4719] = 1'b0;  addr_rom[ 4719]='h00000000;  wr_data_rom[ 4719]='h00000000;
    rd_cycle[ 4720] = 1'b0;  wr_cycle[ 4720] = 1'b0;  addr_rom[ 4720]='h00000000;  wr_data_rom[ 4720]='h00000000;
    rd_cycle[ 4721] = 1'b0;  wr_cycle[ 4721] = 1'b0;  addr_rom[ 4721]='h00000000;  wr_data_rom[ 4721]='h00000000;
    rd_cycle[ 4722] = 1'b0;  wr_cycle[ 4722] = 1'b0;  addr_rom[ 4722]='h00000000;  wr_data_rom[ 4722]='h00000000;
    rd_cycle[ 4723] = 1'b0;  wr_cycle[ 4723] = 1'b0;  addr_rom[ 4723]='h00000000;  wr_data_rom[ 4723]='h00000000;
    rd_cycle[ 4724] = 1'b0;  wr_cycle[ 4724] = 1'b0;  addr_rom[ 4724]='h00000000;  wr_data_rom[ 4724]='h00000000;
    rd_cycle[ 4725] = 1'b0;  wr_cycle[ 4725] = 1'b0;  addr_rom[ 4725]='h00000000;  wr_data_rom[ 4725]='h00000000;
    rd_cycle[ 4726] = 1'b0;  wr_cycle[ 4726] = 1'b0;  addr_rom[ 4726]='h00000000;  wr_data_rom[ 4726]='h00000000;
    rd_cycle[ 4727] = 1'b0;  wr_cycle[ 4727] = 1'b0;  addr_rom[ 4727]='h00000000;  wr_data_rom[ 4727]='h00000000;
    rd_cycle[ 4728] = 1'b0;  wr_cycle[ 4728] = 1'b0;  addr_rom[ 4728]='h00000000;  wr_data_rom[ 4728]='h00000000;
    rd_cycle[ 4729] = 1'b0;  wr_cycle[ 4729] = 1'b0;  addr_rom[ 4729]='h00000000;  wr_data_rom[ 4729]='h00000000;
    rd_cycle[ 4730] = 1'b0;  wr_cycle[ 4730] = 1'b0;  addr_rom[ 4730]='h00000000;  wr_data_rom[ 4730]='h00000000;
    rd_cycle[ 4731] = 1'b0;  wr_cycle[ 4731] = 1'b0;  addr_rom[ 4731]='h00000000;  wr_data_rom[ 4731]='h00000000;
    rd_cycle[ 4732] = 1'b0;  wr_cycle[ 4732] = 1'b0;  addr_rom[ 4732]='h00000000;  wr_data_rom[ 4732]='h00000000;
    rd_cycle[ 4733] = 1'b0;  wr_cycle[ 4733] = 1'b0;  addr_rom[ 4733]='h00000000;  wr_data_rom[ 4733]='h00000000;
    rd_cycle[ 4734] = 1'b0;  wr_cycle[ 4734] = 1'b0;  addr_rom[ 4734]='h00000000;  wr_data_rom[ 4734]='h00000000;
    rd_cycle[ 4735] = 1'b0;  wr_cycle[ 4735] = 1'b0;  addr_rom[ 4735]='h00000000;  wr_data_rom[ 4735]='h00000000;
    rd_cycle[ 4736] = 1'b0;  wr_cycle[ 4736] = 1'b0;  addr_rom[ 4736]='h00000000;  wr_data_rom[ 4736]='h00000000;
    rd_cycle[ 4737] = 1'b0;  wr_cycle[ 4737] = 1'b0;  addr_rom[ 4737]='h00000000;  wr_data_rom[ 4737]='h00000000;
    rd_cycle[ 4738] = 1'b0;  wr_cycle[ 4738] = 1'b0;  addr_rom[ 4738]='h00000000;  wr_data_rom[ 4738]='h00000000;
    rd_cycle[ 4739] = 1'b0;  wr_cycle[ 4739] = 1'b0;  addr_rom[ 4739]='h00000000;  wr_data_rom[ 4739]='h00000000;
    rd_cycle[ 4740] = 1'b0;  wr_cycle[ 4740] = 1'b0;  addr_rom[ 4740]='h00000000;  wr_data_rom[ 4740]='h00000000;
    rd_cycle[ 4741] = 1'b0;  wr_cycle[ 4741] = 1'b0;  addr_rom[ 4741]='h00000000;  wr_data_rom[ 4741]='h00000000;
    rd_cycle[ 4742] = 1'b0;  wr_cycle[ 4742] = 1'b0;  addr_rom[ 4742]='h00000000;  wr_data_rom[ 4742]='h00000000;
    rd_cycle[ 4743] = 1'b0;  wr_cycle[ 4743] = 1'b0;  addr_rom[ 4743]='h00000000;  wr_data_rom[ 4743]='h00000000;
    rd_cycle[ 4744] = 1'b0;  wr_cycle[ 4744] = 1'b0;  addr_rom[ 4744]='h00000000;  wr_data_rom[ 4744]='h00000000;
    rd_cycle[ 4745] = 1'b0;  wr_cycle[ 4745] = 1'b0;  addr_rom[ 4745]='h00000000;  wr_data_rom[ 4745]='h00000000;
    rd_cycle[ 4746] = 1'b0;  wr_cycle[ 4746] = 1'b0;  addr_rom[ 4746]='h00000000;  wr_data_rom[ 4746]='h00000000;
    rd_cycle[ 4747] = 1'b0;  wr_cycle[ 4747] = 1'b0;  addr_rom[ 4747]='h00000000;  wr_data_rom[ 4747]='h00000000;
    rd_cycle[ 4748] = 1'b0;  wr_cycle[ 4748] = 1'b0;  addr_rom[ 4748]='h00000000;  wr_data_rom[ 4748]='h00000000;
    rd_cycle[ 4749] = 1'b0;  wr_cycle[ 4749] = 1'b0;  addr_rom[ 4749]='h00000000;  wr_data_rom[ 4749]='h00000000;
    rd_cycle[ 4750] = 1'b0;  wr_cycle[ 4750] = 1'b0;  addr_rom[ 4750]='h00000000;  wr_data_rom[ 4750]='h00000000;
    rd_cycle[ 4751] = 1'b0;  wr_cycle[ 4751] = 1'b0;  addr_rom[ 4751]='h00000000;  wr_data_rom[ 4751]='h00000000;
    rd_cycle[ 4752] = 1'b0;  wr_cycle[ 4752] = 1'b0;  addr_rom[ 4752]='h00000000;  wr_data_rom[ 4752]='h00000000;
    rd_cycle[ 4753] = 1'b0;  wr_cycle[ 4753] = 1'b0;  addr_rom[ 4753]='h00000000;  wr_data_rom[ 4753]='h00000000;
    rd_cycle[ 4754] = 1'b0;  wr_cycle[ 4754] = 1'b0;  addr_rom[ 4754]='h00000000;  wr_data_rom[ 4754]='h00000000;
    rd_cycle[ 4755] = 1'b0;  wr_cycle[ 4755] = 1'b0;  addr_rom[ 4755]='h00000000;  wr_data_rom[ 4755]='h00000000;
    rd_cycle[ 4756] = 1'b0;  wr_cycle[ 4756] = 1'b0;  addr_rom[ 4756]='h00000000;  wr_data_rom[ 4756]='h00000000;
    rd_cycle[ 4757] = 1'b0;  wr_cycle[ 4757] = 1'b0;  addr_rom[ 4757]='h00000000;  wr_data_rom[ 4757]='h00000000;
    rd_cycle[ 4758] = 1'b0;  wr_cycle[ 4758] = 1'b0;  addr_rom[ 4758]='h00000000;  wr_data_rom[ 4758]='h00000000;
    rd_cycle[ 4759] = 1'b0;  wr_cycle[ 4759] = 1'b0;  addr_rom[ 4759]='h00000000;  wr_data_rom[ 4759]='h00000000;
    rd_cycle[ 4760] = 1'b0;  wr_cycle[ 4760] = 1'b0;  addr_rom[ 4760]='h00000000;  wr_data_rom[ 4760]='h00000000;
    rd_cycle[ 4761] = 1'b0;  wr_cycle[ 4761] = 1'b0;  addr_rom[ 4761]='h00000000;  wr_data_rom[ 4761]='h00000000;
    rd_cycle[ 4762] = 1'b0;  wr_cycle[ 4762] = 1'b0;  addr_rom[ 4762]='h00000000;  wr_data_rom[ 4762]='h00000000;
    rd_cycle[ 4763] = 1'b0;  wr_cycle[ 4763] = 1'b0;  addr_rom[ 4763]='h00000000;  wr_data_rom[ 4763]='h00000000;
    rd_cycle[ 4764] = 1'b0;  wr_cycle[ 4764] = 1'b0;  addr_rom[ 4764]='h00000000;  wr_data_rom[ 4764]='h00000000;
    rd_cycle[ 4765] = 1'b0;  wr_cycle[ 4765] = 1'b0;  addr_rom[ 4765]='h00000000;  wr_data_rom[ 4765]='h00000000;
    rd_cycle[ 4766] = 1'b0;  wr_cycle[ 4766] = 1'b0;  addr_rom[ 4766]='h00000000;  wr_data_rom[ 4766]='h00000000;
    rd_cycle[ 4767] = 1'b0;  wr_cycle[ 4767] = 1'b0;  addr_rom[ 4767]='h00000000;  wr_data_rom[ 4767]='h00000000;
    rd_cycle[ 4768] = 1'b0;  wr_cycle[ 4768] = 1'b0;  addr_rom[ 4768]='h00000000;  wr_data_rom[ 4768]='h00000000;
    rd_cycle[ 4769] = 1'b0;  wr_cycle[ 4769] = 1'b0;  addr_rom[ 4769]='h00000000;  wr_data_rom[ 4769]='h00000000;
    rd_cycle[ 4770] = 1'b0;  wr_cycle[ 4770] = 1'b0;  addr_rom[ 4770]='h00000000;  wr_data_rom[ 4770]='h00000000;
    rd_cycle[ 4771] = 1'b0;  wr_cycle[ 4771] = 1'b0;  addr_rom[ 4771]='h00000000;  wr_data_rom[ 4771]='h00000000;
    rd_cycle[ 4772] = 1'b0;  wr_cycle[ 4772] = 1'b0;  addr_rom[ 4772]='h00000000;  wr_data_rom[ 4772]='h00000000;
    rd_cycle[ 4773] = 1'b0;  wr_cycle[ 4773] = 1'b0;  addr_rom[ 4773]='h00000000;  wr_data_rom[ 4773]='h00000000;
    rd_cycle[ 4774] = 1'b0;  wr_cycle[ 4774] = 1'b0;  addr_rom[ 4774]='h00000000;  wr_data_rom[ 4774]='h00000000;
    rd_cycle[ 4775] = 1'b0;  wr_cycle[ 4775] = 1'b0;  addr_rom[ 4775]='h00000000;  wr_data_rom[ 4775]='h00000000;
    rd_cycle[ 4776] = 1'b0;  wr_cycle[ 4776] = 1'b0;  addr_rom[ 4776]='h00000000;  wr_data_rom[ 4776]='h00000000;
    rd_cycle[ 4777] = 1'b0;  wr_cycle[ 4777] = 1'b0;  addr_rom[ 4777]='h00000000;  wr_data_rom[ 4777]='h00000000;
    rd_cycle[ 4778] = 1'b0;  wr_cycle[ 4778] = 1'b0;  addr_rom[ 4778]='h00000000;  wr_data_rom[ 4778]='h00000000;
    rd_cycle[ 4779] = 1'b0;  wr_cycle[ 4779] = 1'b0;  addr_rom[ 4779]='h00000000;  wr_data_rom[ 4779]='h00000000;
    rd_cycle[ 4780] = 1'b0;  wr_cycle[ 4780] = 1'b0;  addr_rom[ 4780]='h00000000;  wr_data_rom[ 4780]='h00000000;
    rd_cycle[ 4781] = 1'b0;  wr_cycle[ 4781] = 1'b0;  addr_rom[ 4781]='h00000000;  wr_data_rom[ 4781]='h00000000;
    rd_cycle[ 4782] = 1'b0;  wr_cycle[ 4782] = 1'b0;  addr_rom[ 4782]='h00000000;  wr_data_rom[ 4782]='h00000000;
    rd_cycle[ 4783] = 1'b0;  wr_cycle[ 4783] = 1'b0;  addr_rom[ 4783]='h00000000;  wr_data_rom[ 4783]='h00000000;
    rd_cycle[ 4784] = 1'b0;  wr_cycle[ 4784] = 1'b0;  addr_rom[ 4784]='h00000000;  wr_data_rom[ 4784]='h00000000;
    rd_cycle[ 4785] = 1'b0;  wr_cycle[ 4785] = 1'b0;  addr_rom[ 4785]='h00000000;  wr_data_rom[ 4785]='h00000000;
    rd_cycle[ 4786] = 1'b0;  wr_cycle[ 4786] = 1'b0;  addr_rom[ 4786]='h00000000;  wr_data_rom[ 4786]='h00000000;
    rd_cycle[ 4787] = 1'b0;  wr_cycle[ 4787] = 1'b0;  addr_rom[ 4787]='h00000000;  wr_data_rom[ 4787]='h00000000;
    rd_cycle[ 4788] = 1'b0;  wr_cycle[ 4788] = 1'b0;  addr_rom[ 4788]='h00000000;  wr_data_rom[ 4788]='h00000000;
    rd_cycle[ 4789] = 1'b0;  wr_cycle[ 4789] = 1'b0;  addr_rom[ 4789]='h00000000;  wr_data_rom[ 4789]='h00000000;
    rd_cycle[ 4790] = 1'b0;  wr_cycle[ 4790] = 1'b0;  addr_rom[ 4790]='h00000000;  wr_data_rom[ 4790]='h00000000;
    rd_cycle[ 4791] = 1'b0;  wr_cycle[ 4791] = 1'b0;  addr_rom[ 4791]='h00000000;  wr_data_rom[ 4791]='h00000000;
    rd_cycle[ 4792] = 1'b0;  wr_cycle[ 4792] = 1'b0;  addr_rom[ 4792]='h00000000;  wr_data_rom[ 4792]='h00000000;
    rd_cycle[ 4793] = 1'b0;  wr_cycle[ 4793] = 1'b0;  addr_rom[ 4793]='h00000000;  wr_data_rom[ 4793]='h00000000;
    rd_cycle[ 4794] = 1'b0;  wr_cycle[ 4794] = 1'b0;  addr_rom[ 4794]='h00000000;  wr_data_rom[ 4794]='h00000000;
    rd_cycle[ 4795] = 1'b0;  wr_cycle[ 4795] = 1'b0;  addr_rom[ 4795]='h00000000;  wr_data_rom[ 4795]='h00000000;
    rd_cycle[ 4796] = 1'b0;  wr_cycle[ 4796] = 1'b0;  addr_rom[ 4796]='h00000000;  wr_data_rom[ 4796]='h00000000;
    rd_cycle[ 4797] = 1'b0;  wr_cycle[ 4797] = 1'b0;  addr_rom[ 4797]='h00000000;  wr_data_rom[ 4797]='h00000000;
    rd_cycle[ 4798] = 1'b0;  wr_cycle[ 4798] = 1'b0;  addr_rom[ 4798]='h00000000;  wr_data_rom[ 4798]='h00000000;
    rd_cycle[ 4799] = 1'b0;  wr_cycle[ 4799] = 1'b0;  addr_rom[ 4799]='h00000000;  wr_data_rom[ 4799]='h00000000;
    rd_cycle[ 4800] = 1'b0;  wr_cycle[ 4800] = 1'b0;  addr_rom[ 4800]='h00000000;  wr_data_rom[ 4800]='h00000000;
    rd_cycle[ 4801] = 1'b0;  wr_cycle[ 4801] = 1'b0;  addr_rom[ 4801]='h00000000;  wr_data_rom[ 4801]='h00000000;
    rd_cycle[ 4802] = 1'b0;  wr_cycle[ 4802] = 1'b0;  addr_rom[ 4802]='h00000000;  wr_data_rom[ 4802]='h00000000;
    rd_cycle[ 4803] = 1'b0;  wr_cycle[ 4803] = 1'b0;  addr_rom[ 4803]='h00000000;  wr_data_rom[ 4803]='h00000000;
    rd_cycle[ 4804] = 1'b0;  wr_cycle[ 4804] = 1'b0;  addr_rom[ 4804]='h00000000;  wr_data_rom[ 4804]='h00000000;
    rd_cycle[ 4805] = 1'b0;  wr_cycle[ 4805] = 1'b0;  addr_rom[ 4805]='h00000000;  wr_data_rom[ 4805]='h00000000;
    rd_cycle[ 4806] = 1'b0;  wr_cycle[ 4806] = 1'b0;  addr_rom[ 4806]='h00000000;  wr_data_rom[ 4806]='h00000000;
    rd_cycle[ 4807] = 1'b0;  wr_cycle[ 4807] = 1'b0;  addr_rom[ 4807]='h00000000;  wr_data_rom[ 4807]='h00000000;
    rd_cycle[ 4808] = 1'b0;  wr_cycle[ 4808] = 1'b0;  addr_rom[ 4808]='h00000000;  wr_data_rom[ 4808]='h00000000;
    rd_cycle[ 4809] = 1'b0;  wr_cycle[ 4809] = 1'b0;  addr_rom[ 4809]='h00000000;  wr_data_rom[ 4809]='h00000000;
    rd_cycle[ 4810] = 1'b0;  wr_cycle[ 4810] = 1'b0;  addr_rom[ 4810]='h00000000;  wr_data_rom[ 4810]='h00000000;
    rd_cycle[ 4811] = 1'b0;  wr_cycle[ 4811] = 1'b0;  addr_rom[ 4811]='h00000000;  wr_data_rom[ 4811]='h00000000;
    rd_cycle[ 4812] = 1'b0;  wr_cycle[ 4812] = 1'b0;  addr_rom[ 4812]='h00000000;  wr_data_rom[ 4812]='h00000000;
    rd_cycle[ 4813] = 1'b0;  wr_cycle[ 4813] = 1'b0;  addr_rom[ 4813]='h00000000;  wr_data_rom[ 4813]='h00000000;
    rd_cycle[ 4814] = 1'b0;  wr_cycle[ 4814] = 1'b0;  addr_rom[ 4814]='h00000000;  wr_data_rom[ 4814]='h00000000;
    rd_cycle[ 4815] = 1'b0;  wr_cycle[ 4815] = 1'b0;  addr_rom[ 4815]='h00000000;  wr_data_rom[ 4815]='h00000000;
    rd_cycle[ 4816] = 1'b0;  wr_cycle[ 4816] = 1'b0;  addr_rom[ 4816]='h00000000;  wr_data_rom[ 4816]='h00000000;
    rd_cycle[ 4817] = 1'b0;  wr_cycle[ 4817] = 1'b0;  addr_rom[ 4817]='h00000000;  wr_data_rom[ 4817]='h00000000;
    rd_cycle[ 4818] = 1'b0;  wr_cycle[ 4818] = 1'b0;  addr_rom[ 4818]='h00000000;  wr_data_rom[ 4818]='h00000000;
    rd_cycle[ 4819] = 1'b0;  wr_cycle[ 4819] = 1'b0;  addr_rom[ 4819]='h00000000;  wr_data_rom[ 4819]='h00000000;
    rd_cycle[ 4820] = 1'b0;  wr_cycle[ 4820] = 1'b0;  addr_rom[ 4820]='h00000000;  wr_data_rom[ 4820]='h00000000;
    rd_cycle[ 4821] = 1'b0;  wr_cycle[ 4821] = 1'b0;  addr_rom[ 4821]='h00000000;  wr_data_rom[ 4821]='h00000000;
    rd_cycle[ 4822] = 1'b0;  wr_cycle[ 4822] = 1'b0;  addr_rom[ 4822]='h00000000;  wr_data_rom[ 4822]='h00000000;
    rd_cycle[ 4823] = 1'b0;  wr_cycle[ 4823] = 1'b0;  addr_rom[ 4823]='h00000000;  wr_data_rom[ 4823]='h00000000;
    rd_cycle[ 4824] = 1'b0;  wr_cycle[ 4824] = 1'b0;  addr_rom[ 4824]='h00000000;  wr_data_rom[ 4824]='h00000000;
    rd_cycle[ 4825] = 1'b0;  wr_cycle[ 4825] = 1'b0;  addr_rom[ 4825]='h00000000;  wr_data_rom[ 4825]='h00000000;
    rd_cycle[ 4826] = 1'b0;  wr_cycle[ 4826] = 1'b0;  addr_rom[ 4826]='h00000000;  wr_data_rom[ 4826]='h00000000;
    rd_cycle[ 4827] = 1'b0;  wr_cycle[ 4827] = 1'b0;  addr_rom[ 4827]='h00000000;  wr_data_rom[ 4827]='h00000000;
    rd_cycle[ 4828] = 1'b0;  wr_cycle[ 4828] = 1'b0;  addr_rom[ 4828]='h00000000;  wr_data_rom[ 4828]='h00000000;
    rd_cycle[ 4829] = 1'b0;  wr_cycle[ 4829] = 1'b0;  addr_rom[ 4829]='h00000000;  wr_data_rom[ 4829]='h00000000;
    rd_cycle[ 4830] = 1'b0;  wr_cycle[ 4830] = 1'b0;  addr_rom[ 4830]='h00000000;  wr_data_rom[ 4830]='h00000000;
    rd_cycle[ 4831] = 1'b0;  wr_cycle[ 4831] = 1'b0;  addr_rom[ 4831]='h00000000;  wr_data_rom[ 4831]='h00000000;
    rd_cycle[ 4832] = 1'b0;  wr_cycle[ 4832] = 1'b0;  addr_rom[ 4832]='h00000000;  wr_data_rom[ 4832]='h00000000;
    rd_cycle[ 4833] = 1'b0;  wr_cycle[ 4833] = 1'b0;  addr_rom[ 4833]='h00000000;  wr_data_rom[ 4833]='h00000000;
    rd_cycle[ 4834] = 1'b0;  wr_cycle[ 4834] = 1'b0;  addr_rom[ 4834]='h00000000;  wr_data_rom[ 4834]='h00000000;
    rd_cycle[ 4835] = 1'b0;  wr_cycle[ 4835] = 1'b0;  addr_rom[ 4835]='h00000000;  wr_data_rom[ 4835]='h00000000;
    rd_cycle[ 4836] = 1'b0;  wr_cycle[ 4836] = 1'b0;  addr_rom[ 4836]='h00000000;  wr_data_rom[ 4836]='h00000000;
    rd_cycle[ 4837] = 1'b0;  wr_cycle[ 4837] = 1'b0;  addr_rom[ 4837]='h00000000;  wr_data_rom[ 4837]='h00000000;
    rd_cycle[ 4838] = 1'b0;  wr_cycle[ 4838] = 1'b0;  addr_rom[ 4838]='h00000000;  wr_data_rom[ 4838]='h00000000;
    rd_cycle[ 4839] = 1'b0;  wr_cycle[ 4839] = 1'b0;  addr_rom[ 4839]='h00000000;  wr_data_rom[ 4839]='h00000000;
    rd_cycle[ 4840] = 1'b0;  wr_cycle[ 4840] = 1'b0;  addr_rom[ 4840]='h00000000;  wr_data_rom[ 4840]='h00000000;
    rd_cycle[ 4841] = 1'b0;  wr_cycle[ 4841] = 1'b0;  addr_rom[ 4841]='h00000000;  wr_data_rom[ 4841]='h00000000;
    rd_cycle[ 4842] = 1'b0;  wr_cycle[ 4842] = 1'b0;  addr_rom[ 4842]='h00000000;  wr_data_rom[ 4842]='h00000000;
    rd_cycle[ 4843] = 1'b0;  wr_cycle[ 4843] = 1'b0;  addr_rom[ 4843]='h00000000;  wr_data_rom[ 4843]='h00000000;
    rd_cycle[ 4844] = 1'b0;  wr_cycle[ 4844] = 1'b0;  addr_rom[ 4844]='h00000000;  wr_data_rom[ 4844]='h00000000;
    rd_cycle[ 4845] = 1'b0;  wr_cycle[ 4845] = 1'b0;  addr_rom[ 4845]='h00000000;  wr_data_rom[ 4845]='h00000000;
    rd_cycle[ 4846] = 1'b0;  wr_cycle[ 4846] = 1'b0;  addr_rom[ 4846]='h00000000;  wr_data_rom[ 4846]='h00000000;
    rd_cycle[ 4847] = 1'b0;  wr_cycle[ 4847] = 1'b0;  addr_rom[ 4847]='h00000000;  wr_data_rom[ 4847]='h00000000;
    rd_cycle[ 4848] = 1'b0;  wr_cycle[ 4848] = 1'b0;  addr_rom[ 4848]='h00000000;  wr_data_rom[ 4848]='h00000000;
    rd_cycle[ 4849] = 1'b0;  wr_cycle[ 4849] = 1'b0;  addr_rom[ 4849]='h00000000;  wr_data_rom[ 4849]='h00000000;
    rd_cycle[ 4850] = 1'b0;  wr_cycle[ 4850] = 1'b0;  addr_rom[ 4850]='h00000000;  wr_data_rom[ 4850]='h00000000;
    rd_cycle[ 4851] = 1'b0;  wr_cycle[ 4851] = 1'b0;  addr_rom[ 4851]='h00000000;  wr_data_rom[ 4851]='h00000000;
    rd_cycle[ 4852] = 1'b0;  wr_cycle[ 4852] = 1'b0;  addr_rom[ 4852]='h00000000;  wr_data_rom[ 4852]='h00000000;
    rd_cycle[ 4853] = 1'b0;  wr_cycle[ 4853] = 1'b0;  addr_rom[ 4853]='h00000000;  wr_data_rom[ 4853]='h00000000;
    rd_cycle[ 4854] = 1'b0;  wr_cycle[ 4854] = 1'b0;  addr_rom[ 4854]='h00000000;  wr_data_rom[ 4854]='h00000000;
    rd_cycle[ 4855] = 1'b0;  wr_cycle[ 4855] = 1'b0;  addr_rom[ 4855]='h00000000;  wr_data_rom[ 4855]='h00000000;
    rd_cycle[ 4856] = 1'b0;  wr_cycle[ 4856] = 1'b0;  addr_rom[ 4856]='h00000000;  wr_data_rom[ 4856]='h00000000;
    rd_cycle[ 4857] = 1'b0;  wr_cycle[ 4857] = 1'b0;  addr_rom[ 4857]='h00000000;  wr_data_rom[ 4857]='h00000000;
    rd_cycle[ 4858] = 1'b0;  wr_cycle[ 4858] = 1'b0;  addr_rom[ 4858]='h00000000;  wr_data_rom[ 4858]='h00000000;
    rd_cycle[ 4859] = 1'b0;  wr_cycle[ 4859] = 1'b0;  addr_rom[ 4859]='h00000000;  wr_data_rom[ 4859]='h00000000;
    rd_cycle[ 4860] = 1'b0;  wr_cycle[ 4860] = 1'b0;  addr_rom[ 4860]='h00000000;  wr_data_rom[ 4860]='h00000000;
    rd_cycle[ 4861] = 1'b0;  wr_cycle[ 4861] = 1'b0;  addr_rom[ 4861]='h00000000;  wr_data_rom[ 4861]='h00000000;
    rd_cycle[ 4862] = 1'b0;  wr_cycle[ 4862] = 1'b0;  addr_rom[ 4862]='h00000000;  wr_data_rom[ 4862]='h00000000;
    rd_cycle[ 4863] = 1'b0;  wr_cycle[ 4863] = 1'b0;  addr_rom[ 4863]='h00000000;  wr_data_rom[ 4863]='h00000000;
    rd_cycle[ 4864] = 1'b0;  wr_cycle[ 4864] = 1'b0;  addr_rom[ 4864]='h00000000;  wr_data_rom[ 4864]='h00000000;
    rd_cycle[ 4865] = 1'b0;  wr_cycle[ 4865] = 1'b0;  addr_rom[ 4865]='h00000000;  wr_data_rom[ 4865]='h00000000;
    rd_cycle[ 4866] = 1'b0;  wr_cycle[ 4866] = 1'b0;  addr_rom[ 4866]='h00000000;  wr_data_rom[ 4866]='h00000000;
    rd_cycle[ 4867] = 1'b0;  wr_cycle[ 4867] = 1'b0;  addr_rom[ 4867]='h00000000;  wr_data_rom[ 4867]='h00000000;
    rd_cycle[ 4868] = 1'b0;  wr_cycle[ 4868] = 1'b0;  addr_rom[ 4868]='h00000000;  wr_data_rom[ 4868]='h00000000;
    rd_cycle[ 4869] = 1'b0;  wr_cycle[ 4869] = 1'b0;  addr_rom[ 4869]='h00000000;  wr_data_rom[ 4869]='h00000000;
    rd_cycle[ 4870] = 1'b0;  wr_cycle[ 4870] = 1'b0;  addr_rom[ 4870]='h00000000;  wr_data_rom[ 4870]='h00000000;
    rd_cycle[ 4871] = 1'b0;  wr_cycle[ 4871] = 1'b0;  addr_rom[ 4871]='h00000000;  wr_data_rom[ 4871]='h00000000;
    rd_cycle[ 4872] = 1'b0;  wr_cycle[ 4872] = 1'b0;  addr_rom[ 4872]='h00000000;  wr_data_rom[ 4872]='h00000000;
    rd_cycle[ 4873] = 1'b0;  wr_cycle[ 4873] = 1'b0;  addr_rom[ 4873]='h00000000;  wr_data_rom[ 4873]='h00000000;
    rd_cycle[ 4874] = 1'b0;  wr_cycle[ 4874] = 1'b0;  addr_rom[ 4874]='h00000000;  wr_data_rom[ 4874]='h00000000;
    rd_cycle[ 4875] = 1'b0;  wr_cycle[ 4875] = 1'b0;  addr_rom[ 4875]='h00000000;  wr_data_rom[ 4875]='h00000000;
    rd_cycle[ 4876] = 1'b0;  wr_cycle[ 4876] = 1'b0;  addr_rom[ 4876]='h00000000;  wr_data_rom[ 4876]='h00000000;
    rd_cycle[ 4877] = 1'b0;  wr_cycle[ 4877] = 1'b0;  addr_rom[ 4877]='h00000000;  wr_data_rom[ 4877]='h00000000;
    rd_cycle[ 4878] = 1'b0;  wr_cycle[ 4878] = 1'b0;  addr_rom[ 4878]='h00000000;  wr_data_rom[ 4878]='h00000000;
    rd_cycle[ 4879] = 1'b0;  wr_cycle[ 4879] = 1'b0;  addr_rom[ 4879]='h00000000;  wr_data_rom[ 4879]='h00000000;
    rd_cycle[ 4880] = 1'b0;  wr_cycle[ 4880] = 1'b0;  addr_rom[ 4880]='h00000000;  wr_data_rom[ 4880]='h00000000;
    rd_cycle[ 4881] = 1'b0;  wr_cycle[ 4881] = 1'b0;  addr_rom[ 4881]='h00000000;  wr_data_rom[ 4881]='h00000000;
    rd_cycle[ 4882] = 1'b0;  wr_cycle[ 4882] = 1'b0;  addr_rom[ 4882]='h00000000;  wr_data_rom[ 4882]='h00000000;
    rd_cycle[ 4883] = 1'b0;  wr_cycle[ 4883] = 1'b0;  addr_rom[ 4883]='h00000000;  wr_data_rom[ 4883]='h00000000;
    rd_cycle[ 4884] = 1'b0;  wr_cycle[ 4884] = 1'b0;  addr_rom[ 4884]='h00000000;  wr_data_rom[ 4884]='h00000000;
    rd_cycle[ 4885] = 1'b0;  wr_cycle[ 4885] = 1'b0;  addr_rom[ 4885]='h00000000;  wr_data_rom[ 4885]='h00000000;
    rd_cycle[ 4886] = 1'b0;  wr_cycle[ 4886] = 1'b0;  addr_rom[ 4886]='h00000000;  wr_data_rom[ 4886]='h00000000;
    rd_cycle[ 4887] = 1'b0;  wr_cycle[ 4887] = 1'b0;  addr_rom[ 4887]='h00000000;  wr_data_rom[ 4887]='h00000000;
    rd_cycle[ 4888] = 1'b0;  wr_cycle[ 4888] = 1'b0;  addr_rom[ 4888]='h00000000;  wr_data_rom[ 4888]='h00000000;
    rd_cycle[ 4889] = 1'b0;  wr_cycle[ 4889] = 1'b0;  addr_rom[ 4889]='h00000000;  wr_data_rom[ 4889]='h00000000;
    rd_cycle[ 4890] = 1'b0;  wr_cycle[ 4890] = 1'b0;  addr_rom[ 4890]='h00000000;  wr_data_rom[ 4890]='h00000000;
    rd_cycle[ 4891] = 1'b0;  wr_cycle[ 4891] = 1'b0;  addr_rom[ 4891]='h00000000;  wr_data_rom[ 4891]='h00000000;
    rd_cycle[ 4892] = 1'b0;  wr_cycle[ 4892] = 1'b0;  addr_rom[ 4892]='h00000000;  wr_data_rom[ 4892]='h00000000;
    rd_cycle[ 4893] = 1'b0;  wr_cycle[ 4893] = 1'b0;  addr_rom[ 4893]='h00000000;  wr_data_rom[ 4893]='h00000000;
    rd_cycle[ 4894] = 1'b0;  wr_cycle[ 4894] = 1'b0;  addr_rom[ 4894]='h00000000;  wr_data_rom[ 4894]='h00000000;
    rd_cycle[ 4895] = 1'b0;  wr_cycle[ 4895] = 1'b0;  addr_rom[ 4895]='h00000000;  wr_data_rom[ 4895]='h00000000;
    rd_cycle[ 4896] = 1'b0;  wr_cycle[ 4896] = 1'b0;  addr_rom[ 4896]='h00000000;  wr_data_rom[ 4896]='h00000000;
    rd_cycle[ 4897] = 1'b0;  wr_cycle[ 4897] = 1'b0;  addr_rom[ 4897]='h00000000;  wr_data_rom[ 4897]='h00000000;
    rd_cycle[ 4898] = 1'b0;  wr_cycle[ 4898] = 1'b0;  addr_rom[ 4898]='h00000000;  wr_data_rom[ 4898]='h00000000;
    rd_cycle[ 4899] = 1'b0;  wr_cycle[ 4899] = 1'b0;  addr_rom[ 4899]='h00000000;  wr_data_rom[ 4899]='h00000000;
    rd_cycle[ 4900] = 1'b0;  wr_cycle[ 4900] = 1'b0;  addr_rom[ 4900]='h00000000;  wr_data_rom[ 4900]='h00000000;
    rd_cycle[ 4901] = 1'b0;  wr_cycle[ 4901] = 1'b0;  addr_rom[ 4901]='h00000000;  wr_data_rom[ 4901]='h00000000;
    rd_cycle[ 4902] = 1'b0;  wr_cycle[ 4902] = 1'b0;  addr_rom[ 4902]='h00000000;  wr_data_rom[ 4902]='h00000000;
    rd_cycle[ 4903] = 1'b0;  wr_cycle[ 4903] = 1'b0;  addr_rom[ 4903]='h00000000;  wr_data_rom[ 4903]='h00000000;
    rd_cycle[ 4904] = 1'b0;  wr_cycle[ 4904] = 1'b0;  addr_rom[ 4904]='h00000000;  wr_data_rom[ 4904]='h00000000;
    rd_cycle[ 4905] = 1'b0;  wr_cycle[ 4905] = 1'b0;  addr_rom[ 4905]='h00000000;  wr_data_rom[ 4905]='h00000000;
    rd_cycle[ 4906] = 1'b0;  wr_cycle[ 4906] = 1'b0;  addr_rom[ 4906]='h00000000;  wr_data_rom[ 4906]='h00000000;
    rd_cycle[ 4907] = 1'b0;  wr_cycle[ 4907] = 1'b0;  addr_rom[ 4907]='h00000000;  wr_data_rom[ 4907]='h00000000;
    rd_cycle[ 4908] = 1'b0;  wr_cycle[ 4908] = 1'b0;  addr_rom[ 4908]='h00000000;  wr_data_rom[ 4908]='h00000000;
    rd_cycle[ 4909] = 1'b0;  wr_cycle[ 4909] = 1'b0;  addr_rom[ 4909]='h00000000;  wr_data_rom[ 4909]='h00000000;
    rd_cycle[ 4910] = 1'b0;  wr_cycle[ 4910] = 1'b0;  addr_rom[ 4910]='h00000000;  wr_data_rom[ 4910]='h00000000;
    rd_cycle[ 4911] = 1'b0;  wr_cycle[ 4911] = 1'b0;  addr_rom[ 4911]='h00000000;  wr_data_rom[ 4911]='h00000000;
    rd_cycle[ 4912] = 1'b0;  wr_cycle[ 4912] = 1'b0;  addr_rom[ 4912]='h00000000;  wr_data_rom[ 4912]='h00000000;
    rd_cycle[ 4913] = 1'b0;  wr_cycle[ 4913] = 1'b0;  addr_rom[ 4913]='h00000000;  wr_data_rom[ 4913]='h00000000;
    rd_cycle[ 4914] = 1'b0;  wr_cycle[ 4914] = 1'b0;  addr_rom[ 4914]='h00000000;  wr_data_rom[ 4914]='h00000000;
    rd_cycle[ 4915] = 1'b0;  wr_cycle[ 4915] = 1'b0;  addr_rom[ 4915]='h00000000;  wr_data_rom[ 4915]='h00000000;
    rd_cycle[ 4916] = 1'b0;  wr_cycle[ 4916] = 1'b0;  addr_rom[ 4916]='h00000000;  wr_data_rom[ 4916]='h00000000;
    rd_cycle[ 4917] = 1'b0;  wr_cycle[ 4917] = 1'b0;  addr_rom[ 4917]='h00000000;  wr_data_rom[ 4917]='h00000000;
    rd_cycle[ 4918] = 1'b0;  wr_cycle[ 4918] = 1'b0;  addr_rom[ 4918]='h00000000;  wr_data_rom[ 4918]='h00000000;
    rd_cycle[ 4919] = 1'b0;  wr_cycle[ 4919] = 1'b0;  addr_rom[ 4919]='h00000000;  wr_data_rom[ 4919]='h00000000;
    rd_cycle[ 4920] = 1'b0;  wr_cycle[ 4920] = 1'b0;  addr_rom[ 4920]='h00000000;  wr_data_rom[ 4920]='h00000000;
    rd_cycle[ 4921] = 1'b0;  wr_cycle[ 4921] = 1'b0;  addr_rom[ 4921]='h00000000;  wr_data_rom[ 4921]='h00000000;
    rd_cycle[ 4922] = 1'b0;  wr_cycle[ 4922] = 1'b0;  addr_rom[ 4922]='h00000000;  wr_data_rom[ 4922]='h00000000;
    rd_cycle[ 4923] = 1'b0;  wr_cycle[ 4923] = 1'b0;  addr_rom[ 4923]='h00000000;  wr_data_rom[ 4923]='h00000000;
    rd_cycle[ 4924] = 1'b0;  wr_cycle[ 4924] = 1'b0;  addr_rom[ 4924]='h00000000;  wr_data_rom[ 4924]='h00000000;
    rd_cycle[ 4925] = 1'b0;  wr_cycle[ 4925] = 1'b0;  addr_rom[ 4925]='h00000000;  wr_data_rom[ 4925]='h00000000;
    rd_cycle[ 4926] = 1'b0;  wr_cycle[ 4926] = 1'b0;  addr_rom[ 4926]='h00000000;  wr_data_rom[ 4926]='h00000000;
    rd_cycle[ 4927] = 1'b0;  wr_cycle[ 4927] = 1'b0;  addr_rom[ 4927]='h00000000;  wr_data_rom[ 4927]='h00000000;
    rd_cycle[ 4928] = 1'b0;  wr_cycle[ 4928] = 1'b0;  addr_rom[ 4928]='h00000000;  wr_data_rom[ 4928]='h00000000;
    rd_cycle[ 4929] = 1'b0;  wr_cycle[ 4929] = 1'b0;  addr_rom[ 4929]='h00000000;  wr_data_rom[ 4929]='h00000000;
    rd_cycle[ 4930] = 1'b0;  wr_cycle[ 4930] = 1'b0;  addr_rom[ 4930]='h00000000;  wr_data_rom[ 4930]='h00000000;
    rd_cycle[ 4931] = 1'b0;  wr_cycle[ 4931] = 1'b0;  addr_rom[ 4931]='h00000000;  wr_data_rom[ 4931]='h00000000;
    rd_cycle[ 4932] = 1'b0;  wr_cycle[ 4932] = 1'b0;  addr_rom[ 4932]='h00000000;  wr_data_rom[ 4932]='h00000000;
    rd_cycle[ 4933] = 1'b0;  wr_cycle[ 4933] = 1'b0;  addr_rom[ 4933]='h00000000;  wr_data_rom[ 4933]='h00000000;
    rd_cycle[ 4934] = 1'b0;  wr_cycle[ 4934] = 1'b0;  addr_rom[ 4934]='h00000000;  wr_data_rom[ 4934]='h00000000;
    rd_cycle[ 4935] = 1'b0;  wr_cycle[ 4935] = 1'b0;  addr_rom[ 4935]='h00000000;  wr_data_rom[ 4935]='h00000000;
    rd_cycle[ 4936] = 1'b0;  wr_cycle[ 4936] = 1'b0;  addr_rom[ 4936]='h00000000;  wr_data_rom[ 4936]='h00000000;
    rd_cycle[ 4937] = 1'b0;  wr_cycle[ 4937] = 1'b0;  addr_rom[ 4937]='h00000000;  wr_data_rom[ 4937]='h00000000;
    rd_cycle[ 4938] = 1'b0;  wr_cycle[ 4938] = 1'b0;  addr_rom[ 4938]='h00000000;  wr_data_rom[ 4938]='h00000000;
    rd_cycle[ 4939] = 1'b0;  wr_cycle[ 4939] = 1'b0;  addr_rom[ 4939]='h00000000;  wr_data_rom[ 4939]='h00000000;
    rd_cycle[ 4940] = 1'b0;  wr_cycle[ 4940] = 1'b0;  addr_rom[ 4940]='h00000000;  wr_data_rom[ 4940]='h00000000;
    rd_cycle[ 4941] = 1'b0;  wr_cycle[ 4941] = 1'b0;  addr_rom[ 4941]='h00000000;  wr_data_rom[ 4941]='h00000000;
    rd_cycle[ 4942] = 1'b0;  wr_cycle[ 4942] = 1'b0;  addr_rom[ 4942]='h00000000;  wr_data_rom[ 4942]='h00000000;
    rd_cycle[ 4943] = 1'b0;  wr_cycle[ 4943] = 1'b0;  addr_rom[ 4943]='h00000000;  wr_data_rom[ 4943]='h00000000;
    rd_cycle[ 4944] = 1'b0;  wr_cycle[ 4944] = 1'b0;  addr_rom[ 4944]='h00000000;  wr_data_rom[ 4944]='h00000000;
    rd_cycle[ 4945] = 1'b0;  wr_cycle[ 4945] = 1'b0;  addr_rom[ 4945]='h00000000;  wr_data_rom[ 4945]='h00000000;
    rd_cycle[ 4946] = 1'b0;  wr_cycle[ 4946] = 1'b0;  addr_rom[ 4946]='h00000000;  wr_data_rom[ 4946]='h00000000;
    rd_cycle[ 4947] = 1'b0;  wr_cycle[ 4947] = 1'b0;  addr_rom[ 4947]='h00000000;  wr_data_rom[ 4947]='h00000000;
    rd_cycle[ 4948] = 1'b0;  wr_cycle[ 4948] = 1'b0;  addr_rom[ 4948]='h00000000;  wr_data_rom[ 4948]='h00000000;
    rd_cycle[ 4949] = 1'b0;  wr_cycle[ 4949] = 1'b0;  addr_rom[ 4949]='h00000000;  wr_data_rom[ 4949]='h00000000;
    rd_cycle[ 4950] = 1'b0;  wr_cycle[ 4950] = 1'b0;  addr_rom[ 4950]='h00000000;  wr_data_rom[ 4950]='h00000000;
    rd_cycle[ 4951] = 1'b0;  wr_cycle[ 4951] = 1'b0;  addr_rom[ 4951]='h00000000;  wr_data_rom[ 4951]='h00000000;
    rd_cycle[ 4952] = 1'b0;  wr_cycle[ 4952] = 1'b0;  addr_rom[ 4952]='h00000000;  wr_data_rom[ 4952]='h00000000;
    rd_cycle[ 4953] = 1'b0;  wr_cycle[ 4953] = 1'b0;  addr_rom[ 4953]='h00000000;  wr_data_rom[ 4953]='h00000000;
    rd_cycle[ 4954] = 1'b0;  wr_cycle[ 4954] = 1'b0;  addr_rom[ 4954]='h00000000;  wr_data_rom[ 4954]='h00000000;
    rd_cycle[ 4955] = 1'b0;  wr_cycle[ 4955] = 1'b0;  addr_rom[ 4955]='h00000000;  wr_data_rom[ 4955]='h00000000;
    rd_cycle[ 4956] = 1'b0;  wr_cycle[ 4956] = 1'b0;  addr_rom[ 4956]='h00000000;  wr_data_rom[ 4956]='h00000000;
    rd_cycle[ 4957] = 1'b0;  wr_cycle[ 4957] = 1'b0;  addr_rom[ 4957]='h00000000;  wr_data_rom[ 4957]='h00000000;
    rd_cycle[ 4958] = 1'b0;  wr_cycle[ 4958] = 1'b0;  addr_rom[ 4958]='h00000000;  wr_data_rom[ 4958]='h00000000;
    rd_cycle[ 4959] = 1'b0;  wr_cycle[ 4959] = 1'b0;  addr_rom[ 4959]='h00000000;  wr_data_rom[ 4959]='h00000000;
    rd_cycle[ 4960] = 1'b0;  wr_cycle[ 4960] = 1'b0;  addr_rom[ 4960]='h00000000;  wr_data_rom[ 4960]='h00000000;
    rd_cycle[ 4961] = 1'b0;  wr_cycle[ 4961] = 1'b0;  addr_rom[ 4961]='h00000000;  wr_data_rom[ 4961]='h00000000;
    rd_cycle[ 4962] = 1'b0;  wr_cycle[ 4962] = 1'b0;  addr_rom[ 4962]='h00000000;  wr_data_rom[ 4962]='h00000000;
    rd_cycle[ 4963] = 1'b0;  wr_cycle[ 4963] = 1'b0;  addr_rom[ 4963]='h00000000;  wr_data_rom[ 4963]='h00000000;
    rd_cycle[ 4964] = 1'b0;  wr_cycle[ 4964] = 1'b0;  addr_rom[ 4964]='h00000000;  wr_data_rom[ 4964]='h00000000;
    rd_cycle[ 4965] = 1'b0;  wr_cycle[ 4965] = 1'b0;  addr_rom[ 4965]='h00000000;  wr_data_rom[ 4965]='h00000000;
    rd_cycle[ 4966] = 1'b0;  wr_cycle[ 4966] = 1'b0;  addr_rom[ 4966]='h00000000;  wr_data_rom[ 4966]='h00000000;
    rd_cycle[ 4967] = 1'b0;  wr_cycle[ 4967] = 1'b0;  addr_rom[ 4967]='h00000000;  wr_data_rom[ 4967]='h00000000;
    rd_cycle[ 4968] = 1'b0;  wr_cycle[ 4968] = 1'b0;  addr_rom[ 4968]='h00000000;  wr_data_rom[ 4968]='h00000000;
    rd_cycle[ 4969] = 1'b0;  wr_cycle[ 4969] = 1'b0;  addr_rom[ 4969]='h00000000;  wr_data_rom[ 4969]='h00000000;
    rd_cycle[ 4970] = 1'b0;  wr_cycle[ 4970] = 1'b0;  addr_rom[ 4970]='h00000000;  wr_data_rom[ 4970]='h00000000;
    rd_cycle[ 4971] = 1'b0;  wr_cycle[ 4971] = 1'b0;  addr_rom[ 4971]='h00000000;  wr_data_rom[ 4971]='h00000000;
    rd_cycle[ 4972] = 1'b0;  wr_cycle[ 4972] = 1'b0;  addr_rom[ 4972]='h00000000;  wr_data_rom[ 4972]='h00000000;
    rd_cycle[ 4973] = 1'b0;  wr_cycle[ 4973] = 1'b0;  addr_rom[ 4973]='h00000000;  wr_data_rom[ 4973]='h00000000;
    rd_cycle[ 4974] = 1'b0;  wr_cycle[ 4974] = 1'b0;  addr_rom[ 4974]='h00000000;  wr_data_rom[ 4974]='h00000000;
    rd_cycle[ 4975] = 1'b0;  wr_cycle[ 4975] = 1'b0;  addr_rom[ 4975]='h00000000;  wr_data_rom[ 4975]='h00000000;
    rd_cycle[ 4976] = 1'b0;  wr_cycle[ 4976] = 1'b0;  addr_rom[ 4976]='h00000000;  wr_data_rom[ 4976]='h00000000;
    rd_cycle[ 4977] = 1'b0;  wr_cycle[ 4977] = 1'b0;  addr_rom[ 4977]='h00000000;  wr_data_rom[ 4977]='h00000000;
    rd_cycle[ 4978] = 1'b0;  wr_cycle[ 4978] = 1'b0;  addr_rom[ 4978]='h00000000;  wr_data_rom[ 4978]='h00000000;
    rd_cycle[ 4979] = 1'b0;  wr_cycle[ 4979] = 1'b0;  addr_rom[ 4979]='h00000000;  wr_data_rom[ 4979]='h00000000;
    rd_cycle[ 4980] = 1'b0;  wr_cycle[ 4980] = 1'b0;  addr_rom[ 4980]='h00000000;  wr_data_rom[ 4980]='h00000000;
    rd_cycle[ 4981] = 1'b0;  wr_cycle[ 4981] = 1'b0;  addr_rom[ 4981]='h00000000;  wr_data_rom[ 4981]='h00000000;
    rd_cycle[ 4982] = 1'b0;  wr_cycle[ 4982] = 1'b0;  addr_rom[ 4982]='h00000000;  wr_data_rom[ 4982]='h00000000;
    rd_cycle[ 4983] = 1'b0;  wr_cycle[ 4983] = 1'b0;  addr_rom[ 4983]='h00000000;  wr_data_rom[ 4983]='h00000000;
    rd_cycle[ 4984] = 1'b0;  wr_cycle[ 4984] = 1'b0;  addr_rom[ 4984]='h00000000;  wr_data_rom[ 4984]='h00000000;
    rd_cycle[ 4985] = 1'b0;  wr_cycle[ 4985] = 1'b0;  addr_rom[ 4985]='h00000000;  wr_data_rom[ 4985]='h00000000;
    rd_cycle[ 4986] = 1'b0;  wr_cycle[ 4986] = 1'b0;  addr_rom[ 4986]='h00000000;  wr_data_rom[ 4986]='h00000000;
    rd_cycle[ 4987] = 1'b0;  wr_cycle[ 4987] = 1'b0;  addr_rom[ 4987]='h00000000;  wr_data_rom[ 4987]='h00000000;
    rd_cycle[ 4988] = 1'b0;  wr_cycle[ 4988] = 1'b0;  addr_rom[ 4988]='h00000000;  wr_data_rom[ 4988]='h00000000;
    rd_cycle[ 4989] = 1'b0;  wr_cycle[ 4989] = 1'b0;  addr_rom[ 4989]='h00000000;  wr_data_rom[ 4989]='h00000000;
    rd_cycle[ 4990] = 1'b0;  wr_cycle[ 4990] = 1'b0;  addr_rom[ 4990]='h00000000;  wr_data_rom[ 4990]='h00000000;
    rd_cycle[ 4991] = 1'b0;  wr_cycle[ 4991] = 1'b0;  addr_rom[ 4991]='h00000000;  wr_data_rom[ 4991]='h00000000;
    rd_cycle[ 4992] = 1'b0;  wr_cycle[ 4992] = 1'b0;  addr_rom[ 4992]='h00000000;  wr_data_rom[ 4992]='h00000000;
    rd_cycle[ 4993] = 1'b0;  wr_cycle[ 4993] = 1'b0;  addr_rom[ 4993]='h00000000;  wr_data_rom[ 4993]='h00000000;
    rd_cycle[ 4994] = 1'b0;  wr_cycle[ 4994] = 1'b0;  addr_rom[ 4994]='h00000000;  wr_data_rom[ 4994]='h00000000;
    rd_cycle[ 4995] = 1'b0;  wr_cycle[ 4995] = 1'b0;  addr_rom[ 4995]='h00000000;  wr_data_rom[ 4995]='h00000000;
    rd_cycle[ 4996] = 1'b0;  wr_cycle[ 4996] = 1'b0;  addr_rom[ 4996]='h00000000;  wr_data_rom[ 4996]='h00000000;
    rd_cycle[ 4997] = 1'b0;  wr_cycle[ 4997] = 1'b0;  addr_rom[ 4997]='h00000000;  wr_data_rom[ 4997]='h00000000;
    rd_cycle[ 4998] = 1'b0;  wr_cycle[ 4998] = 1'b0;  addr_rom[ 4998]='h00000000;  wr_data_rom[ 4998]='h00000000;
    rd_cycle[ 4999] = 1'b0;  wr_cycle[ 4999] = 1'b0;  addr_rom[ 4999]='h00000000;  wr_data_rom[ 4999]='h00000000;
    // 1000 sequence read cycles
    rd_cycle[ 5000] = 1'b1;  wr_cycle[ 5000] = 1'b0;  addr_rom[ 5000]='h00000000;  wr_data_rom[ 5000]='h00000000;
    rd_cycle[ 5001] = 1'b1;  wr_cycle[ 5001] = 1'b0;  addr_rom[ 5001]='h00000004;  wr_data_rom[ 5001]='h00000000;
    rd_cycle[ 5002] = 1'b1;  wr_cycle[ 5002] = 1'b0;  addr_rom[ 5002]='h00000008;  wr_data_rom[ 5002]='h00000000;
    rd_cycle[ 5003] = 1'b1;  wr_cycle[ 5003] = 1'b0;  addr_rom[ 5003]='h0000000c;  wr_data_rom[ 5003]='h00000000;
    rd_cycle[ 5004] = 1'b1;  wr_cycle[ 5004] = 1'b0;  addr_rom[ 5004]='h00000010;  wr_data_rom[ 5004]='h00000000;
    rd_cycle[ 5005] = 1'b1;  wr_cycle[ 5005] = 1'b0;  addr_rom[ 5005]='h00000014;  wr_data_rom[ 5005]='h00000000;
    rd_cycle[ 5006] = 1'b1;  wr_cycle[ 5006] = 1'b0;  addr_rom[ 5006]='h00000018;  wr_data_rom[ 5006]='h00000000;
    rd_cycle[ 5007] = 1'b1;  wr_cycle[ 5007] = 1'b0;  addr_rom[ 5007]='h0000001c;  wr_data_rom[ 5007]='h00000000;
    rd_cycle[ 5008] = 1'b1;  wr_cycle[ 5008] = 1'b0;  addr_rom[ 5008]='h00000020;  wr_data_rom[ 5008]='h00000000;
    rd_cycle[ 5009] = 1'b1;  wr_cycle[ 5009] = 1'b0;  addr_rom[ 5009]='h00000024;  wr_data_rom[ 5009]='h00000000;
    rd_cycle[ 5010] = 1'b1;  wr_cycle[ 5010] = 1'b0;  addr_rom[ 5010]='h00000028;  wr_data_rom[ 5010]='h00000000;
    rd_cycle[ 5011] = 1'b1;  wr_cycle[ 5011] = 1'b0;  addr_rom[ 5011]='h0000002c;  wr_data_rom[ 5011]='h00000000;
    rd_cycle[ 5012] = 1'b1;  wr_cycle[ 5012] = 1'b0;  addr_rom[ 5012]='h00000030;  wr_data_rom[ 5012]='h00000000;
    rd_cycle[ 5013] = 1'b1;  wr_cycle[ 5013] = 1'b0;  addr_rom[ 5013]='h00000034;  wr_data_rom[ 5013]='h00000000;
    rd_cycle[ 5014] = 1'b1;  wr_cycle[ 5014] = 1'b0;  addr_rom[ 5014]='h00000038;  wr_data_rom[ 5014]='h00000000;
    rd_cycle[ 5015] = 1'b1;  wr_cycle[ 5015] = 1'b0;  addr_rom[ 5015]='h0000003c;  wr_data_rom[ 5015]='h00000000;
    rd_cycle[ 5016] = 1'b1;  wr_cycle[ 5016] = 1'b0;  addr_rom[ 5016]='h00000040;  wr_data_rom[ 5016]='h00000000;
    rd_cycle[ 5017] = 1'b1;  wr_cycle[ 5017] = 1'b0;  addr_rom[ 5017]='h00000044;  wr_data_rom[ 5017]='h00000000;
    rd_cycle[ 5018] = 1'b1;  wr_cycle[ 5018] = 1'b0;  addr_rom[ 5018]='h00000048;  wr_data_rom[ 5018]='h00000000;
    rd_cycle[ 5019] = 1'b1;  wr_cycle[ 5019] = 1'b0;  addr_rom[ 5019]='h0000004c;  wr_data_rom[ 5019]='h00000000;
    rd_cycle[ 5020] = 1'b1;  wr_cycle[ 5020] = 1'b0;  addr_rom[ 5020]='h00000050;  wr_data_rom[ 5020]='h00000000;
    rd_cycle[ 5021] = 1'b1;  wr_cycle[ 5021] = 1'b0;  addr_rom[ 5021]='h00000054;  wr_data_rom[ 5021]='h00000000;
    rd_cycle[ 5022] = 1'b1;  wr_cycle[ 5022] = 1'b0;  addr_rom[ 5022]='h00000058;  wr_data_rom[ 5022]='h00000000;
    rd_cycle[ 5023] = 1'b1;  wr_cycle[ 5023] = 1'b0;  addr_rom[ 5023]='h0000005c;  wr_data_rom[ 5023]='h00000000;
    rd_cycle[ 5024] = 1'b1;  wr_cycle[ 5024] = 1'b0;  addr_rom[ 5024]='h00000060;  wr_data_rom[ 5024]='h00000000;
    rd_cycle[ 5025] = 1'b1;  wr_cycle[ 5025] = 1'b0;  addr_rom[ 5025]='h00000064;  wr_data_rom[ 5025]='h00000000;
    rd_cycle[ 5026] = 1'b1;  wr_cycle[ 5026] = 1'b0;  addr_rom[ 5026]='h00000068;  wr_data_rom[ 5026]='h00000000;
    rd_cycle[ 5027] = 1'b1;  wr_cycle[ 5027] = 1'b0;  addr_rom[ 5027]='h0000006c;  wr_data_rom[ 5027]='h00000000;
    rd_cycle[ 5028] = 1'b1;  wr_cycle[ 5028] = 1'b0;  addr_rom[ 5028]='h00000070;  wr_data_rom[ 5028]='h00000000;
    rd_cycle[ 5029] = 1'b1;  wr_cycle[ 5029] = 1'b0;  addr_rom[ 5029]='h00000074;  wr_data_rom[ 5029]='h00000000;
    rd_cycle[ 5030] = 1'b1;  wr_cycle[ 5030] = 1'b0;  addr_rom[ 5030]='h00000078;  wr_data_rom[ 5030]='h00000000;
    rd_cycle[ 5031] = 1'b1;  wr_cycle[ 5031] = 1'b0;  addr_rom[ 5031]='h0000007c;  wr_data_rom[ 5031]='h00000000;
    rd_cycle[ 5032] = 1'b1;  wr_cycle[ 5032] = 1'b0;  addr_rom[ 5032]='h00000080;  wr_data_rom[ 5032]='h00000000;
    rd_cycle[ 5033] = 1'b1;  wr_cycle[ 5033] = 1'b0;  addr_rom[ 5033]='h00000084;  wr_data_rom[ 5033]='h00000000;
    rd_cycle[ 5034] = 1'b1;  wr_cycle[ 5034] = 1'b0;  addr_rom[ 5034]='h00000088;  wr_data_rom[ 5034]='h00000000;
    rd_cycle[ 5035] = 1'b1;  wr_cycle[ 5035] = 1'b0;  addr_rom[ 5035]='h0000008c;  wr_data_rom[ 5035]='h00000000;
    rd_cycle[ 5036] = 1'b1;  wr_cycle[ 5036] = 1'b0;  addr_rom[ 5036]='h00000090;  wr_data_rom[ 5036]='h00000000;
    rd_cycle[ 5037] = 1'b1;  wr_cycle[ 5037] = 1'b0;  addr_rom[ 5037]='h00000094;  wr_data_rom[ 5037]='h00000000;
    rd_cycle[ 5038] = 1'b1;  wr_cycle[ 5038] = 1'b0;  addr_rom[ 5038]='h00000098;  wr_data_rom[ 5038]='h00000000;
    rd_cycle[ 5039] = 1'b1;  wr_cycle[ 5039] = 1'b0;  addr_rom[ 5039]='h0000009c;  wr_data_rom[ 5039]='h00000000;
    rd_cycle[ 5040] = 1'b1;  wr_cycle[ 5040] = 1'b0;  addr_rom[ 5040]='h000000a0;  wr_data_rom[ 5040]='h00000000;
    rd_cycle[ 5041] = 1'b1;  wr_cycle[ 5041] = 1'b0;  addr_rom[ 5041]='h000000a4;  wr_data_rom[ 5041]='h00000000;
    rd_cycle[ 5042] = 1'b1;  wr_cycle[ 5042] = 1'b0;  addr_rom[ 5042]='h000000a8;  wr_data_rom[ 5042]='h00000000;
    rd_cycle[ 5043] = 1'b1;  wr_cycle[ 5043] = 1'b0;  addr_rom[ 5043]='h000000ac;  wr_data_rom[ 5043]='h00000000;
    rd_cycle[ 5044] = 1'b1;  wr_cycle[ 5044] = 1'b0;  addr_rom[ 5044]='h000000b0;  wr_data_rom[ 5044]='h00000000;
    rd_cycle[ 5045] = 1'b1;  wr_cycle[ 5045] = 1'b0;  addr_rom[ 5045]='h000000b4;  wr_data_rom[ 5045]='h00000000;
    rd_cycle[ 5046] = 1'b1;  wr_cycle[ 5046] = 1'b0;  addr_rom[ 5046]='h000000b8;  wr_data_rom[ 5046]='h00000000;
    rd_cycle[ 5047] = 1'b1;  wr_cycle[ 5047] = 1'b0;  addr_rom[ 5047]='h000000bc;  wr_data_rom[ 5047]='h00000000;
    rd_cycle[ 5048] = 1'b1;  wr_cycle[ 5048] = 1'b0;  addr_rom[ 5048]='h000000c0;  wr_data_rom[ 5048]='h00000000;
    rd_cycle[ 5049] = 1'b1;  wr_cycle[ 5049] = 1'b0;  addr_rom[ 5049]='h000000c4;  wr_data_rom[ 5049]='h00000000;
    rd_cycle[ 5050] = 1'b1;  wr_cycle[ 5050] = 1'b0;  addr_rom[ 5050]='h000000c8;  wr_data_rom[ 5050]='h00000000;
    rd_cycle[ 5051] = 1'b1;  wr_cycle[ 5051] = 1'b0;  addr_rom[ 5051]='h000000cc;  wr_data_rom[ 5051]='h00000000;
    rd_cycle[ 5052] = 1'b1;  wr_cycle[ 5052] = 1'b0;  addr_rom[ 5052]='h000000d0;  wr_data_rom[ 5052]='h00000000;
    rd_cycle[ 5053] = 1'b1;  wr_cycle[ 5053] = 1'b0;  addr_rom[ 5053]='h000000d4;  wr_data_rom[ 5053]='h00000000;
    rd_cycle[ 5054] = 1'b1;  wr_cycle[ 5054] = 1'b0;  addr_rom[ 5054]='h000000d8;  wr_data_rom[ 5054]='h00000000;
    rd_cycle[ 5055] = 1'b1;  wr_cycle[ 5055] = 1'b0;  addr_rom[ 5055]='h000000dc;  wr_data_rom[ 5055]='h00000000;
    rd_cycle[ 5056] = 1'b1;  wr_cycle[ 5056] = 1'b0;  addr_rom[ 5056]='h000000e0;  wr_data_rom[ 5056]='h00000000;
    rd_cycle[ 5057] = 1'b1;  wr_cycle[ 5057] = 1'b0;  addr_rom[ 5057]='h000000e4;  wr_data_rom[ 5057]='h00000000;
    rd_cycle[ 5058] = 1'b1;  wr_cycle[ 5058] = 1'b0;  addr_rom[ 5058]='h000000e8;  wr_data_rom[ 5058]='h00000000;
    rd_cycle[ 5059] = 1'b1;  wr_cycle[ 5059] = 1'b0;  addr_rom[ 5059]='h000000ec;  wr_data_rom[ 5059]='h00000000;
    rd_cycle[ 5060] = 1'b1;  wr_cycle[ 5060] = 1'b0;  addr_rom[ 5060]='h000000f0;  wr_data_rom[ 5060]='h00000000;
    rd_cycle[ 5061] = 1'b1;  wr_cycle[ 5061] = 1'b0;  addr_rom[ 5061]='h000000f4;  wr_data_rom[ 5061]='h00000000;
    rd_cycle[ 5062] = 1'b1;  wr_cycle[ 5062] = 1'b0;  addr_rom[ 5062]='h000000f8;  wr_data_rom[ 5062]='h00000000;
    rd_cycle[ 5063] = 1'b1;  wr_cycle[ 5063] = 1'b0;  addr_rom[ 5063]='h000000fc;  wr_data_rom[ 5063]='h00000000;
    rd_cycle[ 5064] = 1'b1;  wr_cycle[ 5064] = 1'b0;  addr_rom[ 5064]='h00000100;  wr_data_rom[ 5064]='h00000000;
    rd_cycle[ 5065] = 1'b1;  wr_cycle[ 5065] = 1'b0;  addr_rom[ 5065]='h00000104;  wr_data_rom[ 5065]='h00000000;
    rd_cycle[ 5066] = 1'b1;  wr_cycle[ 5066] = 1'b0;  addr_rom[ 5066]='h00000108;  wr_data_rom[ 5066]='h00000000;
    rd_cycle[ 5067] = 1'b1;  wr_cycle[ 5067] = 1'b0;  addr_rom[ 5067]='h0000010c;  wr_data_rom[ 5067]='h00000000;
    rd_cycle[ 5068] = 1'b1;  wr_cycle[ 5068] = 1'b0;  addr_rom[ 5068]='h00000110;  wr_data_rom[ 5068]='h00000000;
    rd_cycle[ 5069] = 1'b1;  wr_cycle[ 5069] = 1'b0;  addr_rom[ 5069]='h00000114;  wr_data_rom[ 5069]='h00000000;
    rd_cycle[ 5070] = 1'b1;  wr_cycle[ 5070] = 1'b0;  addr_rom[ 5070]='h00000118;  wr_data_rom[ 5070]='h00000000;
    rd_cycle[ 5071] = 1'b1;  wr_cycle[ 5071] = 1'b0;  addr_rom[ 5071]='h0000011c;  wr_data_rom[ 5071]='h00000000;
    rd_cycle[ 5072] = 1'b1;  wr_cycle[ 5072] = 1'b0;  addr_rom[ 5072]='h00000120;  wr_data_rom[ 5072]='h00000000;
    rd_cycle[ 5073] = 1'b1;  wr_cycle[ 5073] = 1'b0;  addr_rom[ 5073]='h00000124;  wr_data_rom[ 5073]='h00000000;
    rd_cycle[ 5074] = 1'b1;  wr_cycle[ 5074] = 1'b0;  addr_rom[ 5074]='h00000128;  wr_data_rom[ 5074]='h00000000;
    rd_cycle[ 5075] = 1'b1;  wr_cycle[ 5075] = 1'b0;  addr_rom[ 5075]='h0000012c;  wr_data_rom[ 5075]='h00000000;
    rd_cycle[ 5076] = 1'b1;  wr_cycle[ 5076] = 1'b0;  addr_rom[ 5076]='h00000130;  wr_data_rom[ 5076]='h00000000;
    rd_cycle[ 5077] = 1'b1;  wr_cycle[ 5077] = 1'b0;  addr_rom[ 5077]='h00000134;  wr_data_rom[ 5077]='h00000000;
    rd_cycle[ 5078] = 1'b1;  wr_cycle[ 5078] = 1'b0;  addr_rom[ 5078]='h00000138;  wr_data_rom[ 5078]='h00000000;
    rd_cycle[ 5079] = 1'b1;  wr_cycle[ 5079] = 1'b0;  addr_rom[ 5079]='h0000013c;  wr_data_rom[ 5079]='h00000000;
    rd_cycle[ 5080] = 1'b1;  wr_cycle[ 5080] = 1'b0;  addr_rom[ 5080]='h00000140;  wr_data_rom[ 5080]='h00000000;
    rd_cycle[ 5081] = 1'b1;  wr_cycle[ 5081] = 1'b0;  addr_rom[ 5081]='h00000144;  wr_data_rom[ 5081]='h00000000;
    rd_cycle[ 5082] = 1'b1;  wr_cycle[ 5082] = 1'b0;  addr_rom[ 5082]='h00000148;  wr_data_rom[ 5082]='h00000000;
    rd_cycle[ 5083] = 1'b1;  wr_cycle[ 5083] = 1'b0;  addr_rom[ 5083]='h0000014c;  wr_data_rom[ 5083]='h00000000;
    rd_cycle[ 5084] = 1'b1;  wr_cycle[ 5084] = 1'b0;  addr_rom[ 5084]='h00000150;  wr_data_rom[ 5084]='h00000000;
    rd_cycle[ 5085] = 1'b1;  wr_cycle[ 5085] = 1'b0;  addr_rom[ 5085]='h00000154;  wr_data_rom[ 5085]='h00000000;
    rd_cycle[ 5086] = 1'b1;  wr_cycle[ 5086] = 1'b0;  addr_rom[ 5086]='h00000158;  wr_data_rom[ 5086]='h00000000;
    rd_cycle[ 5087] = 1'b1;  wr_cycle[ 5087] = 1'b0;  addr_rom[ 5087]='h0000015c;  wr_data_rom[ 5087]='h00000000;
    rd_cycle[ 5088] = 1'b1;  wr_cycle[ 5088] = 1'b0;  addr_rom[ 5088]='h00000160;  wr_data_rom[ 5088]='h00000000;
    rd_cycle[ 5089] = 1'b1;  wr_cycle[ 5089] = 1'b0;  addr_rom[ 5089]='h00000164;  wr_data_rom[ 5089]='h00000000;
    rd_cycle[ 5090] = 1'b1;  wr_cycle[ 5090] = 1'b0;  addr_rom[ 5090]='h00000168;  wr_data_rom[ 5090]='h00000000;
    rd_cycle[ 5091] = 1'b1;  wr_cycle[ 5091] = 1'b0;  addr_rom[ 5091]='h0000016c;  wr_data_rom[ 5091]='h00000000;
    rd_cycle[ 5092] = 1'b1;  wr_cycle[ 5092] = 1'b0;  addr_rom[ 5092]='h00000170;  wr_data_rom[ 5092]='h00000000;
    rd_cycle[ 5093] = 1'b1;  wr_cycle[ 5093] = 1'b0;  addr_rom[ 5093]='h00000174;  wr_data_rom[ 5093]='h00000000;
    rd_cycle[ 5094] = 1'b1;  wr_cycle[ 5094] = 1'b0;  addr_rom[ 5094]='h00000178;  wr_data_rom[ 5094]='h00000000;
    rd_cycle[ 5095] = 1'b1;  wr_cycle[ 5095] = 1'b0;  addr_rom[ 5095]='h0000017c;  wr_data_rom[ 5095]='h00000000;
    rd_cycle[ 5096] = 1'b1;  wr_cycle[ 5096] = 1'b0;  addr_rom[ 5096]='h00000180;  wr_data_rom[ 5096]='h00000000;
    rd_cycle[ 5097] = 1'b1;  wr_cycle[ 5097] = 1'b0;  addr_rom[ 5097]='h00000184;  wr_data_rom[ 5097]='h00000000;
    rd_cycle[ 5098] = 1'b1;  wr_cycle[ 5098] = 1'b0;  addr_rom[ 5098]='h00000188;  wr_data_rom[ 5098]='h00000000;
    rd_cycle[ 5099] = 1'b1;  wr_cycle[ 5099] = 1'b0;  addr_rom[ 5099]='h0000018c;  wr_data_rom[ 5099]='h00000000;
    rd_cycle[ 5100] = 1'b1;  wr_cycle[ 5100] = 1'b0;  addr_rom[ 5100]='h00000190;  wr_data_rom[ 5100]='h00000000;
    rd_cycle[ 5101] = 1'b1;  wr_cycle[ 5101] = 1'b0;  addr_rom[ 5101]='h00000194;  wr_data_rom[ 5101]='h00000000;
    rd_cycle[ 5102] = 1'b1;  wr_cycle[ 5102] = 1'b0;  addr_rom[ 5102]='h00000198;  wr_data_rom[ 5102]='h00000000;
    rd_cycle[ 5103] = 1'b1;  wr_cycle[ 5103] = 1'b0;  addr_rom[ 5103]='h0000019c;  wr_data_rom[ 5103]='h00000000;
    rd_cycle[ 5104] = 1'b1;  wr_cycle[ 5104] = 1'b0;  addr_rom[ 5104]='h000001a0;  wr_data_rom[ 5104]='h00000000;
    rd_cycle[ 5105] = 1'b1;  wr_cycle[ 5105] = 1'b0;  addr_rom[ 5105]='h000001a4;  wr_data_rom[ 5105]='h00000000;
    rd_cycle[ 5106] = 1'b1;  wr_cycle[ 5106] = 1'b0;  addr_rom[ 5106]='h000001a8;  wr_data_rom[ 5106]='h00000000;
    rd_cycle[ 5107] = 1'b1;  wr_cycle[ 5107] = 1'b0;  addr_rom[ 5107]='h000001ac;  wr_data_rom[ 5107]='h00000000;
    rd_cycle[ 5108] = 1'b1;  wr_cycle[ 5108] = 1'b0;  addr_rom[ 5108]='h000001b0;  wr_data_rom[ 5108]='h00000000;
    rd_cycle[ 5109] = 1'b1;  wr_cycle[ 5109] = 1'b0;  addr_rom[ 5109]='h000001b4;  wr_data_rom[ 5109]='h00000000;
    rd_cycle[ 5110] = 1'b1;  wr_cycle[ 5110] = 1'b0;  addr_rom[ 5110]='h000001b8;  wr_data_rom[ 5110]='h00000000;
    rd_cycle[ 5111] = 1'b1;  wr_cycle[ 5111] = 1'b0;  addr_rom[ 5111]='h000001bc;  wr_data_rom[ 5111]='h00000000;
    rd_cycle[ 5112] = 1'b1;  wr_cycle[ 5112] = 1'b0;  addr_rom[ 5112]='h000001c0;  wr_data_rom[ 5112]='h00000000;
    rd_cycle[ 5113] = 1'b1;  wr_cycle[ 5113] = 1'b0;  addr_rom[ 5113]='h000001c4;  wr_data_rom[ 5113]='h00000000;
    rd_cycle[ 5114] = 1'b1;  wr_cycle[ 5114] = 1'b0;  addr_rom[ 5114]='h000001c8;  wr_data_rom[ 5114]='h00000000;
    rd_cycle[ 5115] = 1'b1;  wr_cycle[ 5115] = 1'b0;  addr_rom[ 5115]='h000001cc;  wr_data_rom[ 5115]='h00000000;
    rd_cycle[ 5116] = 1'b1;  wr_cycle[ 5116] = 1'b0;  addr_rom[ 5116]='h000001d0;  wr_data_rom[ 5116]='h00000000;
    rd_cycle[ 5117] = 1'b1;  wr_cycle[ 5117] = 1'b0;  addr_rom[ 5117]='h000001d4;  wr_data_rom[ 5117]='h00000000;
    rd_cycle[ 5118] = 1'b1;  wr_cycle[ 5118] = 1'b0;  addr_rom[ 5118]='h000001d8;  wr_data_rom[ 5118]='h00000000;
    rd_cycle[ 5119] = 1'b1;  wr_cycle[ 5119] = 1'b0;  addr_rom[ 5119]='h000001dc;  wr_data_rom[ 5119]='h00000000;
    rd_cycle[ 5120] = 1'b1;  wr_cycle[ 5120] = 1'b0;  addr_rom[ 5120]='h000001e0;  wr_data_rom[ 5120]='h00000000;
    rd_cycle[ 5121] = 1'b1;  wr_cycle[ 5121] = 1'b0;  addr_rom[ 5121]='h000001e4;  wr_data_rom[ 5121]='h00000000;
    rd_cycle[ 5122] = 1'b1;  wr_cycle[ 5122] = 1'b0;  addr_rom[ 5122]='h000001e8;  wr_data_rom[ 5122]='h00000000;
    rd_cycle[ 5123] = 1'b1;  wr_cycle[ 5123] = 1'b0;  addr_rom[ 5123]='h000001ec;  wr_data_rom[ 5123]='h00000000;
    rd_cycle[ 5124] = 1'b1;  wr_cycle[ 5124] = 1'b0;  addr_rom[ 5124]='h000001f0;  wr_data_rom[ 5124]='h00000000;
    rd_cycle[ 5125] = 1'b1;  wr_cycle[ 5125] = 1'b0;  addr_rom[ 5125]='h000001f4;  wr_data_rom[ 5125]='h00000000;
    rd_cycle[ 5126] = 1'b1;  wr_cycle[ 5126] = 1'b0;  addr_rom[ 5126]='h000001f8;  wr_data_rom[ 5126]='h00000000;
    rd_cycle[ 5127] = 1'b1;  wr_cycle[ 5127] = 1'b0;  addr_rom[ 5127]='h000001fc;  wr_data_rom[ 5127]='h00000000;
    rd_cycle[ 5128] = 1'b1;  wr_cycle[ 5128] = 1'b0;  addr_rom[ 5128]='h00000200;  wr_data_rom[ 5128]='h00000000;
    rd_cycle[ 5129] = 1'b1;  wr_cycle[ 5129] = 1'b0;  addr_rom[ 5129]='h00000204;  wr_data_rom[ 5129]='h00000000;
    rd_cycle[ 5130] = 1'b1;  wr_cycle[ 5130] = 1'b0;  addr_rom[ 5130]='h00000208;  wr_data_rom[ 5130]='h00000000;
    rd_cycle[ 5131] = 1'b1;  wr_cycle[ 5131] = 1'b0;  addr_rom[ 5131]='h0000020c;  wr_data_rom[ 5131]='h00000000;
    rd_cycle[ 5132] = 1'b1;  wr_cycle[ 5132] = 1'b0;  addr_rom[ 5132]='h00000210;  wr_data_rom[ 5132]='h00000000;
    rd_cycle[ 5133] = 1'b1;  wr_cycle[ 5133] = 1'b0;  addr_rom[ 5133]='h00000214;  wr_data_rom[ 5133]='h00000000;
    rd_cycle[ 5134] = 1'b1;  wr_cycle[ 5134] = 1'b0;  addr_rom[ 5134]='h00000218;  wr_data_rom[ 5134]='h00000000;
    rd_cycle[ 5135] = 1'b1;  wr_cycle[ 5135] = 1'b0;  addr_rom[ 5135]='h0000021c;  wr_data_rom[ 5135]='h00000000;
    rd_cycle[ 5136] = 1'b1;  wr_cycle[ 5136] = 1'b0;  addr_rom[ 5136]='h00000220;  wr_data_rom[ 5136]='h00000000;
    rd_cycle[ 5137] = 1'b1;  wr_cycle[ 5137] = 1'b0;  addr_rom[ 5137]='h00000224;  wr_data_rom[ 5137]='h00000000;
    rd_cycle[ 5138] = 1'b1;  wr_cycle[ 5138] = 1'b0;  addr_rom[ 5138]='h00000228;  wr_data_rom[ 5138]='h00000000;
    rd_cycle[ 5139] = 1'b1;  wr_cycle[ 5139] = 1'b0;  addr_rom[ 5139]='h0000022c;  wr_data_rom[ 5139]='h00000000;
    rd_cycle[ 5140] = 1'b1;  wr_cycle[ 5140] = 1'b0;  addr_rom[ 5140]='h00000230;  wr_data_rom[ 5140]='h00000000;
    rd_cycle[ 5141] = 1'b1;  wr_cycle[ 5141] = 1'b0;  addr_rom[ 5141]='h00000234;  wr_data_rom[ 5141]='h00000000;
    rd_cycle[ 5142] = 1'b1;  wr_cycle[ 5142] = 1'b0;  addr_rom[ 5142]='h00000238;  wr_data_rom[ 5142]='h00000000;
    rd_cycle[ 5143] = 1'b1;  wr_cycle[ 5143] = 1'b0;  addr_rom[ 5143]='h0000023c;  wr_data_rom[ 5143]='h00000000;
    rd_cycle[ 5144] = 1'b1;  wr_cycle[ 5144] = 1'b0;  addr_rom[ 5144]='h00000240;  wr_data_rom[ 5144]='h00000000;
    rd_cycle[ 5145] = 1'b1;  wr_cycle[ 5145] = 1'b0;  addr_rom[ 5145]='h00000244;  wr_data_rom[ 5145]='h00000000;
    rd_cycle[ 5146] = 1'b1;  wr_cycle[ 5146] = 1'b0;  addr_rom[ 5146]='h00000248;  wr_data_rom[ 5146]='h00000000;
    rd_cycle[ 5147] = 1'b1;  wr_cycle[ 5147] = 1'b0;  addr_rom[ 5147]='h0000024c;  wr_data_rom[ 5147]='h00000000;
    rd_cycle[ 5148] = 1'b1;  wr_cycle[ 5148] = 1'b0;  addr_rom[ 5148]='h00000250;  wr_data_rom[ 5148]='h00000000;
    rd_cycle[ 5149] = 1'b1;  wr_cycle[ 5149] = 1'b0;  addr_rom[ 5149]='h00000254;  wr_data_rom[ 5149]='h00000000;
    rd_cycle[ 5150] = 1'b1;  wr_cycle[ 5150] = 1'b0;  addr_rom[ 5150]='h00000258;  wr_data_rom[ 5150]='h00000000;
    rd_cycle[ 5151] = 1'b1;  wr_cycle[ 5151] = 1'b0;  addr_rom[ 5151]='h0000025c;  wr_data_rom[ 5151]='h00000000;
    rd_cycle[ 5152] = 1'b1;  wr_cycle[ 5152] = 1'b0;  addr_rom[ 5152]='h00000260;  wr_data_rom[ 5152]='h00000000;
    rd_cycle[ 5153] = 1'b1;  wr_cycle[ 5153] = 1'b0;  addr_rom[ 5153]='h00000264;  wr_data_rom[ 5153]='h00000000;
    rd_cycle[ 5154] = 1'b1;  wr_cycle[ 5154] = 1'b0;  addr_rom[ 5154]='h00000268;  wr_data_rom[ 5154]='h00000000;
    rd_cycle[ 5155] = 1'b1;  wr_cycle[ 5155] = 1'b0;  addr_rom[ 5155]='h0000026c;  wr_data_rom[ 5155]='h00000000;
    rd_cycle[ 5156] = 1'b1;  wr_cycle[ 5156] = 1'b0;  addr_rom[ 5156]='h00000270;  wr_data_rom[ 5156]='h00000000;
    rd_cycle[ 5157] = 1'b1;  wr_cycle[ 5157] = 1'b0;  addr_rom[ 5157]='h00000274;  wr_data_rom[ 5157]='h00000000;
    rd_cycle[ 5158] = 1'b1;  wr_cycle[ 5158] = 1'b0;  addr_rom[ 5158]='h00000278;  wr_data_rom[ 5158]='h00000000;
    rd_cycle[ 5159] = 1'b1;  wr_cycle[ 5159] = 1'b0;  addr_rom[ 5159]='h0000027c;  wr_data_rom[ 5159]='h00000000;
    rd_cycle[ 5160] = 1'b1;  wr_cycle[ 5160] = 1'b0;  addr_rom[ 5160]='h00000280;  wr_data_rom[ 5160]='h00000000;
    rd_cycle[ 5161] = 1'b1;  wr_cycle[ 5161] = 1'b0;  addr_rom[ 5161]='h00000284;  wr_data_rom[ 5161]='h00000000;
    rd_cycle[ 5162] = 1'b1;  wr_cycle[ 5162] = 1'b0;  addr_rom[ 5162]='h00000288;  wr_data_rom[ 5162]='h00000000;
    rd_cycle[ 5163] = 1'b1;  wr_cycle[ 5163] = 1'b0;  addr_rom[ 5163]='h0000028c;  wr_data_rom[ 5163]='h00000000;
    rd_cycle[ 5164] = 1'b1;  wr_cycle[ 5164] = 1'b0;  addr_rom[ 5164]='h00000290;  wr_data_rom[ 5164]='h00000000;
    rd_cycle[ 5165] = 1'b1;  wr_cycle[ 5165] = 1'b0;  addr_rom[ 5165]='h00000294;  wr_data_rom[ 5165]='h00000000;
    rd_cycle[ 5166] = 1'b1;  wr_cycle[ 5166] = 1'b0;  addr_rom[ 5166]='h00000298;  wr_data_rom[ 5166]='h00000000;
    rd_cycle[ 5167] = 1'b1;  wr_cycle[ 5167] = 1'b0;  addr_rom[ 5167]='h0000029c;  wr_data_rom[ 5167]='h00000000;
    rd_cycle[ 5168] = 1'b1;  wr_cycle[ 5168] = 1'b0;  addr_rom[ 5168]='h000002a0;  wr_data_rom[ 5168]='h00000000;
    rd_cycle[ 5169] = 1'b1;  wr_cycle[ 5169] = 1'b0;  addr_rom[ 5169]='h000002a4;  wr_data_rom[ 5169]='h00000000;
    rd_cycle[ 5170] = 1'b1;  wr_cycle[ 5170] = 1'b0;  addr_rom[ 5170]='h000002a8;  wr_data_rom[ 5170]='h00000000;
    rd_cycle[ 5171] = 1'b1;  wr_cycle[ 5171] = 1'b0;  addr_rom[ 5171]='h000002ac;  wr_data_rom[ 5171]='h00000000;
    rd_cycle[ 5172] = 1'b1;  wr_cycle[ 5172] = 1'b0;  addr_rom[ 5172]='h000002b0;  wr_data_rom[ 5172]='h00000000;
    rd_cycle[ 5173] = 1'b1;  wr_cycle[ 5173] = 1'b0;  addr_rom[ 5173]='h000002b4;  wr_data_rom[ 5173]='h00000000;
    rd_cycle[ 5174] = 1'b1;  wr_cycle[ 5174] = 1'b0;  addr_rom[ 5174]='h000002b8;  wr_data_rom[ 5174]='h00000000;
    rd_cycle[ 5175] = 1'b1;  wr_cycle[ 5175] = 1'b0;  addr_rom[ 5175]='h000002bc;  wr_data_rom[ 5175]='h00000000;
    rd_cycle[ 5176] = 1'b1;  wr_cycle[ 5176] = 1'b0;  addr_rom[ 5176]='h000002c0;  wr_data_rom[ 5176]='h00000000;
    rd_cycle[ 5177] = 1'b1;  wr_cycle[ 5177] = 1'b0;  addr_rom[ 5177]='h000002c4;  wr_data_rom[ 5177]='h00000000;
    rd_cycle[ 5178] = 1'b1;  wr_cycle[ 5178] = 1'b0;  addr_rom[ 5178]='h000002c8;  wr_data_rom[ 5178]='h00000000;
    rd_cycle[ 5179] = 1'b1;  wr_cycle[ 5179] = 1'b0;  addr_rom[ 5179]='h000002cc;  wr_data_rom[ 5179]='h00000000;
    rd_cycle[ 5180] = 1'b1;  wr_cycle[ 5180] = 1'b0;  addr_rom[ 5180]='h000002d0;  wr_data_rom[ 5180]='h00000000;
    rd_cycle[ 5181] = 1'b1;  wr_cycle[ 5181] = 1'b0;  addr_rom[ 5181]='h000002d4;  wr_data_rom[ 5181]='h00000000;
    rd_cycle[ 5182] = 1'b1;  wr_cycle[ 5182] = 1'b0;  addr_rom[ 5182]='h000002d8;  wr_data_rom[ 5182]='h00000000;
    rd_cycle[ 5183] = 1'b1;  wr_cycle[ 5183] = 1'b0;  addr_rom[ 5183]='h000002dc;  wr_data_rom[ 5183]='h00000000;
    rd_cycle[ 5184] = 1'b1;  wr_cycle[ 5184] = 1'b0;  addr_rom[ 5184]='h000002e0;  wr_data_rom[ 5184]='h00000000;
    rd_cycle[ 5185] = 1'b1;  wr_cycle[ 5185] = 1'b0;  addr_rom[ 5185]='h000002e4;  wr_data_rom[ 5185]='h00000000;
    rd_cycle[ 5186] = 1'b1;  wr_cycle[ 5186] = 1'b0;  addr_rom[ 5186]='h000002e8;  wr_data_rom[ 5186]='h00000000;
    rd_cycle[ 5187] = 1'b1;  wr_cycle[ 5187] = 1'b0;  addr_rom[ 5187]='h000002ec;  wr_data_rom[ 5187]='h00000000;
    rd_cycle[ 5188] = 1'b1;  wr_cycle[ 5188] = 1'b0;  addr_rom[ 5188]='h000002f0;  wr_data_rom[ 5188]='h00000000;
    rd_cycle[ 5189] = 1'b1;  wr_cycle[ 5189] = 1'b0;  addr_rom[ 5189]='h000002f4;  wr_data_rom[ 5189]='h00000000;
    rd_cycle[ 5190] = 1'b1;  wr_cycle[ 5190] = 1'b0;  addr_rom[ 5190]='h000002f8;  wr_data_rom[ 5190]='h00000000;
    rd_cycle[ 5191] = 1'b1;  wr_cycle[ 5191] = 1'b0;  addr_rom[ 5191]='h000002fc;  wr_data_rom[ 5191]='h00000000;
    rd_cycle[ 5192] = 1'b1;  wr_cycle[ 5192] = 1'b0;  addr_rom[ 5192]='h00000300;  wr_data_rom[ 5192]='h00000000;
    rd_cycle[ 5193] = 1'b1;  wr_cycle[ 5193] = 1'b0;  addr_rom[ 5193]='h00000304;  wr_data_rom[ 5193]='h00000000;
    rd_cycle[ 5194] = 1'b1;  wr_cycle[ 5194] = 1'b0;  addr_rom[ 5194]='h00000308;  wr_data_rom[ 5194]='h00000000;
    rd_cycle[ 5195] = 1'b1;  wr_cycle[ 5195] = 1'b0;  addr_rom[ 5195]='h0000030c;  wr_data_rom[ 5195]='h00000000;
    rd_cycle[ 5196] = 1'b1;  wr_cycle[ 5196] = 1'b0;  addr_rom[ 5196]='h00000310;  wr_data_rom[ 5196]='h00000000;
    rd_cycle[ 5197] = 1'b1;  wr_cycle[ 5197] = 1'b0;  addr_rom[ 5197]='h00000314;  wr_data_rom[ 5197]='h00000000;
    rd_cycle[ 5198] = 1'b1;  wr_cycle[ 5198] = 1'b0;  addr_rom[ 5198]='h00000318;  wr_data_rom[ 5198]='h00000000;
    rd_cycle[ 5199] = 1'b1;  wr_cycle[ 5199] = 1'b0;  addr_rom[ 5199]='h0000031c;  wr_data_rom[ 5199]='h00000000;
    rd_cycle[ 5200] = 1'b1;  wr_cycle[ 5200] = 1'b0;  addr_rom[ 5200]='h00000320;  wr_data_rom[ 5200]='h00000000;
    rd_cycle[ 5201] = 1'b1;  wr_cycle[ 5201] = 1'b0;  addr_rom[ 5201]='h00000324;  wr_data_rom[ 5201]='h00000000;
    rd_cycle[ 5202] = 1'b1;  wr_cycle[ 5202] = 1'b0;  addr_rom[ 5202]='h00000328;  wr_data_rom[ 5202]='h00000000;
    rd_cycle[ 5203] = 1'b1;  wr_cycle[ 5203] = 1'b0;  addr_rom[ 5203]='h0000032c;  wr_data_rom[ 5203]='h00000000;
    rd_cycle[ 5204] = 1'b1;  wr_cycle[ 5204] = 1'b0;  addr_rom[ 5204]='h00000330;  wr_data_rom[ 5204]='h00000000;
    rd_cycle[ 5205] = 1'b1;  wr_cycle[ 5205] = 1'b0;  addr_rom[ 5205]='h00000334;  wr_data_rom[ 5205]='h00000000;
    rd_cycle[ 5206] = 1'b1;  wr_cycle[ 5206] = 1'b0;  addr_rom[ 5206]='h00000338;  wr_data_rom[ 5206]='h00000000;
    rd_cycle[ 5207] = 1'b1;  wr_cycle[ 5207] = 1'b0;  addr_rom[ 5207]='h0000033c;  wr_data_rom[ 5207]='h00000000;
    rd_cycle[ 5208] = 1'b1;  wr_cycle[ 5208] = 1'b0;  addr_rom[ 5208]='h00000340;  wr_data_rom[ 5208]='h00000000;
    rd_cycle[ 5209] = 1'b1;  wr_cycle[ 5209] = 1'b0;  addr_rom[ 5209]='h00000344;  wr_data_rom[ 5209]='h00000000;
    rd_cycle[ 5210] = 1'b1;  wr_cycle[ 5210] = 1'b0;  addr_rom[ 5210]='h00000348;  wr_data_rom[ 5210]='h00000000;
    rd_cycle[ 5211] = 1'b1;  wr_cycle[ 5211] = 1'b0;  addr_rom[ 5211]='h0000034c;  wr_data_rom[ 5211]='h00000000;
    rd_cycle[ 5212] = 1'b1;  wr_cycle[ 5212] = 1'b0;  addr_rom[ 5212]='h00000350;  wr_data_rom[ 5212]='h00000000;
    rd_cycle[ 5213] = 1'b1;  wr_cycle[ 5213] = 1'b0;  addr_rom[ 5213]='h00000354;  wr_data_rom[ 5213]='h00000000;
    rd_cycle[ 5214] = 1'b1;  wr_cycle[ 5214] = 1'b0;  addr_rom[ 5214]='h00000358;  wr_data_rom[ 5214]='h00000000;
    rd_cycle[ 5215] = 1'b1;  wr_cycle[ 5215] = 1'b0;  addr_rom[ 5215]='h0000035c;  wr_data_rom[ 5215]='h00000000;
    rd_cycle[ 5216] = 1'b1;  wr_cycle[ 5216] = 1'b0;  addr_rom[ 5216]='h00000360;  wr_data_rom[ 5216]='h00000000;
    rd_cycle[ 5217] = 1'b1;  wr_cycle[ 5217] = 1'b0;  addr_rom[ 5217]='h00000364;  wr_data_rom[ 5217]='h00000000;
    rd_cycle[ 5218] = 1'b1;  wr_cycle[ 5218] = 1'b0;  addr_rom[ 5218]='h00000368;  wr_data_rom[ 5218]='h00000000;
    rd_cycle[ 5219] = 1'b1;  wr_cycle[ 5219] = 1'b0;  addr_rom[ 5219]='h0000036c;  wr_data_rom[ 5219]='h00000000;
    rd_cycle[ 5220] = 1'b1;  wr_cycle[ 5220] = 1'b0;  addr_rom[ 5220]='h00000370;  wr_data_rom[ 5220]='h00000000;
    rd_cycle[ 5221] = 1'b1;  wr_cycle[ 5221] = 1'b0;  addr_rom[ 5221]='h00000374;  wr_data_rom[ 5221]='h00000000;
    rd_cycle[ 5222] = 1'b1;  wr_cycle[ 5222] = 1'b0;  addr_rom[ 5222]='h00000378;  wr_data_rom[ 5222]='h00000000;
    rd_cycle[ 5223] = 1'b1;  wr_cycle[ 5223] = 1'b0;  addr_rom[ 5223]='h0000037c;  wr_data_rom[ 5223]='h00000000;
    rd_cycle[ 5224] = 1'b1;  wr_cycle[ 5224] = 1'b0;  addr_rom[ 5224]='h00000380;  wr_data_rom[ 5224]='h00000000;
    rd_cycle[ 5225] = 1'b1;  wr_cycle[ 5225] = 1'b0;  addr_rom[ 5225]='h00000384;  wr_data_rom[ 5225]='h00000000;
    rd_cycle[ 5226] = 1'b1;  wr_cycle[ 5226] = 1'b0;  addr_rom[ 5226]='h00000388;  wr_data_rom[ 5226]='h00000000;
    rd_cycle[ 5227] = 1'b1;  wr_cycle[ 5227] = 1'b0;  addr_rom[ 5227]='h0000038c;  wr_data_rom[ 5227]='h00000000;
    rd_cycle[ 5228] = 1'b1;  wr_cycle[ 5228] = 1'b0;  addr_rom[ 5228]='h00000390;  wr_data_rom[ 5228]='h00000000;
    rd_cycle[ 5229] = 1'b1;  wr_cycle[ 5229] = 1'b0;  addr_rom[ 5229]='h00000394;  wr_data_rom[ 5229]='h00000000;
    rd_cycle[ 5230] = 1'b1;  wr_cycle[ 5230] = 1'b0;  addr_rom[ 5230]='h00000398;  wr_data_rom[ 5230]='h00000000;
    rd_cycle[ 5231] = 1'b1;  wr_cycle[ 5231] = 1'b0;  addr_rom[ 5231]='h0000039c;  wr_data_rom[ 5231]='h00000000;
    rd_cycle[ 5232] = 1'b1;  wr_cycle[ 5232] = 1'b0;  addr_rom[ 5232]='h000003a0;  wr_data_rom[ 5232]='h00000000;
    rd_cycle[ 5233] = 1'b1;  wr_cycle[ 5233] = 1'b0;  addr_rom[ 5233]='h000003a4;  wr_data_rom[ 5233]='h00000000;
    rd_cycle[ 5234] = 1'b1;  wr_cycle[ 5234] = 1'b0;  addr_rom[ 5234]='h000003a8;  wr_data_rom[ 5234]='h00000000;
    rd_cycle[ 5235] = 1'b1;  wr_cycle[ 5235] = 1'b0;  addr_rom[ 5235]='h000003ac;  wr_data_rom[ 5235]='h00000000;
    rd_cycle[ 5236] = 1'b1;  wr_cycle[ 5236] = 1'b0;  addr_rom[ 5236]='h000003b0;  wr_data_rom[ 5236]='h00000000;
    rd_cycle[ 5237] = 1'b1;  wr_cycle[ 5237] = 1'b0;  addr_rom[ 5237]='h000003b4;  wr_data_rom[ 5237]='h00000000;
    rd_cycle[ 5238] = 1'b1;  wr_cycle[ 5238] = 1'b0;  addr_rom[ 5238]='h000003b8;  wr_data_rom[ 5238]='h00000000;
    rd_cycle[ 5239] = 1'b1;  wr_cycle[ 5239] = 1'b0;  addr_rom[ 5239]='h000003bc;  wr_data_rom[ 5239]='h00000000;
    rd_cycle[ 5240] = 1'b1;  wr_cycle[ 5240] = 1'b0;  addr_rom[ 5240]='h000003c0;  wr_data_rom[ 5240]='h00000000;
    rd_cycle[ 5241] = 1'b1;  wr_cycle[ 5241] = 1'b0;  addr_rom[ 5241]='h000003c4;  wr_data_rom[ 5241]='h00000000;
    rd_cycle[ 5242] = 1'b1;  wr_cycle[ 5242] = 1'b0;  addr_rom[ 5242]='h000003c8;  wr_data_rom[ 5242]='h00000000;
    rd_cycle[ 5243] = 1'b1;  wr_cycle[ 5243] = 1'b0;  addr_rom[ 5243]='h000003cc;  wr_data_rom[ 5243]='h00000000;
    rd_cycle[ 5244] = 1'b1;  wr_cycle[ 5244] = 1'b0;  addr_rom[ 5244]='h000003d0;  wr_data_rom[ 5244]='h00000000;
    rd_cycle[ 5245] = 1'b1;  wr_cycle[ 5245] = 1'b0;  addr_rom[ 5245]='h000003d4;  wr_data_rom[ 5245]='h00000000;
    rd_cycle[ 5246] = 1'b1;  wr_cycle[ 5246] = 1'b0;  addr_rom[ 5246]='h000003d8;  wr_data_rom[ 5246]='h00000000;
    rd_cycle[ 5247] = 1'b1;  wr_cycle[ 5247] = 1'b0;  addr_rom[ 5247]='h000003dc;  wr_data_rom[ 5247]='h00000000;
    rd_cycle[ 5248] = 1'b1;  wr_cycle[ 5248] = 1'b0;  addr_rom[ 5248]='h000003e0;  wr_data_rom[ 5248]='h00000000;
    rd_cycle[ 5249] = 1'b1;  wr_cycle[ 5249] = 1'b0;  addr_rom[ 5249]='h000003e4;  wr_data_rom[ 5249]='h00000000;
    rd_cycle[ 5250] = 1'b1;  wr_cycle[ 5250] = 1'b0;  addr_rom[ 5250]='h000003e8;  wr_data_rom[ 5250]='h00000000;
    rd_cycle[ 5251] = 1'b1;  wr_cycle[ 5251] = 1'b0;  addr_rom[ 5251]='h000003ec;  wr_data_rom[ 5251]='h00000000;
    rd_cycle[ 5252] = 1'b1;  wr_cycle[ 5252] = 1'b0;  addr_rom[ 5252]='h000003f0;  wr_data_rom[ 5252]='h00000000;
    rd_cycle[ 5253] = 1'b1;  wr_cycle[ 5253] = 1'b0;  addr_rom[ 5253]='h000003f4;  wr_data_rom[ 5253]='h00000000;
    rd_cycle[ 5254] = 1'b1;  wr_cycle[ 5254] = 1'b0;  addr_rom[ 5254]='h000003f8;  wr_data_rom[ 5254]='h00000000;
    rd_cycle[ 5255] = 1'b1;  wr_cycle[ 5255] = 1'b0;  addr_rom[ 5255]='h000003fc;  wr_data_rom[ 5255]='h00000000;
    rd_cycle[ 5256] = 1'b1;  wr_cycle[ 5256] = 1'b0;  addr_rom[ 5256]='h00000400;  wr_data_rom[ 5256]='h00000000;
    rd_cycle[ 5257] = 1'b1;  wr_cycle[ 5257] = 1'b0;  addr_rom[ 5257]='h00000404;  wr_data_rom[ 5257]='h00000000;
    rd_cycle[ 5258] = 1'b1;  wr_cycle[ 5258] = 1'b0;  addr_rom[ 5258]='h00000408;  wr_data_rom[ 5258]='h00000000;
    rd_cycle[ 5259] = 1'b1;  wr_cycle[ 5259] = 1'b0;  addr_rom[ 5259]='h0000040c;  wr_data_rom[ 5259]='h00000000;
    rd_cycle[ 5260] = 1'b1;  wr_cycle[ 5260] = 1'b0;  addr_rom[ 5260]='h00000410;  wr_data_rom[ 5260]='h00000000;
    rd_cycle[ 5261] = 1'b1;  wr_cycle[ 5261] = 1'b0;  addr_rom[ 5261]='h00000414;  wr_data_rom[ 5261]='h00000000;
    rd_cycle[ 5262] = 1'b1;  wr_cycle[ 5262] = 1'b0;  addr_rom[ 5262]='h00000418;  wr_data_rom[ 5262]='h00000000;
    rd_cycle[ 5263] = 1'b1;  wr_cycle[ 5263] = 1'b0;  addr_rom[ 5263]='h0000041c;  wr_data_rom[ 5263]='h00000000;
    rd_cycle[ 5264] = 1'b1;  wr_cycle[ 5264] = 1'b0;  addr_rom[ 5264]='h00000420;  wr_data_rom[ 5264]='h00000000;
    rd_cycle[ 5265] = 1'b1;  wr_cycle[ 5265] = 1'b0;  addr_rom[ 5265]='h00000424;  wr_data_rom[ 5265]='h00000000;
    rd_cycle[ 5266] = 1'b1;  wr_cycle[ 5266] = 1'b0;  addr_rom[ 5266]='h00000428;  wr_data_rom[ 5266]='h00000000;
    rd_cycle[ 5267] = 1'b1;  wr_cycle[ 5267] = 1'b0;  addr_rom[ 5267]='h0000042c;  wr_data_rom[ 5267]='h00000000;
    rd_cycle[ 5268] = 1'b1;  wr_cycle[ 5268] = 1'b0;  addr_rom[ 5268]='h00000430;  wr_data_rom[ 5268]='h00000000;
    rd_cycle[ 5269] = 1'b1;  wr_cycle[ 5269] = 1'b0;  addr_rom[ 5269]='h00000434;  wr_data_rom[ 5269]='h00000000;
    rd_cycle[ 5270] = 1'b1;  wr_cycle[ 5270] = 1'b0;  addr_rom[ 5270]='h00000438;  wr_data_rom[ 5270]='h00000000;
    rd_cycle[ 5271] = 1'b1;  wr_cycle[ 5271] = 1'b0;  addr_rom[ 5271]='h0000043c;  wr_data_rom[ 5271]='h00000000;
    rd_cycle[ 5272] = 1'b1;  wr_cycle[ 5272] = 1'b0;  addr_rom[ 5272]='h00000440;  wr_data_rom[ 5272]='h00000000;
    rd_cycle[ 5273] = 1'b1;  wr_cycle[ 5273] = 1'b0;  addr_rom[ 5273]='h00000444;  wr_data_rom[ 5273]='h00000000;
    rd_cycle[ 5274] = 1'b1;  wr_cycle[ 5274] = 1'b0;  addr_rom[ 5274]='h00000448;  wr_data_rom[ 5274]='h00000000;
    rd_cycle[ 5275] = 1'b1;  wr_cycle[ 5275] = 1'b0;  addr_rom[ 5275]='h0000044c;  wr_data_rom[ 5275]='h00000000;
    rd_cycle[ 5276] = 1'b1;  wr_cycle[ 5276] = 1'b0;  addr_rom[ 5276]='h00000450;  wr_data_rom[ 5276]='h00000000;
    rd_cycle[ 5277] = 1'b1;  wr_cycle[ 5277] = 1'b0;  addr_rom[ 5277]='h00000454;  wr_data_rom[ 5277]='h00000000;
    rd_cycle[ 5278] = 1'b1;  wr_cycle[ 5278] = 1'b0;  addr_rom[ 5278]='h00000458;  wr_data_rom[ 5278]='h00000000;
    rd_cycle[ 5279] = 1'b1;  wr_cycle[ 5279] = 1'b0;  addr_rom[ 5279]='h0000045c;  wr_data_rom[ 5279]='h00000000;
    rd_cycle[ 5280] = 1'b1;  wr_cycle[ 5280] = 1'b0;  addr_rom[ 5280]='h00000460;  wr_data_rom[ 5280]='h00000000;
    rd_cycle[ 5281] = 1'b1;  wr_cycle[ 5281] = 1'b0;  addr_rom[ 5281]='h00000464;  wr_data_rom[ 5281]='h00000000;
    rd_cycle[ 5282] = 1'b1;  wr_cycle[ 5282] = 1'b0;  addr_rom[ 5282]='h00000468;  wr_data_rom[ 5282]='h00000000;
    rd_cycle[ 5283] = 1'b1;  wr_cycle[ 5283] = 1'b0;  addr_rom[ 5283]='h0000046c;  wr_data_rom[ 5283]='h00000000;
    rd_cycle[ 5284] = 1'b1;  wr_cycle[ 5284] = 1'b0;  addr_rom[ 5284]='h00000470;  wr_data_rom[ 5284]='h00000000;
    rd_cycle[ 5285] = 1'b1;  wr_cycle[ 5285] = 1'b0;  addr_rom[ 5285]='h00000474;  wr_data_rom[ 5285]='h00000000;
    rd_cycle[ 5286] = 1'b1;  wr_cycle[ 5286] = 1'b0;  addr_rom[ 5286]='h00000478;  wr_data_rom[ 5286]='h00000000;
    rd_cycle[ 5287] = 1'b1;  wr_cycle[ 5287] = 1'b0;  addr_rom[ 5287]='h0000047c;  wr_data_rom[ 5287]='h00000000;
    rd_cycle[ 5288] = 1'b1;  wr_cycle[ 5288] = 1'b0;  addr_rom[ 5288]='h00000480;  wr_data_rom[ 5288]='h00000000;
    rd_cycle[ 5289] = 1'b1;  wr_cycle[ 5289] = 1'b0;  addr_rom[ 5289]='h00000484;  wr_data_rom[ 5289]='h00000000;
    rd_cycle[ 5290] = 1'b1;  wr_cycle[ 5290] = 1'b0;  addr_rom[ 5290]='h00000488;  wr_data_rom[ 5290]='h00000000;
    rd_cycle[ 5291] = 1'b1;  wr_cycle[ 5291] = 1'b0;  addr_rom[ 5291]='h0000048c;  wr_data_rom[ 5291]='h00000000;
    rd_cycle[ 5292] = 1'b1;  wr_cycle[ 5292] = 1'b0;  addr_rom[ 5292]='h00000490;  wr_data_rom[ 5292]='h00000000;
    rd_cycle[ 5293] = 1'b1;  wr_cycle[ 5293] = 1'b0;  addr_rom[ 5293]='h00000494;  wr_data_rom[ 5293]='h00000000;
    rd_cycle[ 5294] = 1'b1;  wr_cycle[ 5294] = 1'b0;  addr_rom[ 5294]='h00000498;  wr_data_rom[ 5294]='h00000000;
    rd_cycle[ 5295] = 1'b1;  wr_cycle[ 5295] = 1'b0;  addr_rom[ 5295]='h0000049c;  wr_data_rom[ 5295]='h00000000;
    rd_cycle[ 5296] = 1'b1;  wr_cycle[ 5296] = 1'b0;  addr_rom[ 5296]='h000004a0;  wr_data_rom[ 5296]='h00000000;
    rd_cycle[ 5297] = 1'b1;  wr_cycle[ 5297] = 1'b0;  addr_rom[ 5297]='h000004a4;  wr_data_rom[ 5297]='h00000000;
    rd_cycle[ 5298] = 1'b1;  wr_cycle[ 5298] = 1'b0;  addr_rom[ 5298]='h000004a8;  wr_data_rom[ 5298]='h00000000;
    rd_cycle[ 5299] = 1'b1;  wr_cycle[ 5299] = 1'b0;  addr_rom[ 5299]='h000004ac;  wr_data_rom[ 5299]='h00000000;
    rd_cycle[ 5300] = 1'b1;  wr_cycle[ 5300] = 1'b0;  addr_rom[ 5300]='h000004b0;  wr_data_rom[ 5300]='h00000000;
    rd_cycle[ 5301] = 1'b1;  wr_cycle[ 5301] = 1'b0;  addr_rom[ 5301]='h000004b4;  wr_data_rom[ 5301]='h00000000;
    rd_cycle[ 5302] = 1'b1;  wr_cycle[ 5302] = 1'b0;  addr_rom[ 5302]='h000004b8;  wr_data_rom[ 5302]='h00000000;
    rd_cycle[ 5303] = 1'b1;  wr_cycle[ 5303] = 1'b0;  addr_rom[ 5303]='h000004bc;  wr_data_rom[ 5303]='h00000000;
    rd_cycle[ 5304] = 1'b1;  wr_cycle[ 5304] = 1'b0;  addr_rom[ 5304]='h000004c0;  wr_data_rom[ 5304]='h00000000;
    rd_cycle[ 5305] = 1'b1;  wr_cycle[ 5305] = 1'b0;  addr_rom[ 5305]='h000004c4;  wr_data_rom[ 5305]='h00000000;
    rd_cycle[ 5306] = 1'b1;  wr_cycle[ 5306] = 1'b0;  addr_rom[ 5306]='h000004c8;  wr_data_rom[ 5306]='h00000000;
    rd_cycle[ 5307] = 1'b1;  wr_cycle[ 5307] = 1'b0;  addr_rom[ 5307]='h000004cc;  wr_data_rom[ 5307]='h00000000;
    rd_cycle[ 5308] = 1'b1;  wr_cycle[ 5308] = 1'b0;  addr_rom[ 5308]='h000004d0;  wr_data_rom[ 5308]='h00000000;
    rd_cycle[ 5309] = 1'b1;  wr_cycle[ 5309] = 1'b0;  addr_rom[ 5309]='h000004d4;  wr_data_rom[ 5309]='h00000000;
    rd_cycle[ 5310] = 1'b1;  wr_cycle[ 5310] = 1'b0;  addr_rom[ 5310]='h000004d8;  wr_data_rom[ 5310]='h00000000;
    rd_cycle[ 5311] = 1'b1;  wr_cycle[ 5311] = 1'b0;  addr_rom[ 5311]='h000004dc;  wr_data_rom[ 5311]='h00000000;
    rd_cycle[ 5312] = 1'b1;  wr_cycle[ 5312] = 1'b0;  addr_rom[ 5312]='h000004e0;  wr_data_rom[ 5312]='h00000000;
    rd_cycle[ 5313] = 1'b1;  wr_cycle[ 5313] = 1'b0;  addr_rom[ 5313]='h000004e4;  wr_data_rom[ 5313]='h00000000;
    rd_cycle[ 5314] = 1'b1;  wr_cycle[ 5314] = 1'b0;  addr_rom[ 5314]='h000004e8;  wr_data_rom[ 5314]='h00000000;
    rd_cycle[ 5315] = 1'b1;  wr_cycle[ 5315] = 1'b0;  addr_rom[ 5315]='h000004ec;  wr_data_rom[ 5315]='h00000000;
    rd_cycle[ 5316] = 1'b1;  wr_cycle[ 5316] = 1'b0;  addr_rom[ 5316]='h000004f0;  wr_data_rom[ 5316]='h00000000;
    rd_cycle[ 5317] = 1'b1;  wr_cycle[ 5317] = 1'b0;  addr_rom[ 5317]='h000004f4;  wr_data_rom[ 5317]='h00000000;
    rd_cycle[ 5318] = 1'b1;  wr_cycle[ 5318] = 1'b0;  addr_rom[ 5318]='h000004f8;  wr_data_rom[ 5318]='h00000000;
    rd_cycle[ 5319] = 1'b1;  wr_cycle[ 5319] = 1'b0;  addr_rom[ 5319]='h000004fc;  wr_data_rom[ 5319]='h00000000;
    rd_cycle[ 5320] = 1'b1;  wr_cycle[ 5320] = 1'b0;  addr_rom[ 5320]='h00000500;  wr_data_rom[ 5320]='h00000000;
    rd_cycle[ 5321] = 1'b1;  wr_cycle[ 5321] = 1'b0;  addr_rom[ 5321]='h00000504;  wr_data_rom[ 5321]='h00000000;
    rd_cycle[ 5322] = 1'b1;  wr_cycle[ 5322] = 1'b0;  addr_rom[ 5322]='h00000508;  wr_data_rom[ 5322]='h00000000;
    rd_cycle[ 5323] = 1'b1;  wr_cycle[ 5323] = 1'b0;  addr_rom[ 5323]='h0000050c;  wr_data_rom[ 5323]='h00000000;
    rd_cycle[ 5324] = 1'b1;  wr_cycle[ 5324] = 1'b0;  addr_rom[ 5324]='h00000510;  wr_data_rom[ 5324]='h00000000;
    rd_cycle[ 5325] = 1'b1;  wr_cycle[ 5325] = 1'b0;  addr_rom[ 5325]='h00000514;  wr_data_rom[ 5325]='h00000000;
    rd_cycle[ 5326] = 1'b1;  wr_cycle[ 5326] = 1'b0;  addr_rom[ 5326]='h00000518;  wr_data_rom[ 5326]='h00000000;
    rd_cycle[ 5327] = 1'b1;  wr_cycle[ 5327] = 1'b0;  addr_rom[ 5327]='h0000051c;  wr_data_rom[ 5327]='h00000000;
    rd_cycle[ 5328] = 1'b1;  wr_cycle[ 5328] = 1'b0;  addr_rom[ 5328]='h00000520;  wr_data_rom[ 5328]='h00000000;
    rd_cycle[ 5329] = 1'b1;  wr_cycle[ 5329] = 1'b0;  addr_rom[ 5329]='h00000524;  wr_data_rom[ 5329]='h00000000;
    rd_cycle[ 5330] = 1'b1;  wr_cycle[ 5330] = 1'b0;  addr_rom[ 5330]='h00000528;  wr_data_rom[ 5330]='h00000000;
    rd_cycle[ 5331] = 1'b1;  wr_cycle[ 5331] = 1'b0;  addr_rom[ 5331]='h0000052c;  wr_data_rom[ 5331]='h00000000;
    rd_cycle[ 5332] = 1'b1;  wr_cycle[ 5332] = 1'b0;  addr_rom[ 5332]='h00000530;  wr_data_rom[ 5332]='h00000000;
    rd_cycle[ 5333] = 1'b1;  wr_cycle[ 5333] = 1'b0;  addr_rom[ 5333]='h00000534;  wr_data_rom[ 5333]='h00000000;
    rd_cycle[ 5334] = 1'b1;  wr_cycle[ 5334] = 1'b0;  addr_rom[ 5334]='h00000538;  wr_data_rom[ 5334]='h00000000;
    rd_cycle[ 5335] = 1'b1;  wr_cycle[ 5335] = 1'b0;  addr_rom[ 5335]='h0000053c;  wr_data_rom[ 5335]='h00000000;
    rd_cycle[ 5336] = 1'b1;  wr_cycle[ 5336] = 1'b0;  addr_rom[ 5336]='h00000540;  wr_data_rom[ 5336]='h00000000;
    rd_cycle[ 5337] = 1'b1;  wr_cycle[ 5337] = 1'b0;  addr_rom[ 5337]='h00000544;  wr_data_rom[ 5337]='h00000000;
    rd_cycle[ 5338] = 1'b1;  wr_cycle[ 5338] = 1'b0;  addr_rom[ 5338]='h00000548;  wr_data_rom[ 5338]='h00000000;
    rd_cycle[ 5339] = 1'b1;  wr_cycle[ 5339] = 1'b0;  addr_rom[ 5339]='h0000054c;  wr_data_rom[ 5339]='h00000000;
    rd_cycle[ 5340] = 1'b1;  wr_cycle[ 5340] = 1'b0;  addr_rom[ 5340]='h00000550;  wr_data_rom[ 5340]='h00000000;
    rd_cycle[ 5341] = 1'b1;  wr_cycle[ 5341] = 1'b0;  addr_rom[ 5341]='h00000554;  wr_data_rom[ 5341]='h00000000;
    rd_cycle[ 5342] = 1'b1;  wr_cycle[ 5342] = 1'b0;  addr_rom[ 5342]='h00000558;  wr_data_rom[ 5342]='h00000000;
    rd_cycle[ 5343] = 1'b1;  wr_cycle[ 5343] = 1'b0;  addr_rom[ 5343]='h0000055c;  wr_data_rom[ 5343]='h00000000;
    rd_cycle[ 5344] = 1'b1;  wr_cycle[ 5344] = 1'b0;  addr_rom[ 5344]='h00000560;  wr_data_rom[ 5344]='h00000000;
    rd_cycle[ 5345] = 1'b1;  wr_cycle[ 5345] = 1'b0;  addr_rom[ 5345]='h00000564;  wr_data_rom[ 5345]='h00000000;
    rd_cycle[ 5346] = 1'b1;  wr_cycle[ 5346] = 1'b0;  addr_rom[ 5346]='h00000568;  wr_data_rom[ 5346]='h00000000;
    rd_cycle[ 5347] = 1'b1;  wr_cycle[ 5347] = 1'b0;  addr_rom[ 5347]='h0000056c;  wr_data_rom[ 5347]='h00000000;
    rd_cycle[ 5348] = 1'b1;  wr_cycle[ 5348] = 1'b0;  addr_rom[ 5348]='h00000570;  wr_data_rom[ 5348]='h00000000;
    rd_cycle[ 5349] = 1'b1;  wr_cycle[ 5349] = 1'b0;  addr_rom[ 5349]='h00000574;  wr_data_rom[ 5349]='h00000000;
    rd_cycle[ 5350] = 1'b1;  wr_cycle[ 5350] = 1'b0;  addr_rom[ 5350]='h00000578;  wr_data_rom[ 5350]='h00000000;
    rd_cycle[ 5351] = 1'b1;  wr_cycle[ 5351] = 1'b0;  addr_rom[ 5351]='h0000057c;  wr_data_rom[ 5351]='h00000000;
    rd_cycle[ 5352] = 1'b1;  wr_cycle[ 5352] = 1'b0;  addr_rom[ 5352]='h00000580;  wr_data_rom[ 5352]='h00000000;
    rd_cycle[ 5353] = 1'b1;  wr_cycle[ 5353] = 1'b0;  addr_rom[ 5353]='h00000584;  wr_data_rom[ 5353]='h00000000;
    rd_cycle[ 5354] = 1'b1;  wr_cycle[ 5354] = 1'b0;  addr_rom[ 5354]='h00000588;  wr_data_rom[ 5354]='h00000000;
    rd_cycle[ 5355] = 1'b1;  wr_cycle[ 5355] = 1'b0;  addr_rom[ 5355]='h0000058c;  wr_data_rom[ 5355]='h00000000;
    rd_cycle[ 5356] = 1'b1;  wr_cycle[ 5356] = 1'b0;  addr_rom[ 5356]='h00000590;  wr_data_rom[ 5356]='h00000000;
    rd_cycle[ 5357] = 1'b1;  wr_cycle[ 5357] = 1'b0;  addr_rom[ 5357]='h00000594;  wr_data_rom[ 5357]='h00000000;
    rd_cycle[ 5358] = 1'b1;  wr_cycle[ 5358] = 1'b0;  addr_rom[ 5358]='h00000598;  wr_data_rom[ 5358]='h00000000;
    rd_cycle[ 5359] = 1'b1;  wr_cycle[ 5359] = 1'b0;  addr_rom[ 5359]='h0000059c;  wr_data_rom[ 5359]='h00000000;
    rd_cycle[ 5360] = 1'b1;  wr_cycle[ 5360] = 1'b0;  addr_rom[ 5360]='h000005a0;  wr_data_rom[ 5360]='h00000000;
    rd_cycle[ 5361] = 1'b1;  wr_cycle[ 5361] = 1'b0;  addr_rom[ 5361]='h000005a4;  wr_data_rom[ 5361]='h00000000;
    rd_cycle[ 5362] = 1'b1;  wr_cycle[ 5362] = 1'b0;  addr_rom[ 5362]='h000005a8;  wr_data_rom[ 5362]='h00000000;
    rd_cycle[ 5363] = 1'b1;  wr_cycle[ 5363] = 1'b0;  addr_rom[ 5363]='h000005ac;  wr_data_rom[ 5363]='h00000000;
    rd_cycle[ 5364] = 1'b1;  wr_cycle[ 5364] = 1'b0;  addr_rom[ 5364]='h000005b0;  wr_data_rom[ 5364]='h00000000;
    rd_cycle[ 5365] = 1'b1;  wr_cycle[ 5365] = 1'b0;  addr_rom[ 5365]='h000005b4;  wr_data_rom[ 5365]='h00000000;
    rd_cycle[ 5366] = 1'b1;  wr_cycle[ 5366] = 1'b0;  addr_rom[ 5366]='h000005b8;  wr_data_rom[ 5366]='h00000000;
    rd_cycle[ 5367] = 1'b1;  wr_cycle[ 5367] = 1'b0;  addr_rom[ 5367]='h000005bc;  wr_data_rom[ 5367]='h00000000;
    rd_cycle[ 5368] = 1'b1;  wr_cycle[ 5368] = 1'b0;  addr_rom[ 5368]='h000005c0;  wr_data_rom[ 5368]='h00000000;
    rd_cycle[ 5369] = 1'b1;  wr_cycle[ 5369] = 1'b0;  addr_rom[ 5369]='h000005c4;  wr_data_rom[ 5369]='h00000000;
    rd_cycle[ 5370] = 1'b1;  wr_cycle[ 5370] = 1'b0;  addr_rom[ 5370]='h000005c8;  wr_data_rom[ 5370]='h00000000;
    rd_cycle[ 5371] = 1'b1;  wr_cycle[ 5371] = 1'b0;  addr_rom[ 5371]='h000005cc;  wr_data_rom[ 5371]='h00000000;
    rd_cycle[ 5372] = 1'b1;  wr_cycle[ 5372] = 1'b0;  addr_rom[ 5372]='h000005d0;  wr_data_rom[ 5372]='h00000000;
    rd_cycle[ 5373] = 1'b1;  wr_cycle[ 5373] = 1'b0;  addr_rom[ 5373]='h000005d4;  wr_data_rom[ 5373]='h00000000;
    rd_cycle[ 5374] = 1'b1;  wr_cycle[ 5374] = 1'b0;  addr_rom[ 5374]='h000005d8;  wr_data_rom[ 5374]='h00000000;
    rd_cycle[ 5375] = 1'b1;  wr_cycle[ 5375] = 1'b0;  addr_rom[ 5375]='h000005dc;  wr_data_rom[ 5375]='h00000000;
    rd_cycle[ 5376] = 1'b1;  wr_cycle[ 5376] = 1'b0;  addr_rom[ 5376]='h000005e0;  wr_data_rom[ 5376]='h00000000;
    rd_cycle[ 5377] = 1'b1;  wr_cycle[ 5377] = 1'b0;  addr_rom[ 5377]='h000005e4;  wr_data_rom[ 5377]='h00000000;
    rd_cycle[ 5378] = 1'b1;  wr_cycle[ 5378] = 1'b0;  addr_rom[ 5378]='h000005e8;  wr_data_rom[ 5378]='h00000000;
    rd_cycle[ 5379] = 1'b1;  wr_cycle[ 5379] = 1'b0;  addr_rom[ 5379]='h000005ec;  wr_data_rom[ 5379]='h00000000;
    rd_cycle[ 5380] = 1'b1;  wr_cycle[ 5380] = 1'b0;  addr_rom[ 5380]='h000005f0;  wr_data_rom[ 5380]='h00000000;
    rd_cycle[ 5381] = 1'b1;  wr_cycle[ 5381] = 1'b0;  addr_rom[ 5381]='h000005f4;  wr_data_rom[ 5381]='h00000000;
    rd_cycle[ 5382] = 1'b1;  wr_cycle[ 5382] = 1'b0;  addr_rom[ 5382]='h000005f8;  wr_data_rom[ 5382]='h00000000;
    rd_cycle[ 5383] = 1'b1;  wr_cycle[ 5383] = 1'b0;  addr_rom[ 5383]='h000005fc;  wr_data_rom[ 5383]='h00000000;
    rd_cycle[ 5384] = 1'b1;  wr_cycle[ 5384] = 1'b0;  addr_rom[ 5384]='h00000600;  wr_data_rom[ 5384]='h00000000;
    rd_cycle[ 5385] = 1'b1;  wr_cycle[ 5385] = 1'b0;  addr_rom[ 5385]='h00000604;  wr_data_rom[ 5385]='h00000000;
    rd_cycle[ 5386] = 1'b1;  wr_cycle[ 5386] = 1'b0;  addr_rom[ 5386]='h00000608;  wr_data_rom[ 5386]='h00000000;
    rd_cycle[ 5387] = 1'b1;  wr_cycle[ 5387] = 1'b0;  addr_rom[ 5387]='h0000060c;  wr_data_rom[ 5387]='h00000000;
    rd_cycle[ 5388] = 1'b1;  wr_cycle[ 5388] = 1'b0;  addr_rom[ 5388]='h00000610;  wr_data_rom[ 5388]='h00000000;
    rd_cycle[ 5389] = 1'b1;  wr_cycle[ 5389] = 1'b0;  addr_rom[ 5389]='h00000614;  wr_data_rom[ 5389]='h00000000;
    rd_cycle[ 5390] = 1'b1;  wr_cycle[ 5390] = 1'b0;  addr_rom[ 5390]='h00000618;  wr_data_rom[ 5390]='h00000000;
    rd_cycle[ 5391] = 1'b1;  wr_cycle[ 5391] = 1'b0;  addr_rom[ 5391]='h0000061c;  wr_data_rom[ 5391]='h00000000;
    rd_cycle[ 5392] = 1'b1;  wr_cycle[ 5392] = 1'b0;  addr_rom[ 5392]='h00000620;  wr_data_rom[ 5392]='h00000000;
    rd_cycle[ 5393] = 1'b1;  wr_cycle[ 5393] = 1'b0;  addr_rom[ 5393]='h00000624;  wr_data_rom[ 5393]='h00000000;
    rd_cycle[ 5394] = 1'b1;  wr_cycle[ 5394] = 1'b0;  addr_rom[ 5394]='h00000628;  wr_data_rom[ 5394]='h00000000;
    rd_cycle[ 5395] = 1'b1;  wr_cycle[ 5395] = 1'b0;  addr_rom[ 5395]='h0000062c;  wr_data_rom[ 5395]='h00000000;
    rd_cycle[ 5396] = 1'b1;  wr_cycle[ 5396] = 1'b0;  addr_rom[ 5396]='h00000630;  wr_data_rom[ 5396]='h00000000;
    rd_cycle[ 5397] = 1'b1;  wr_cycle[ 5397] = 1'b0;  addr_rom[ 5397]='h00000634;  wr_data_rom[ 5397]='h00000000;
    rd_cycle[ 5398] = 1'b1;  wr_cycle[ 5398] = 1'b0;  addr_rom[ 5398]='h00000638;  wr_data_rom[ 5398]='h00000000;
    rd_cycle[ 5399] = 1'b1;  wr_cycle[ 5399] = 1'b0;  addr_rom[ 5399]='h0000063c;  wr_data_rom[ 5399]='h00000000;
    rd_cycle[ 5400] = 1'b1;  wr_cycle[ 5400] = 1'b0;  addr_rom[ 5400]='h00000640;  wr_data_rom[ 5400]='h00000000;
    rd_cycle[ 5401] = 1'b1;  wr_cycle[ 5401] = 1'b0;  addr_rom[ 5401]='h00000644;  wr_data_rom[ 5401]='h00000000;
    rd_cycle[ 5402] = 1'b1;  wr_cycle[ 5402] = 1'b0;  addr_rom[ 5402]='h00000648;  wr_data_rom[ 5402]='h00000000;
    rd_cycle[ 5403] = 1'b1;  wr_cycle[ 5403] = 1'b0;  addr_rom[ 5403]='h0000064c;  wr_data_rom[ 5403]='h00000000;
    rd_cycle[ 5404] = 1'b1;  wr_cycle[ 5404] = 1'b0;  addr_rom[ 5404]='h00000650;  wr_data_rom[ 5404]='h00000000;
    rd_cycle[ 5405] = 1'b1;  wr_cycle[ 5405] = 1'b0;  addr_rom[ 5405]='h00000654;  wr_data_rom[ 5405]='h00000000;
    rd_cycle[ 5406] = 1'b1;  wr_cycle[ 5406] = 1'b0;  addr_rom[ 5406]='h00000658;  wr_data_rom[ 5406]='h00000000;
    rd_cycle[ 5407] = 1'b1;  wr_cycle[ 5407] = 1'b0;  addr_rom[ 5407]='h0000065c;  wr_data_rom[ 5407]='h00000000;
    rd_cycle[ 5408] = 1'b1;  wr_cycle[ 5408] = 1'b0;  addr_rom[ 5408]='h00000660;  wr_data_rom[ 5408]='h00000000;
    rd_cycle[ 5409] = 1'b1;  wr_cycle[ 5409] = 1'b0;  addr_rom[ 5409]='h00000664;  wr_data_rom[ 5409]='h00000000;
    rd_cycle[ 5410] = 1'b1;  wr_cycle[ 5410] = 1'b0;  addr_rom[ 5410]='h00000668;  wr_data_rom[ 5410]='h00000000;
    rd_cycle[ 5411] = 1'b1;  wr_cycle[ 5411] = 1'b0;  addr_rom[ 5411]='h0000066c;  wr_data_rom[ 5411]='h00000000;
    rd_cycle[ 5412] = 1'b1;  wr_cycle[ 5412] = 1'b0;  addr_rom[ 5412]='h00000670;  wr_data_rom[ 5412]='h00000000;
    rd_cycle[ 5413] = 1'b1;  wr_cycle[ 5413] = 1'b0;  addr_rom[ 5413]='h00000674;  wr_data_rom[ 5413]='h00000000;
    rd_cycle[ 5414] = 1'b1;  wr_cycle[ 5414] = 1'b0;  addr_rom[ 5414]='h00000678;  wr_data_rom[ 5414]='h00000000;
    rd_cycle[ 5415] = 1'b1;  wr_cycle[ 5415] = 1'b0;  addr_rom[ 5415]='h0000067c;  wr_data_rom[ 5415]='h00000000;
    rd_cycle[ 5416] = 1'b1;  wr_cycle[ 5416] = 1'b0;  addr_rom[ 5416]='h00000680;  wr_data_rom[ 5416]='h00000000;
    rd_cycle[ 5417] = 1'b1;  wr_cycle[ 5417] = 1'b0;  addr_rom[ 5417]='h00000684;  wr_data_rom[ 5417]='h00000000;
    rd_cycle[ 5418] = 1'b1;  wr_cycle[ 5418] = 1'b0;  addr_rom[ 5418]='h00000688;  wr_data_rom[ 5418]='h00000000;
    rd_cycle[ 5419] = 1'b1;  wr_cycle[ 5419] = 1'b0;  addr_rom[ 5419]='h0000068c;  wr_data_rom[ 5419]='h00000000;
    rd_cycle[ 5420] = 1'b1;  wr_cycle[ 5420] = 1'b0;  addr_rom[ 5420]='h00000690;  wr_data_rom[ 5420]='h00000000;
    rd_cycle[ 5421] = 1'b1;  wr_cycle[ 5421] = 1'b0;  addr_rom[ 5421]='h00000694;  wr_data_rom[ 5421]='h00000000;
    rd_cycle[ 5422] = 1'b1;  wr_cycle[ 5422] = 1'b0;  addr_rom[ 5422]='h00000698;  wr_data_rom[ 5422]='h00000000;
    rd_cycle[ 5423] = 1'b1;  wr_cycle[ 5423] = 1'b0;  addr_rom[ 5423]='h0000069c;  wr_data_rom[ 5423]='h00000000;
    rd_cycle[ 5424] = 1'b1;  wr_cycle[ 5424] = 1'b0;  addr_rom[ 5424]='h000006a0;  wr_data_rom[ 5424]='h00000000;
    rd_cycle[ 5425] = 1'b1;  wr_cycle[ 5425] = 1'b0;  addr_rom[ 5425]='h000006a4;  wr_data_rom[ 5425]='h00000000;
    rd_cycle[ 5426] = 1'b1;  wr_cycle[ 5426] = 1'b0;  addr_rom[ 5426]='h000006a8;  wr_data_rom[ 5426]='h00000000;
    rd_cycle[ 5427] = 1'b1;  wr_cycle[ 5427] = 1'b0;  addr_rom[ 5427]='h000006ac;  wr_data_rom[ 5427]='h00000000;
    rd_cycle[ 5428] = 1'b1;  wr_cycle[ 5428] = 1'b0;  addr_rom[ 5428]='h000006b0;  wr_data_rom[ 5428]='h00000000;
    rd_cycle[ 5429] = 1'b1;  wr_cycle[ 5429] = 1'b0;  addr_rom[ 5429]='h000006b4;  wr_data_rom[ 5429]='h00000000;
    rd_cycle[ 5430] = 1'b1;  wr_cycle[ 5430] = 1'b0;  addr_rom[ 5430]='h000006b8;  wr_data_rom[ 5430]='h00000000;
    rd_cycle[ 5431] = 1'b1;  wr_cycle[ 5431] = 1'b0;  addr_rom[ 5431]='h000006bc;  wr_data_rom[ 5431]='h00000000;
    rd_cycle[ 5432] = 1'b1;  wr_cycle[ 5432] = 1'b0;  addr_rom[ 5432]='h000006c0;  wr_data_rom[ 5432]='h00000000;
    rd_cycle[ 5433] = 1'b1;  wr_cycle[ 5433] = 1'b0;  addr_rom[ 5433]='h000006c4;  wr_data_rom[ 5433]='h00000000;
    rd_cycle[ 5434] = 1'b1;  wr_cycle[ 5434] = 1'b0;  addr_rom[ 5434]='h000006c8;  wr_data_rom[ 5434]='h00000000;
    rd_cycle[ 5435] = 1'b1;  wr_cycle[ 5435] = 1'b0;  addr_rom[ 5435]='h000006cc;  wr_data_rom[ 5435]='h00000000;
    rd_cycle[ 5436] = 1'b1;  wr_cycle[ 5436] = 1'b0;  addr_rom[ 5436]='h000006d0;  wr_data_rom[ 5436]='h00000000;
    rd_cycle[ 5437] = 1'b1;  wr_cycle[ 5437] = 1'b0;  addr_rom[ 5437]='h000006d4;  wr_data_rom[ 5437]='h00000000;
    rd_cycle[ 5438] = 1'b1;  wr_cycle[ 5438] = 1'b0;  addr_rom[ 5438]='h000006d8;  wr_data_rom[ 5438]='h00000000;
    rd_cycle[ 5439] = 1'b1;  wr_cycle[ 5439] = 1'b0;  addr_rom[ 5439]='h000006dc;  wr_data_rom[ 5439]='h00000000;
    rd_cycle[ 5440] = 1'b1;  wr_cycle[ 5440] = 1'b0;  addr_rom[ 5440]='h000006e0;  wr_data_rom[ 5440]='h00000000;
    rd_cycle[ 5441] = 1'b1;  wr_cycle[ 5441] = 1'b0;  addr_rom[ 5441]='h000006e4;  wr_data_rom[ 5441]='h00000000;
    rd_cycle[ 5442] = 1'b1;  wr_cycle[ 5442] = 1'b0;  addr_rom[ 5442]='h000006e8;  wr_data_rom[ 5442]='h00000000;
    rd_cycle[ 5443] = 1'b1;  wr_cycle[ 5443] = 1'b0;  addr_rom[ 5443]='h000006ec;  wr_data_rom[ 5443]='h00000000;
    rd_cycle[ 5444] = 1'b1;  wr_cycle[ 5444] = 1'b0;  addr_rom[ 5444]='h000006f0;  wr_data_rom[ 5444]='h00000000;
    rd_cycle[ 5445] = 1'b1;  wr_cycle[ 5445] = 1'b0;  addr_rom[ 5445]='h000006f4;  wr_data_rom[ 5445]='h00000000;
    rd_cycle[ 5446] = 1'b1;  wr_cycle[ 5446] = 1'b0;  addr_rom[ 5446]='h000006f8;  wr_data_rom[ 5446]='h00000000;
    rd_cycle[ 5447] = 1'b1;  wr_cycle[ 5447] = 1'b0;  addr_rom[ 5447]='h000006fc;  wr_data_rom[ 5447]='h00000000;
    rd_cycle[ 5448] = 1'b1;  wr_cycle[ 5448] = 1'b0;  addr_rom[ 5448]='h00000700;  wr_data_rom[ 5448]='h00000000;
    rd_cycle[ 5449] = 1'b1;  wr_cycle[ 5449] = 1'b0;  addr_rom[ 5449]='h00000704;  wr_data_rom[ 5449]='h00000000;
    rd_cycle[ 5450] = 1'b1;  wr_cycle[ 5450] = 1'b0;  addr_rom[ 5450]='h00000708;  wr_data_rom[ 5450]='h00000000;
    rd_cycle[ 5451] = 1'b1;  wr_cycle[ 5451] = 1'b0;  addr_rom[ 5451]='h0000070c;  wr_data_rom[ 5451]='h00000000;
    rd_cycle[ 5452] = 1'b1;  wr_cycle[ 5452] = 1'b0;  addr_rom[ 5452]='h00000710;  wr_data_rom[ 5452]='h00000000;
    rd_cycle[ 5453] = 1'b1;  wr_cycle[ 5453] = 1'b0;  addr_rom[ 5453]='h00000714;  wr_data_rom[ 5453]='h00000000;
    rd_cycle[ 5454] = 1'b1;  wr_cycle[ 5454] = 1'b0;  addr_rom[ 5454]='h00000718;  wr_data_rom[ 5454]='h00000000;
    rd_cycle[ 5455] = 1'b1;  wr_cycle[ 5455] = 1'b0;  addr_rom[ 5455]='h0000071c;  wr_data_rom[ 5455]='h00000000;
    rd_cycle[ 5456] = 1'b1;  wr_cycle[ 5456] = 1'b0;  addr_rom[ 5456]='h00000720;  wr_data_rom[ 5456]='h00000000;
    rd_cycle[ 5457] = 1'b1;  wr_cycle[ 5457] = 1'b0;  addr_rom[ 5457]='h00000724;  wr_data_rom[ 5457]='h00000000;
    rd_cycle[ 5458] = 1'b1;  wr_cycle[ 5458] = 1'b0;  addr_rom[ 5458]='h00000728;  wr_data_rom[ 5458]='h00000000;
    rd_cycle[ 5459] = 1'b1;  wr_cycle[ 5459] = 1'b0;  addr_rom[ 5459]='h0000072c;  wr_data_rom[ 5459]='h00000000;
    rd_cycle[ 5460] = 1'b1;  wr_cycle[ 5460] = 1'b0;  addr_rom[ 5460]='h00000730;  wr_data_rom[ 5460]='h00000000;
    rd_cycle[ 5461] = 1'b1;  wr_cycle[ 5461] = 1'b0;  addr_rom[ 5461]='h00000734;  wr_data_rom[ 5461]='h00000000;
    rd_cycle[ 5462] = 1'b1;  wr_cycle[ 5462] = 1'b0;  addr_rom[ 5462]='h00000738;  wr_data_rom[ 5462]='h00000000;
    rd_cycle[ 5463] = 1'b1;  wr_cycle[ 5463] = 1'b0;  addr_rom[ 5463]='h0000073c;  wr_data_rom[ 5463]='h00000000;
    rd_cycle[ 5464] = 1'b1;  wr_cycle[ 5464] = 1'b0;  addr_rom[ 5464]='h00000740;  wr_data_rom[ 5464]='h00000000;
    rd_cycle[ 5465] = 1'b1;  wr_cycle[ 5465] = 1'b0;  addr_rom[ 5465]='h00000744;  wr_data_rom[ 5465]='h00000000;
    rd_cycle[ 5466] = 1'b1;  wr_cycle[ 5466] = 1'b0;  addr_rom[ 5466]='h00000748;  wr_data_rom[ 5466]='h00000000;
    rd_cycle[ 5467] = 1'b1;  wr_cycle[ 5467] = 1'b0;  addr_rom[ 5467]='h0000074c;  wr_data_rom[ 5467]='h00000000;
    rd_cycle[ 5468] = 1'b1;  wr_cycle[ 5468] = 1'b0;  addr_rom[ 5468]='h00000750;  wr_data_rom[ 5468]='h00000000;
    rd_cycle[ 5469] = 1'b1;  wr_cycle[ 5469] = 1'b0;  addr_rom[ 5469]='h00000754;  wr_data_rom[ 5469]='h00000000;
    rd_cycle[ 5470] = 1'b1;  wr_cycle[ 5470] = 1'b0;  addr_rom[ 5470]='h00000758;  wr_data_rom[ 5470]='h00000000;
    rd_cycle[ 5471] = 1'b1;  wr_cycle[ 5471] = 1'b0;  addr_rom[ 5471]='h0000075c;  wr_data_rom[ 5471]='h00000000;
    rd_cycle[ 5472] = 1'b1;  wr_cycle[ 5472] = 1'b0;  addr_rom[ 5472]='h00000760;  wr_data_rom[ 5472]='h00000000;
    rd_cycle[ 5473] = 1'b1;  wr_cycle[ 5473] = 1'b0;  addr_rom[ 5473]='h00000764;  wr_data_rom[ 5473]='h00000000;
    rd_cycle[ 5474] = 1'b1;  wr_cycle[ 5474] = 1'b0;  addr_rom[ 5474]='h00000768;  wr_data_rom[ 5474]='h00000000;
    rd_cycle[ 5475] = 1'b1;  wr_cycle[ 5475] = 1'b0;  addr_rom[ 5475]='h0000076c;  wr_data_rom[ 5475]='h00000000;
    rd_cycle[ 5476] = 1'b1;  wr_cycle[ 5476] = 1'b0;  addr_rom[ 5476]='h00000770;  wr_data_rom[ 5476]='h00000000;
    rd_cycle[ 5477] = 1'b1;  wr_cycle[ 5477] = 1'b0;  addr_rom[ 5477]='h00000774;  wr_data_rom[ 5477]='h00000000;
    rd_cycle[ 5478] = 1'b1;  wr_cycle[ 5478] = 1'b0;  addr_rom[ 5478]='h00000778;  wr_data_rom[ 5478]='h00000000;
    rd_cycle[ 5479] = 1'b1;  wr_cycle[ 5479] = 1'b0;  addr_rom[ 5479]='h0000077c;  wr_data_rom[ 5479]='h00000000;
    rd_cycle[ 5480] = 1'b1;  wr_cycle[ 5480] = 1'b0;  addr_rom[ 5480]='h00000780;  wr_data_rom[ 5480]='h00000000;
    rd_cycle[ 5481] = 1'b1;  wr_cycle[ 5481] = 1'b0;  addr_rom[ 5481]='h00000784;  wr_data_rom[ 5481]='h00000000;
    rd_cycle[ 5482] = 1'b1;  wr_cycle[ 5482] = 1'b0;  addr_rom[ 5482]='h00000788;  wr_data_rom[ 5482]='h00000000;
    rd_cycle[ 5483] = 1'b1;  wr_cycle[ 5483] = 1'b0;  addr_rom[ 5483]='h0000078c;  wr_data_rom[ 5483]='h00000000;
    rd_cycle[ 5484] = 1'b1;  wr_cycle[ 5484] = 1'b0;  addr_rom[ 5484]='h00000790;  wr_data_rom[ 5484]='h00000000;
    rd_cycle[ 5485] = 1'b1;  wr_cycle[ 5485] = 1'b0;  addr_rom[ 5485]='h00000794;  wr_data_rom[ 5485]='h00000000;
    rd_cycle[ 5486] = 1'b1;  wr_cycle[ 5486] = 1'b0;  addr_rom[ 5486]='h00000798;  wr_data_rom[ 5486]='h00000000;
    rd_cycle[ 5487] = 1'b1;  wr_cycle[ 5487] = 1'b0;  addr_rom[ 5487]='h0000079c;  wr_data_rom[ 5487]='h00000000;
    rd_cycle[ 5488] = 1'b1;  wr_cycle[ 5488] = 1'b0;  addr_rom[ 5488]='h000007a0;  wr_data_rom[ 5488]='h00000000;
    rd_cycle[ 5489] = 1'b1;  wr_cycle[ 5489] = 1'b0;  addr_rom[ 5489]='h000007a4;  wr_data_rom[ 5489]='h00000000;
    rd_cycle[ 5490] = 1'b1;  wr_cycle[ 5490] = 1'b0;  addr_rom[ 5490]='h000007a8;  wr_data_rom[ 5490]='h00000000;
    rd_cycle[ 5491] = 1'b1;  wr_cycle[ 5491] = 1'b0;  addr_rom[ 5491]='h000007ac;  wr_data_rom[ 5491]='h00000000;
    rd_cycle[ 5492] = 1'b1;  wr_cycle[ 5492] = 1'b0;  addr_rom[ 5492]='h000007b0;  wr_data_rom[ 5492]='h00000000;
    rd_cycle[ 5493] = 1'b1;  wr_cycle[ 5493] = 1'b0;  addr_rom[ 5493]='h000007b4;  wr_data_rom[ 5493]='h00000000;
    rd_cycle[ 5494] = 1'b1;  wr_cycle[ 5494] = 1'b0;  addr_rom[ 5494]='h000007b8;  wr_data_rom[ 5494]='h00000000;
    rd_cycle[ 5495] = 1'b1;  wr_cycle[ 5495] = 1'b0;  addr_rom[ 5495]='h000007bc;  wr_data_rom[ 5495]='h00000000;
    rd_cycle[ 5496] = 1'b1;  wr_cycle[ 5496] = 1'b0;  addr_rom[ 5496]='h000007c0;  wr_data_rom[ 5496]='h00000000;
    rd_cycle[ 5497] = 1'b1;  wr_cycle[ 5497] = 1'b0;  addr_rom[ 5497]='h000007c4;  wr_data_rom[ 5497]='h00000000;
    rd_cycle[ 5498] = 1'b1;  wr_cycle[ 5498] = 1'b0;  addr_rom[ 5498]='h000007c8;  wr_data_rom[ 5498]='h00000000;
    rd_cycle[ 5499] = 1'b1;  wr_cycle[ 5499] = 1'b0;  addr_rom[ 5499]='h000007cc;  wr_data_rom[ 5499]='h00000000;
    rd_cycle[ 5500] = 1'b1;  wr_cycle[ 5500] = 1'b0;  addr_rom[ 5500]='h000007d0;  wr_data_rom[ 5500]='h00000000;
    rd_cycle[ 5501] = 1'b1;  wr_cycle[ 5501] = 1'b0;  addr_rom[ 5501]='h000007d4;  wr_data_rom[ 5501]='h00000000;
    rd_cycle[ 5502] = 1'b1;  wr_cycle[ 5502] = 1'b0;  addr_rom[ 5502]='h000007d8;  wr_data_rom[ 5502]='h00000000;
    rd_cycle[ 5503] = 1'b1;  wr_cycle[ 5503] = 1'b0;  addr_rom[ 5503]='h000007dc;  wr_data_rom[ 5503]='h00000000;
    rd_cycle[ 5504] = 1'b1;  wr_cycle[ 5504] = 1'b0;  addr_rom[ 5504]='h000007e0;  wr_data_rom[ 5504]='h00000000;
    rd_cycle[ 5505] = 1'b1;  wr_cycle[ 5505] = 1'b0;  addr_rom[ 5505]='h000007e4;  wr_data_rom[ 5505]='h00000000;
    rd_cycle[ 5506] = 1'b1;  wr_cycle[ 5506] = 1'b0;  addr_rom[ 5506]='h000007e8;  wr_data_rom[ 5506]='h00000000;
    rd_cycle[ 5507] = 1'b1;  wr_cycle[ 5507] = 1'b0;  addr_rom[ 5507]='h000007ec;  wr_data_rom[ 5507]='h00000000;
    rd_cycle[ 5508] = 1'b1;  wr_cycle[ 5508] = 1'b0;  addr_rom[ 5508]='h000007f0;  wr_data_rom[ 5508]='h00000000;
    rd_cycle[ 5509] = 1'b1;  wr_cycle[ 5509] = 1'b0;  addr_rom[ 5509]='h000007f4;  wr_data_rom[ 5509]='h00000000;
    rd_cycle[ 5510] = 1'b1;  wr_cycle[ 5510] = 1'b0;  addr_rom[ 5510]='h000007f8;  wr_data_rom[ 5510]='h00000000;
    rd_cycle[ 5511] = 1'b1;  wr_cycle[ 5511] = 1'b0;  addr_rom[ 5511]='h000007fc;  wr_data_rom[ 5511]='h00000000;
    rd_cycle[ 5512] = 1'b1;  wr_cycle[ 5512] = 1'b0;  addr_rom[ 5512]='h00000800;  wr_data_rom[ 5512]='h00000000;
    rd_cycle[ 5513] = 1'b1;  wr_cycle[ 5513] = 1'b0;  addr_rom[ 5513]='h00000804;  wr_data_rom[ 5513]='h00000000;
    rd_cycle[ 5514] = 1'b1;  wr_cycle[ 5514] = 1'b0;  addr_rom[ 5514]='h00000808;  wr_data_rom[ 5514]='h00000000;
    rd_cycle[ 5515] = 1'b1;  wr_cycle[ 5515] = 1'b0;  addr_rom[ 5515]='h0000080c;  wr_data_rom[ 5515]='h00000000;
    rd_cycle[ 5516] = 1'b1;  wr_cycle[ 5516] = 1'b0;  addr_rom[ 5516]='h00000810;  wr_data_rom[ 5516]='h00000000;
    rd_cycle[ 5517] = 1'b1;  wr_cycle[ 5517] = 1'b0;  addr_rom[ 5517]='h00000814;  wr_data_rom[ 5517]='h00000000;
    rd_cycle[ 5518] = 1'b1;  wr_cycle[ 5518] = 1'b0;  addr_rom[ 5518]='h00000818;  wr_data_rom[ 5518]='h00000000;
    rd_cycle[ 5519] = 1'b1;  wr_cycle[ 5519] = 1'b0;  addr_rom[ 5519]='h0000081c;  wr_data_rom[ 5519]='h00000000;
    rd_cycle[ 5520] = 1'b1;  wr_cycle[ 5520] = 1'b0;  addr_rom[ 5520]='h00000820;  wr_data_rom[ 5520]='h00000000;
    rd_cycle[ 5521] = 1'b1;  wr_cycle[ 5521] = 1'b0;  addr_rom[ 5521]='h00000824;  wr_data_rom[ 5521]='h00000000;
    rd_cycle[ 5522] = 1'b1;  wr_cycle[ 5522] = 1'b0;  addr_rom[ 5522]='h00000828;  wr_data_rom[ 5522]='h00000000;
    rd_cycle[ 5523] = 1'b1;  wr_cycle[ 5523] = 1'b0;  addr_rom[ 5523]='h0000082c;  wr_data_rom[ 5523]='h00000000;
    rd_cycle[ 5524] = 1'b1;  wr_cycle[ 5524] = 1'b0;  addr_rom[ 5524]='h00000830;  wr_data_rom[ 5524]='h00000000;
    rd_cycle[ 5525] = 1'b1;  wr_cycle[ 5525] = 1'b0;  addr_rom[ 5525]='h00000834;  wr_data_rom[ 5525]='h00000000;
    rd_cycle[ 5526] = 1'b1;  wr_cycle[ 5526] = 1'b0;  addr_rom[ 5526]='h00000838;  wr_data_rom[ 5526]='h00000000;
    rd_cycle[ 5527] = 1'b1;  wr_cycle[ 5527] = 1'b0;  addr_rom[ 5527]='h0000083c;  wr_data_rom[ 5527]='h00000000;
    rd_cycle[ 5528] = 1'b1;  wr_cycle[ 5528] = 1'b0;  addr_rom[ 5528]='h00000840;  wr_data_rom[ 5528]='h00000000;
    rd_cycle[ 5529] = 1'b1;  wr_cycle[ 5529] = 1'b0;  addr_rom[ 5529]='h00000844;  wr_data_rom[ 5529]='h00000000;
    rd_cycle[ 5530] = 1'b1;  wr_cycle[ 5530] = 1'b0;  addr_rom[ 5530]='h00000848;  wr_data_rom[ 5530]='h00000000;
    rd_cycle[ 5531] = 1'b1;  wr_cycle[ 5531] = 1'b0;  addr_rom[ 5531]='h0000084c;  wr_data_rom[ 5531]='h00000000;
    rd_cycle[ 5532] = 1'b1;  wr_cycle[ 5532] = 1'b0;  addr_rom[ 5532]='h00000850;  wr_data_rom[ 5532]='h00000000;
    rd_cycle[ 5533] = 1'b1;  wr_cycle[ 5533] = 1'b0;  addr_rom[ 5533]='h00000854;  wr_data_rom[ 5533]='h00000000;
    rd_cycle[ 5534] = 1'b1;  wr_cycle[ 5534] = 1'b0;  addr_rom[ 5534]='h00000858;  wr_data_rom[ 5534]='h00000000;
    rd_cycle[ 5535] = 1'b1;  wr_cycle[ 5535] = 1'b0;  addr_rom[ 5535]='h0000085c;  wr_data_rom[ 5535]='h00000000;
    rd_cycle[ 5536] = 1'b1;  wr_cycle[ 5536] = 1'b0;  addr_rom[ 5536]='h00000860;  wr_data_rom[ 5536]='h00000000;
    rd_cycle[ 5537] = 1'b1;  wr_cycle[ 5537] = 1'b0;  addr_rom[ 5537]='h00000864;  wr_data_rom[ 5537]='h00000000;
    rd_cycle[ 5538] = 1'b1;  wr_cycle[ 5538] = 1'b0;  addr_rom[ 5538]='h00000868;  wr_data_rom[ 5538]='h00000000;
    rd_cycle[ 5539] = 1'b1;  wr_cycle[ 5539] = 1'b0;  addr_rom[ 5539]='h0000086c;  wr_data_rom[ 5539]='h00000000;
    rd_cycle[ 5540] = 1'b1;  wr_cycle[ 5540] = 1'b0;  addr_rom[ 5540]='h00000870;  wr_data_rom[ 5540]='h00000000;
    rd_cycle[ 5541] = 1'b1;  wr_cycle[ 5541] = 1'b0;  addr_rom[ 5541]='h00000874;  wr_data_rom[ 5541]='h00000000;
    rd_cycle[ 5542] = 1'b1;  wr_cycle[ 5542] = 1'b0;  addr_rom[ 5542]='h00000878;  wr_data_rom[ 5542]='h00000000;
    rd_cycle[ 5543] = 1'b1;  wr_cycle[ 5543] = 1'b0;  addr_rom[ 5543]='h0000087c;  wr_data_rom[ 5543]='h00000000;
    rd_cycle[ 5544] = 1'b1;  wr_cycle[ 5544] = 1'b0;  addr_rom[ 5544]='h00000880;  wr_data_rom[ 5544]='h00000000;
    rd_cycle[ 5545] = 1'b1;  wr_cycle[ 5545] = 1'b0;  addr_rom[ 5545]='h00000884;  wr_data_rom[ 5545]='h00000000;
    rd_cycle[ 5546] = 1'b1;  wr_cycle[ 5546] = 1'b0;  addr_rom[ 5546]='h00000888;  wr_data_rom[ 5546]='h00000000;
    rd_cycle[ 5547] = 1'b1;  wr_cycle[ 5547] = 1'b0;  addr_rom[ 5547]='h0000088c;  wr_data_rom[ 5547]='h00000000;
    rd_cycle[ 5548] = 1'b1;  wr_cycle[ 5548] = 1'b0;  addr_rom[ 5548]='h00000890;  wr_data_rom[ 5548]='h00000000;
    rd_cycle[ 5549] = 1'b1;  wr_cycle[ 5549] = 1'b0;  addr_rom[ 5549]='h00000894;  wr_data_rom[ 5549]='h00000000;
    rd_cycle[ 5550] = 1'b1;  wr_cycle[ 5550] = 1'b0;  addr_rom[ 5550]='h00000898;  wr_data_rom[ 5550]='h00000000;
    rd_cycle[ 5551] = 1'b1;  wr_cycle[ 5551] = 1'b0;  addr_rom[ 5551]='h0000089c;  wr_data_rom[ 5551]='h00000000;
    rd_cycle[ 5552] = 1'b1;  wr_cycle[ 5552] = 1'b0;  addr_rom[ 5552]='h000008a0;  wr_data_rom[ 5552]='h00000000;
    rd_cycle[ 5553] = 1'b1;  wr_cycle[ 5553] = 1'b0;  addr_rom[ 5553]='h000008a4;  wr_data_rom[ 5553]='h00000000;
    rd_cycle[ 5554] = 1'b1;  wr_cycle[ 5554] = 1'b0;  addr_rom[ 5554]='h000008a8;  wr_data_rom[ 5554]='h00000000;
    rd_cycle[ 5555] = 1'b1;  wr_cycle[ 5555] = 1'b0;  addr_rom[ 5555]='h000008ac;  wr_data_rom[ 5555]='h00000000;
    rd_cycle[ 5556] = 1'b1;  wr_cycle[ 5556] = 1'b0;  addr_rom[ 5556]='h000008b0;  wr_data_rom[ 5556]='h00000000;
    rd_cycle[ 5557] = 1'b1;  wr_cycle[ 5557] = 1'b0;  addr_rom[ 5557]='h000008b4;  wr_data_rom[ 5557]='h00000000;
    rd_cycle[ 5558] = 1'b1;  wr_cycle[ 5558] = 1'b0;  addr_rom[ 5558]='h000008b8;  wr_data_rom[ 5558]='h00000000;
    rd_cycle[ 5559] = 1'b1;  wr_cycle[ 5559] = 1'b0;  addr_rom[ 5559]='h000008bc;  wr_data_rom[ 5559]='h00000000;
    rd_cycle[ 5560] = 1'b1;  wr_cycle[ 5560] = 1'b0;  addr_rom[ 5560]='h000008c0;  wr_data_rom[ 5560]='h00000000;
    rd_cycle[ 5561] = 1'b1;  wr_cycle[ 5561] = 1'b0;  addr_rom[ 5561]='h000008c4;  wr_data_rom[ 5561]='h00000000;
    rd_cycle[ 5562] = 1'b1;  wr_cycle[ 5562] = 1'b0;  addr_rom[ 5562]='h000008c8;  wr_data_rom[ 5562]='h00000000;
    rd_cycle[ 5563] = 1'b1;  wr_cycle[ 5563] = 1'b0;  addr_rom[ 5563]='h000008cc;  wr_data_rom[ 5563]='h00000000;
    rd_cycle[ 5564] = 1'b1;  wr_cycle[ 5564] = 1'b0;  addr_rom[ 5564]='h000008d0;  wr_data_rom[ 5564]='h00000000;
    rd_cycle[ 5565] = 1'b1;  wr_cycle[ 5565] = 1'b0;  addr_rom[ 5565]='h000008d4;  wr_data_rom[ 5565]='h00000000;
    rd_cycle[ 5566] = 1'b1;  wr_cycle[ 5566] = 1'b0;  addr_rom[ 5566]='h000008d8;  wr_data_rom[ 5566]='h00000000;
    rd_cycle[ 5567] = 1'b1;  wr_cycle[ 5567] = 1'b0;  addr_rom[ 5567]='h000008dc;  wr_data_rom[ 5567]='h00000000;
    rd_cycle[ 5568] = 1'b1;  wr_cycle[ 5568] = 1'b0;  addr_rom[ 5568]='h000008e0;  wr_data_rom[ 5568]='h00000000;
    rd_cycle[ 5569] = 1'b1;  wr_cycle[ 5569] = 1'b0;  addr_rom[ 5569]='h000008e4;  wr_data_rom[ 5569]='h00000000;
    rd_cycle[ 5570] = 1'b1;  wr_cycle[ 5570] = 1'b0;  addr_rom[ 5570]='h000008e8;  wr_data_rom[ 5570]='h00000000;
    rd_cycle[ 5571] = 1'b1;  wr_cycle[ 5571] = 1'b0;  addr_rom[ 5571]='h000008ec;  wr_data_rom[ 5571]='h00000000;
    rd_cycle[ 5572] = 1'b1;  wr_cycle[ 5572] = 1'b0;  addr_rom[ 5572]='h000008f0;  wr_data_rom[ 5572]='h00000000;
    rd_cycle[ 5573] = 1'b1;  wr_cycle[ 5573] = 1'b0;  addr_rom[ 5573]='h000008f4;  wr_data_rom[ 5573]='h00000000;
    rd_cycle[ 5574] = 1'b1;  wr_cycle[ 5574] = 1'b0;  addr_rom[ 5574]='h000008f8;  wr_data_rom[ 5574]='h00000000;
    rd_cycle[ 5575] = 1'b1;  wr_cycle[ 5575] = 1'b0;  addr_rom[ 5575]='h000008fc;  wr_data_rom[ 5575]='h00000000;
    rd_cycle[ 5576] = 1'b1;  wr_cycle[ 5576] = 1'b0;  addr_rom[ 5576]='h00000900;  wr_data_rom[ 5576]='h00000000;
    rd_cycle[ 5577] = 1'b1;  wr_cycle[ 5577] = 1'b0;  addr_rom[ 5577]='h00000904;  wr_data_rom[ 5577]='h00000000;
    rd_cycle[ 5578] = 1'b1;  wr_cycle[ 5578] = 1'b0;  addr_rom[ 5578]='h00000908;  wr_data_rom[ 5578]='h00000000;
    rd_cycle[ 5579] = 1'b1;  wr_cycle[ 5579] = 1'b0;  addr_rom[ 5579]='h0000090c;  wr_data_rom[ 5579]='h00000000;
    rd_cycle[ 5580] = 1'b1;  wr_cycle[ 5580] = 1'b0;  addr_rom[ 5580]='h00000910;  wr_data_rom[ 5580]='h00000000;
    rd_cycle[ 5581] = 1'b1;  wr_cycle[ 5581] = 1'b0;  addr_rom[ 5581]='h00000914;  wr_data_rom[ 5581]='h00000000;
    rd_cycle[ 5582] = 1'b1;  wr_cycle[ 5582] = 1'b0;  addr_rom[ 5582]='h00000918;  wr_data_rom[ 5582]='h00000000;
    rd_cycle[ 5583] = 1'b1;  wr_cycle[ 5583] = 1'b0;  addr_rom[ 5583]='h0000091c;  wr_data_rom[ 5583]='h00000000;
    rd_cycle[ 5584] = 1'b1;  wr_cycle[ 5584] = 1'b0;  addr_rom[ 5584]='h00000920;  wr_data_rom[ 5584]='h00000000;
    rd_cycle[ 5585] = 1'b1;  wr_cycle[ 5585] = 1'b0;  addr_rom[ 5585]='h00000924;  wr_data_rom[ 5585]='h00000000;
    rd_cycle[ 5586] = 1'b1;  wr_cycle[ 5586] = 1'b0;  addr_rom[ 5586]='h00000928;  wr_data_rom[ 5586]='h00000000;
    rd_cycle[ 5587] = 1'b1;  wr_cycle[ 5587] = 1'b0;  addr_rom[ 5587]='h0000092c;  wr_data_rom[ 5587]='h00000000;
    rd_cycle[ 5588] = 1'b1;  wr_cycle[ 5588] = 1'b0;  addr_rom[ 5588]='h00000930;  wr_data_rom[ 5588]='h00000000;
    rd_cycle[ 5589] = 1'b1;  wr_cycle[ 5589] = 1'b0;  addr_rom[ 5589]='h00000934;  wr_data_rom[ 5589]='h00000000;
    rd_cycle[ 5590] = 1'b1;  wr_cycle[ 5590] = 1'b0;  addr_rom[ 5590]='h00000938;  wr_data_rom[ 5590]='h00000000;
    rd_cycle[ 5591] = 1'b1;  wr_cycle[ 5591] = 1'b0;  addr_rom[ 5591]='h0000093c;  wr_data_rom[ 5591]='h00000000;
    rd_cycle[ 5592] = 1'b1;  wr_cycle[ 5592] = 1'b0;  addr_rom[ 5592]='h00000940;  wr_data_rom[ 5592]='h00000000;
    rd_cycle[ 5593] = 1'b1;  wr_cycle[ 5593] = 1'b0;  addr_rom[ 5593]='h00000944;  wr_data_rom[ 5593]='h00000000;
    rd_cycle[ 5594] = 1'b1;  wr_cycle[ 5594] = 1'b0;  addr_rom[ 5594]='h00000948;  wr_data_rom[ 5594]='h00000000;
    rd_cycle[ 5595] = 1'b1;  wr_cycle[ 5595] = 1'b0;  addr_rom[ 5595]='h0000094c;  wr_data_rom[ 5595]='h00000000;
    rd_cycle[ 5596] = 1'b1;  wr_cycle[ 5596] = 1'b0;  addr_rom[ 5596]='h00000950;  wr_data_rom[ 5596]='h00000000;
    rd_cycle[ 5597] = 1'b1;  wr_cycle[ 5597] = 1'b0;  addr_rom[ 5597]='h00000954;  wr_data_rom[ 5597]='h00000000;
    rd_cycle[ 5598] = 1'b1;  wr_cycle[ 5598] = 1'b0;  addr_rom[ 5598]='h00000958;  wr_data_rom[ 5598]='h00000000;
    rd_cycle[ 5599] = 1'b1;  wr_cycle[ 5599] = 1'b0;  addr_rom[ 5599]='h0000095c;  wr_data_rom[ 5599]='h00000000;
    rd_cycle[ 5600] = 1'b1;  wr_cycle[ 5600] = 1'b0;  addr_rom[ 5600]='h00000960;  wr_data_rom[ 5600]='h00000000;
    rd_cycle[ 5601] = 1'b1;  wr_cycle[ 5601] = 1'b0;  addr_rom[ 5601]='h00000964;  wr_data_rom[ 5601]='h00000000;
    rd_cycle[ 5602] = 1'b1;  wr_cycle[ 5602] = 1'b0;  addr_rom[ 5602]='h00000968;  wr_data_rom[ 5602]='h00000000;
    rd_cycle[ 5603] = 1'b1;  wr_cycle[ 5603] = 1'b0;  addr_rom[ 5603]='h0000096c;  wr_data_rom[ 5603]='h00000000;
    rd_cycle[ 5604] = 1'b1;  wr_cycle[ 5604] = 1'b0;  addr_rom[ 5604]='h00000970;  wr_data_rom[ 5604]='h00000000;
    rd_cycle[ 5605] = 1'b1;  wr_cycle[ 5605] = 1'b0;  addr_rom[ 5605]='h00000974;  wr_data_rom[ 5605]='h00000000;
    rd_cycle[ 5606] = 1'b1;  wr_cycle[ 5606] = 1'b0;  addr_rom[ 5606]='h00000978;  wr_data_rom[ 5606]='h00000000;
    rd_cycle[ 5607] = 1'b1;  wr_cycle[ 5607] = 1'b0;  addr_rom[ 5607]='h0000097c;  wr_data_rom[ 5607]='h00000000;
    rd_cycle[ 5608] = 1'b1;  wr_cycle[ 5608] = 1'b0;  addr_rom[ 5608]='h00000980;  wr_data_rom[ 5608]='h00000000;
    rd_cycle[ 5609] = 1'b1;  wr_cycle[ 5609] = 1'b0;  addr_rom[ 5609]='h00000984;  wr_data_rom[ 5609]='h00000000;
    rd_cycle[ 5610] = 1'b1;  wr_cycle[ 5610] = 1'b0;  addr_rom[ 5610]='h00000988;  wr_data_rom[ 5610]='h00000000;
    rd_cycle[ 5611] = 1'b1;  wr_cycle[ 5611] = 1'b0;  addr_rom[ 5611]='h0000098c;  wr_data_rom[ 5611]='h00000000;
    rd_cycle[ 5612] = 1'b1;  wr_cycle[ 5612] = 1'b0;  addr_rom[ 5612]='h00000990;  wr_data_rom[ 5612]='h00000000;
    rd_cycle[ 5613] = 1'b1;  wr_cycle[ 5613] = 1'b0;  addr_rom[ 5613]='h00000994;  wr_data_rom[ 5613]='h00000000;
    rd_cycle[ 5614] = 1'b1;  wr_cycle[ 5614] = 1'b0;  addr_rom[ 5614]='h00000998;  wr_data_rom[ 5614]='h00000000;
    rd_cycle[ 5615] = 1'b1;  wr_cycle[ 5615] = 1'b0;  addr_rom[ 5615]='h0000099c;  wr_data_rom[ 5615]='h00000000;
    rd_cycle[ 5616] = 1'b1;  wr_cycle[ 5616] = 1'b0;  addr_rom[ 5616]='h000009a0;  wr_data_rom[ 5616]='h00000000;
    rd_cycle[ 5617] = 1'b1;  wr_cycle[ 5617] = 1'b0;  addr_rom[ 5617]='h000009a4;  wr_data_rom[ 5617]='h00000000;
    rd_cycle[ 5618] = 1'b1;  wr_cycle[ 5618] = 1'b0;  addr_rom[ 5618]='h000009a8;  wr_data_rom[ 5618]='h00000000;
    rd_cycle[ 5619] = 1'b1;  wr_cycle[ 5619] = 1'b0;  addr_rom[ 5619]='h000009ac;  wr_data_rom[ 5619]='h00000000;
    rd_cycle[ 5620] = 1'b1;  wr_cycle[ 5620] = 1'b0;  addr_rom[ 5620]='h000009b0;  wr_data_rom[ 5620]='h00000000;
    rd_cycle[ 5621] = 1'b1;  wr_cycle[ 5621] = 1'b0;  addr_rom[ 5621]='h000009b4;  wr_data_rom[ 5621]='h00000000;
    rd_cycle[ 5622] = 1'b1;  wr_cycle[ 5622] = 1'b0;  addr_rom[ 5622]='h000009b8;  wr_data_rom[ 5622]='h00000000;
    rd_cycle[ 5623] = 1'b1;  wr_cycle[ 5623] = 1'b0;  addr_rom[ 5623]='h000009bc;  wr_data_rom[ 5623]='h00000000;
    rd_cycle[ 5624] = 1'b1;  wr_cycle[ 5624] = 1'b0;  addr_rom[ 5624]='h000009c0;  wr_data_rom[ 5624]='h00000000;
    rd_cycle[ 5625] = 1'b1;  wr_cycle[ 5625] = 1'b0;  addr_rom[ 5625]='h000009c4;  wr_data_rom[ 5625]='h00000000;
    rd_cycle[ 5626] = 1'b1;  wr_cycle[ 5626] = 1'b0;  addr_rom[ 5626]='h000009c8;  wr_data_rom[ 5626]='h00000000;
    rd_cycle[ 5627] = 1'b1;  wr_cycle[ 5627] = 1'b0;  addr_rom[ 5627]='h000009cc;  wr_data_rom[ 5627]='h00000000;
    rd_cycle[ 5628] = 1'b1;  wr_cycle[ 5628] = 1'b0;  addr_rom[ 5628]='h000009d0;  wr_data_rom[ 5628]='h00000000;
    rd_cycle[ 5629] = 1'b1;  wr_cycle[ 5629] = 1'b0;  addr_rom[ 5629]='h000009d4;  wr_data_rom[ 5629]='h00000000;
    rd_cycle[ 5630] = 1'b1;  wr_cycle[ 5630] = 1'b0;  addr_rom[ 5630]='h000009d8;  wr_data_rom[ 5630]='h00000000;
    rd_cycle[ 5631] = 1'b1;  wr_cycle[ 5631] = 1'b0;  addr_rom[ 5631]='h000009dc;  wr_data_rom[ 5631]='h00000000;
    rd_cycle[ 5632] = 1'b1;  wr_cycle[ 5632] = 1'b0;  addr_rom[ 5632]='h000009e0;  wr_data_rom[ 5632]='h00000000;
    rd_cycle[ 5633] = 1'b1;  wr_cycle[ 5633] = 1'b0;  addr_rom[ 5633]='h000009e4;  wr_data_rom[ 5633]='h00000000;
    rd_cycle[ 5634] = 1'b1;  wr_cycle[ 5634] = 1'b0;  addr_rom[ 5634]='h000009e8;  wr_data_rom[ 5634]='h00000000;
    rd_cycle[ 5635] = 1'b1;  wr_cycle[ 5635] = 1'b0;  addr_rom[ 5635]='h000009ec;  wr_data_rom[ 5635]='h00000000;
    rd_cycle[ 5636] = 1'b1;  wr_cycle[ 5636] = 1'b0;  addr_rom[ 5636]='h000009f0;  wr_data_rom[ 5636]='h00000000;
    rd_cycle[ 5637] = 1'b1;  wr_cycle[ 5637] = 1'b0;  addr_rom[ 5637]='h000009f4;  wr_data_rom[ 5637]='h00000000;
    rd_cycle[ 5638] = 1'b1;  wr_cycle[ 5638] = 1'b0;  addr_rom[ 5638]='h000009f8;  wr_data_rom[ 5638]='h00000000;
    rd_cycle[ 5639] = 1'b1;  wr_cycle[ 5639] = 1'b0;  addr_rom[ 5639]='h000009fc;  wr_data_rom[ 5639]='h00000000;
    rd_cycle[ 5640] = 1'b1;  wr_cycle[ 5640] = 1'b0;  addr_rom[ 5640]='h00000a00;  wr_data_rom[ 5640]='h00000000;
    rd_cycle[ 5641] = 1'b1;  wr_cycle[ 5641] = 1'b0;  addr_rom[ 5641]='h00000a04;  wr_data_rom[ 5641]='h00000000;
    rd_cycle[ 5642] = 1'b1;  wr_cycle[ 5642] = 1'b0;  addr_rom[ 5642]='h00000a08;  wr_data_rom[ 5642]='h00000000;
    rd_cycle[ 5643] = 1'b1;  wr_cycle[ 5643] = 1'b0;  addr_rom[ 5643]='h00000a0c;  wr_data_rom[ 5643]='h00000000;
    rd_cycle[ 5644] = 1'b1;  wr_cycle[ 5644] = 1'b0;  addr_rom[ 5644]='h00000a10;  wr_data_rom[ 5644]='h00000000;
    rd_cycle[ 5645] = 1'b1;  wr_cycle[ 5645] = 1'b0;  addr_rom[ 5645]='h00000a14;  wr_data_rom[ 5645]='h00000000;
    rd_cycle[ 5646] = 1'b1;  wr_cycle[ 5646] = 1'b0;  addr_rom[ 5646]='h00000a18;  wr_data_rom[ 5646]='h00000000;
    rd_cycle[ 5647] = 1'b1;  wr_cycle[ 5647] = 1'b0;  addr_rom[ 5647]='h00000a1c;  wr_data_rom[ 5647]='h00000000;
    rd_cycle[ 5648] = 1'b1;  wr_cycle[ 5648] = 1'b0;  addr_rom[ 5648]='h00000a20;  wr_data_rom[ 5648]='h00000000;
    rd_cycle[ 5649] = 1'b1;  wr_cycle[ 5649] = 1'b0;  addr_rom[ 5649]='h00000a24;  wr_data_rom[ 5649]='h00000000;
    rd_cycle[ 5650] = 1'b1;  wr_cycle[ 5650] = 1'b0;  addr_rom[ 5650]='h00000a28;  wr_data_rom[ 5650]='h00000000;
    rd_cycle[ 5651] = 1'b1;  wr_cycle[ 5651] = 1'b0;  addr_rom[ 5651]='h00000a2c;  wr_data_rom[ 5651]='h00000000;
    rd_cycle[ 5652] = 1'b1;  wr_cycle[ 5652] = 1'b0;  addr_rom[ 5652]='h00000a30;  wr_data_rom[ 5652]='h00000000;
    rd_cycle[ 5653] = 1'b1;  wr_cycle[ 5653] = 1'b0;  addr_rom[ 5653]='h00000a34;  wr_data_rom[ 5653]='h00000000;
    rd_cycle[ 5654] = 1'b1;  wr_cycle[ 5654] = 1'b0;  addr_rom[ 5654]='h00000a38;  wr_data_rom[ 5654]='h00000000;
    rd_cycle[ 5655] = 1'b1;  wr_cycle[ 5655] = 1'b0;  addr_rom[ 5655]='h00000a3c;  wr_data_rom[ 5655]='h00000000;
    rd_cycle[ 5656] = 1'b1;  wr_cycle[ 5656] = 1'b0;  addr_rom[ 5656]='h00000a40;  wr_data_rom[ 5656]='h00000000;
    rd_cycle[ 5657] = 1'b1;  wr_cycle[ 5657] = 1'b0;  addr_rom[ 5657]='h00000a44;  wr_data_rom[ 5657]='h00000000;
    rd_cycle[ 5658] = 1'b1;  wr_cycle[ 5658] = 1'b0;  addr_rom[ 5658]='h00000a48;  wr_data_rom[ 5658]='h00000000;
    rd_cycle[ 5659] = 1'b1;  wr_cycle[ 5659] = 1'b0;  addr_rom[ 5659]='h00000a4c;  wr_data_rom[ 5659]='h00000000;
    rd_cycle[ 5660] = 1'b1;  wr_cycle[ 5660] = 1'b0;  addr_rom[ 5660]='h00000a50;  wr_data_rom[ 5660]='h00000000;
    rd_cycle[ 5661] = 1'b1;  wr_cycle[ 5661] = 1'b0;  addr_rom[ 5661]='h00000a54;  wr_data_rom[ 5661]='h00000000;
    rd_cycle[ 5662] = 1'b1;  wr_cycle[ 5662] = 1'b0;  addr_rom[ 5662]='h00000a58;  wr_data_rom[ 5662]='h00000000;
    rd_cycle[ 5663] = 1'b1;  wr_cycle[ 5663] = 1'b0;  addr_rom[ 5663]='h00000a5c;  wr_data_rom[ 5663]='h00000000;
    rd_cycle[ 5664] = 1'b1;  wr_cycle[ 5664] = 1'b0;  addr_rom[ 5664]='h00000a60;  wr_data_rom[ 5664]='h00000000;
    rd_cycle[ 5665] = 1'b1;  wr_cycle[ 5665] = 1'b0;  addr_rom[ 5665]='h00000a64;  wr_data_rom[ 5665]='h00000000;
    rd_cycle[ 5666] = 1'b1;  wr_cycle[ 5666] = 1'b0;  addr_rom[ 5666]='h00000a68;  wr_data_rom[ 5666]='h00000000;
    rd_cycle[ 5667] = 1'b1;  wr_cycle[ 5667] = 1'b0;  addr_rom[ 5667]='h00000a6c;  wr_data_rom[ 5667]='h00000000;
    rd_cycle[ 5668] = 1'b1;  wr_cycle[ 5668] = 1'b0;  addr_rom[ 5668]='h00000a70;  wr_data_rom[ 5668]='h00000000;
    rd_cycle[ 5669] = 1'b1;  wr_cycle[ 5669] = 1'b0;  addr_rom[ 5669]='h00000a74;  wr_data_rom[ 5669]='h00000000;
    rd_cycle[ 5670] = 1'b1;  wr_cycle[ 5670] = 1'b0;  addr_rom[ 5670]='h00000a78;  wr_data_rom[ 5670]='h00000000;
    rd_cycle[ 5671] = 1'b1;  wr_cycle[ 5671] = 1'b0;  addr_rom[ 5671]='h00000a7c;  wr_data_rom[ 5671]='h00000000;
    rd_cycle[ 5672] = 1'b1;  wr_cycle[ 5672] = 1'b0;  addr_rom[ 5672]='h00000a80;  wr_data_rom[ 5672]='h00000000;
    rd_cycle[ 5673] = 1'b1;  wr_cycle[ 5673] = 1'b0;  addr_rom[ 5673]='h00000a84;  wr_data_rom[ 5673]='h00000000;
    rd_cycle[ 5674] = 1'b1;  wr_cycle[ 5674] = 1'b0;  addr_rom[ 5674]='h00000a88;  wr_data_rom[ 5674]='h00000000;
    rd_cycle[ 5675] = 1'b1;  wr_cycle[ 5675] = 1'b0;  addr_rom[ 5675]='h00000a8c;  wr_data_rom[ 5675]='h00000000;
    rd_cycle[ 5676] = 1'b1;  wr_cycle[ 5676] = 1'b0;  addr_rom[ 5676]='h00000a90;  wr_data_rom[ 5676]='h00000000;
    rd_cycle[ 5677] = 1'b1;  wr_cycle[ 5677] = 1'b0;  addr_rom[ 5677]='h00000a94;  wr_data_rom[ 5677]='h00000000;
    rd_cycle[ 5678] = 1'b1;  wr_cycle[ 5678] = 1'b0;  addr_rom[ 5678]='h00000a98;  wr_data_rom[ 5678]='h00000000;
    rd_cycle[ 5679] = 1'b1;  wr_cycle[ 5679] = 1'b0;  addr_rom[ 5679]='h00000a9c;  wr_data_rom[ 5679]='h00000000;
    rd_cycle[ 5680] = 1'b1;  wr_cycle[ 5680] = 1'b0;  addr_rom[ 5680]='h00000aa0;  wr_data_rom[ 5680]='h00000000;
    rd_cycle[ 5681] = 1'b1;  wr_cycle[ 5681] = 1'b0;  addr_rom[ 5681]='h00000aa4;  wr_data_rom[ 5681]='h00000000;
    rd_cycle[ 5682] = 1'b1;  wr_cycle[ 5682] = 1'b0;  addr_rom[ 5682]='h00000aa8;  wr_data_rom[ 5682]='h00000000;
    rd_cycle[ 5683] = 1'b1;  wr_cycle[ 5683] = 1'b0;  addr_rom[ 5683]='h00000aac;  wr_data_rom[ 5683]='h00000000;
    rd_cycle[ 5684] = 1'b1;  wr_cycle[ 5684] = 1'b0;  addr_rom[ 5684]='h00000ab0;  wr_data_rom[ 5684]='h00000000;
    rd_cycle[ 5685] = 1'b1;  wr_cycle[ 5685] = 1'b0;  addr_rom[ 5685]='h00000ab4;  wr_data_rom[ 5685]='h00000000;
    rd_cycle[ 5686] = 1'b1;  wr_cycle[ 5686] = 1'b0;  addr_rom[ 5686]='h00000ab8;  wr_data_rom[ 5686]='h00000000;
    rd_cycle[ 5687] = 1'b1;  wr_cycle[ 5687] = 1'b0;  addr_rom[ 5687]='h00000abc;  wr_data_rom[ 5687]='h00000000;
    rd_cycle[ 5688] = 1'b1;  wr_cycle[ 5688] = 1'b0;  addr_rom[ 5688]='h00000ac0;  wr_data_rom[ 5688]='h00000000;
    rd_cycle[ 5689] = 1'b1;  wr_cycle[ 5689] = 1'b0;  addr_rom[ 5689]='h00000ac4;  wr_data_rom[ 5689]='h00000000;
    rd_cycle[ 5690] = 1'b1;  wr_cycle[ 5690] = 1'b0;  addr_rom[ 5690]='h00000ac8;  wr_data_rom[ 5690]='h00000000;
    rd_cycle[ 5691] = 1'b1;  wr_cycle[ 5691] = 1'b0;  addr_rom[ 5691]='h00000acc;  wr_data_rom[ 5691]='h00000000;
    rd_cycle[ 5692] = 1'b1;  wr_cycle[ 5692] = 1'b0;  addr_rom[ 5692]='h00000ad0;  wr_data_rom[ 5692]='h00000000;
    rd_cycle[ 5693] = 1'b1;  wr_cycle[ 5693] = 1'b0;  addr_rom[ 5693]='h00000ad4;  wr_data_rom[ 5693]='h00000000;
    rd_cycle[ 5694] = 1'b1;  wr_cycle[ 5694] = 1'b0;  addr_rom[ 5694]='h00000ad8;  wr_data_rom[ 5694]='h00000000;
    rd_cycle[ 5695] = 1'b1;  wr_cycle[ 5695] = 1'b0;  addr_rom[ 5695]='h00000adc;  wr_data_rom[ 5695]='h00000000;
    rd_cycle[ 5696] = 1'b1;  wr_cycle[ 5696] = 1'b0;  addr_rom[ 5696]='h00000ae0;  wr_data_rom[ 5696]='h00000000;
    rd_cycle[ 5697] = 1'b1;  wr_cycle[ 5697] = 1'b0;  addr_rom[ 5697]='h00000ae4;  wr_data_rom[ 5697]='h00000000;
    rd_cycle[ 5698] = 1'b1;  wr_cycle[ 5698] = 1'b0;  addr_rom[ 5698]='h00000ae8;  wr_data_rom[ 5698]='h00000000;
    rd_cycle[ 5699] = 1'b1;  wr_cycle[ 5699] = 1'b0;  addr_rom[ 5699]='h00000aec;  wr_data_rom[ 5699]='h00000000;
    rd_cycle[ 5700] = 1'b1;  wr_cycle[ 5700] = 1'b0;  addr_rom[ 5700]='h00000af0;  wr_data_rom[ 5700]='h00000000;
    rd_cycle[ 5701] = 1'b1;  wr_cycle[ 5701] = 1'b0;  addr_rom[ 5701]='h00000af4;  wr_data_rom[ 5701]='h00000000;
    rd_cycle[ 5702] = 1'b1;  wr_cycle[ 5702] = 1'b0;  addr_rom[ 5702]='h00000af8;  wr_data_rom[ 5702]='h00000000;
    rd_cycle[ 5703] = 1'b1;  wr_cycle[ 5703] = 1'b0;  addr_rom[ 5703]='h00000afc;  wr_data_rom[ 5703]='h00000000;
    rd_cycle[ 5704] = 1'b1;  wr_cycle[ 5704] = 1'b0;  addr_rom[ 5704]='h00000b00;  wr_data_rom[ 5704]='h00000000;
    rd_cycle[ 5705] = 1'b1;  wr_cycle[ 5705] = 1'b0;  addr_rom[ 5705]='h00000b04;  wr_data_rom[ 5705]='h00000000;
    rd_cycle[ 5706] = 1'b1;  wr_cycle[ 5706] = 1'b0;  addr_rom[ 5706]='h00000b08;  wr_data_rom[ 5706]='h00000000;
    rd_cycle[ 5707] = 1'b1;  wr_cycle[ 5707] = 1'b0;  addr_rom[ 5707]='h00000b0c;  wr_data_rom[ 5707]='h00000000;
    rd_cycle[ 5708] = 1'b1;  wr_cycle[ 5708] = 1'b0;  addr_rom[ 5708]='h00000b10;  wr_data_rom[ 5708]='h00000000;
    rd_cycle[ 5709] = 1'b1;  wr_cycle[ 5709] = 1'b0;  addr_rom[ 5709]='h00000b14;  wr_data_rom[ 5709]='h00000000;
    rd_cycle[ 5710] = 1'b1;  wr_cycle[ 5710] = 1'b0;  addr_rom[ 5710]='h00000b18;  wr_data_rom[ 5710]='h00000000;
    rd_cycle[ 5711] = 1'b1;  wr_cycle[ 5711] = 1'b0;  addr_rom[ 5711]='h00000b1c;  wr_data_rom[ 5711]='h00000000;
    rd_cycle[ 5712] = 1'b1;  wr_cycle[ 5712] = 1'b0;  addr_rom[ 5712]='h00000b20;  wr_data_rom[ 5712]='h00000000;
    rd_cycle[ 5713] = 1'b1;  wr_cycle[ 5713] = 1'b0;  addr_rom[ 5713]='h00000b24;  wr_data_rom[ 5713]='h00000000;
    rd_cycle[ 5714] = 1'b1;  wr_cycle[ 5714] = 1'b0;  addr_rom[ 5714]='h00000b28;  wr_data_rom[ 5714]='h00000000;
    rd_cycle[ 5715] = 1'b1;  wr_cycle[ 5715] = 1'b0;  addr_rom[ 5715]='h00000b2c;  wr_data_rom[ 5715]='h00000000;
    rd_cycle[ 5716] = 1'b1;  wr_cycle[ 5716] = 1'b0;  addr_rom[ 5716]='h00000b30;  wr_data_rom[ 5716]='h00000000;
    rd_cycle[ 5717] = 1'b1;  wr_cycle[ 5717] = 1'b0;  addr_rom[ 5717]='h00000b34;  wr_data_rom[ 5717]='h00000000;
    rd_cycle[ 5718] = 1'b1;  wr_cycle[ 5718] = 1'b0;  addr_rom[ 5718]='h00000b38;  wr_data_rom[ 5718]='h00000000;
    rd_cycle[ 5719] = 1'b1;  wr_cycle[ 5719] = 1'b0;  addr_rom[ 5719]='h00000b3c;  wr_data_rom[ 5719]='h00000000;
    rd_cycle[ 5720] = 1'b1;  wr_cycle[ 5720] = 1'b0;  addr_rom[ 5720]='h00000b40;  wr_data_rom[ 5720]='h00000000;
    rd_cycle[ 5721] = 1'b1;  wr_cycle[ 5721] = 1'b0;  addr_rom[ 5721]='h00000b44;  wr_data_rom[ 5721]='h00000000;
    rd_cycle[ 5722] = 1'b1;  wr_cycle[ 5722] = 1'b0;  addr_rom[ 5722]='h00000b48;  wr_data_rom[ 5722]='h00000000;
    rd_cycle[ 5723] = 1'b1;  wr_cycle[ 5723] = 1'b0;  addr_rom[ 5723]='h00000b4c;  wr_data_rom[ 5723]='h00000000;
    rd_cycle[ 5724] = 1'b1;  wr_cycle[ 5724] = 1'b0;  addr_rom[ 5724]='h00000b50;  wr_data_rom[ 5724]='h00000000;
    rd_cycle[ 5725] = 1'b1;  wr_cycle[ 5725] = 1'b0;  addr_rom[ 5725]='h00000b54;  wr_data_rom[ 5725]='h00000000;
    rd_cycle[ 5726] = 1'b1;  wr_cycle[ 5726] = 1'b0;  addr_rom[ 5726]='h00000b58;  wr_data_rom[ 5726]='h00000000;
    rd_cycle[ 5727] = 1'b1;  wr_cycle[ 5727] = 1'b0;  addr_rom[ 5727]='h00000b5c;  wr_data_rom[ 5727]='h00000000;
    rd_cycle[ 5728] = 1'b1;  wr_cycle[ 5728] = 1'b0;  addr_rom[ 5728]='h00000b60;  wr_data_rom[ 5728]='h00000000;
    rd_cycle[ 5729] = 1'b1;  wr_cycle[ 5729] = 1'b0;  addr_rom[ 5729]='h00000b64;  wr_data_rom[ 5729]='h00000000;
    rd_cycle[ 5730] = 1'b1;  wr_cycle[ 5730] = 1'b0;  addr_rom[ 5730]='h00000b68;  wr_data_rom[ 5730]='h00000000;
    rd_cycle[ 5731] = 1'b1;  wr_cycle[ 5731] = 1'b0;  addr_rom[ 5731]='h00000b6c;  wr_data_rom[ 5731]='h00000000;
    rd_cycle[ 5732] = 1'b1;  wr_cycle[ 5732] = 1'b0;  addr_rom[ 5732]='h00000b70;  wr_data_rom[ 5732]='h00000000;
    rd_cycle[ 5733] = 1'b1;  wr_cycle[ 5733] = 1'b0;  addr_rom[ 5733]='h00000b74;  wr_data_rom[ 5733]='h00000000;
    rd_cycle[ 5734] = 1'b1;  wr_cycle[ 5734] = 1'b0;  addr_rom[ 5734]='h00000b78;  wr_data_rom[ 5734]='h00000000;
    rd_cycle[ 5735] = 1'b1;  wr_cycle[ 5735] = 1'b0;  addr_rom[ 5735]='h00000b7c;  wr_data_rom[ 5735]='h00000000;
    rd_cycle[ 5736] = 1'b1;  wr_cycle[ 5736] = 1'b0;  addr_rom[ 5736]='h00000b80;  wr_data_rom[ 5736]='h00000000;
    rd_cycle[ 5737] = 1'b1;  wr_cycle[ 5737] = 1'b0;  addr_rom[ 5737]='h00000b84;  wr_data_rom[ 5737]='h00000000;
    rd_cycle[ 5738] = 1'b1;  wr_cycle[ 5738] = 1'b0;  addr_rom[ 5738]='h00000b88;  wr_data_rom[ 5738]='h00000000;
    rd_cycle[ 5739] = 1'b1;  wr_cycle[ 5739] = 1'b0;  addr_rom[ 5739]='h00000b8c;  wr_data_rom[ 5739]='h00000000;
    rd_cycle[ 5740] = 1'b1;  wr_cycle[ 5740] = 1'b0;  addr_rom[ 5740]='h00000b90;  wr_data_rom[ 5740]='h00000000;
    rd_cycle[ 5741] = 1'b1;  wr_cycle[ 5741] = 1'b0;  addr_rom[ 5741]='h00000b94;  wr_data_rom[ 5741]='h00000000;
    rd_cycle[ 5742] = 1'b1;  wr_cycle[ 5742] = 1'b0;  addr_rom[ 5742]='h00000b98;  wr_data_rom[ 5742]='h00000000;
    rd_cycle[ 5743] = 1'b1;  wr_cycle[ 5743] = 1'b0;  addr_rom[ 5743]='h00000b9c;  wr_data_rom[ 5743]='h00000000;
    rd_cycle[ 5744] = 1'b1;  wr_cycle[ 5744] = 1'b0;  addr_rom[ 5744]='h00000ba0;  wr_data_rom[ 5744]='h00000000;
    rd_cycle[ 5745] = 1'b1;  wr_cycle[ 5745] = 1'b0;  addr_rom[ 5745]='h00000ba4;  wr_data_rom[ 5745]='h00000000;
    rd_cycle[ 5746] = 1'b1;  wr_cycle[ 5746] = 1'b0;  addr_rom[ 5746]='h00000ba8;  wr_data_rom[ 5746]='h00000000;
    rd_cycle[ 5747] = 1'b1;  wr_cycle[ 5747] = 1'b0;  addr_rom[ 5747]='h00000bac;  wr_data_rom[ 5747]='h00000000;
    rd_cycle[ 5748] = 1'b1;  wr_cycle[ 5748] = 1'b0;  addr_rom[ 5748]='h00000bb0;  wr_data_rom[ 5748]='h00000000;
    rd_cycle[ 5749] = 1'b1;  wr_cycle[ 5749] = 1'b0;  addr_rom[ 5749]='h00000bb4;  wr_data_rom[ 5749]='h00000000;
    rd_cycle[ 5750] = 1'b1;  wr_cycle[ 5750] = 1'b0;  addr_rom[ 5750]='h00000bb8;  wr_data_rom[ 5750]='h00000000;
    rd_cycle[ 5751] = 1'b1;  wr_cycle[ 5751] = 1'b0;  addr_rom[ 5751]='h00000bbc;  wr_data_rom[ 5751]='h00000000;
    rd_cycle[ 5752] = 1'b1;  wr_cycle[ 5752] = 1'b0;  addr_rom[ 5752]='h00000bc0;  wr_data_rom[ 5752]='h00000000;
    rd_cycle[ 5753] = 1'b1;  wr_cycle[ 5753] = 1'b0;  addr_rom[ 5753]='h00000bc4;  wr_data_rom[ 5753]='h00000000;
    rd_cycle[ 5754] = 1'b1;  wr_cycle[ 5754] = 1'b0;  addr_rom[ 5754]='h00000bc8;  wr_data_rom[ 5754]='h00000000;
    rd_cycle[ 5755] = 1'b1;  wr_cycle[ 5755] = 1'b0;  addr_rom[ 5755]='h00000bcc;  wr_data_rom[ 5755]='h00000000;
    rd_cycle[ 5756] = 1'b1;  wr_cycle[ 5756] = 1'b0;  addr_rom[ 5756]='h00000bd0;  wr_data_rom[ 5756]='h00000000;
    rd_cycle[ 5757] = 1'b1;  wr_cycle[ 5757] = 1'b0;  addr_rom[ 5757]='h00000bd4;  wr_data_rom[ 5757]='h00000000;
    rd_cycle[ 5758] = 1'b1;  wr_cycle[ 5758] = 1'b0;  addr_rom[ 5758]='h00000bd8;  wr_data_rom[ 5758]='h00000000;
    rd_cycle[ 5759] = 1'b1;  wr_cycle[ 5759] = 1'b0;  addr_rom[ 5759]='h00000bdc;  wr_data_rom[ 5759]='h00000000;
    rd_cycle[ 5760] = 1'b1;  wr_cycle[ 5760] = 1'b0;  addr_rom[ 5760]='h00000be0;  wr_data_rom[ 5760]='h00000000;
    rd_cycle[ 5761] = 1'b1;  wr_cycle[ 5761] = 1'b0;  addr_rom[ 5761]='h00000be4;  wr_data_rom[ 5761]='h00000000;
    rd_cycle[ 5762] = 1'b1;  wr_cycle[ 5762] = 1'b0;  addr_rom[ 5762]='h00000be8;  wr_data_rom[ 5762]='h00000000;
    rd_cycle[ 5763] = 1'b1;  wr_cycle[ 5763] = 1'b0;  addr_rom[ 5763]='h00000bec;  wr_data_rom[ 5763]='h00000000;
    rd_cycle[ 5764] = 1'b1;  wr_cycle[ 5764] = 1'b0;  addr_rom[ 5764]='h00000bf0;  wr_data_rom[ 5764]='h00000000;
    rd_cycle[ 5765] = 1'b1;  wr_cycle[ 5765] = 1'b0;  addr_rom[ 5765]='h00000bf4;  wr_data_rom[ 5765]='h00000000;
    rd_cycle[ 5766] = 1'b1;  wr_cycle[ 5766] = 1'b0;  addr_rom[ 5766]='h00000bf8;  wr_data_rom[ 5766]='h00000000;
    rd_cycle[ 5767] = 1'b1;  wr_cycle[ 5767] = 1'b0;  addr_rom[ 5767]='h00000bfc;  wr_data_rom[ 5767]='h00000000;
    rd_cycle[ 5768] = 1'b1;  wr_cycle[ 5768] = 1'b0;  addr_rom[ 5768]='h00000c00;  wr_data_rom[ 5768]='h00000000;
    rd_cycle[ 5769] = 1'b1;  wr_cycle[ 5769] = 1'b0;  addr_rom[ 5769]='h00000c04;  wr_data_rom[ 5769]='h00000000;
    rd_cycle[ 5770] = 1'b1;  wr_cycle[ 5770] = 1'b0;  addr_rom[ 5770]='h00000c08;  wr_data_rom[ 5770]='h00000000;
    rd_cycle[ 5771] = 1'b1;  wr_cycle[ 5771] = 1'b0;  addr_rom[ 5771]='h00000c0c;  wr_data_rom[ 5771]='h00000000;
    rd_cycle[ 5772] = 1'b1;  wr_cycle[ 5772] = 1'b0;  addr_rom[ 5772]='h00000c10;  wr_data_rom[ 5772]='h00000000;
    rd_cycle[ 5773] = 1'b1;  wr_cycle[ 5773] = 1'b0;  addr_rom[ 5773]='h00000c14;  wr_data_rom[ 5773]='h00000000;
    rd_cycle[ 5774] = 1'b1;  wr_cycle[ 5774] = 1'b0;  addr_rom[ 5774]='h00000c18;  wr_data_rom[ 5774]='h00000000;
    rd_cycle[ 5775] = 1'b1;  wr_cycle[ 5775] = 1'b0;  addr_rom[ 5775]='h00000c1c;  wr_data_rom[ 5775]='h00000000;
    rd_cycle[ 5776] = 1'b1;  wr_cycle[ 5776] = 1'b0;  addr_rom[ 5776]='h00000c20;  wr_data_rom[ 5776]='h00000000;
    rd_cycle[ 5777] = 1'b1;  wr_cycle[ 5777] = 1'b0;  addr_rom[ 5777]='h00000c24;  wr_data_rom[ 5777]='h00000000;
    rd_cycle[ 5778] = 1'b1;  wr_cycle[ 5778] = 1'b0;  addr_rom[ 5778]='h00000c28;  wr_data_rom[ 5778]='h00000000;
    rd_cycle[ 5779] = 1'b1;  wr_cycle[ 5779] = 1'b0;  addr_rom[ 5779]='h00000c2c;  wr_data_rom[ 5779]='h00000000;
    rd_cycle[ 5780] = 1'b1;  wr_cycle[ 5780] = 1'b0;  addr_rom[ 5780]='h00000c30;  wr_data_rom[ 5780]='h00000000;
    rd_cycle[ 5781] = 1'b1;  wr_cycle[ 5781] = 1'b0;  addr_rom[ 5781]='h00000c34;  wr_data_rom[ 5781]='h00000000;
    rd_cycle[ 5782] = 1'b1;  wr_cycle[ 5782] = 1'b0;  addr_rom[ 5782]='h00000c38;  wr_data_rom[ 5782]='h00000000;
    rd_cycle[ 5783] = 1'b1;  wr_cycle[ 5783] = 1'b0;  addr_rom[ 5783]='h00000c3c;  wr_data_rom[ 5783]='h00000000;
    rd_cycle[ 5784] = 1'b1;  wr_cycle[ 5784] = 1'b0;  addr_rom[ 5784]='h00000c40;  wr_data_rom[ 5784]='h00000000;
    rd_cycle[ 5785] = 1'b1;  wr_cycle[ 5785] = 1'b0;  addr_rom[ 5785]='h00000c44;  wr_data_rom[ 5785]='h00000000;
    rd_cycle[ 5786] = 1'b1;  wr_cycle[ 5786] = 1'b0;  addr_rom[ 5786]='h00000c48;  wr_data_rom[ 5786]='h00000000;
    rd_cycle[ 5787] = 1'b1;  wr_cycle[ 5787] = 1'b0;  addr_rom[ 5787]='h00000c4c;  wr_data_rom[ 5787]='h00000000;
    rd_cycle[ 5788] = 1'b1;  wr_cycle[ 5788] = 1'b0;  addr_rom[ 5788]='h00000c50;  wr_data_rom[ 5788]='h00000000;
    rd_cycle[ 5789] = 1'b1;  wr_cycle[ 5789] = 1'b0;  addr_rom[ 5789]='h00000c54;  wr_data_rom[ 5789]='h00000000;
    rd_cycle[ 5790] = 1'b1;  wr_cycle[ 5790] = 1'b0;  addr_rom[ 5790]='h00000c58;  wr_data_rom[ 5790]='h00000000;
    rd_cycle[ 5791] = 1'b1;  wr_cycle[ 5791] = 1'b0;  addr_rom[ 5791]='h00000c5c;  wr_data_rom[ 5791]='h00000000;
    rd_cycle[ 5792] = 1'b1;  wr_cycle[ 5792] = 1'b0;  addr_rom[ 5792]='h00000c60;  wr_data_rom[ 5792]='h00000000;
    rd_cycle[ 5793] = 1'b1;  wr_cycle[ 5793] = 1'b0;  addr_rom[ 5793]='h00000c64;  wr_data_rom[ 5793]='h00000000;
    rd_cycle[ 5794] = 1'b1;  wr_cycle[ 5794] = 1'b0;  addr_rom[ 5794]='h00000c68;  wr_data_rom[ 5794]='h00000000;
    rd_cycle[ 5795] = 1'b1;  wr_cycle[ 5795] = 1'b0;  addr_rom[ 5795]='h00000c6c;  wr_data_rom[ 5795]='h00000000;
    rd_cycle[ 5796] = 1'b1;  wr_cycle[ 5796] = 1'b0;  addr_rom[ 5796]='h00000c70;  wr_data_rom[ 5796]='h00000000;
    rd_cycle[ 5797] = 1'b1;  wr_cycle[ 5797] = 1'b0;  addr_rom[ 5797]='h00000c74;  wr_data_rom[ 5797]='h00000000;
    rd_cycle[ 5798] = 1'b1;  wr_cycle[ 5798] = 1'b0;  addr_rom[ 5798]='h00000c78;  wr_data_rom[ 5798]='h00000000;
    rd_cycle[ 5799] = 1'b1;  wr_cycle[ 5799] = 1'b0;  addr_rom[ 5799]='h00000c7c;  wr_data_rom[ 5799]='h00000000;
    rd_cycle[ 5800] = 1'b1;  wr_cycle[ 5800] = 1'b0;  addr_rom[ 5800]='h00000c80;  wr_data_rom[ 5800]='h00000000;
    rd_cycle[ 5801] = 1'b1;  wr_cycle[ 5801] = 1'b0;  addr_rom[ 5801]='h00000c84;  wr_data_rom[ 5801]='h00000000;
    rd_cycle[ 5802] = 1'b1;  wr_cycle[ 5802] = 1'b0;  addr_rom[ 5802]='h00000c88;  wr_data_rom[ 5802]='h00000000;
    rd_cycle[ 5803] = 1'b1;  wr_cycle[ 5803] = 1'b0;  addr_rom[ 5803]='h00000c8c;  wr_data_rom[ 5803]='h00000000;
    rd_cycle[ 5804] = 1'b1;  wr_cycle[ 5804] = 1'b0;  addr_rom[ 5804]='h00000c90;  wr_data_rom[ 5804]='h00000000;
    rd_cycle[ 5805] = 1'b1;  wr_cycle[ 5805] = 1'b0;  addr_rom[ 5805]='h00000c94;  wr_data_rom[ 5805]='h00000000;
    rd_cycle[ 5806] = 1'b1;  wr_cycle[ 5806] = 1'b0;  addr_rom[ 5806]='h00000c98;  wr_data_rom[ 5806]='h00000000;
    rd_cycle[ 5807] = 1'b1;  wr_cycle[ 5807] = 1'b0;  addr_rom[ 5807]='h00000c9c;  wr_data_rom[ 5807]='h00000000;
    rd_cycle[ 5808] = 1'b1;  wr_cycle[ 5808] = 1'b0;  addr_rom[ 5808]='h00000ca0;  wr_data_rom[ 5808]='h00000000;
    rd_cycle[ 5809] = 1'b1;  wr_cycle[ 5809] = 1'b0;  addr_rom[ 5809]='h00000ca4;  wr_data_rom[ 5809]='h00000000;
    rd_cycle[ 5810] = 1'b1;  wr_cycle[ 5810] = 1'b0;  addr_rom[ 5810]='h00000ca8;  wr_data_rom[ 5810]='h00000000;
    rd_cycle[ 5811] = 1'b1;  wr_cycle[ 5811] = 1'b0;  addr_rom[ 5811]='h00000cac;  wr_data_rom[ 5811]='h00000000;
    rd_cycle[ 5812] = 1'b1;  wr_cycle[ 5812] = 1'b0;  addr_rom[ 5812]='h00000cb0;  wr_data_rom[ 5812]='h00000000;
    rd_cycle[ 5813] = 1'b1;  wr_cycle[ 5813] = 1'b0;  addr_rom[ 5813]='h00000cb4;  wr_data_rom[ 5813]='h00000000;
    rd_cycle[ 5814] = 1'b1;  wr_cycle[ 5814] = 1'b0;  addr_rom[ 5814]='h00000cb8;  wr_data_rom[ 5814]='h00000000;
    rd_cycle[ 5815] = 1'b1;  wr_cycle[ 5815] = 1'b0;  addr_rom[ 5815]='h00000cbc;  wr_data_rom[ 5815]='h00000000;
    rd_cycle[ 5816] = 1'b1;  wr_cycle[ 5816] = 1'b0;  addr_rom[ 5816]='h00000cc0;  wr_data_rom[ 5816]='h00000000;
    rd_cycle[ 5817] = 1'b1;  wr_cycle[ 5817] = 1'b0;  addr_rom[ 5817]='h00000cc4;  wr_data_rom[ 5817]='h00000000;
    rd_cycle[ 5818] = 1'b1;  wr_cycle[ 5818] = 1'b0;  addr_rom[ 5818]='h00000cc8;  wr_data_rom[ 5818]='h00000000;
    rd_cycle[ 5819] = 1'b1;  wr_cycle[ 5819] = 1'b0;  addr_rom[ 5819]='h00000ccc;  wr_data_rom[ 5819]='h00000000;
    rd_cycle[ 5820] = 1'b1;  wr_cycle[ 5820] = 1'b0;  addr_rom[ 5820]='h00000cd0;  wr_data_rom[ 5820]='h00000000;
    rd_cycle[ 5821] = 1'b1;  wr_cycle[ 5821] = 1'b0;  addr_rom[ 5821]='h00000cd4;  wr_data_rom[ 5821]='h00000000;
    rd_cycle[ 5822] = 1'b1;  wr_cycle[ 5822] = 1'b0;  addr_rom[ 5822]='h00000cd8;  wr_data_rom[ 5822]='h00000000;
    rd_cycle[ 5823] = 1'b1;  wr_cycle[ 5823] = 1'b0;  addr_rom[ 5823]='h00000cdc;  wr_data_rom[ 5823]='h00000000;
    rd_cycle[ 5824] = 1'b1;  wr_cycle[ 5824] = 1'b0;  addr_rom[ 5824]='h00000ce0;  wr_data_rom[ 5824]='h00000000;
    rd_cycle[ 5825] = 1'b1;  wr_cycle[ 5825] = 1'b0;  addr_rom[ 5825]='h00000ce4;  wr_data_rom[ 5825]='h00000000;
    rd_cycle[ 5826] = 1'b1;  wr_cycle[ 5826] = 1'b0;  addr_rom[ 5826]='h00000ce8;  wr_data_rom[ 5826]='h00000000;
    rd_cycle[ 5827] = 1'b1;  wr_cycle[ 5827] = 1'b0;  addr_rom[ 5827]='h00000cec;  wr_data_rom[ 5827]='h00000000;
    rd_cycle[ 5828] = 1'b1;  wr_cycle[ 5828] = 1'b0;  addr_rom[ 5828]='h00000cf0;  wr_data_rom[ 5828]='h00000000;
    rd_cycle[ 5829] = 1'b1;  wr_cycle[ 5829] = 1'b0;  addr_rom[ 5829]='h00000cf4;  wr_data_rom[ 5829]='h00000000;
    rd_cycle[ 5830] = 1'b1;  wr_cycle[ 5830] = 1'b0;  addr_rom[ 5830]='h00000cf8;  wr_data_rom[ 5830]='h00000000;
    rd_cycle[ 5831] = 1'b1;  wr_cycle[ 5831] = 1'b0;  addr_rom[ 5831]='h00000cfc;  wr_data_rom[ 5831]='h00000000;
    rd_cycle[ 5832] = 1'b1;  wr_cycle[ 5832] = 1'b0;  addr_rom[ 5832]='h00000d00;  wr_data_rom[ 5832]='h00000000;
    rd_cycle[ 5833] = 1'b1;  wr_cycle[ 5833] = 1'b0;  addr_rom[ 5833]='h00000d04;  wr_data_rom[ 5833]='h00000000;
    rd_cycle[ 5834] = 1'b1;  wr_cycle[ 5834] = 1'b0;  addr_rom[ 5834]='h00000d08;  wr_data_rom[ 5834]='h00000000;
    rd_cycle[ 5835] = 1'b1;  wr_cycle[ 5835] = 1'b0;  addr_rom[ 5835]='h00000d0c;  wr_data_rom[ 5835]='h00000000;
    rd_cycle[ 5836] = 1'b1;  wr_cycle[ 5836] = 1'b0;  addr_rom[ 5836]='h00000d10;  wr_data_rom[ 5836]='h00000000;
    rd_cycle[ 5837] = 1'b1;  wr_cycle[ 5837] = 1'b0;  addr_rom[ 5837]='h00000d14;  wr_data_rom[ 5837]='h00000000;
    rd_cycle[ 5838] = 1'b1;  wr_cycle[ 5838] = 1'b0;  addr_rom[ 5838]='h00000d18;  wr_data_rom[ 5838]='h00000000;
    rd_cycle[ 5839] = 1'b1;  wr_cycle[ 5839] = 1'b0;  addr_rom[ 5839]='h00000d1c;  wr_data_rom[ 5839]='h00000000;
    rd_cycle[ 5840] = 1'b1;  wr_cycle[ 5840] = 1'b0;  addr_rom[ 5840]='h00000d20;  wr_data_rom[ 5840]='h00000000;
    rd_cycle[ 5841] = 1'b1;  wr_cycle[ 5841] = 1'b0;  addr_rom[ 5841]='h00000d24;  wr_data_rom[ 5841]='h00000000;
    rd_cycle[ 5842] = 1'b1;  wr_cycle[ 5842] = 1'b0;  addr_rom[ 5842]='h00000d28;  wr_data_rom[ 5842]='h00000000;
    rd_cycle[ 5843] = 1'b1;  wr_cycle[ 5843] = 1'b0;  addr_rom[ 5843]='h00000d2c;  wr_data_rom[ 5843]='h00000000;
    rd_cycle[ 5844] = 1'b1;  wr_cycle[ 5844] = 1'b0;  addr_rom[ 5844]='h00000d30;  wr_data_rom[ 5844]='h00000000;
    rd_cycle[ 5845] = 1'b1;  wr_cycle[ 5845] = 1'b0;  addr_rom[ 5845]='h00000d34;  wr_data_rom[ 5845]='h00000000;
    rd_cycle[ 5846] = 1'b1;  wr_cycle[ 5846] = 1'b0;  addr_rom[ 5846]='h00000d38;  wr_data_rom[ 5846]='h00000000;
    rd_cycle[ 5847] = 1'b1;  wr_cycle[ 5847] = 1'b0;  addr_rom[ 5847]='h00000d3c;  wr_data_rom[ 5847]='h00000000;
    rd_cycle[ 5848] = 1'b1;  wr_cycle[ 5848] = 1'b0;  addr_rom[ 5848]='h00000d40;  wr_data_rom[ 5848]='h00000000;
    rd_cycle[ 5849] = 1'b1;  wr_cycle[ 5849] = 1'b0;  addr_rom[ 5849]='h00000d44;  wr_data_rom[ 5849]='h00000000;
    rd_cycle[ 5850] = 1'b1;  wr_cycle[ 5850] = 1'b0;  addr_rom[ 5850]='h00000d48;  wr_data_rom[ 5850]='h00000000;
    rd_cycle[ 5851] = 1'b1;  wr_cycle[ 5851] = 1'b0;  addr_rom[ 5851]='h00000d4c;  wr_data_rom[ 5851]='h00000000;
    rd_cycle[ 5852] = 1'b1;  wr_cycle[ 5852] = 1'b0;  addr_rom[ 5852]='h00000d50;  wr_data_rom[ 5852]='h00000000;
    rd_cycle[ 5853] = 1'b1;  wr_cycle[ 5853] = 1'b0;  addr_rom[ 5853]='h00000d54;  wr_data_rom[ 5853]='h00000000;
    rd_cycle[ 5854] = 1'b1;  wr_cycle[ 5854] = 1'b0;  addr_rom[ 5854]='h00000d58;  wr_data_rom[ 5854]='h00000000;
    rd_cycle[ 5855] = 1'b1;  wr_cycle[ 5855] = 1'b0;  addr_rom[ 5855]='h00000d5c;  wr_data_rom[ 5855]='h00000000;
    rd_cycle[ 5856] = 1'b1;  wr_cycle[ 5856] = 1'b0;  addr_rom[ 5856]='h00000d60;  wr_data_rom[ 5856]='h00000000;
    rd_cycle[ 5857] = 1'b1;  wr_cycle[ 5857] = 1'b0;  addr_rom[ 5857]='h00000d64;  wr_data_rom[ 5857]='h00000000;
    rd_cycle[ 5858] = 1'b1;  wr_cycle[ 5858] = 1'b0;  addr_rom[ 5858]='h00000d68;  wr_data_rom[ 5858]='h00000000;
    rd_cycle[ 5859] = 1'b1;  wr_cycle[ 5859] = 1'b0;  addr_rom[ 5859]='h00000d6c;  wr_data_rom[ 5859]='h00000000;
    rd_cycle[ 5860] = 1'b1;  wr_cycle[ 5860] = 1'b0;  addr_rom[ 5860]='h00000d70;  wr_data_rom[ 5860]='h00000000;
    rd_cycle[ 5861] = 1'b1;  wr_cycle[ 5861] = 1'b0;  addr_rom[ 5861]='h00000d74;  wr_data_rom[ 5861]='h00000000;
    rd_cycle[ 5862] = 1'b1;  wr_cycle[ 5862] = 1'b0;  addr_rom[ 5862]='h00000d78;  wr_data_rom[ 5862]='h00000000;
    rd_cycle[ 5863] = 1'b1;  wr_cycle[ 5863] = 1'b0;  addr_rom[ 5863]='h00000d7c;  wr_data_rom[ 5863]='h00000000;
    rd_cycle[ 5864] = 1'b1;  wr_cycle[ 5864] = 1'b0;  addr_rom[ 5864]='h00000d80;  wr_data_rom[ 5864]='h00000000;
    rd_cycle[ 5865] = 1'b1;  wr_cycle[ 5865] = 1'b0;  addr_rom[ 5865]='h00000d84;  wr_data_rom[ 5865]='h00000000;
    rd_cycle[ 5866] = 1'b1;  wr_cycle[ 5866] = 1'b0;  addr_rom[ 5866]='h00000d88;  wr_data_rom[ 5866]='h00000000;
    rd_cycle[ 5867] = 1'b1;  wr_cycle[ 5867] = 1'b0;  addr_rom[ 5867]='h00000d8c;  wr_data_rom[ 5867]='h00000000;
    rd_cycle[ 5868] = 1'b1;  wr_cycle[ 5868] = 1'b0;  addr_rom[ 5868]='h00000d90;  wr_data_rom[ 5868]='h00000000;
    rd_cycle[ 5869] = 1'b1;  wr_cycle[ 5869] = 1'b0;  addr_rom[ 5869]='h00000d94;  wr_data_rom[ 5869]='h00000000;
    rd_cycle[ 5870] = 1'b1;  wr_cycle[ 5870] = 1'b0;  addr_rom[ 5870]='h00000d98;  wr_data_rom[ 5870]='h00000000;
    rd_cycle[ 5871] = 1'b1;  wr_cycle[ 5871] = 1'b0;  addr_rom[ 5871]='h00000d9c;  wr_data_rom[ 5871]='h00000000;
    rd_cycle[ 5872] = 1'b1;  wr_cycle[ 5872] = 1'b0;  addr_rom[ 5872]='h00000da0;  wr_data_rom[ 5872]='h00000000;
    rd_cycle[ 5873] = 1'b1;  wr_cycle[ 5873] = 1'b0;  addr_rom[ 5873]='h00000da4;  wr_data_rom[ 5873]='h00000000;
    rd_cycle[ 5874] = 1'b1;  wr_cycle[ 5874] = 1'b0;  addr_rom[ 5874]='h00000da8;  wr_data_rom[ 5874]='h00000000;
    rd_cycle[ 5875] = 1'b1;  wr_cycle[ 5875] = 1'b0;  addr_rom[ 5875]='h00000dac;  wr_data_rom[ 5875]='h00000000;
    rd_cycle[ 5876] = 1'b1;  wr_cycle[ 5876] = 1'b0;  addr_rom[ 5876]='h00000db0;  wr_data_rom[ 5876]='h00000000;
    rd_cycle[ 5877] = 1'b1;  wr_cycle[ 5877] = 1'b0;  addr_rom[ 5877]='h00000db4;  wr_data_rom[ 5877]='h00000000;
    rd_cycle[ 5878] = 1'b1;  wr_cycle[ 5878] = 1'b0;  addr_rom[ 5878]='h00000db8;  wr_data_rom[ 5878]='h00000000;
    rd_cycle[ 5879] = 1'b1;  wr_cycle[ 5879] = 1'b0;  addr_rom[ 5879]='h00000dbc;  wr_data_rom[ 5879]='h00000000;
    rd_cycle[ 5880] = 1'b1;  wr_cycle[ 5880] = 1'b0;  addr_rom[ 5880]='h00000dc0;  wr_data_rom[ 5880]='h00000000;
    rd_cycle[ 5881] = 1'b1;  wr_cycle[ 5881] = 1'b0;  addr_rom[ 5881]='h00000dc4;  wr_data_rom[ 5881]='h00000000;
    rd_cycle[ 5882] = 1'b1;  wr_cycle[ 5882] = 1'b0;  addr_rom[ 5882]='h00000dc8;  wr_data_rom[ 5882]='h00000000;
    rd_cycle[ 5883] = 1'b1;  wr_cycle[ 5883] = 1'b0;  addr_rom[ 5883]='h00000dcc;  wr_data_rom[ 5883]='h00000000;
    rd_cycle[ 5884] = 1'b1;  wr_cycle[ 5884] = 1'b0;  addr_rom[ 5884]='h00000dd0;  wr_data_rom[ 5884]='h00000000;
    rd_cycle[ 5885] = 1'b1;  wr_cycle[ 5885] = 1'b0;  addr_rom[ 5885]='h00000dd4;  wr_data_rom[ 5885]='h00000000;
    rd_cycle[ 5886] = 1'b1;  wr_cycle[ 5886] = 1'b0;  addr_rom[ 5886]='h00000dd8;  wr_data_rom[ 5886]='h00000000;
    rd_cycle[ 5887] = 1'b1;  wr_cycle[ 5887] = 1'b0;  addr_rom[ 5887]='h00000ddc;  wr_data_rom[ 5887]='h00000000;
    rd_cycle[ 5888] = 1'b1;  wr_cycle[ 5888] = 1'b0;  addr_rom[ 5888]='h00000de0;  wr_data_rom[ 5888]='h00000000;
    rd_cycle[ 5889] = 1'b1;  wr_cycle[ 5889] = 1'b0;  addr_rom[ 5889]='h00000de4;  wr_data_rom[ 5889]='h00000000;
    rd_cycle[ 5890] = 1'b1;  wr_cycle[ 5890] = 1'b0;  addr_rom[ 5890]='h00000de8;  wr_data_rom[ 5890]='h00000000;
    rd_cycle[ 5891] = 1'b1;  wr_cycle[ 5891] = 1'b0;  addr_rom[ 5891]='h00000dec;  wr_data_rom[ 5891]='h00000000;
    rd_cycle[ 5892] = 1'b1;  wr_cycle[ 5892] = 1'b0;  addr_rom[ 5892]='h00000df0;  wr_data_rom[ 5892]='h00000000;
    rd_cycle[ 5893] = 1'b1;  wr_cycle[ 5893] = 1'b0;  addr_rom[ 5893]='h00000df4;  wr_data_rom[ 5893]='h00000000;
    rd_cycle[ 5894] = 1'b1;  wr_cycle[ 5894] = 1'b0;  addr_rom[ 5894]='h00000df8;  wr_data_rom[ 5894]='h00000000;
    rd_cycle[ 5895] = 1'b1;  wr_cycle[ 5895] = 1'b0;  addr_rom[ 5895]='h00000dfc;  wr_data_rom[ 5895]='h00000000;
    rd_cycle[ 5896] = 1'b1;  wr_cycle[ 5896] = 1'b0;  addr_rom[ 5896]='h00000e00;  wr_data_rom[ 5896]='h00000000;
    rd_cycle[ 5897] = 1'b1;  wr_cycle[ 5897] = 1'b0;  addr_rom[ 5897]='h00000e04;  wr_data_rom[ 5897]='h00000000;
    rd_cycle[ 5898] = 1'b1;  wr_cycle[ 5898] = 1'b0;  addr_rom[ 5898]='h00000e08;  wr_data_rom[ 5898]='h00000000;
    rd_cycle[ 5899] = 1'b1;  wr_cycle[ 5899] = 1'b0;  addr_rom[ 5899]='h00000e0c;  wr_data_rom[ 5899]='h00000000;
    rd_cycle[ 5900] = 1'b1;  wr_cycle[ 5900] = 1'b0;  addr_rom[ 5900]='h00000e10;  wr_data_rom[ 5900]='h00000000;
    rd_cycle[ 5901] = 1'b1;  wr_cycle[ 5901] = 1'b0;  addr_rom[ 5901]='h00000e14;  wr_data_rom[ 5901]='h00000000;
    rd_cycle[ 5902] = 1'b1;  wr_cycle[ 5902] = 1'b0;  addr_rom[ 5902]='h00000e18;  wr_data_rom[ 5902]='h00000000;
    rd_cycle[ 5903] = 1'b1;  wr_cycle[ 5903] = 1'b0;  addr_rom[ 5903]='h00000e1c;  wr_data_rom[ 5903]='h00000000;
    rd_cycle[ 5904] = 1'b1;  wr_cycle[ 5904] = 1'b0;  addr_rom[ 5904]='h00000e20;  wr_data_rom[ 5904]='h00000000;
    rd_cycle[ 5905] = 1'b1;  wr_cycle[ 5905] = 1'b0;  addr_rom[ 5905]='h00000e24;  wr_data_rom[ 5905]='h00000000;
    rd_cycle[ 5906] = 1'b1;  wr_cycle[ 5906] = 1'b0;  addr_rom[ 5906]='h00000e28;  wr_data_rom[ 5906]='h00000000;
    rd_cycle[ 5907] = 1'b1;  wr_cycle[ 5907] = 1'b0;  addr_rom[ 5907]='h00000e2c;  wr_data_rom[ 5907]='h00000000;
    rd_cycle[ 5908] = 1'b1;  wr_cycle[ 5908] = 1'b0;  addr_rom[ 5908]='h00000e30;  wr_data_rom[ 5908]='h00000000;
    rd_cycle[ 5909] = 1'b1;  wr_cycle[ 5909] = 1'b0;  addr_rom[ 5909]='h00000e34;  wr_data_rom[ 5909]='h00000000;
    rd_cycle[ 5910] = 1'b1;  wr_cycle[ 5910] = 1'b0;  addr_rom[ 5910]='h00000e38;  wr_data_rom[ 5910]='h00000000;
    rd_cycle[ 5911] = 1'b1;  wr_cycle[ 5911] = 1'b0;  addr_rom[ 5911]='h00000e3c;  wr_data_rom[ 5911]='h00000000;
    rd_cycle[ 5912] = 1'b1;  wr_cycle[ 5912] = 1'b0;  addr_rom[ 5912]='h00000e40;  wr_data_rom[ 5912]='h00000000;
    rd_cycle[ 5913] = 1'b1;  wr_cycle[ 5913] = 1'b0;  addr_rom[ 5913]='h00000e44;  wr_data_rom[ 5913]='h00000000;
    rd_cycle[ 5914] = 1'b1;  wr_cycle[ 5914] = 1'b0;  addr_rom[ 5914]='h00000e48;  wr_data_rom[ 5914]='h00000000;
    rd_cycle[ 5915] = 1'b1;  wr_cycle[ 5915] = 1'b0;  addr_rom[ 5915]='h00000e4c;  wr_data_rom[ 5915]='h00000000;
    rd_cycle[ 5916] = 1'b1;  wr_cycle[ 5916] = 1'b0;  addr_rom[ 5916]='h00000e50;  wr_data_rom[ 5916]='h00000000;
    rd_cycle[ 5917] = 1'b1;  wr_cycle[ 5917] = 1'b0;  addr_rom[ 5917]='h00000e54;  wr_data_rom[ 5917]='h00000000;
    rd_cycle[ 5918] = 1'b1;  wr_cycle[ 5918] = 1'b0;  addr_rom[ 5918]='h00000e58;  wr_data_rom[ 5918]='h00000000;
    rd_cycle[ 5919] = 1'b1;  wr_cycle[ 5919] = 1'b0;  addr_rom[ 5919]='h00000e5c;  wr_data_rom[ 5919]='h00000000;
    rd_cycle[ 5920] = 1'b1;  wr_cycle[ 5920] = 1'b0;  addr_rom[ 5920]='h00000e60;  wr_data_rom[ 5920]='h00000000;
    rd_cycle[ 5921] = 1'b1;  wr_cycle[ 5921] = 1'b0;  addr_rom[ 5921]='h00000e64;  wr_data_rom[ 5921]='h00000000;
    rd_cycle[ 5922] = 1'b1;  wr_cycle[ 5922] = 1'b0;  addr_rom[ 5922]='h00000e68;  wr_data_rom[ 5922]='h00000000;
    rd_cycle[ 5923] = 1'b1;  wr_cycle[ 5923] = 1'b0;  addr_rom[ 5923]='h00000e6c;  wr_data_rom[ 5923]='h00000000;
    rd_cycle[ 5924] = 1'b1;  wr_cycle[ 5924] = 1'b0;  addr_rom[ 5924]='h00000e70;  wr_data_rom[ 5924]='h00000000;
    rd_cycle[ 5925] = 1'b1;  wr_cycle[ 5925] = 1'b0;  addr_rom[ 5925]='h00000e74;  wr_data_rom[ 5925]='h00000000;
    rd_cycle[ 5926] = 1'b1;  wr_cycle[ 5926] = 1'b0;  addr_rom[ 5926]='h00000e78;  wr_data_rom[ 5926]='h00000000;
    rd_cycle[ 5927] = 1'b1;  wr_cycle[ 5927] = 1'b0;  addr_rom[ 5927]='h00000e7c;  wr_data_rom[ 5927]='h00000000;
    rd_cycle[ 5928] = 1'b1;  wr_cycle[ 5928] = 1'b0;  addr_rom[ 5928]='h00000e80;  wr_data_rom[ 5928]='h00000000;
    rd_cycle[ 5929] = 1'b1;  wr_cycle[ 5929] = 1'b0;  addr_rom[ 5929]='h00000e84;  wr_data_rom[ 5929]='h00000000;
    rd_cycle[ 5930] = 1'b1;  wr_cycle[ 5930] = 1'b0;  addr_rom[ 5930]='h00000e88;  wr_data_rom[ 5930]='h00000000;
    rd_cycle[ 5931] = 1'b1;  wr_cycle[ 5931] = 1'b0;  addr_rom[ 5931]='h00000e8c;  wr_data_rom[ 5931]='h00000000;
    rd_cycle[ 5932] = 1'b1;  wr_cycle[ 5932] = 1'b0;  addr_rom[ 5932]='h00000e90;  wr_data_rom[ 5932]='h00000000;
    rd_cycle[ 5933] = 1'b1;  wr_cycle[ 5933] = 1'b0;  addr_rom[ 5933]='h00000e94;  wr_data_rom[ 5933]='h00000000;
    rd_cycle[ 5934] = 1'b1;  wr_cycle[ 5934] = 1'b0;  addr_rom[ 5934]='h00000e98;  wr_data_rom[ 5934]='h00000000;
    rd_cycle[ 5935] = 1'b1;  wr_cycle[ 5935] = 1'b0;  addr_rom[ 5935]='h00000e9c;  wr_data_rom[ 5935]='h00000000;
    rd_cycle[ 5936] = 1'b1;  wr_cycle[ 5936] = 1'b0;  addr_rom[ 5936]='h00000ea0;  wr_data_rom[ 5936]='h00000000;
    rd_cycle[ 5937] = 1'b1;  wr_cycle[ 5937] = 1'b0;  addr_rom[ 5937]='h00000ea4;  wr_data_rom[ 5937]='h00000000;
    rd_cycle[ 5938] = 1'b1;  wr_cycle[ 5938] = 1'b0;  addr_rom[ 5938]='h00000ea8;  wr_data_rom[ 5938]='h00000000;
    rd_cycle[ 5939] = 1'b1;  wr_cycle[ 5939] = 1'b0;  addr_rom[ 5939]='h00000eac;  wr_data_rom[ 5939]='h00000000;
    rd_cycle[ 5940] = 1'b1;  wr_cycle[ 5940] = 1'b0;  addr_rom[ 5940]='h00000eb0;  wr_data_rom[ 5940]='h00000000;
    rd_cycle[ 5941] = 1'b1;  wr_cycle[ 5941] = 1'b0;  addr_rom[ 5941]='h00000eb4;  wr_data_rom[ 5941]='h00000000;
    rd_cycle[ 5942] = 1'b1;  wr_cycle[ 5942] = 1'b0;  addr_rom[ 5942]='h00000eb8;  wr_data_rom[ 5942]='h00000000;
    rd_cycle[ 5943] = 1'b1;  wr_cycle[ 5943] = 1'b0;  addr_rom[ 5943]='h00000ebc;  wr_data_rom[ 5943]='h00000000;
    rd_cycle[ 5944] = 1'b1;  wr_cycle[ 5944] = 1'b0;  addr_rom[ 5944]='h00000ec0;  wr_data_rom[ 5944]='h00000000;
    rd_cycle[ 5945] = 1'b1;  wr_cycle[ 5945] = 1'b0;  addr_rom[ 5945]='h00000ec4;  wr_data_rom[ 5945]='h00000000;
    rd_cycle[ 5946] = 1'b1;  wr_cycle[ 5946] = 1'b0;  addr_rom[ 5946]='h00000ec8;  wr_data_rom[ 5946]='h00000000;
    rd_cycle[ 5947] = 1'b1;  wr_cycle[ 5947] = 1'b0;  addr_rom[ 5947]='h00000ecc;  wr_data_rom[ 5947]='h00000000;
    rd_cycle[ 5948] = 1'b1;  wr_cycle[ 5948] = 1'b0;  addr_rom[ 5948]='h00000ed0;  wr_data_rom[ 5948]='h00000000;
    rd_cycle[ 5949] = 1'b1;  wr_cycle[ 5949] = 1'b0;  addr_rom[ 5949]='h00000ed4;  wr_data_rom[ 5949]='h00000000;
    rd_cycle[ 5950] = 1'b1;  wr_cycle[ 5950] = 1'b0;  addr_rom[ 5950]='h00000ed8;  wr_data_rom[ 5950]='h00000000;
    rd_cycle[ 5951] = 1'b1;  wr_cycle[ 5951] = 1'b0;  addr_rom[ 5951]='h00000edc;  wr_data_rom[ 5951]='h00000000;
    rd_cycle[ 5952] = 1'b1;  wr_cycle[ 5952] = 1'b0;  addr_rom[ 5952]='h00000ee0;  wr_data_rom[ 5952]='h00000000;
    rd_cycle[ 5953] = 1'b1;  wr_cycle[ 5953] = 1'b0;  addr_rom[ 5953]='h00000ee4;  wr_data_rom[ 5953]='h00000000;
    rd_cycle[ 5954] = 1'b1;  wr_cycle[ 5954] = 1'b0;  addr_rom[ 5954]='h00000ee8;  wr_data_rom[ 5954]='h00000000;
    rd_cycle[ 5955] = 1'b1;  wr_cycle[ 5955] = 1'b0;  addr_rom[ 5955]='h00000eec;  wr_data_rom[ 5955]='h00000000;
    rd_cycle[ 5956] = 1'b1;  wr_cycle[ 5956] = 1'b0;  addr_rom[ 5956]='h00000ef0;  wr_data_rom[ 5956]='h00000000;
    rd_cycle[ 5957] = 1'b1;  wr_cycle[ 5957] = 1'b0;  addr_rom[ 5957]='h00000ef4;  wr_data_rom[ 5957]='h00000000;
    rd_cycle[ 5958] = 1'b1;  wr_cycle[ 5958] = 1'b0;  addr_rom[ 5958]='h00000ef8;  wr_data_rom[ 5958]='h00000000;
    rd_cycle[ 5959] = 1'b1;  wr_cycle[ 5959] = 1'b0;  addr_rom[ 5959]='h00000efc;  wr_data_rom[ 5959]='h00000000;
    rd_cycle[ 5960] = 1'b1;  wr_cycle[ 5960] = 1'b0;  addr_rom[ 5960]='h00000f00;  wr_data_rom[ 5960]='h00000000;
    rd_cycle[ 5961] = 1'b1;  wr_cycle[ 5961] = 1'b0;  addr_rom[ 5961]='h00000f04;  wr_data_rom[ 5961]='h00000000;
    rd_cycle[ 5962] = 1'b1;  wr_cycle[ 5962] = 1'b0;  addr_rom[ 5962]='h00000f08;  wr_data_rom[ 5962]='h00000000;
    rd_cycle[ 5963] = 1'b1;  wr_cycle[ 5963] = 1'b0;  addr_rom[ 5963]='h00000f0c;  wr_data_rom[ 5963]='h00000000;
    rd_cycle[ 5964] = 1'b1;  wr_cycle[ 5964] = 1'b0;  addr_rom[ 5964]='h00000f10;  wr_data_rom[ 5964]='h00000000;
    rd_cycle[ 5965] = 1'b1;  wr_cycle[ 5965] = 1'b0;  addr_rom[ 5965]='h00000f14;  wr_data_rom[ 5965]='h00000000;
    rd_cycle[ 5966] = 1'b1;  wr_cycle[ 5966] = 1'b0;  addr_rom[ 5966]='h00000f18;  wr_data_rom[ 5966]='h00000000;
    rd_cycle[ 5967] = 1'b1;  wr_cycle[ 5967] = 1'b0;  addr_rom[ 5967]='h00000f1c;  wr_data_rom[ 5967]='h00000000;
    rd_cycle[ 5968] = 1'b1;  wr_cycle[ 5968] = 1'b0;  addr_rom[ 5968]='h00000f20;  wr_data_rom[ 5968]='h00000000;
    rd_cycle[ 5969] = 1'b1;  wr_cycle[ 5969] = 1'b0;  addr_rom[ 5969]='h00000f24;  wr_data_rom[ 5969]='h00000000;
    rd_cycle[ 5970] = 1'b1;  wr_cycle[ 5970] = 1'b0;  addr_rom[ 5970]='h00000f28;  wr_data_rom[ 5970]='h00000000;
    rd_cycle[ 5971] = 1'b1;  wr_cycle[ 5971] = 1'b0;  addr_rom[ 5971]='h00000f2c;  wr_data_rom[ 5971]='h00000000;
    rd_cycle[ 5972] = 1'b1;  wr_cycle[ 5972] = 1'b0;  addr_rom[ 5972]='h00000f30;  wr_data_rom[ 5972]='h00000000;
    rd_cycle[ 5973] = 1'b1;  wr_cycle[ 5973] = 1'b0;  addr_rom[ 5973]='h00000f34;  wr_data_rom[ 5973]='h00000000;
    rd_cycle[ 5974] = 1'b1;  wr_cycle[ 5974] = 1'b0;  addr_rom[ 5974]='h00000f38;  wr_data_rom[ 5974]='h00000000;
    rd_cycle[ 5975] = 1'b1;  wr_cycle[ 5975] = 1'b0;  addr_rom[ 5975]='h00000f3c;  wr_data_rom[ 5975]='h00000000;
    rd_cycle[ 5976] = 1'b1;  wr_cycle[ 5976] = 1'b0;  addr_rom[ 5976]='h00000f40;  wr_data_rom[ 5976]='h00000000;
    rd_cycle[ 5977] = 1'b1;  wr_cycle[ 5977] = 1'b0;  addr_rom[ 5977]='h00000f44;  wr_data_rom[ 5977]='h00000000;
    rd_cycle[ 5978] = 1'b1;  wr_cycle[ 5978] = 1'b0;  addr_rom[ 5978]='h00000f48;  wr_data_rom[ 5978]='h00000000;
    rd_cycle[ 5979] = 1'b1;  wr_cycle[ 5979] = 1'b0;  addr_rom[ 5979]='h00000f4c;  wr_data_rom[ 5979]='h00000000;
    rd_cycle[ 5980] = 1'b1;  wr_cycle[ 5980] = 1'b0;  addr_rom[ 5980]='h00000f50;  wr_data_rom[ 5980]='h00000000;
    rd_cycle[ 5981] = 1'b1;  wr_cycle[ 5981] = 1'b0;  addr_rom[ 5981]='h00000f54;  wr_data_rom[ 5981]='h00000000;
    rd_cycle[ 5982] = 1'b1;  wr_cycle[ 5982] = 1'b0;  addr_rom[ 5982]='h00000f58;  wr_data_rom[ 5982]='h00000000;
    rd_cycle[ 5983] = 1'b1;  wr_cycle[ 5983] = 1'b0;  addr_rom[ 5983]='h00000f5c;  wr_data_rom[ 5983]='h00000000;
    rd_cycle[ 5984] = 1'b1;  wr_cycle[ 5984] = 1'b0;  addr_rom[ 5984]='h00000f60;  wr_data_rom[ 5984]='h00000000;
    rd_cycle[ 5985] = 1'b1;  wr_cycle[ 5985] = 1'b0;  addr_rom[ 5985]='h00000f64;  wr_data_rom[ 5985]='h00000000;
    rd_cycle[ 5986] = 1'b1;  wr_cycle[ 5986] = 1'b0;  addr_rom[ 5986]='h00000f68;  wr_data_rom[ 5986]='h00000000;
    rd_cycle[ 5987] = 1'b1;  wr_cycle[ 5987] = 1'b0;  addr_rom[ 5987]='h00000f6c;  wr_data_rom[ 5987]='h00000000;
    rd_cycle[ 5988] = 1'b1;  wr_cycle[ 5988] = 1'b0;  addr_rom[ 5988]='h00000f70;  wr_data_rom[ 5988]='h00000000;
    rd_cycle[ 5989] = 1'b1;  wr_cycle[ 5989] = 1'b0;  addr_rom[ 5989]='h00000f74;  wr_data_rom[ 5989]='h00000000;
    rd_cycle[ 5990] = 1'b1;  wr_cycle[ 5990] = 1'b0;  addr_rom[ 5990]='h00000f78;  wr_data_rom[ 5990]='h00000000;
    rd_cycle[ 5991] = 1'b1;  wr_cycle[ 5991] = 1'b0;  addr_rom[ 5991]='h00000f7c;  wr_data_rom[ 5991]='h00000000;
    rd_cycle[ 5992] = 1'b1;  wr_cycle[ 5992] = 1'b0;  addr_rom[ 5992]='h00000f80;  wr_data_rom[ 5992]='h00000000;
    rd_cycle[ 5993] = 1'b1;  wr_cycle[ 5993] = 1'b0;  addr_rom[ 5993]='h00000f84;  wr_data_rom[ 5993]='h00000000;
    rd_cycle[ 5994] = 1'b1;  wr_cycle[ 5994] = 1'b0;  addr_rom[ 5994]='h00000f88;  wr_data_rom[ 5994]='h00000000;
    rd_cycle[ 5995] = 1'b1;  wr_cycle[ 5995] = 1'b0;  addr_rom[ 5995]='h00000f8c;  wr_data_rom[ 5995]='h00000000;
    rd_cycle[ 5996] = 1'b1;  wr_cycle[ 5996] = 1'b0;  addr_rom[ 5996]='h00000f90;  wr_data_rom[ 5996]='h00000000;
    rd_cycle[ 5997] = 1'b1;  wr_cycle[ 5997] = 1'b0;  addr_rom[ 5997]='h00000f94;  wr_data_rom[ 5997]='h00000000;
    rd_cycle[ 5998] = 1'b1;  wr_cycle[ 5998] = 1'b0;  addr_rom[ 5998]='h00000f98;  wr_data_rom[ 5998]='h00000000;
    rd_cycle[ 5999] = 1'b1;  wr_cycle[ 5999] = 1'b0;  addr_rom[ 5999]='h00000f9c;  wr_data_rom[ 5999]='h00000000;
end

initial begin
    validation_data[    0] = 'h00000cc5; 
    validation_data[    1] = 'h00000421; 
    validation_data[    2] = 'h00000221; 
    validation_data[    3] = 'h00000a99; 
    validation_data[    4] = 'h00000030; 
    validation_data[    5] = 'h00000963; 
    validation_data[    6] = 'h000004e5; 
    validation_data[    7] = 'h000007c0; 
    validation_data[    8] = 'h00000503; 
    validation_data[    9] = 'h00000731; 
    validation_data[   10] = 'h0000090a; 
    validation_data[   11] = 'h00000b6e; 
    validation_data[   12] = 'h00000645; 
    validation_data[   13] = 'h0000088c; 
    validation_data[   14] = 'h00000a7e; 
    validation_data[   15] = 'h000008f5; 
    validation_data[   16] = 'h0000031f; 
    validation_data[   17] = 'h00000251; 
    validation_data[   18] = 'h00000c3b; 
    validation_data[   19] = 'h00000c1e; 
    validation_data[   20] = 'h00000d8a; 
    validation_data[   21] = 'h00000946; 
    validation_data[   22] = 'h00000d40; 
    validation_data[   23] = 'h00000e7a; 
    validation_data[   24] = 'h000004bf; 
    validation_data[   25] = 'h00000f34; 
    validation_data[   26] = 'h00000907; 
    validation_data[   27] = 'h0000011b; 
    validation_data[   28] = 'h000008ce; 
    validation_data[   29] = 'h000001c8; 
    validation_data[   30] = 'h000008f1; 
    validation_data[   31] = 'h00000f88; 
    validation_data[   32] = 'h00000ddc; 
    validation_data[   33] = 'h00000a22; 
    validation_data[   34] = 'h00000a79; 
    validation_data[   35] = 'h00000c68; 
    validation_data[   36] = 'h00000cca; 
    validation_data[   37] = 'h0000073d; 
    validation_data[   38] = 'h00000bb1; 
    validation_data[   39] = 'h00000e24; 
    validation_data[   40] = 'h00000241; 
    validation_data[   41] = 'h00000108; 
    validation_data[   42] = 'h00000257; 
    validation_data[   43] = 'h000009a3; 
    validation_data[   44] = 'h00000bdc; 
    validation_data[   45] = 'h000009bd; 
    validation_data[   46] = 'h000004b8; 
    validation_data[   47] = 'h000006d8; 
    validation_data[   48] = 'h000007a0; 
    validation_data[   49] = 'h00000472; 
    validation_data[   50] = 'h000006b6; 
    validation_data[   51] = 'h00000ddf; 
    validation_data[   52] = 'h00000607; 
    validation_data[   53] = 'h00000f70; 
    validation_data[   54] = 'h0000058b; 
    validation_data[   55] = 'h000006ce; 
    validation_data[   56] = 'h0000039e; 
    validation_data[   57] = 'h0000017f; 
    validation_data[   58] = 'h000000de; 
    validation_data[   59] = 'h00000b73; 
    validation_data[   60] = 'h00000126; 
    validation_data[   61] = 'h00000867; 
    validation_data[   62] = 'h0000086d; 
    validation_data[   63] = 'h000002c1; 
    validation_data[   64] = 'h00000ee8; 
    validation_data[   65] = 'h00000276; 
    validation_data[   66] = 'h00000f21; 
    validation_data[   67] = 'h00000bbb; 
    validation_data[   68] = 'h00000831; 
    validation_data[   69] = 'h000006d8; 
    validation_data[   70] = 'h00000e89; 
    validation_data[   71] = 'h00000e4b; 
    validation_data[   72] = 'h00000cd5; 
    validation_data[   73] = 'h000001a3; 
    validation_data[   74] = 'h00000cd7; 
    validation_data[   75] = 'h00000f99; 
    validation_data[   76] = 'h00000d00; 
    validation_data[   77] = 'h000000e1; 
    validation_data[   78] = 'h00000e15; 
    validation_data[   79] = 'h00000c17; 
    validation_data[   80] = 'h0000094c; 
    validation_data[   81] = 'h00000ed0; 
    validation_data[   82] = 'h00000e88; 
    validation_data[   83] = 'h00000267; 
    validation_data[   84] = 'h00000411; 
    validation_data[   85] = 'h00000aa9; 
    validation_data[   86] = 'h00000eb7; 
    validation_data[   87] = 'h0000031d; 
    validation_data[   88] = 'h00000c5e; 
    validation_data[   89] = 'h00000c7f; 
    validation_data[   90] = 'h000003a2; 
    validation_data[   91] = 'h00000358; 
    validation_data[   92] = 'h000009d8; 
    validation_data[   93] = 'h000005ac; 
    validation_data[   94] = 'h0000004f; 
    validation_data[   95] = 'h00000b42; 
    validation_data[   96] = 'h000001c8; 
    validation_data[   97] = 'h0000091f; 
    validation_data[   98] = 'h00000d4a; 
    validation_data[   99] = 'h000006ad; 
    validation_data[  100] = 'h000007b1; 
    validation_data[  101] = 'h0000062e; 
    validation_data[  102] = 'h0000071b; 
    validation_data[  103] = 'h00000b3f; 
    validation_data[  104] = 'h000003dd; 
    validation_data[  105] = 'h00000f3a; 
    validation_data[  106] = 'h00000203; 
    validation_data[  107] = 'h000008b7; 
    validation_data[  108] = 'h000008f5; 
    validation_data[  109] = 'h0000036e; 
    validation_data[  110] = 'h00000763; 
    validation_data[  111] = 'h0000028f; 
    validation_data[  112] = 'h000009ad; 
    validation_data[  113] = 'h00000611; 
    validation_data[  114] = 'h000008c2; 
    validation_data[  115] = 'h00000730; 
    validation_data[  116] = 'h000001ad; 
    validation_data[  117] = 'h000004b6; 
    validation_data[  118] = 'h0000028c; 
    validation_data[  119] = 'h00000628; 
    validation_data[  120] = 'h00000c8d; 
    validation_data[  121] = 'h000008f2; 
    validation_data[  122] = 'h00000a1e; 
    validation_data[  123] = 'h00000758; 
    validation_data[  124] = 'h00000ba3; 
    validation_data[  125] = 'h00000750; 
    validation_data[  126] = 'h00000ea5; 
    validation_data[  127] = 'h000003fc; 
    validation_data[  128] = 'h00000884; 
    validation_data[  129] = 'h0000082a; 
    validation_data[  130] = 'h00000ad3; 
    validation_data[  131] = 'h000007c8; 
    validation_data[  132] = 'h00000f81; 
    validation_data[  133] = 'h00000121; 
    validation_data[  134] = 'h00000476; 
    validation_data[  135] = 'h000005e5; 
    validation_data[  136] = 'h000009db; 
    validation_data[  137] = 'h000000d6; 
    validation_data[  138] = 'h00000749; 
    validation_data[  139] = 'h00000ef3; 
    validation_data[  140] = 'h00000c25; 
    validation_data[  141] = 'h00000158; 
    validation_data[  142] = 'h0000044e; 
    validation_data[  143] = 'h00000d23; 
    validation_data[  144] = 'h000008db; 
    validation_data[  145] = 'h0000085d; 
    validation_data[  146] = 'h00000c99; 
    validation_data[  147] = 'h00000f13; 
    validation_data[  148] = 'h000007e0; 
    validation_data[  149] = 'h00000057; 
    validation_data[  150] = 'h00000670; 
    validation_data[  151] = 'h00000376; 
    validation_data[  152] = 'h00000443; 
    validation_data[  153] = 'h00000e05; 
    validation_data[  154] = 'h000006df; 
    validation_data[  155] = 'h00000b54; 
    validation_data[  156] = 'h00000604; 
    validation_data[  157] = 'h000004d9; 
    validation_data[  158] = 'h000003d4; 
    validation_data[  159] = 'h00000f8a; 
    validation_data[  160] = 'h00000829; 
    validation_data[  161] = 'h00000ce3; 
    validation_data[  162] = 'h0000094c; 
    validation_data[  163] = 'h00000e7a; 
    validation_data[  164] = 'h00000157; 
    validation_data[  165] = 'h00000835; 
    validation_data[  166] = 'h00000926; 
    validation_data[  167] = 'h00000af4; 
    validation_data[  168] = 'h00000918; 
    validation_data[  169] = 'h000007e5; 
    validation_data[  170] = 'h000009ce; 
    validation_data[  171] = 'h00000a7a; 
    validation_data[  172] = 'h000009d9; 
    validation_data[  173] = 'h000007de; 
    validation_data[  174] = 'h00000bd3; 
    validation_data[  175] = 'h00000530; 
    validation_data[  176] = 'h000009b7; 
    validation_data[  177] = 'h00000ce5; 
    validation_data[  178] = 'h00000a50; 
    validation_data[  179] = 'h00000a4b; 
    validation_data[  180] = 'h00000056; 
    validation_data[  181] = 'h0000084d; 
    validation_data[  182] = 'h00000c56; 
    validation_data[  183] = 'h000002cf; 
    validation_data[  184] = 'h0000080e; 
    validation_data[  185] = 'h00000c79; 
    validation_data[  186] = 'h00000c71; 
    validation_data[  187] = 'h000007cf; 
    validation_data[  188] = 'h0000093b; 
    validation_data[  189] = 'h00000038; 
    validation_data[  190] = 'h00000609; 
    validation_data[  191] = 'h00000b83; 
    validation_data[  192] = 'h000001d1; 
    validation_data[  193] = 'h00000c6e; 
    validation_data[  194] = 'h00000217; 
    validation_data[  195] = 'h00000e3a; 
    validation_data[  196] = 'h00000b94; 
    validation_data[  197] = 'h0000065d; 
    validation_data[  198] = 'h00000359; 
    validation_data[  199] = 'h00000cdf; 
    validation_data[  200] = 'h00000f3f; 
    validation_data[  201] = 'h00000131; 
    validation_data[  202] = 'h00000338; 
    validation_data[  203] = 'h00000080; 
    validation_data[  204] = 'h0000051c; 
    validation_data[  205] = 'h000006e9; 
    validation_data[  206] = 'h00000133; 
    validation_data[  207] = 'h00000351; 
    validation_data[  208] = 'h000004a6; 
    validation_data[  209] = 'h0000027e; 
    validation_data[  210] = 'h00000992; 
    validation_data[  211] = 'h00000bf7; 
    validation_data[  212] = 'h00000307; 
    validation_data[  213] = 'h000003e8; 
    validation_data[  214] = 'h00000317; 
    validation_data[  215] = 'h000003c4; 
    validation_data[  216] = 'h00000d9d; 
    validation_data[  217] = 'h00000e56; 
    validation_data[  218] = 'h00000117; 
    validation_data[  219] = 'h00000719; 
    validation_data[  220] = 'h00000d32; 
    validation_data[  221] = 'h00000d7d; 
    validation_data[  222] = 'h00000195; 
    validation_data[  223] = 'h000003cc; 
    validation_data[  224] = 'h00000233; 
    validation_data[  225] = 'h00000212; 
    validation_data[  226] = 'h00000124; 
    validation_data[  227] = 'h00000b1f; 
    validation_data[  228] = 'h00000f63; 
    validation_data[  229] = 'h000007b2; 
    validation_data[  230] = 'h00000447; 
    validation_data[  231] = 'h00000b69; 
    validation_data[  232] = 'h000001df; 
    validation_data[  233] = 'h00000b7d; 
    validation_data[  234] = 'h00000d12; 
    validation_data[  235] = 'h00000b4a; 
    validation_data[  236] = 'h000007f6; 
    validation_data[  237] = 'h000008fc; 
    validation_data[  238] = 'h00000289; 
    validation_data[  239] = 'h00000080; 
    validation_data[  240] = 'h00000f33; 
    validation_data[  241] = 'h0000028d; 
    validation_data[  242] = 'h00000d2c; 
    validation_data[  243] = 'h000009f2; 
    validation_data[  244] = 'h00000df5; 
    validation_data[  245] = 'h000008b2; 
    validation_data[  246] = 'h00000e76; 
    validation_data[  247] = 'h00000653; 
    validation_data[  248] = 'h0000011c; 
    validation_data[  249] = 'h00000097; 
    validation_data[  250] = 'h00000660; 
    validation_data[  251] = 'h0000000e; 
    validation_data[  252] = 'h000005c0; 
    validation_data[  253] = 'h0000011d; 
    validation_data[  254] = 'h00000489; 
    validation_data[  255] = 'h00000431; 
    validation_data[  256] = 'h0000012e; 
    validation_data[  257] = 'h00000786; 
    validation_data[  258] = 'h00000614; 
    validation_data[  259] = 'h000006f8; 
    validation_data[  260] = 'h000000d9; 
    validation_data[  261] = 'h000005c3; 
    validation_data[  262] = 'h00000e48; 
    validation_data[  263] = 'h00000d52; 
    validation_data[  264] = 'h00000118; 
    validation_data[  265] = 'h000004a6; 
    validation_data[  266] = 'h00000766; 
    validation_data[  267] = 'h00000473; 
    validation_data[  268] = 'h00000d6c; 
    validation_data[  269] = 'h00000c13; 
    validation_data[  270] = 'h00000ab0; 
    validation_data[  271] = 'h00000e34; 
    validation_data[  272] = 'h000006be; 
    validation_data[  273] = 'h00000690; 
    validation_data[  274] = 'h0000055f; 
    validation_data[  275] = 'h00000017; 
    validation_data[  276] = 'h00000f31; 
    validation_data[  277] = 'h000001e2; 
    validation_data[  278] = 'h00000439; 
    validation_data[  279] = 'h000006c8; 
    validation_data[  280] = 'h00000c9b; 
    validation_data[  281] = 'h00000a93; 
    validation_data[  282] = 'h00000e5d; 
    validation_data[  283] = 'h00000549; 
    validation_data[  284] = 'h000000c0; 
    validation_data[  285] = 'h000000b6; 
    validation_data[  286] = 'h00000017; 
    validation_data[  287] = 'h000003c6; 
    validation_data[  288] = 'h000004da; 
    validation_data[  289] = 'h00000635; 
    validation_data[  290] = 'h0000077a; 
    validation_data[  291] = 'h00000973; 
    validation_data[  292] = 'h000006d5; 
    validation_data[  293] = 'h00000c15; 
    validation_data[  294] = 'h00000a12; 
    validation_data[  295] = 'h00000ad4; 
    validation_data[  296] = 'h00000b12; 
    validation_data[  297] = 'h0000065e; 
    validation_data[  298] = 'h00000620; 
    validation_data[  299] = 'h00000564; 
    validation_data[  300] = 'h00000b43; 
    validation_data[  301] = 'h00000457; 
    validation_data[  302] = 'h000001b1; 
    validation_data[  303] = 'h00000ae6; 
    validation_data[  304] = 'h00000cc0; 
    validation_data[  305] = 'h000005a1; 
    validation_data[  306] = 'h00000959; 
    validation_data[  307] = 'h0000068f; 
    validation_data[  308] = 'h000006bf; 
    validation_data[  309] = 'h00000563; 
    validation_data[  310] = 'h00000edf; 
    validation_data[  311] = 'h00000919; 
    validation_data[  312] = 'h000008fd; 
    validation_data[  313] = 'h00000f65; 
    validation_data[  314] = 'h0000000a; 
    validation_data[  315] = 'h000004b8; 
    validation_data[  316] = 'h00000637; 
    validation_data[  317] = 'h000003a0; 
    validation_data[  318] = 'h00000e2b; 
    validation_data[  319] = 'h00000f40; 
    validation_data[  320] = 'h00000123; 
    validation_data[  321] = 'h00000f2b; 
    validation_data[  322] = 'h0000025f; 
    validation_data[  323] = 'h00000e7b; 
    validation_data[  324] = 'h00000d9d; 
    validation_data[  325] = 'h00000d8e; 
    validation_data[  326] = 'h000005de; 
    validation_data[  327] = 'h000000c9; 
    validation_data[  328] = 'h00000903; 
    validation_data[  329] = 'h00000238; 
    validation_data[  330] = 'h00000405; 
    validation_data[  331] = 'h0000027f; 
    validation_data[  332] = 'h000002fa; 
    validation_data[  333] = 'h00000bdc; 
    validation_data[  334] = 'h00000ed2; 
    validation_data[  335] = 'h00000a61; 
    validation_data[  336] = 'h0000061c; 
    validation_data[  337] = 'h00000a7f; 
    validation_data[  338] = 'h00000b44; 
    validation_data[  339] = 'h000005c6; 
    validation_data[  340] = 'h00000551; 
    validation_data[  341] = 'h000007ab; 
    validation_data[  342] = 'h000000f6; 
    validation_data[  343] = 'h000004ca; 
    validation_data[  344] = 'h00000228; 
    validation_data[  345] = 'h000007a7; 
    validation_data[  346] = 'h0000023f; 
    validation_data[  347] = 'h000006a0; 
    validation_data[  348] = 'h00000323; 
    validation_data[  349] = 'h000007f0; 
    validation_data[  350] = 'h00000bfb; 
    validation_data[  351] = 'h00000e1b; 
    validation_data[  352] = 'h00000554; 
    validation_data[  353] = 'h00000add; 
    validation_data[  354] = 'h0000056a; 
    validation_data[  355] = 'h00000287; 
    validation_data[  356] = 'h00000540; 
    validation_data[  357] = 'h00000a9a; 
    validation_data[  358] = 'h0000079e; 
    validation_data[  359] = 'h000000f9; 
    validation_data[  360] = 'h00000e8c; 
    validation_data[  361] = 'h000008cd; 
    validation_data[  362] = 'h00000af9; 
    validation_data[  363] = 'h00000677; 
    validation_data[  364] = 'h000006a1; 
    validation_data[  365] = 'h00000a04; 
    validation_data[  366] = 'h00000820; 
    validation_data[  367] = 'h0000023a; 
    validation_data[  368] = 'h00000cb8; 
    validation_data[  369] = 'h00000128; 
    validation_data[  370] = 'h0000055d; 
    validation_data[  371] = 'h00000f79; 
    validation_data[  372] = 'h000001c5; 
    validation_data[  373] = 'h0000020c; 
    validation_data[  374] = 'h00000552; 
    validation_data[  375] = 'h00000659; 
    validation_data[  376] = 'h0000070e; 
    validation_data[  377] = 'h000005be; 
    validation_data[  378] = 'h00000cec; 
    validation_data[  379] = 'h0000063e; 
    validation_data[  380] = 'h0000049b; 
    validation_data[  381] = 'h00000f9b; 
    validation_data[  382] = 'h000009ef; 
    validation_data[  383] = 'h00000199; 
    validation_data[  384] = 'h00000e07; 
    validation_data[  385] = 'h00000839; 
    validation_data[  386] = 'h000008e8; 
    validation_data[  387] = 'h00000477; 
    validation_data[  388] = 'h00000897; 
    validation_data[  389] = 'h00000421; 
    validation_data[  390] = 'h000009c1; 
    validation_data[  391] = 'h00000ecc; 
    validation_data[  392] = 'h0000008c; 
    validation_data[  393] = 'h00000d0c; 
    validation_data[  394] = 'h0000021f; 
    validation_data[  395] = 'h00000a64; 
    validation_data[  396] = 'h00000f93; 
    validation_data[  397] = 'h00000513; 
    validation_data[  398] = 'h000003f3; 
    validation_data[  399] = 'h00000f3d; 
    validation_data[  400] = 'h000005d7; 
    validation_data[  401] = 'h00000c12; 
    validation_data[  402] = 'h000005c7; 
    validation_data[  403] = 'h0000042c; 
    validation_data[  404] = 'h00000487; 
    validation_data[  405] = 'h0000007f; 
    validation_data[  406] = 'h00000309; 
    validation_data[  407] = 'h00000f13; 
    validation_data[  408] = 'h000008b0; 
    validation_data[  409] = 'h00000a36; 
    validation_data[  410] = 'h00000b7c; 
    validation_data[  411] = 'h00000ef0; 
    validation_data[  412] = 'h00000cf8; 
    validation_data[  413] = 'h00000400; 
    validation_data[  414] = 'h000006d7; 
    validation_data[  415] = 'h00000a3c; 
    validation_data[  416] = 'h00000899; 
    validation_data[  417] = 'h000007f7; 
    validation_data[  418] = 'h00000f1f; 
    validation_data[  419] = 'h00000741; 
    validation_data[  420] = 'h0000083c; 
    validation_data[  421] = 'h000007e2; 
    validation_data[  422] = 'h0000098b; 
    validation_data[  423] = 'h000004c7; 
    validation_data[  424] = 'h0000069f; 
    validation_data[  425] = 'h00000a81; 
    validation_data[  426] = 'h00000502; 
    validation_data[  427] = 'h0000029f; 
    validation_data[  428] = 'h00000f62; 
    validation_data[  429] = 'h000004d1; 
    validation_data[  430] = 'h00000f1d; 
    validation_data[  431] = 'h00000d81; 
    validation_data[  432] = 'h0000070c; 
    validation_data[  433] = 'h000003b7; 
    validation_data[  434] = 'h00000a62; 
    validation_data[  435] = 'h00000036; 
    validation_data[  436] = 'h00000e0d; 
    validation_data[  437] = 'h0000064d; 
    validation_data[  438] = 'h00000295; 
    validation_data[  439] = 'h00000115; 
    validation_data[  440] = 'h00000e81; 
    validation_data[  441] = 'h00000c0a; 
    validation_data[  442] = 'h00000421; 
    validation_data[  443] = 'h00000347; 
    validation_data[  444] = 'h000006db; 
    validation_data[  445] = 'h00000568; 
    validation_data[  446] = 'h00000c0a; 
    validation_data[  447] = 'h00000011; 
    validation_data[  448] = 'h00000b4e; 
    validation_data[  449] = 'h00000197; 
    validation_data[  450] = 'h000000e9; 
    validation_data[  451] = 'h000000c1; 
    validation_data[  452] = 'h0000056d; 
    validation_data[  453] = 'h00000cad; 
    validation_data[  454] = 'h00000080; 
    validation_data[  455] = 'h00000b54; 
    validation_data[  456] = 'h00000107; 
    validation_data[  457] = 'h00000598; 
    validation_data[  458] = 'h0000084f; 
    validation_data[  459] = 'h0000016c; 
    validation_data[  460] = 'h00000dc8; 
    validation_data[  461] = 'h000007c7; 
    validation_data[  462] = 'h00000af2; 
    validation_data[  463] = 'h00000414; 
    validation_data[  464] = 'h00000aad; 
    validation_data[  465] = 'h000003bf; 
    validation_data[  466] = 'h000007d4; 
    validation_data[  467] = 'h00000d4c; 
    validation_data[  468] = 'h00000571; 
    validation_data[  469] = 'h00000ee4; 
    validation_data[  470] = 'h00000eaf; 
    validation_data[  471] = 'h00000f1d; 
    validation_data[  472] = 'h00000aa0; 
    validation_data[  473] = 'h00000911; 
    validation_data[  474] = 'h00000945; 
    validation_data[  475] = 'h00000c25; 
    validation_data[  476] = 'h00000be4; 
    validation_data[  477] = 'h00000e3e; 
    validation_data[  478] = 'h00000bf4; 
    validation_data[  479] = 'h00000352; 
    validation_data[  480] = 'h00000704; 
    validation_data[  481] = 'h000004cb; 
    validation_data[  482] = 'h000004b1; 
    validation_data[  483] = 'h00000f67; 
    validation_data[  484] = 'h000003de; 
    validation_data[  485] = 'h0000015a; 
    validation_data[  486] = 'h00000e6b; 
    validation_data[  487] = 'h00000a5e; 
    validation_data[  488] = 'h00000994; 
    validation_data[  489] = 'h00000738; 
    validation_data[  490] = 'h0000017c; 
    validation_data[  491] = 'h00000ad1; 
    validation_data[  492] = 'h0000094b; 
    validation_data[  493] = 'h000001c2; 
    validation_data[  494] = 'h00000a99; 
    validation_data[  495] = 'h000006fb; 
    validation_data[  496] = 'h0000035b; 
    validation_data[  497] = 'h00000ceb; 
    validation_data[  498] = 'h00000ea2; 
    validation_data[  499] = 'h00000709; 
    validation_data[  500] = 'h00000559; 
    validation_data[  501] = 'h00000264; 
    validation_data[  502] = 'h00000ab1; 
    validation_data[  503] = 'h00000495; 
    validation_data[  504] = 'h000007c8; 
    validation_data[  505] = 'h000005ad; 
    validation_data[  506] = 'h00000086; 
    validation_data[  507] = 'h000003f1; 
    validation_data[  508] = 'h00000f7d; 
    validation_data[  509] = 'h00000445; 
    validation_data[  510] = 'h00000ad9; 
    validation_data[  511] = 'h00000331; 
    validation_data[  512] = 'h000005a3; 
    validation_data[  513] = 'h000009fb; 
    validation_data[  514] = 'h0000038d; 
    validation_data[  515] = 'h00000969; 
    validation_data[  516] = 'h00000877; 
    validation_data[  517] = 'h00000782; 
    validation_data[  518] = 'h0000004a; 
    validation_data[  519] = 'h00000187; 
    validation_data[  520] = 'h000002b9; 
    validation_data[  521] = 'h00000a46; 
    validation_data[  522] = 'h00000541; 
    validation_data[  523] = 'h000000af; 
    validation_data[  524] = 'h00000c3c; 
    validation_data[  525] = 'h00000779; 
    validation_data[  526] = 'h00000b4b; 
    validation_data[  527] = 'h00000371; 
    validation_data[  528] = 'h000004ec; 
    validation_data[  529] = 'h00000ad6; 
    validation_data[  530] = 'h00000e8a; 
    validation_data[  531] = 'h00000d4f; 
    validation_data[  532] = 'h00000a0d; 
    validation_data[  533] = 'h00000b36; 
    validation_data[  534] = 'h000001e7; 
    validation_data[  535] = 'h0000045a; 
    validation_data[  536] = 'h000004a0; 
    validation_data[  537] = 'h00000e79; 
    validation_data[  538] = 'h000002a1; 
    validation_data[  539] = 'h00000180; 
    validation_data[  540] = 'h000007a6; 
    validation_data[  541] = 'h0000052d; 
    validation_data[  542] = 'h000000c5; 
    validation_data[  543] = 'h00000614; 
    validation_data[  544] = 'h00000786; 
    validation_data[  545] = 'h00000678; 
    validation_data[  546] = 'h00000e65; 
    validation_data[  547] = 'h0000096e; 
    validation_data[  548] = 'h0000063f; 
    validation_data[  549] = 'h00000bd6; 
    validation_data[  550] = 'h00000748; 
    validation_data[  551] = 'h000001e5; 
    validation_data[  552] = 'h00000970; 
    validation_data[  553] = 'h000002cd; 
    validation_data[  554] = 'h00000dbd; 
    validation_data[  555] = 'h000004c9; 
    validation_data[  556] = 'h000005c5; 
    validation_data[  557] = 'h0000084d; 
    validation_data[  558] = 'h00000552; 
    validation_data[  559] = 'h00000186; 
    validation_data[  560] = 'h0000011c; 
    validation_data[  561] = 'h00000708; 
    validation_data[  562] = 'h00000875; 
    validation_data[  563] = 'h000001a9; 
    validation_data[  564] = 'h0000027b; 
    validation_data[  565] = 'h000002f8; 
    validation_data[  566] = 'h00000c42; 
    validation_data[  567] = 'h00000a0a; 
    validation_data[  568] = 'h00000438; 
    validation_data[  569] = 'h0000048d; 
    validation_data[  570] = 'h00000e5f; 
    validation_data[  571] = 'h00000609; 
    validation_data[  572] = 'h00000334; 
    validation_data[  573] = 'h000006be; 
    validation_data[  574] = 'h00000bec; 
    validation_data[  575] = 'h000006f1; 
    validation_data[  576] = 'h00000a61; 
    validation_data[  577] = 'h00000461; 
    validation_data[  578] = 'h0000065e; 
    validation_data[  579] = 'h00000b0e; 
    validation_data[  580] = 'h00000870; 
    validation_data[  581] = 'h00000ef4; 
    validation_data[  582] = 'h00000dcb; 
    validation_data[  583] = 'h000001f7; 
    validation_data[  584] = 'h0000052d; 
    validation_data[  585] = 'h00000b03; 
    validation_data[  586] = 'h00000685; 
    validation_data[  587] = 'h00000f91; 
    validation_data[  588] = 'h00000250; 
    validation_data[  589] = 'h00000153; 
    validation_data[  590] = 'h000008af; 
    validation_data[  591] = 'h000007f5; 
    validation_data[  592] = 'h00000c28; 
    validation_data[  593] = 'h00000dd3; 
    validation_data[  594] = 'h00000bf9; 
    validation_data[  595] = 'h00000176; 
    validation_data[  596] = 'h00000205; 
    validation_data[  597] = 'h0000075c; 
    validation_data[  598] = 'h00000113; 
    validation_data[  599] = 'h00000f41; 
    validation_data[  600] = 'h00000c9a; 
    validation_data[  601] = 'h0000075c; 
    validation_data[  602] = 'h000002c1; 
    validation_data[  603] = 'h0000032d; 
    validation_data[  604] = 'h00000e46; 
    validation_data[  605] = 'h00000357; 
    validation_data[  606] = 'h00000ae1; 
    validation_data[  607] = 'h00000bab; 
    validation_data[  608] = 'h00000ab8; 
    validation_data[  609] = 'h0000071a; 
    validation_data[  610] = 'h0000095e; 
    validation_data[  611] = 'h0000077b; 
    validation_data[  612] = 'h00000017; 
    validation_data[  613] = 'h000003da; 
    validation_data[  614] = 'h00000670; 
    validation_data[  615] = 'h00000a1c; 
    validation_data[  616] = 'h000007a9; 
    validation_data[  617] = 'h00000565; 
    validation_data[  618] = 'h00000233; 
    validation_data[  619] = 'h00000c15; 
    validation_data[  620] = 'h000009b5; 
    validation_data[  621] = 'h00000990; 
    validation_data[  622] = 'h00000a50; 
    validation_data[  623] = 'h00000ed3; 
    validation_data[  624] = 'h000009bd; 
    validation_data[  625] = 'h00000524; 
    validation_data[  626] = 'h00000543; 
    validation_data[  627] = 'h00000e89; 
    validation_data[  628] = 'h000008fc; 
    validation_data[  629] = 'h000008aa; 
    validation_data[  630] = 'h0000096b; 
    validation_data[  631] = 'h000008f2; 
    validation_data[  632] = 'h00000257; 
    validation_data[  633] = 'h00000047; 
    validation_data[  634] = 'h0000053b; 
    validation_data[  635] = 'h000008d3; 
    validation_data[  636] = 'h00000932; 
    validation_data[  637] = 'h0000038b; 
    validation_data[  638] = 'h00000774; 
    validation_data[  639] = 'h00000751; 
    validation_data[  640] = 'h00000c3c; 
    validation_data[  641] = 'h00000a9a; 
    validation_data[  642] = 'h00000a98; 
    validation_data[  643] = 'h0000024f; 
    validation_data[  644] = 'h0000078f; 
    validation_data[  645] = 'h00000a51; 
    validation_data[  646] = 'h000007db; 
    validation_data[  647] = 'h00000d22; 
    validation_data[  648] = 'h000003bd; 
    validation_data[  649] = 'h00000b72; 
    validation_data[  650] = 'h000007ec; 
    validation_data[  651] = 'h0000030f; 
    validation_data[  652] = 'h00000453; 
    validation_data[  653] = 'h000004ec; 
    validation_data[  654] = 'h00000870; 
    validation_data[  655] = 'h00000a79; 
    validation_data[  656] = 'h00000792; 
    validation_data[  657] = 'h00000b90; 
    validation_data[  658] = 'h00000686; 
    validation_data[  659] = 'h00000a23; 
    validation_data[  660] = 'h000002eb; 
    validation_data[  661] = 'h00000d57; 
    validation_data[  662] = 'h00000b5e; 
    validation_data[  663] = 'h0000028a; 
    validation_data[  664] = 'h000004cd; 
    validation_data[  665] = 'h00000cc3; 
    validation_data[  666] = 'h0000071f; 
    validation_data[  667] = 'h00000d5b; 
    validation_data[  668] = 'h00000e55; 
    validation_data[  669] = 'h00000e20; 
    validation_data[  670] = 'h0000096b; 
    validation_data[  671] = 'h0000096f; 
    validation_data[  672] = 'h00000194; 
    validation_data[  673] = 'h00000959; 
    validation_data[  674] = 'h00000401; 
    validation_data[  675] = 'h00000edb; 
    validation_data[  676] = 'h00000ee5; 
    validation_data[  677] = 'h00000eb7; 
    validation_data[  678] = 'h00000bcd; 
    validation_data[  679] = 'h00000c4b; 
    validation_data[  680] = 'h000000f2; 
    validation_data[  681] = 'h0000008f; 
    validation_data[  682] = 'h00000383; 
    validation_data[  683] = 'h0000084c; 
    validation_data[  684] = 'h00000570; 
    validation_data[  685] = 'h0000077f; 
    validation_data[  686] = 'h00000c41; 
    validation_data[  687] = 'h000001f0; 
    validation_data[  688] = 'h000001f9; 
    validation_data[  689] = 'h00000d3e; 
    validation_data[  690] = 'h00000160; 
    validation_data[  691] = 'h00000f92; 
    validation_data[  692] = 'h000000c6; 
    validation_data[  693] = 'h00000836; 
    validation_data[  694] = 'h00000bfd; 
    validation_data[  695] = 'h00000ee7; 
    validation_data[  696] = 'h00000d64; 
    validation_data[  697] = 'h00000074; 
    validation_data[  698] = 'h00000cb4; 
    validation_data[  699] = 'h00000362; 
    validation_data[  700] = 'h00000065; 
    validation_data[  701] = 'h00000c50; 
    validation_data[  702] = 'h00000d02; 
    validation_data[  703] = 'h00000865; 
    validation_data[  704] = 'h000003cd; 
    validation_data[  705] = 'h00000a00; 
    validation_data[  706] = 'h00000a70; 
    validation_data[  707] = 'h00000a0c; 
    validation_data[  708] = 'h000008ea; 
    validation_data[  709] = 'h00000cab; 
    validation_data[  710] = 'h00000edd; 
    validation_data[  711] = 'h00000f7a; 
    validation_data[  712] = 'h00000219; 
    validation_data[  713] = 'h00000652; 
    validation_data[  714] = 'h0000063b; 
    validation_data[  715] = 'h00000d93; 
    validation_data[  716] = 'h0000024e; 
    validation_data[  717] = 'h00000f9f; 
    validation_data[  718] = 'h00000350; 
    validation_data[  719] = 'h0000000a; 
    validation_data[  720] = 'h000008d5; 
    validation_data[  721] = 'h000000e4; 
    validation_data[  722] = 'h000003fc; 
    validation_data[  723] = 'h00000cea; 
    validation_data[  724] = 'h00000d49; 
    validation_data[  725] = 'h00000dc6; 
    validation_data[  726] = 'h00000aba; 
    validation_data[  727] = 'h00000ae7; 
    validation_data[  728] = 'h00000431; 
    validation_data[  729] = 'h00000ce9; 
    validation_data[  730] = 'h000009e8; 
    validation_data[  731] = 'h000008e4; 
    validation_data[  732] = 'h00000137; 
    validation_data[  733] = 'h00000133; 
    validation_data[  734] = 'h00000072; 
    validation_data[  735] = 'h00000a1d; 
    validation_data[  736] = 'h00000dc3; 
    validation_data[  737] = 'h000004a8; 
    validation_data[  738] = 'h00000563; 
    validation_data[  739] = 'h00000862; 
    validation_data[  740] = 'h00000f10; 
    validation_data[  741] = 'h000007be; 
    validation_data[  742] = 'h00000be0; 
    validation_data[  743] = 'h00000082; 
    validation_data[  744] = 'h00000383; 
    validation_data[  745] = 'h00000882; 
    validation_data[  746] = 'h000006a0; 
    validation_data[  747] = 'h0000004f; 
    validation_data[  748] = 'h000001f6; 
    validation_data[  749] = 'h00000886; 
    validation_data[  750] = 'h0000073b; 
    validation_data[  751] = 'h00000b85; 
    validation_data[  752] = 'h00000978; 
    validation_data[  753] = 'h00000516; 
    validation_data[  754] = 'h000009c2; 
    validation_data[  755] = 'h0000069d; 
    validation_data[  756] = 'h00000d51; 
    validation_data[  757] = 'h00000f87; 
    validation_data[  758] = 'h000005dc; 
    validation_data[  759] = 'h00000c40; 
    validation_data[  760] = 'h00000a31; 
    validation_data[  761] = 'h0000003e; 
    validation_data[  762] = 'h00000860; 
    validation_data[  763] = 'h000009c9; 
    validation_data[  764] = 'h00000b7d; 
    validation_data[  765] = 'h00000f78; 
    validation_data[  766] = 'h00000a30; 
    validation_data[  767] = 'h00000a99; 
    validation_data[  768] = 'h0000046a; 
    validation_data[  769] = 'h000009f2; 
    validation_data[  770] = 'h00000a3c; 
    validation_data[  771] = 'h000008fb; 
    validation_data[  772] = 'h00000f60; 
    validation_data[  773] = 'h00000049; 
    validation_data[  774] = 'h000009ad; 
    validation_data[  775] = 'h000006db; 
    validation_data[  776] = 'h000003da; 
    validation_data[  777] = 'h00000579; 
    validation_data[  778] = 'h00000549; 
    validation_data[  779] = 'h000002f3; 
    validation_data[  780] = 'h000008ea; 
    validation_data[  781] = 'h00000418; 
    validation_data[  782] = 'h00000734; 
    validation_data[  783] = 'h00000269; 
    validation_data[  784] = 'h00000867; 
    validation_data[  785] = 'h00000253; 
    validation_data[  786] = 'h00000711; 
    validation_data[  787] = 'h00000cd7; 
    validation_data[  788] = 'h000004e5; 
    validation_data[  789] = 'h000004e2; 
    validation_data[  790] = 'h0000019c; 
    validation_data[  791] = 'h00000b5d; 
    validation_data[  792] = 'h0000085f; 
    validation_data[  793] = 'h000007c0; 
    validation_data[  794] = 'h00000501; 
    validation_data[  795] = 'h00000cc9; 
    validation_data[  796] = 'h0000049f; 
    validation_data[  797] = 'h00000e8a; 
    validation_data[  798] = 'h00000d03; 
    validation_data[  799] = 'h000007c3; 
    validation_data[  800] = 'h00000439; 
    validation_data[  801] = 'h00000657; 
    validation_data[  802] = 'h00000401; 
    validation_data[  803] = 'h0000084e; 
    validation_data[  804] = 'h00000eec; 
    validation_data[  805] = 'h000004bc; 
    validation_data[  806] = 'h0000035b; 
    validation_data[  807] = 'h000001ca; 
    validation_data[  808] = 'h00000111; 
    validation_data[  809] = 'h00000335; 
    validation_data[  810] = 'h00000dd1; 
    validation_data[  811] = 'h000003cd; 
    validation_data[  812] = 'h00000c7a; 
    validation_data[  813] = 'h00000c61; 
    validation_data[  814] = 'h00000af5; 
    validation_data[  815] = 'h00000878; 
    validation_data[  816] = 'h00000384; 
    validation_data[  817] = 'h00000ed4; 
    validation_data[  818] = 'h00000296; 
    validation_data[  819] = 'h000007b2; 
    validation_data[  820] = 'h000009bf; 
    validation_data[  821] = 'h00000cef; 
    validation_data[  822] = 'h00000d95; 
    validation_data[  823] = 'h00000c96; 
    validation_data[  824] = 'h00000488; 
    validation_data[  825] = 'h000008f9; 
    validation_data[  826] = 'h00000926; 
    validation_data[  827] = 'h00000a7c; 
    validation_data[  828] = 'h000000f3; 
    validation_data[  829] = 'h00000415; 
    validation_data[  830] = 'h00000946; 
    validation_data[  831] = 'h00000a24; 
    validation_data[  832] = 'h0000095b; 
    validation_data[  833] = 'h0000011e; 
    validation_data[  834] = 'h00000f74; 
    validation_data[  835] = 'h000002e4; 
    validation_data[  836] = 'h00000eed; 
    validation_data[  837] = 'h0000072c; 
    validation_data[  838] = 'h00000f52; 
    validation_data[  839] = 'h000007f4; 
    validation_data[  840] = 'h000001b5; 
    validation_data[  841] = 'h00000261; 
    validation_data[  842] = 'h000005c4; 
    validation_data[  843] = 'h00000276; 
    validation_data[  844] = 'h000003f5; 
    validation_data[  845] = 'h00000c44; 
    validation_data[  846] = 'h00000a1d; 
    validation_data[  847] = 'h00000306; 
    validation_data[  848] = 'h00000448; 
    validation_data[  849] = 'h00000c13; 
    validation_data[  850] = 'h00000ea0; 
    validation_data[  851] = 'h00000186; 
    validation_data[  852] = 'h00000f93; 
    validation_data[  853] = 'h00000d8a; 
    validation_data[  854] = 'h00000d1e; 
    validation_data[  855] = 'h0000007f; 
    validation_data[  856] = 'h000008d0; 
    validation_data[  857] = 'h00000eac; 
    validation_data[  858] = 'h00000d6e; 
    validation_data[  859] = 'h00000a57; 
    validation_data[  860] = 'h0000097a; 
    validation_data[  861] = 'h00000c5e; 
    validation_data[  862] = 'h0000069a; 
    validation_data[  863] = 'h00000c73; 
    validation_data[  864] = 'h00000b0b; 
    validation_data[  865] = 'h00000b6a; 
    validation_data[  866] = 'h00000212; 
    validation_data[  867] = 'h0000008e; 
    validation_data[  868] = 'h00000a7c; 
    validation_data[  869] = 'h00000118; 
    validation_data[  870] = 'h00000f8c; 
    validation_data[  871] = 'h00000338; 
    validation_data[  872] = 'h000005a6; 
    validation_data[  873] = 'h00000034; 
    validation_data[  874] = 'h00000078; 
    validation_data[  875] = 'h00000af4; 
    validation_data[  876] = 'h000002dc; 
    validation_data[  877] = 'h00000a85; 
    validation_data[  878] = 'h00000f20; 
    validation_data[  879] = 'h0000047c; 
    validation_data[  880] = 'h00000065; 
    validation_data[  881] = 'h00000d5c; 
    validation_data[  882] = 'h00000051; 
    validation_data[  883] = 'h00000419; 
    validation_data[  884] = 'h000000f1; 
    validation_data[  885] = 'h0000064f; 
    validation_data[  886] = 'h00000eef; 
    validation_data[  887] = 'h00000e27; 
    validation_data[  888] = 'h00000ee6; 
    validation_data[  889] = 'h00000102; 
    validation_data[  890] = 'h000007f3; 
    validation_data[  891] = 'h0000041f; 
    validation_data[  892] = 'h00000cef; 
    validation_data[  893] = 'h000003c0; 
    validation_data[  894] = 'h00000ca7; 
    validation_data[  895] = 'h00000623; 
    validation_data[  896] = 'h000002f8; 
    validation_data[  897] = 'h0000026d; 
    validation_data[  898] = 'h000007f4; 
    validation_data[  899] = 'h0000011e; 
    validation_data[  900] = 'h00000312; 
    validation_data[  901] = 'h000006bf; 
    validation_data[  902] = 'h00000bcf; 
    validation_data[  903] = 'h00000926; 
    validation_data[  904] = 'h00000654; 
    validation_data[  905] = 'h00000686; 
    validation_data[  906] = 'h000008e5; 
    validation_data[  907] = 'h000009b9; 
    validation_data[  908] = 'h0000032b; 
    validation_data[  909] = 'h00000d2e; 
    validation_data[  910] = 'h00000186; 
    validation_data[  911] = 'h00000823; 
    validation_data[  912] = 'h00000266; 
    validation_data[  913] = 'h0000098f; 
    validation_data[  914] = 'h000005b0; 
    validation_data[  915] = 'h00000b91; 
    validation_data[  916] = 'h00000acc; 
    validation_data[  917] = 'h000003bf; 
    validation_data[  918] = 'h00000c0a; 
    validation_data[  919] = 'h00000a96; 
    validation_data[  920] = 'h00000d68; 
    validation_data[  921] = 'h000009a4; 
    validation_data[  922] = 'h00000cf3; 
    validation_data[  923] = 'h000004b0; 
    validation_data[  924] = 'h00000519; 
    validation_data[  925] = 'h00000bb3; 
    validation_data[  926] = 'h000001b3; 
    validation_data[  927] = 'h00000069; 
    validation_data[  928] = 'h00000884; 
    validation_data[  929] = 'h0000099c; 
    validation_data[  930] = 'h0000003b; 
    validation_data[  931] = 'h00000f7f; 
    validation_data[  932] = 'h00000294; 
    validation_data[  933] = 'h000007e7; 
    validation_data[  934] = 'h0000058f; 
    validation_data[  935] = 'h00000b58; 
    validation_data[  936] = 'h00000352; 
    validation_data[  937] = 'h00000ba0; 
    validation_data[  938] = 'h00000330; 
    validation_data[  939] = 'h000000c1; 
    validation_data[  940] = 'h0000060f; 
    validation_data[  941] = 'h000009be; 
    validation_data[  942] = 'h00000317; 
    validation_data[  943] = 'h000001be; 
    validation_data[  944] = 'h0000052e; 
    validation_data[  945] = 'h0000023f; 
    validation_data[  946] = 'h00000442; 
    validation_data[  947] = 'h00000c5a; 
    validation_data[  948] = 'h000005e8; 
    validation_data[  949] = 'h000005a1; 
    validation_data[  950] = 'h00000cc8; 
    validation_data[  951] = 'h00000ef0; 
    validation_data[  952] = 'h000008a3; 
    validation_data[  953] = 'h000006b5; 
    validation_data[  954] = 'h00000dfb; 
    validation_data[  955] = 'h00000111; 
    validation_data[  956] = 'h00000c51; 
    validation_data[  957] = 'h00000f35; 
    validation_data[  958] = 'h00000f7c; 
    validation_data[  959] = 'h000006bc; 
    validation_data[  960] = 'h000009a6; 
    validation_data[  961] = 'h000006f3; 
    validation_data[  962] = 'h0000012f; 
    validation_data[  963] = 'h00000ace; 
    validation_data[  964] = 'h00000b62; 
    validation_data[  965] = 'h00000840; 
    validation_data[  966] = 'h000005ea; 
    validation_data[  967] = 'h00000236; 
    validation_data[  968] = 'h00000e64; 
    validation_data[  969] = 'h00000392; 
    validation_data[  970] = 'h00000c19; 
    validation_data[  971] = 'h0000062f; 
    validation_data[  972] = 'h00000e92; 
    validation_data[  973] = 'h00000623; 
    validation_data[  974] = 'h0000062c; 
    validation_data[  975] = 'h00000433; 
    validation_data[  976] = 'h00000bcd; 
    validation_data[  977] = 'h00000b7a; 
    validation_data[  978] = 'h000001c0; 
    validation_data[  979] = 'h00000133; 
    validation_data[  980] = 'h0000058d; 
    validation_data[  981] = 'h000008e6; 
    validation_data[  982] = 'h00000802; 
    validation_data[  983] = 'h000003f8; 
    validation_data[  984] = 'h00000f6e; 
    validation_data[  985] = 'h00000512; 
    validation_data[  986] = 'h00000b8e; 
    validation_data[  987] = 'h00000bc0; 
    validation_data[  988] = 'h00000a23; 
    validation_data[  989] = 'h0000099b; 
    validation_data[  990] = 'h00000c84; 
    validation_data[  991] = 'h00000e93; 
    validation_data[  992] = 'h000005e8; 
    validation_data[  993] = 'h0000049c; 
    validation_data[  994] = 'h00000b8c; 
    validation_data[  995] = 'h00000a0e; 
    validation_data[  996] = 'h0000076f; 
    validation_data[  997] = 'h00000609; 
    validation_data[  998] = 'h0000076b; 
    validation_data[  999] = 'h00000e29; 

end


reg clk = 1'b1, rst = 1'b1;
initial #4 rst = 1'b0;
always  #1 clk = ~clk;

wire  miss;
wire [31:0] rd_data;
reg  [31:0] index = 0, wr_data = 0, addr = 0;
reg  rd_req = 1'b0, wr_req = 1'b0;
reg rd_req_ff = 1'b0, miss_ff = 1'b0;
reg [31:0] validation_count = 0;

always @ (posedge clk or posedge rst)
    if(rst) begin
        rd_req_ff <= 1'b0;
        miss_ff   <= 1'b0;
    end else begin
        rd_req_ff <= rd_req;
        miss_ff   <= miss;
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        validation_count <= 0;
    end else begin
        if(validation_count>=`DATA_COUNT) begin
            validation_count <= 'hffffffff;
        end else if(rd_req_ff && (index>(4*`DATA_COUNT))) begin
            if(~miss_ff) begin
                if(validation_data[validation_count]==rd_data)
                    validation_count <= validation_count+1;
                else
                    validation_count <= 0;
            end
        end else begin
            validation_count <= 0;
        end
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        index   <= 0;
        wr_data <= 0;
        addr    <= 0;
        rd_req  <= 1'b0;
        wr_req  <= 1'b0;
    end else begin
        if(~miss) begin
            if(index<`RDWR_COUNT) begin
                if(wr_cycle[index]) begin
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b1;
                end else if(rd_cycle[index]) begin
                    wr_data <= 0;
                    rd_req  <= 1'b1;
                    wr_req  <= 1'b0;
                end else begin
                    wr_data <= 0;
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b0;
                end
                wr_data <= wr_data_rom[index];
                addr    <= addr_rom[index];
                index <= index + 1;
            end else begin
                wr_data <= 0;
                addr    <= 0;
                rd_req  <= 1'b0;
                wr_req  <= 1'b0;
            end
        end
    end

cache #(
    .LINE_ADDR_LEN  ( 3             ),
    .SET_ADDR_LEN   ( 2             ),
    .TAG_ADDR_LEN   ( 12            ),
    .WAY_CNT        ( 3             )
) cache_test_instance (
    .clk            ( clk           ),
    .rst            ( rst           ),
    .miss           ( miss          ),
    .addr           ( addr          ),
    .rd_req         ( rd_req        ),
    .rd_data        ( rd_data       ),
    .wr_req         ( wr_req        ),
    .wr_data        ( wr_data       )
);

endmodule

