
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    ram_cell[       0] = 32'h00000313;
    ram_cell[       1] = 32'h00000223;
    ram_cell[       2] = 32'h000003e8;
    ram_cell[       3] = 32'h00000707;
    ram_cell[       4] = 32'h0000001f;
    ram_cell[       5] = 32'h00000219;
    ram_cell[       6] = 32'h00000066;
    ram_cell[       7] = 32'h0000036d;
    ram_cell[       8] = 32'h00000731;
    ram_cell[       9] = 32'h000001f8;
    ram_cell[      10] = 32'h0000056e;
    ram_cell[      11] = 32'h00000229;
    ram_cell[      12] = 32'h00000358;
    ram_cell[      13] = 32'h00000757;
    ram_cell[      14] = 32'h00000328;
    ram_cell[      15] = 32'h000001be;
    ram_cell[      16] = 32'h0000012c;
    ram_cell[      17] = 32'h0000017c;
    ram_cell[      18] = 32'h000002be;
    ram_cell[      19] = 32'h000001fd;
    ram_cell[      20] = 32'h00000260;
    ram_cell[      21] = 32'h00000720;
    ram_cell[      22] = 32'h00000362;
    ram_cell[      23] = 32'h00000735;
    ram_cell[      24] = 32'h0000001c;
    ram_cell[      25] = 32'h00000704;
    ram_cell[      26] = 32'h0000052a;
    ram_cell[      27] = 32'h000000ac;
    ram_cell[      28] = 32'h00000538;
    ram_cell[      29] = 32'h00000025;
    ram_cell[      30] = 32'h0000051c;
    ram_cell[      31] = 32'h0000069a;
    ram_cell[      32] = 32'h00000288;
    ram_cell[      33] = 32'h0000057a;
    ram_cell[      34] = 32'h00000257;
    ram_cell[      35] = 32'h00000081;
    ram_cell[      36] = 32'h000004e9;
    ram_cell[      37] = 32'h00000621;
    ram_cell[      38] = 32'h0000029f;
    ram_cell[      39] = 32'h00000447;
    ram_cell[      40] = 32'h0000007a;
    ram_cell[      41] = 32'h00000387;
    ram_cell[      42] = 32'h000006fa;
    ram_cell[      43] = 32'h00000171;
    ram_cell[      44] = 32'h00000695;
    ram_cell[      45] = 32'h000002d8;
    ram_cell[      46] = 32'h0000016e;
    ram_cell[      47] = 32'h000001c4;
    ram_cell[      48] = 32'h0000001b;
    ram_cell[      49] = 32'h000005a6;
    ram_cell[      50] = 32'h000003e9;
    ram_cell[      51] = 32'h00000099;
    ram_cell[      52] = 32'h00000446;
    ram_cell[      53] = 32'h00000356;
    ram_cell[      54] = 32'h000004a3;
    ram_cell[      55] = 32'h000007ab;
    ram_cell[      56] = 32'h00000239;
    ram_cell[      57] = 32'h000000f1;
    ram_cell[      58] = 32'h00000625;
    ram_cell[      59] = 32'h00000200;
    ram_cell[      60] = 32'h000003ea;
    ram_cell[      61] = 32'h00000398;
    ram_cell[      62] = 32'h0000013b;
    ram_cell[      63] = 32'h00000372;
    ram_cell[      64] = 32'h000002c9;
    ram_cell[      65] = 32'h000005f8;
    ram_cell[      66] = 32'h000000dc;
    ram_cell[      67] = 32'h00000561;
    ram_cell[      68] = 32'h000001b6;
    ram_cell[      69] = 32'h000004ee;
    ram_cell[      70] = 32'h00000598;
    ram_cell[      71] = 32'h000005d1;
    ram_cell[      72] = 32'h000005b4;
    ram_cell[      73] = 32'h00000578;
    ram_cell[      74] = 32'h000003fd;
    ram_cell[      75] = 32'h0000079c;
    ram_cell[      76] = 32'h00000037;
    ram_cell[      77] = 32'h0000018f;
    ram_cell[      78] = 32'h00000271;
    ram_cell[      79] = 32'h000000bc;
    ram_cell[      80] = 32'h00000485;
    ram_cell[      81] = 32'h000007f9;
    ram_cell[      82] = 32'h00000541;
    ram_cell[      83] = 32'h00000090;
    ram_cell[      84] = 32'h000007ce;
    ram_cell[      85] = 32'h0000012a;
    ram_cell[      86] = 32'h000007c8;
    ram_cell[      87] = 32'h000006ef;
    ram_cell[      88] = 32'h0000025d;
    ram_cell[      89] = 32'h0000008b;
    ram_cell[      90] = 32'h000003cf;
    ram_cell[      91] = 32'h000005b9;
    ram_cell[      92] = 32'h0000076d;
    ram_cell[      93] = 32'h0000013a;
    ram_cell[      94] = 32'h0000058c;
    ram_cell[      95] = 32'h0000003b;
    ram_cell[      96] = 32'h000006f8;
    ram_cell[      97] = 32'h0000017d;
    ram_cell[      98] = 32'h0000052d;
    ram_cell[      99] = 32'h0000077d;
    ram_cell[     100] = 32'h000001d2;
    ram_cell[     101] = 32'h000006bf;
    ram_cell[     102] = 32'h00000027;
    ram_cell[     103] = 32'h000005a7;
    ram_cell[     104] = 32'h00000196;
    ram_cell[     105] = 32'h000002c6;
    ram_cell[     106] = 32'h000002d6;
    ram_cell[     107] = 32'h0000044e;
    ram_cell[     108] = 32'h00000031;
    ram_cell[     109] = 32'h0000032b;
    ram_cell[     110] = 32'h0000024b;
    ram_cell[     111] = 32'h000000d6;
    ram_cell[     112] = 32'h000006a8;
    ram_cell[     113] = 32'h0000079b;
    ram_cell[     114] = 32'h000004c7;
    ram_cell[     115] = 32'h0000049b;
    ram_cell[     116] = 32'h00000415;
    ram_cell[     117] = 32'h00000267;
    ram_cell[     118] = 32'h0000063d;
    ram_cell[     119] = 32'h0000076f;
    ram_cell[     120] = 32'h000002d4;
    ram_cell[     121] = 32'h000001ba;
    ram_cell[     122] = 32'h0000051f;
    ram_cell[     123] = 32'h00000304;
    ram_cell[     124] = 32'h000000e9;
    ram_cell[     125] = 32'h000005a9;
    ram_cell[     126] = 32'h0000072b;
    ram_cell[     127] = 32'h00000098;
    ram_cell[     128] = 32'h00000575;
    ram_cell[     129] = 32'h00000792;
    ram_cell[     130] = 32'h000006a3;
    ram_cell[     131] = 32'h000001af;
    ram_cell[     132] = 32'h00000773;
    ram_cell[     133] = 32'h000006df;
    ram_cell[     134] = 32'h00000301;
    ram_cell[     135] = 32'h0000034a;
    ram_cell[     136] = 32'h000000b6;
    ram_cell[     137] = 32'h00000445;
    ram_cell[     138] = 32'h0000012f;
    ram_cell[     139] = 32'h0000034b;
    ram_cell[     140] = 32'h00000365;
    ram_cell[     141] = 32'h000006b8;
    ram_cell[     142] = 32'h000001ca;
    ram_cell[     143] = 32'h000007b1;
    ram_cell[     144] = 32'h000002d3;
    ram_cell[     145] = 32'h000001fb;
    ram_cell[     146] = 32'h00000230;
    ram_cell[     147] = 32'h000004e2;
    ram_cell[     148] = 32'h000006cf;
    ram_cell[     149] = 32'h000005ba;
    ram_cell[     150] = 32'h00000608;
    ram_cell[     151] = 32'h00000282;
    ram_cell[     152] = 32'h000005f9;
    ram_cell[     153] = 32'h0000005b;
    ram_cell[     154] = 32'h00000787;
    ram_cell[     155] = 32'h000001df;
    ram_cell[     156] = 32'h00000124;
    ram_cell[     157] = 32'h00000484;
    ram_cell[     158] = 32'h000006d1;
    ram_cell[     159] = 32'h00000011;
    ram_cell[     160] = 32'h000001c3;
    ram_cell[     161] = 32'h0000068c;
    ram_cell[     162] = 32'h0000072d;
    ram_cell[     163] = 32'h000006e5;
    ram_cell[     164] = 32'h0000058f;
    ram_cell[     165] = 32'h000004ff;
    ram_cell[     166] = 32'h0000035b;
    ram_cell[     167] = 32'h00000318;
    ram_cell[     168] = 32'h000000e3;
    ram_cell[     169] = 32'h000002cf;
    ram_cell[     170] = 32'h000003e4;
    ram_cell[     171] = 32'h000002e0;
    ram_cell[     172] = 32'h000002fc;
    ram_cell[     173] = 32'h0000064b;
    ram_cell[     174] = 32'h00000283;
    ram_cell[     175] = 32'h00000004;
    ram_cell[     176] = 32'h00000771;
    ram_cell[     177] = 32'h00000281;
    ram_cell[     178] = 32'h00000573;
    ram_cell[     179] = 32'h000000d7;
    ram_cell[     180] = 32'h0000065c;
    ram_cell[     181] = 32'h0000016c;
    ram_cell[     182] = 32'h00000501;
    ram_cell[     183] = 32'h000001d8;
    ram_cell[     184] = 32'h00000245;
    ram_cell[     185] = 32'h00000084;
    ram_cell[     186] = 32'h000004fa;
    ram_cell[     187] = 32'h00000559;
    ram_cell[     188] = 32'h000007f0;
    ram_cell[     189] = 32'h000007f6;
    ram_cell[     190] = 32'h000003c7;
    ram_cell[     191] = 32'h000003cc;
    ram_cell[     192] = 32'h00000606;
    ram_cell[     193] = 32'h000006a5;
    ram_cell[     194] = 32'h0000058e;
    ram_cell[     195] = 32'h0000018e;
    ram_cell[     196] = 32'h000005a2;
    ram_cell[     197] = 32'h00000308;
    ram_cell[     198] = 32'h0000011c;
    ram_cell[     199] = 32'h0000038d;
    ram_cell[     200] = 32'h00000333;
    ram_cell[     201] = 32'h000004d2;
    ram_cell[     202] = 32'h000005da;
    ram_cell[     203] = 32'h000001a4;
    ram_cell[     204] = 32'h00000264;
    ram_cell[     205] = 32'h000000f6;
    ram_cell[     206] = 32'h000002e7;
    ram_cell[     207] = 32'h000002bc;
    ram_cell[     208] = 32'h0000032a;
    ram_cell[     209] = 32'h0000069f;
    ram_cell[     210] = 32'h000005be;
    ram_cell[     211] = 32'h00000554;
    ram_cell[     212] = 32'h000002e6;
    ram_cell[     213] = 32'h0000048e;
    ram_cell[     214] = 32'h00000545;
    ram_cell[     215] = 32'h000000e0;
    ram_cell[     216] = 32'h00000166;
    ram_cell[     217] = 32'h000002d1;
    ram_cell[     218] = 32'h0000037b;
    ram_cell[     219] = 32'h00000464;
    ram_cell[     220] = 32'h0000062a;
    ram_cell[     221] = 32'h0000067a;
    ram_cell[     222] = 32'h000007f3;
    ram_cell[     223] = 32'h0000036e;
    ram_cell[     224] = 32'h0000065f;
    ram_cell[     225] = 32'h000001f6;
    ram_cell[     226] = 32'h0000026e;
    ram_cell[     227] = 32'h000004f0;
    ram_cell[     228] = 32'h000001cd;
    ram_cell[     229] = 32'h00000576;
    ram_cell[     230] = 32'h000005c4;
    ram_cell[     231] = 32'h0000045d;
    ram_cell[     232] = 32'h000005fe;
    ram_cell[     233] = 32'h000007d3;
    ram_cell[     234] = 32'h0000029b;
    ram_cell[     235] = 32'h00000389;
    ram_cell[     236] = 32'h000007ca;
    ram_cell[     237] = 32'h00000647;
    ram_cell[     238] = 32'h00000513;
    ram_cell[     239] = 32'h0000057b;
    ram_cell[     240] = 32'h000007d6;
    ram_cell[     241] = 32'h000004d9;
    ram_cell[     242] = 32'h00000146;
    ram_cell[     243] = 32'h000007e5;
    ram_cell[     244] = 32'h0000073f;
    ram_cell[     245] = 32'h000002d9;
    ram_cell[     246] = 32'h00000607;
    ram_cell[     247] = 32'h00000499;
    ram_cell[     248] = 32'h00000320;
    ram_cell[     249] = 32'h0000032f;
    ram_cell[     250] = 32'h00000491;
    ram_cell[     251] = 32'h000001c8;
    ram_cell[     252] = 32'h000005f5;
    ram_cell[     253] = 32'h00000178;
    ram_cell[     254] = 32'h000004c8;
    ram_cell[     255] = 32'h000000c4;
    ram_cell[     256] = 32'h0000056a;
    ram_cell[     257] = 32'h00000193;
    ram_cell[     258] = 32'h00000537;
    ram_cell[     259] = 32'h00000630;
    ram_cell[     260] = 32'h00000174;
    ram_cell[     261] = 32'h000000da;
    ram_cell[     262] = 32'h00000247;
    ram_cell[     263] = 32'h0000035d;
    ram_cell[     264] = 32'h0000054b;
    ram_cell[     265] = 32'h000004ce;
    ram_cell[     266] = 32'h000003c4;
    ram_cell[     267] = 32'h000001c2;
    ram_cell[     268] = 32'h000007ee;
    ram_cell[     269] = 32'h000007dc;
    ram_cell[     270] = 32'h00000199;
    ram_cell[     271] = 32'h000005d0;
    ram_cell[     272] = 32'h0000065d;
    ram_cell[     273] = 32'h0000012d;
    ram_cell[     274] = 32'h00000185;
    ram_cell[     275] = 32'h00000409;
    ram_cell[     276] = 32'h000006b9;
    ram_cell[     277] = 32'h000000a0;
    ram_cell[     278] = 32'h00000189;
    ram_cell[     279] = 32'h00000074;
    ram_cell[     280] = 32'h0000041e;
    ram_cell[     281] = 32'h000000db;
    ram_cell[     282] = 32'h00000046;
    ram_cell[     283] = 32'h00000068;
    ram_cell[     284] = 32'h0000050f;
    ram_cell[     285] = 32'h000001de;
    ram_cell[     286] = 32'h0000023e;
    ram_cell[     287] = 32'h000003ad;
    ram_cell[     288] = 32'h000003fc;
    ram_cell[     289] = 32'h00000684;
    ram_cell[     290] = 32'h000006a2;
    ram_cell[     291] = 32'h00000548;
    ram_cell[     292] = 32'h00000427;
    ram_cell[     293] = 32'h00000095;
    ram_cell[     294] = 32'h00000224;
    ram_cell[     295] = 32'h000001d1;
    ram_cell[     296] = 32'h00000547;
    ram_cell[     297] = 32'h00000092;
    ram_cell[     298] = 32'h00000688;
    ram_cell[     299] = 32'h000000d2;
    ram_cell[     300] = 32'h0000045f;
    ram_cell[     301] = 32'h000003ac;
    ram_cell[     302] = 32'h000000fd;
    ram_cell[     303] = 32'h000000d3;
    ram_cell[     304] = 32'h000006f2;
    ram_cell[     305] = 32'h0000068e;
    ram_cell[     306] = 32'h0000028e;
    ram_cell[     307] = 32'h0000006c;
    ram_cell[     308] = 32'h000004b5;
    ram_cell[     309] = 32'h000005ed;
    ram_cell[     310] = 32'h000000d5;
    ram_cell[     311] = 32'h00000293;
    ram_cell[     312] = 32'h00000651;
    ram_cell[     313] = 32'h0000053d;
    ram_cell[     314] = 32'h00000776;
    ram_cell[     315] = 32'h000000a8;
    ram_cell[     316] = 32'h0000072e;
    ram_cell[     317] = 32'h000003ca;
    ram_cell[     318] = 32'h000005dd;
    ram_cell[     319] = 32'h00000531;
    ram_cell[     320] = 32'h0000027b;
    ram_cell[     321] = 32'h00000798;
    ram_cell[     322] = 32'h000001ee;
    ram_cell[     323] = 32'h0000029c;
    ram_cell[     324] = 32'h00000233;
    ram_cell[     325] = 32'h000007d9;
    ram_cell[     326] = 32'h000006a4;
    ram_cell[     327] = 32'h0000003c;
    ram_cell[     328] = 32'h000007cb;
    ram_cell[     329] = 32'h0000070d;
    ram_cell[     330] = 32'h00000034;
    ram_cell[     331] = 32'h000001b2;
    ram_cell[     332] = 32'h00000593;
    ram_cell[     333] = 32'h00000634;
    ram_cell[     334] = 32'h00000108;
    ram_cell[     335] = 32'h000005de;
    ram_cell[     336] = 32'h00000136;
    ram_cell[     337] = 32'h000000aa;
    ram_cell[     338] = 32'h00000154;
    ram_cell[     339] = 32'h0000043a;
    ram_cell[     340] = 32'h0000034f;
    ram_cell[     341] = 32'h00000131;
    ram_cell[     342] = 32'h00000770;
    ram_cell[     343] = 32'h000007db;
    ram_cell[     344] = 32'h000001c5;
    ram_cell[     345] = 32'h00000518;
    ram_cell[     346] = 32'h0000023f;
    ram_cell[     347] = 32'h000004c5;
    ram_cell[     348] = 32'h000003c8;
    ram_cell[     349] = 32'h00000552;
    ram_cell[     350] = 32'h00000015;
    ram_cell[     351] = 32'h00000057;
    ram_cell[     352] = 32'h000000a6;
    ram_cell[     353] = 32'h00000567;
    ram_cell[     354] = 32'h000000e2;
    ram_cell[     355] = 32'h000003a1;
    ram_cell[     356] = 32'h000006e0;
    ram_cell[     357] = 32'h000006b7;
    ram_cell[     358] = 32'h00000622;
    ram_cell[     359] = 32'h00000306;
    ram_cell[     360] = 32'h00000003;
    ram_cell[     361] = 32'h000002ac;
    ram_cell[     362] = 32'h00000611;
    ram_cell[     363] = 32'h000006b1;
    ram_cell[     364] = 32'h0000034c;
    ram_cell[     365] = 32'h000006e2;
    ram_cell[     366] = 32'h000006ca;
    ram_cell[     367] = 32'h000001fa;
    ram_cell[     368] = 32'h00000311;
    ram_cell[     369] = 32'h0000014f;
    ram_cell[     370] = 32'h000004b7;
    ram_cell[     371] = 32'h0000030a;
    ram_cell[     372] = 32'h000005b1;
    ram_cell[     373] = 32'h000007a2;
    ram_cell[     374] = 32'h00000657;
    ram_cell[     375] = 32'h000004a9;
    ram_cell[     376] = 32'h0000023a;
    ram_cell[     377] = 32'h00000546;
    ram_cell[     378] = 32'h00000643;
    ram_cell[     379] = 32'h00000734;
    ram_cell[     380] = 32'h000004f9;
    ram_cell[     381] = 32'h00000403;
    ram_cell[     382] = 32'h00000117;
    ram_cell[     383] = 32'h00000187;
    ram_cell[     384] = 32'h00000483;
    ram_cell[     385] = 32'h00000201;
    ram_cell[     386] = 32'h0000008e;
    ram_cell[     387] = 32'h000004da;
    ram_cell[     388] = 32'h000006f0;
    ram_cell[     389] = 32'h00000203;
    ram_cell[     390] = 32'h0000055e;
    ram_cell[     391] = 32'h000007e4;
    ram_cell[     392] = 32'h00000580;
    ram_cell[     393] = 32'h00000054;
    ram_cell[     394] = 32'h000006c1;
    ram_cell[     395] = 32'h00000624;
    ram_cell[     396] = 32'h000000ea;
    ram_cell[     397] = 32'h00000597;
    ram_cell[     398] = 32'h0000031f;
    ram_cell[     399] = 32'h000006ed;
    ram_cell[     400] = 32'h00000749;
    ram_cell[     401] = 32'h000002e5;
    ram_cell[     402] = 32'h00000036;
    ram_cell[     403] = 32'h000000ef;
    ram_cell[     404] = 32'h000005ce;
    ram_cell[     405] = 32'h00000571;
    ram_cell[     406] = 32'h000004f5;
    ram_cell[     407] = 32'h000001cf;
    ram_cell[     408] = 32'h000005c1;
    ram_cell[     409] = 32'h00000148;
    ram_cell[     410] = 32'h0000007d;
    ram_cell[     411] = 32'h00000275;
    ram_cell[     412] = 32'h00000699;
    ram_cell[     413] = 32'h0000035f;
    ram_cell[     414] = 32'h00000118;
    ram_cell[     415] = 32'h00000646;
    ram_cell[     416] = 32'h00000041;
    ram_cell[     417] = 32'h00000243;
    ram_cell[     418] = 32'h000004d8;
    ram_cell[     419] = 32'h0000048f;
    ram_cell[     420] = 32'h0000001e;
    ram_cell[     421] = 32'h00000300;
    ram_cell[     422] = 32'h0000042a;
    ram_cell[     423] = 32'h000005fd;
    ram_cell[     424] = 32'h00000125;
    ram_cell[     425] = 32'h00000682;
    ram_cell[     426] = 32'h0000028b;
    ram_cell[     427] = 32'h000006b5;
    ram_cell[     428] = 32'h00000238;
    ram_cell[     429] = 32'h000005e1;
    ram_cell[     430] = 32'h00000059;
    ram_cell[     431] = 32'h000004ac;
    ram_cell[     432] = 32'h000001c1;
    ram_cell[     433] = 32'h00000420;
    ram_cell[     434] = 32'h00000708;
    ram_cell[     435] = 32'h000002e4;
    ram_cell[     436] = 32'h00000198;
    ram_cell[     437] = 32'h0000011e;
    ram_cell[     438] = 32'h000001ac;
    ram_cell[     439] = 32'h000004a0;
    ram_cell[     440] = 32'h000006db;
    ram_cell[     441] = 32'h000006f1;
    ram_cell[     442] = 32'h00000432;
    ram_cell[     443] = 32'h0000046d;
    ram_cell[     444] = 32'h0000053b;
    ram_cell[     445] = 32'h00000106;
    ram_cell[     446] = 32'h00000780;
    ram_cell[     447] = 32'h00000299;
    ram_cell[     448] = 32'h000004cd;
    ram_cell[     449] = 32'h0000070e;
    ram_cell[     450] = 32'h00000658;
    ram_cell[     451] = 32'h000007b9;
    ram_cell[     452] = 32'h00000570;
    ram_cell[     453] = 32'h00000709;
    ram_cell[     454] = 32'h000005c7;
    ram_cell[     455] = 32'h00000550;
    ram_cell[     456] = 32'h0000045e;
    ram_cell[     457] = 32'h000007b5;
    ram_cell[     458] = 32'h000005c8;
    ram_cell[     459] = 32'h0000038b;
    ram_cell[     460] = 32'h00000493;
    ram_cell[     461] = 32'h000005d6;
    ram_cell[     462] = 32'h0000003d;
    ram_cell[     463] = 32'h0000019e;
    ram_cell[     464] = 32'h000005ea;
    ram_cell[     465] = 32'h00000693;
    ram_cell[     466] = 32'h00000490;
    ram_cell[     467] = 32'h00000505;
    ram_cell[     468] = 32'h00000370;
    ram_cell[     469] = 32'h00000412;
    ram_cell[     470] = 32'h00000449;
    ram_cell[     471] = 32'h00000553;
    ram_cell[     472] = 32'h0000042f;
    ram_cell[     473] = 32'h00000424;
    ram_cell[     474] = 32'h00000116;
    ram_cell[     475] = 32'h000000f9;
    ram_cell[     476] = 32'h0000023d;
    ram_cell[     477] = 32'h000002ce;
    ram_cell[     478] = 32'h00000182;
    ram_cell[     479] = 32'h000001ae;
    ram_cell[     480] = 32'h000002d2;
    ram_cell[     481] = 32'h00000279;
    ram_cell[     482] = 32'h0000062f;
    ram_cell[     483] = 32'h000006f5;
    ram_cell[     484] = 32'h000007f7;
    ram_cell[     485] = 32'h00000235;
    ram_cell[     486] = 32'h00000324;
    ram_cell[     487] = 32'h00000246;
    ram_cell[     488] = 32'h0000022b;
    ram_cell[     489] = 32'h000005b8;
    ram_cell[     490] = 32'h000007ec;
    ram_cell[     491] = 32'h00000322;
    ram_cell[     492] = 32'h00000316;
    ram_cell[     493] = 32'h00000014;
    ram_cell[     494] = 32'h00000794;
    ram_cell[     495] = 32'h000007d2;
    ram_cell[     496] = 32'h00000228;
    ram_cell[     497] = 32'h0000021f;
    ram_cell[     498] = 32'h00000411;
    ram_cell[     499] = 32'h000005ab;
    ram_cell[     500] = 32'h000004b4;
    ram_cell[     501] = 32'h00000509;
    ram_cell[     502] = 32'h00000120;
    ram_cell[     503] = 32'h00000609;
    ram_cell[     504] = 32'h000001e2;
    ram_cell[     505] = 32'h0000010e;
    ram_cell[     506] = 32'h000007a4;
    ram_cell[     507] = 32'h000002c5;
    ram_cell[     508] = 32'h0000053f;
    ram_cell[     509] = 32'h000000f2;
    ram_cell[     510] = 32'h000002c4;
    ram_cell[     511] = 32'h000005d8;
    ram_cell[     512] = 32'h000000fb;
    ram_cell[     513] = 32'h000006c8;
    ram_cell[     514] = 32'h0000051e;
    ram_cell[     515] = 32'h000000a2;
    ram_cell[     516] = 32'h000000f0;
    ram_cell[     517] = 32'h00000507;
    ram_cell[     518] = 32'h00000173;
    ram_cell[     519] = 32'h0000004a;
    ram_cell[     520] = 32'h00000331;
    ram_cell[     521] = 32'h00000022;
    ram_cell[     522] = 32'h00000453;
    ram_cell[     523] = 32'h0000059a;
    ram_cell[     524] = 32'h000002dc;
    ram_cell[     525] = 32'h0000015c;
    ram_cell[     526] = 32'h0000068f;
    ram_cell[     527] = 32'h00000681;
    ram_cell[     528] = 32'h00000539;
    ram_cell[     529] = 32'h0000017f;
    ram_cell[     530] = 32'h00000184;
    ram_cell[     531] = 32'h00000728;
    ram_cell[     532] = 32'h0000025a;
    ram_cell[     533] = 32'h0000033a;
    ram_cell[     534] = 32'h00000048;
    ram_cell[     535] = 32'h0000045c;
    ram_cell[     536] = 32'h0000036a;
    ram_cell[     537] = 32'h000004a4;
    ram_cell[     538] = 32'h000004c9;
    ram_cell[     539] = 32'h000005fa;
    ram_cell[     540] = 32'h0000038c;
    ram_cell[     541] = 32'h0000078d;
    ram_cell[     542] = 32'h00000417;
    ram_cell[     543] = 32'h00000347;
    ram_cell[     544] = 32'h000005cc;
    ram_cell[     545] = 32'h0000071d;
    ram_cell[     546] = 32'h000005c2;
    ram_cell[     547] = 32'h000005c9;
    ram_cell[     548] = 32'h00000747;
    ram_cell[     549] = 32'h000003bf;
    ram_cell[     550] = 32'h000004c2;
    ram_cell[     551] = 32'h0000014e;
    ram_cell[     552] = 32'h0000050a;
    ram_cell[     553] = 32'h00000482;
    ram_cell[     554] = 32'h00000056;
    ram_cell[     555] = 32'h00000438;
    ram_cell[     556] = 32'h000005c6;
    ram_cell[     557] = 32'h00000678;
    ram_cell[     558] = 32'h000003e2;
    ram_cell[     559] = 32'h00000186;
    ram_cell[     560] = 32'h0000073d;
    ram_cell[     561] = 32'h00000100;
    ram_cell[     562] = 32'h00000364;
    ram_cell[     563] = 32'h000005cf;
    ram_cell[     564] = 32'h000001e5;
    ram_cell[     565] = 32'h000004ca;
    ram_cell[     566] = 32'h000000f3;
    ram_cell[     567] = 32'h0000066e;
    ram_cell[     568] = 32'h0000052f;
    ram_cell[     569] = 32'h000006ad;
    ram_cell[     570] = 32'h000003f5;
    ram_cell[     571] = 32'h000003bb;
    ram_cell[     572] = 32'h0000007e;
    ram_cell[     573] = 32'h000006fe;
    ram_cell[     574] = 32'h000002a7;
    ram_cell[     575] = 32'h000004df;
    ram_cell[     576] = 32'h00000591;
    ram_cell[     577] = 32'h00000062;
    ram_cell[     578] = 32'h0000028d;
    ram_cell[     579] = 32'h000007d0;
    ram_cell[     580] = 32'h000003b8;
    ram_cell[     581] = 32'h0000041a;
    ram_cell[     582] = 32'h0000017a;
    ram_cell[     583] = 32'h0000020f;
    ram_cell[     584] = 32'h000003e7;
    ram_cell[     585] = 32'h00000564;
    ram_cell[     586] = 32'h00000206;
    ram_cell[     587] = 32'h00000526;
    ram_cell[     588] = 32'h000005ef;
    ram_cell[     589] = 32'h0000002b;
    ram_cell[     590] = 32'h000007f5;
    ram_cell[     591] = 32'h000003f9;
    ram_cell[     592] = 32'h00000305;
    ram_cell[     593] = 32'h000001ef;
    ram_cell[     594] = 32'h0000025b;
    ram_cell[     595] = 32'h00000722;
    ram_cell[     596] = 32'h000007d7;
    ram_cell[     597] = 32'h00000729;
    ram_cell[     598] = 32'h00000326;
    ram_cell[     599] = 32'h00000703;
    ram_cell[     600] = 32'h0000043c;
    ram_cell[     601] = 32'h000003eb;
    ram_cell[     602] = 32'h000002d5;
    ram_cell[     603] = 32'h000000ce;
    ram_cell[     604] = 32'h0000057e;
    ram_cell[     605] = 32'h00000498;
    ram_cell[     606] = 32'h000006e4;
    ram_cell[     607] = 32'h00000249;
    ram_cell[     608] = 32'h00000751;
    ram_cell[     609] = 32'h000007c5;
    ram_cell[     610] = 32'h000005a3;
    ram_cell[     611] = 32'h0000027e;
    ram_cell[     612] = 32'h000002a6;
    ram_cell[     613] = 32'h00000127;
    ram_cell[     614] = 32'h000007f4;
    ram_cell[     615] = 32'h000005ca;
    ram_cell[     616] = 32'h00000335;
    ram_cell[     617] = 32'h000000a9;
    ram_cell[     618] = 32'h000002de;
    ram_cell[     619] = 32'h000005ac;
    ram_cell[     620] = 32'h0000060f;
    ram_cell[     621] = 32'h00000515;
    ram_cell[     622] = 32'h0000019d;
    ram_cell[     623] = 32'h00000237;
    ram_cell[     624] = 32'h0000076c;
    ram_cell[     625] = 32'h00000130;
    ram_cell[     626] = 32'h00000476;
    ram_cell[     627] = 32'h00000745;
    ram_cell[     628] = 32'h0000071a;
    ram_cell[     629] = 32'h0000077a;
    ram_cell[     630] = 32'h000003af;
    ram_cell[     631] = 32'h000007fe;
    ram_cell[     632] = 32'h000006b4;
    ram_cell[     633] = 32'h00000291;
    ram_cell[     634] = 32'h00000103;
    ram_cell[     635] = 32'h00000151;
    ram_cell[     636] = 32'h0000051b;
    ram_cell[     637] = 32'h0000040d;
    ram_cell[     638] = 32'h00000137;
    ram_cell[     639] = 32'h00000702;
    ram_cell[     640] = 32'h0000021b;
    ram_cell[     641] = 32'h000004fb;
    ram_cell[     642] = 32'h0000047d;
    ram_cell[     643] = 32'h0000078f;
    ram_cell[     644] = 32'h00000407;
    ram_cell[     645] = 32'h000005db;
    ram_cell[     646] = 32'h00000314;
    ram_cell[     647] = 32'h0000075a;
    ram_cell[     648] = 32'h0000049f;
    ram_cell[     649] = 32'h00000673;
    ram_cell[     650] = 32'h000000f5;
    ram_cell[     651] = 32'h0000067e;
    ram_cell[     652] = 32'h000003e6;
    ram_cell[     653] = 32'h0000006e;
    ram_cell[     654] = 32'h000003d6;
    ram_cell[     655] = 32'h000004d6;
    ram_cell[     656] = 32'h000001b0;
    ram_cell[     657] = 32'h00000399;
    ram_cell[     658] = 32'h0000051d;
    ram_cell[     659] = 32'h0000061a;
    ram_cell[     660] = 32'h00000467;
    ram_cell[     661] = 32'h000004ba;
    ram_cell[     662] = 32'h0000015f;
    ram_cell[     663] = 32'h0000033e;
    ram_cell[     664] = 32'h000001d9;
    ram_cell[     665] = 32'h0000019a;
    ram_cell[     666] = 32'h0000062c;
    ram_cell[     667] = 32'h0000033c;
    ram_cell[     668] = 32'h0000071b;
    ram_cell[     669] = 32'h00000018;
    ram_cell[     670] = 32'h000001f0;
    ram_cell[     671] = 32'h000006c6;
    ram_cell[     672] = 32'h0000071c;
    ram_cell[     673] = 32'h000000df;
    ram_cell[     674] = 32'h00000510;
    ram_cell[     675] = 32'h0000067d;
    ram_cell[     676] = 32'h00000435;
    ram_cell[     677] = 32'h000006f9;
    ram_cell[     678] = 32'h00000502;
    ram_cell[     679] = 32'h000007c7;
    ram_cell[     680] = 32'h000003aa;
    ram_cell[     681] = 32'h000005d3;
    ram_cell[     682] = 32'h000004ed;
    ram_cell[     683] = 32'h00000087;
    ram_cell[     684] = 32'h00000053;
    ram_cell[     685] = 32'h000006c4;
    ram_cell[     686] = 32'h000005ec;
    ram_cell[     687] = 32'h00000506;
    ram_cell[     688] = 32'h000006d4;
    ram_cell[     689] = 32'h000005af;
    ram_cell[     690] = 32'h000002df;
    ram_cell[     691] = 32'h00000500;
    ram_cell[     692] = 32'h0000018d;
    ram_cell[     693] = 32'h000003ee;
    ram_cell[     694] = 32'h000005fc;
    ram_cell[     695] = 32'h00000157;
    ram_cell[     696] = 32'h00000002;
    ram_cell[     697] = 32'h00000534;
    ram_cell[     698] = 32'h000002dd;
    ram_cell[     699] = 32'h000005d7;
    ram_cell[     700] = 32'h00000172;
    ram_cell[     701] = 32'h000004ec;
    ram_cell[     702] = 32'h000004dd;
    ram_cell[     703] = 32'h000000b5;
    ram_cell[     704] = 32'h00000793;
    ram_cell[     705] = 32'h000005a0;
    ram_cell[     706] = 32'h00000461;
    ram_cell[     707] = 32'h00000177;
    ram_cell[     708] = 32'h000000ba;
    ram_cell[     709] = 32'h000001fe;
    ram_cell[     710] = 32'h0000020b;
    ram_cell[     711] = 32'h0000032e;
    ram_cell[     712] = 32'h00000252;
    ram_cell[     713] = 32'h00000760;
    ram_cell[     714] = 32'h0000021c;
    ram_cell[     715] = 32'h000006b3;
    ram_cell[     716] = 32'h00000278;
    ram_cell[     717] = 32'h00000270;
    ram_cell[     718] = 32'h00000263;
    ram_cell[     719] = 32'h000007e7;
    ram_cell[     720] = 32'h0000054d;
    ram_cell[     721] = 32'h000005b7;
    ram_cell[     722] = 32'h0000078a;
    ram_cell[     723] = 32'h00000440;
    ram_cell[     724] = 32'h0000029a;
    ram_cell[     725] = 32'h0000075c;
    ram_cell[     726] = 32'h00000089;
    ram_cell[     727] = 32'h00000330;
    ram_cell[     728] = 32'h00000715;
    ram_cell[     729] = 32'h000002f4;
    ram_cell[     730] = 32'h000000b9;
    ram_cell[     731] = 32'h000000ec;
    ram_cell[     732] = 32'h00000010;
    ram_cell[     733] = 32'h0000027c;
    ram_cell[     734] = 32'h00000139;
    ram_cell[     735] = 32'h00000082;
    ram_cell[     736] = 32'h0000018c;
    ram_cell[     737] = 32'h00000191;
    ram_cell[     738] = 32'h00000661;
    ram_cell[     739] = 32'h0000002c;
    ram_cell[     740] = 32'h0000019f;
    ram_cell[     741] = 32'h0000074c;
    ram_cell[     742] = 32'h00000225;
    ram_cell[     743] = 32'h00000414;
    ram_cell[     744] = 32'h00000710;
    ram_cell[     745] = 32'h000006bb;
    ram_cell[     746] = 32'h00000696;
    ram_cell[     747] = 32'h00000044;
    ram_cell[     748] = 32'h0000035c;
    ram_cell[     749] = 32'h000007b8;
    ram_cell[     750] = 32'h0000065a;
    ram_cell[     751] = 32'h00000351;
    ram_cell[     752] = 32'h0000000a;
    ram_cell[     753] = 32'h0000031a;
    ram_cell[     754] = 32'h00000401;
    ram_cell[     755] = 32'h0000012e;
    ram_cell[     756] = 32'h0000066b;
    ram_cell[     757] = 32'h000007d8;
    ram_cell[     758] = 32'h00000114;
    ram_cell[     759] = 32'h0000009f;
    ram_cell[     760] = 32'h00000462;
    ram_cell[     761] = 32'h00000527;
    ram_cell[     762] = 32'h00000102;
    ram_cell[     763] = 32'h00000503;
    ram_cell[     764] = 32'h00000636;
    ram_cell[     765] = 32'h000004a2;
    ram_cell[     766] = 32'h000006a0;
    ram_cell[     767] = 32'h00000723;
    ram_cell[     768] = 32'h0000060a;
    ram_cell[     769] = 32'h00000775;
    ram_cell[     770] = 32'h000005ff;
    ram_cell[     771] = 32'h0000026a;
    ram_cell[     772] = 32'h0000055b;
    ram_cell[     773] = 32'h00000549;
    ram_cell[     774] = 32'h000006dd;
    ram_cell[     775] = 32'h000003d8;
    ram_cell[     776] = 32'h000006bc;
    ram_cell[     777] = 32'h0000004d;
    ram_cell[     778] = 32'h000001bc;
    ram_cell[     779] = 32'h000007a7;
    ram_cell[     780] = 32'h00000746;
    ram_cell[     781] = 32'h00000522;
    ram_cell[     782] = 32'h000002cb;
    ram_cell[     783] = 32'h00000743;
    ram_cell[     784] = 32'h00000376;
    ram_cell[     785] = 32'h00000668;
    ram_cell[     786] = 32'h00000342;
    ram_cell[     787] = 32'h000000a3;
    ram_cell[     788] = 32'h00000155;
    ram_cell[     789] = 32'h000001a5;
    ram_cell[     790] = 32'h000005df;
    ram_cell[     791] = 32'h0000046b;
    ram_cell[     792] = 32'h0000079a;
    ram_cell[     793] = 32'h0000078e;
    ram_cell[     794] = 32'h000006ff;
    ram_cell[     795] = 32'h00000632;
    ram_cell[     796] = 32'h00000023;
    ram_cell[     797] = 32'h0000062b;
    ram_cell[     798] = 32'h000002a3;
    ram_cell[     799] = 32'h0000063a;
    ram_cell[     800] = 32'h00000321;
    ram_cell[     801] = 32'h00000119;
    ram_cell[     802] = 32'h000006c0;
    ram_cell[     803] = 32'h00000251;
    ram_cell[     804] = 32'h00000652;
    ram_cell[     805] = 32'h00000685;
    ram_cell[     806] = 32'h00000380;
    ram_cell[     807] = 32'h00000212;
    ram_cell[     808] = 32'h000007ac;
    ram_cell[     809] = 32'h00000329;
    ram_cell[     810] = 32'h000000b0;
    ram_cell[     811] = 32'h00000222;
    ram_cell[     812] = 32'h00000748;
    ram_cell[     813] = 32'h00000754;
    ram_cell[     814] = 32'h00000273;
    ram_cell[     815] = 32'h00000394;
    ram_cell[     816] = 32'h000004e6;
    ram_cell[     817] = 32'h0000070f;
    ram_cell[     818] = 32'h000001b1;
    ram_cell[     819] = 32'h00000227;
    ram_cell[     820] = 32'h00000663;
    ram_cell[     821] = 32'h0000034d;
    ram_cell[     822] = 32'h00000788;
    ram_cell[     823] = 32'h000002b9;
    ram_cell[     824] = 32'h00000088;
    ram_cell[     825] = 32'h00000373;
    ram_cell[     826] = 32'h000006e6;
    ram_cell[     827] = 32'h000005bc;
    ram_cell[     828] = 32'h0000059f;
    ram_cell[     829] = 32'h000007f8;
    ram_cell[     830] = 32'h00000544;
    ram_cell[     831] = 32'h00000413;
    ram_cell[     832] = 32'h0000021d;
    ram_cell[     833] = 32'h000002bf;
    ram_cell[     834] = 32'h00000012;
    ram_cell[     835] = 32'h00000176;
    ram_cell[     836] = 32'h0000041d;
    ram_cell[     837] = 32'h000002b8;
    ram_cell[     838] = 32'h00000039;
    ram_cell[     839] = 32'h0000049a;
    ram_cell[     840] = 32'h000005dc;
    ram_cell[     841] = 32'h000001a8;
    ram_cell[     842] = 32'h000001cc;
    ram_cell[     843] = 32'h000000d4;
    ram_cell[     844] = 32'h000007e2;
    ram_cell[     845] = 32'h00000452;
    ram_cell[     846] = 32'h00000369;
    ram_cell[     847] = 32'h0000066d;
    ram_cell[     848] = 32'h000005cd;
    ram_cell[     849] = 32'h0000010b;
    ram_cell[     850] = 32'h00000676;
    ram_cell[     851] = 32'h000005a5;
    ram_cell[     852] = 32'h00000135;
    ram_cell[     853] = 32'h0000018b;
    ram_cell[     854] = 32'h000007a3;
    ram_cell[     855] = 32'h0000077b;
    ram_cell[     856] = 32'h0000075d;
    ram_cell[     857] = 32'h00000079;
    ram_cell[     858] = 32'h00000379;
    ram_cell[     859] = 32'h00000542;
    ram_cell[     860] = 32'h00000315;
    ram_cell[     861] = 32'h00000671;
    ram_cell[     862] = 32'h0000079f;
    ram_cell[     863] = 32'h000001e4;
    ram_cell[     864] = 32'h00000215;
    ram_cell[     865] = 32'h0000033f;
    ram_cell[     866] = 32'h0000016a;
    ram_cell[     867] = 32'h00000289;
    ram_cell[     868] = 32'h0000052e;
    ram_cell[     869] = 32'h000003ef;
    ram_cell[     870] = 32'h0000014a;
    ram_cell[     871] = 32'h000007bf;
    ram_cell[     872] = 32'h00000586;
    ram_cell[     873] = 32'h000000ae;
    ram_cell[     874] = 32'h0000060e;
    ram_cell[     875] = 32'h000001bf;
    ram_cell[     876] = 32'h00000338;
    ram_cell[     877] = 32'h0000056c;
    ram_cell[     878] = 32'h000002a1;
    ram_cell[     879] = 32'h00000782;
    ram_cell[     880] = 32'h00000258;
    ram_cell[     881] = 32'h0000078b;
    ram_cell[     882] = 32'h000006c7;
    ram_cell[     883] = 32'h0000058d;
    ram_cell[     884] = 32'h000005f4;
    ram_cell[     885] = 32'h000004c3;
    ram_cell[     886] = 32'h0000046c;
    ram_cell[     887] = 32'h000006d3;
    ram_cell[     888] = 32'h0000064c;
    ram_cell[     889] = 32'h000006c2;
    ram_cell[     890] = 32'h000003b4;
    ram_cell[     891] = 32'h0000014c;
    ram_cell[     892] = 32'h00000013;
    ram_cell[     893] = 32'h0000061d;
    ram_cell[     894] = 32'h000002b7;
    ram_cell[     895] = 32'h000001ed;
    ram_cell[     896] = 32'h00000296;
    ram_cell[     897] = 32'h000004af;
    ram_cell[     898] = 32'h0000004e;
    ram_cell[     899] = 32'h00000637;
    ram_cell[     900] = 32'h000003a3;
    ram_cell[     901] = 32'h00000418;
    ram_cell[     902] = 32'h0000065e;
    ram_cell[     903] = 32'h0000007b;
    ram_cell[     904] = 32'h00000517;
    ram_cell[     905] = 32'h000000ad;
    ram_cell[     906] = 32'h0000047e;
    ram_cell[     907] = 32'h0000053a;
    ram_cell[     908] = 32'h00000006;
    ram_cell[     909] = 32'h00000644;
    ram_cell[     910] = 32'h0000073c;
    ram_cell[     911] = 32'h000001d6;
    ram_cell[     912] = 32'h00000094;
    ram_cell[     913] = 32'h00000473;
    ram_cell[     914] = 32'h00000111;
    ram_cell[     915] = 32'h000003d9;
    ram_cell[     916] = 32'h000002c2;
    ram_cell[     917] = 32'h00000618;
    ram_cell[     918] = 32'h000001ad;
    ram_cell[     919] = 32'h00000242;
    ram_cell[     920] = 32'h00000303;
    ram_cell[     921] = 32'h0000048d;
    ram_cell[     922] = 32'h00000560;
    ram_cell[     923] = 32'h00000126;
    ram_cell[     924] = 32'h000004c1;
    ram_cell[     925] = 32'h00000442;
    ram_cell[     926] = 32'h000003a9;
    ram_cell[     927] = 32'h0000039a;
    ram_cell[     928] = 32'h0000009e;
    ram_cell[     929] = 32'h00000566;
    ram_cell[     930] = 32'h0000056b;
    ram_cell[     931] = 32'h00000648;
    ram_cell[     932] = 32'h000004fc;
    ram_cell[     933] = 32'h000004cb;
    ram_cell[     934] = 32'h000004de;
    ram_cell[     935] = 32'h000002a9;
    ram_cell[     936] = 32'h00000605;
    ram_cell[     937] = 32'h0000056d;
    ram_cell[     938] = 32'h000000b1;
    ram_cell[     939] = 32'h000007c6;
    ram_cell[     940] = 32'h0000061f;
    ram_cell[     941] = 32'h00000689;
    ram_cell[     942] = 32'h000000fa;
    ram_cell[     943] = 32'h00000486;
    ram_cell[     944] = 32'h000000a7;
    ram_cell[     945] = 32'h00000456;
    ram_cell[     946] = 32'h00000471;
    ram_cell[     947] = 32'h0000064e;
    ram_cell[     948] = 32'h00000603;
    ram_cell[     949] = 32'h00000298;
    ram_cell[     950] = 32'h00000188;
    ram_cell[     951] = 32'h0000059b;
    ram_cell[     952] = 32'h000000f4;
    ram_cell[     953] = 32'h00000562;
    ram_cell[     954] = 32'h00000774;
    ram_cell[     955] = 32'h000007d1;
    ram_cell[     956] = 32'h00000017;
    ram_cell[     957] = 32'h00000392;
    ram_cell[     958] = 32'h00000348;
    ram_cell[     959] = 32'h0000038a;
    ram_cell[     960] = 32'h00000650;
    ram_cell[     961] = 32'h000004a1;
    ram_cell[     962] = 32'h000003dc;
    ram_cell[     963] = 32'h0000012b;
    ram_cell[     964] = 32'h0000061e;
    ram_cell[     965] = 32'h0000027d;
    ram_cell[     966] = 32'h0000017e;
    ram_cell[     967] = 32'h00000790;
    ram_cell[     968] = 32'h0000002d;
    ram_cell[     969] = 32'h000000f7;
    ram_cell[     970] = 32'h00000724;
    ram_cell[     971] = 32'h000003de;
    ram_cell[     972] = 32'h000007cd;
    ram_cell[     973] = 32'h000003d0;
    ram_cell[     974] = 32'h00000721;
    ram_cell[     975] = 32'h000001b8;
    ram_cell[     976] = 32'h00000286;
    ram_cell[     977] = 32'h0000024d;
    ram_cell[     978] = 32'h00000028;
    ram_cell[     979] = 32'h000006d8;
    ram_cell[     980] = 32'h0000048a;
    ram_cell[     981] = 32'h00000769;
    ram_cell[     982] = 32'h00000582;
    ram_cell[     983] = 32'h00000368;
    ram_cell[     984] = 32'h000004d5;
    ram_cell[     985] = 32'h0000022c;
    ram_cell[     986] = 32'h00000156;
    ram_cell[     987] = 32'h0000036f;
    ram_cell[     988] = 32'h00000343;
    ram_cell[     989] = 32'h00000210;
    ram_cell[     990] = 32'h000001c0;
    ram_cell[     991] = 32'h000003c9;
    ram_cell[     992] = 32'h000007fd;
    ram_cell[     993] = 32'h000002e2;
    ram_cell[     994] = 32'h0000030e;
    ram_cell[     995] = 32'h00000457;
    ram_cell[     996] = 32'h00000444;
    ram_cell[     997] = 32'h000001f2;
    ram_cell[     998] = 32'h00000353;
    ram_cell[     999] = 32'h0000016b;
    ram_cell[    1000] = 32'h00000677;
    ram_cell[    1001] = 32'h00000133;
    ram_cell[    1002] = 32'h00000613;
    ram_cell[    1003] = 32'h00000352;
    ram_cell[    1004] = 32'h00000334;
    ram_cell[    1005] = 32'h000004aa;
    ram_cell[    1006] = 32'h000001f3;
    ram_cell[    1007] = 32'h00000221;
    ram_cell[    1008] = 32'h0000037c;
    ram_cell[    1009] = 32'h000007cf;
    ram_cell[    1010] = 32'h000001aa;
    ram_cell[    1011] = 32'h0000033d;
    ram_cell[    1012] = 32'h000005d5;
    ram_cell[    1013] = 32'h000003d2;
    ram_cell[    1014] = 32'h0000040b;
    ram_cell[    1015] = 32'h0000010c;
    ram_cell[    1016] = 32'h0000046a;
    ram_cell[    1017] = 32'h00000297;
    ram_cell[    1018] = 32'h00000478;
    ram_cell[    1019] = 32'h0000055f;
    ram_cell[    1020] = 32'h00000595;
    ram_cell[    1021] = 32'h000004a7;
    ram_cell[    1022] = 32'h0000024f;
    ram_cell[    1023] = 32'h0000073e;
    ram_cell[    1024] = 32'h000004f4;
    ram_cell[    1025] = 32'h000001a7;
    ram_cell[    1026] = 32'h0000005f;
    ram_cell[    1027] = 32'h000007fa;
    ram_cell[    1028] = 32'h00000397;
    ram_cell[    1029] = 32'h00000585;
    ram_cell[    1030] = 32'h0000020a;
    ram_cell[    1031] = 32'h000004f2;
    ram_cell[    1032] = 32'h000000c3;
    ram_cell[    1033] = 32'h00000783;
    ram_cell[    1034] = 32'h000005f3;
    ram_cell[    1035] = 32'h000002a2;
    ram_cell[    1036] = 32'h00000055;
    ram_cell[    1037] = 32'h00000393;
    ram_cell[    1038] = 32'h00000007;
    ram_cell[    1039] = 32'h00000451;
    ram_cell[    1040] = 32'h00000113;
    ram_cell[    1041] = 32'h000006d5;
    ram_cell[    1042] = 32'h000006cb;
    ram_cell[    1043] = 32'h000005fb;
    ram_cell[    1044] = 32'h00000645;
    ram_cell[    1045] = 32'h000004d1;
    ram_cell[    1046] = 32'h000002f7;
    ram_cell[    1047] = 32'h0000060c;
    ram_cell[    1048] = 32'h0000054c;
    ram_cell[    1049] = 32'h00000323;
    ram_cell[    1050] = 32'h000005e5;
    ram_cell[    1051] = 32'h000004f8;
    ram_cell[    1052] = 32'h00000638;
    ram_cell[    1053] = 32'h0000013d;
    ram_cell[    1054] = 32'h000000c7;
    ram_cell[    1055] = 32'h00000052;
    ram_cell[    1056] = 32'h0000070b;
    ram_cell[    1057] = 32'h000000a1;
    ram_cell[    1058] = 32'h0000050c;
    ram_cell[    1059] = 32'h00000468;
    ram_cell[    1060] = 32'h00000083;
    ram_cell[    1061] = 32'h00000061;
    ram_cell[    1062] = 32'h000007fb;
    ram_cell[    1063] = 32'h0000011d;
    ram_cell[    1064] = 32'h000002ea;
    ram_cell[    1065] = 32'h00000123;
    ram_cell[    1066] = 32'h000003fb;
    ram_cell[    1067] = 32'h00000525;
    ram_cell[    1068] = 32'h000001d4;
    ram_cell[    1069] = 32'h0000024e;
    ram_cell[    1070] = 32'h00000572;
    ram_cell[    1071] = 32'h0000031c;
    ram_cell[    1072] = 32'h000003b7;
    ram_cell[    1073] = 32'h000002d7;
    ram_cell[    1074] = 32'h00000284;
    ram_cell[    1075] = 32'h0000001d;
    ram_cell[    1076] = 32'h000005e8;
    ram_cell[    1077] = 32'h0000013f;
    ram_cell[    1078] = 32'h00000529;
    ram_cell[    1079] = 32'h000000f8;
    ram_cell[    1080] = 32'h000002e1;
    ram_cell[    1081] = 32'h0000005c;
    ram_cell[    1082] = 32'h000004b1;
    ram_cell[    1083] = 32'h000001d5;
    ram_cell[    1084] = 32'h000004ad;
    ram_cell[    1085] = 32'h00000426;
    ram_cell[    1086] = 32'h000007c9;
    ram_cell[    1087] = 32'h000002a8;
    ram_cell[    1088] = 32'h00000205;
    ram_cell[    1089] = 32'h000002ae;
    ram_cell[    1090] = 32'h000002b4;
    ram_cell[    1091] = 32'h00000755;
    ram_cell[    1092] = 32'h0000041f;
    ram_cell[    1093] = 32'h000003cd;
    ram_cell[    1094] = 32'h000002eb;
    ram_cell[    1095] = 32'h000001a6;
    ram_cell[    1096] = 32'h00000248;
    ram_cell[    1097] = 32'h000003a5;
    ram_cell[    1098] = 32'h0000044d;
    ram_cell[    1099] = 32'h0000031b;
    ram_cell[    1100] = 32'h00000590;
    ram_cell[    1101] = 32'h0000055d;
    ram_cell[    1102] = 32'h000003b5;
    ram_cell[    1103] = 32'h00000294;
    ram_cell[    1104] = 32'h00000234;
    ram_cell[    1105] = 32'h0000016f;
    ram_cell[    1106] = 32'h000000cc;
    ram_cell[    1107] = 32'h000002cd;
    ram_cell[    1108] = 32'h00000795;
    ram_cell[    1109] = 32'h0000022e;
    ram_cell[    1110] = 32'h0000032d;
    ram_cell[    1111] = 32'h000000d8;
    ram_cell[    1112] = 32'h00000049;
    ram_cell[    1113] = 32'h00000268;
    ram_cell[    1114] = 32'h00000051;
    ram_cell[    1115] = 32'h0000001a;
    ram_cell[    1116] = 32'h00000487;
    ram_cell[    1117] = 32'h000002ec;
    ram_cell[    1118] = 32'h000002f6;
    ram_cell[    1119] = 32'h0000000e;
    ram_cell[    1120] = 32'h000000bb;
    ram_cell[    1121] = 32'h000003c6;
    ram_cell[    1122] = 32'h00000739;
    ram_cell[    1123] = 32'h0000011f;
    ram_cell[    1124] = 32'h000006e1;
    ram_cell[    1125] = 32'h000006a1;
    ram_cell[    1126] = 32'h00000665;
    ram_cell[    1127] = 32'h00000312;
    ram_cell[    1128] = 32'h00000786;
    ram_cell[    1129] = 32'h0000013e;
    ram_cell[    1130] = 32'h000007e8;
    ram_cell[    1131] = 32'h000002e3;
    ram_cell[    1132] = 32'h00000259;
    ram_cell[    1133] = 32'h00000767;
    ram_cell[    1134] = 32'h000004b6;
    ram_cell[    1135] = 32'h00000168;
    ram_cell[    1136] = 32'h0000059c;
    ram_cell[    1137] = 32'h0000000f;
    ram_cell[    1138] = 32'h00000516;
    ram_cell[    1139] = 32'h00000143;
    ram_cell[    1140] = 32'h000006af;
    ram_cell[    1141] = 32'h000002db;
    ram_cell[    1142] = 32'h00000016;
    ram_cell[    1143] = 32'h00000378;
    ram_cell[    1144] = 32'h000002fb;
    ram_cell[    1145] = 32'h000000e6;
    ram_cell[    1146] = 32'h0000036c;
    ram_cell[    1147] = 32'h00000627;
    ram_cell[    1148] = 32'h0000076a;
    ram_cell[    1149] = 32'h000003f1;
    ram_cell[    1150] = 32'h0000039d;
    ram_cell[    1151] = 32'h0000050b;
    ram_cell[    1152] = 32'h00000272;
    ram_cell[    1153] = 32'h00000360;
    ram_cell[    1154] = 32'h000007c3;
    ram_cell[    1155] = 32'h00000705;
    ram_cell[    1156] = 32'h00000692;
    ram_cell[    1157] = 32'h000006b0;
    ram_cell[    1158] = 32'h000001f7;
    ram_cell[    1159] = 32'h00000063;
    ram_cell[    1160] = 32'h0000050d;
    ram_cell[    1161] = 32'h0000072a;
    ram_cell[    1162] = 32'h00000045;
    ram_cell[    1163] = 32'h000007e9;
    ram_cell[    1164] = 32'h000000ed;
    ram_cell[    1165] = 32'h000000e1;
    ram_cell[    1166] = 32'h0000025f;
    ram_cell[    1167] = 32'h000005f1;
    ram_cell[    1168] = 32'h000002ba;
    ram_cell[    1169] = 32'h000004b8;
    ram_cell[    1170] = 32'h00000032;
    ram_cell[    1171] = 32'h000000c6;
    ram_cell[    1172] = 32'h00000640;
    ram_cell[    1173] = 32'h00000772;
    ram_cell[    1174] = 32'h0000010f;
    ram_cell[    1175] = 32'h00000085;
    ram_cell[    1176] = 32'h000007a8;
    ram_cell[    1177] = 32'h00000429;
    ram_cell[    1178] = 32'h000001a9;
    ram_cell[    1179] = 32'h00000107;
    ram_cell[    1180] = 32'h000001c7;
    ram_cell[    1181] = 32'h000004db;
    ram_cell[    1182] = 32'h000004eb;
    ram_cell[    1183] = 32'h00000374;
    ram_cell[    1184] = 32'h00000524;
    ram_cell[    1185] = 32'h000007bd;
    ram_cell[    1186] = 32'h0000026f;
    ram_cell[    1187] = 32'h000001e6;
    ram_cell[    1188] = 32'h00000163;
    ram_cell[    1189] = 32'h00000466;
    ram_cell[    1190] = 32'h0000035e;
    ram_cell[    1191] = 32'h0000030c;
    ram_cell[    1192] = 32'h00000690;
    ram_cell[    1193] = 32'h0000049c;
    ram_cell[    1194] = 32'h000003ae;
    ram_cell[    1195] = 32'h000002f3;
    ram_cell[    1196] = 32'h0000066c;
    ram_cell[    1197] = 32'h000003ce;
    ram_cell[    1198] = 32'h000003c3;
    ram_cell[    1199] = 32'h000003f7;
    ram_cell[    1200] = 32'h000007ba;
    ram_cell[    1201] = 32'h00000344;
    ram_cell[    1202] = 32'h000002fa;
    ram_cell[    1203] = 32'h00000402;
    ram_cell[    1204] = 32'h0000054e;
    ram_cell[    1205] = 32'h0000004f;
    ram_cell[    1206] = 32'h00000614;
    ram_cell[    1207] = 32'h0000033b;
    ram_cell[    1208] = 32'h00000153;
    ram_cell[    1209] = 32'h00000207;
    ram_cell[    1210] = 32'h00000520;
    ram_cell[    1211] = 32'h000006b2;
    ram_cell[    1212] = 32'h0000042c;
    ram_cell[    1213] = 32'h0000037a;
    ram_cell[    1214] = 32'h0000010a;
    ram_cell[    1215] = 32'h000007ef;
    ram_cell[    1216] = 32'h000001a3;
    ram_cell[    1217] = 32'h0000046e;
    ram_cell[    1218] = 32'h000001ab;
    ram_cell[    1219] = 32'h00000202;
    ram_cell[    1220] = 32'h000005b6;
    ram_cell[    1221] = 32'h000004bc;
    ram_cell[    1222] = 32'h00000616;
    ram_cell[    1223] = 32'h00000744;
    ram_cell[    1224] = 32'h0000040e;
    ram_cell[    1225] = 32'h00000396;
    ram_cell[    1226] = 32'h000003ff;
    ram_cell[    1227] = 32'h000002ab;
    ram_cell[    1228] = 32'h000002c3;
    ram_cell[    1229] = 32'h000003ec;
    ram_cell[    1230] = 32'h000004e4;
    ram_cell[    1231] = 32'h000004c6;
    ram_cell[    1232] = 32'h000004cc;
    ram_cell[    1233] = 32'h0000040f;
    ram_cell[    1234] = 32'h00000654;
    ram_cell[    1235] = 32'h000000c9;
    ram_cell[    1236] = 32'h00000226;
    ram_cell[    1237] = 32'h00000763;
    ram_cell[    1238] = 32'h0000058a;
    ram_cell[    1239] = 32'h0000075e;
    ram_cell[    1240] = 32'h0000063c;
    ram_cell[    1241] = 32'h000007e1;
    ram_cell[    1242] = 32'h0000071e;
    ram_cell[    1243] = 32'h0000030b;
    ram_cell[    1244] = 32'h000001d0;
    ram_cell[    1245] = 32'h000000a4;
    ram_cell[    1246] = 32'h000006be;
    ram_cell[    1247] = 32'h00000631;
    ram_cell[    1248] = 32'h00000346;
    ram_cell[    1249] = 32'h000003d1;
    ram_cell[    1250] = 32'h00000254;
    ram_cell[    1251] = 32'h000002fd;
    ram_cell[    1252] = 32'h000005f2;
    ram_cell[    1253] = 32'h000006e9;
    ram_cell[    1254] = 32'h00000469;
    ram_cell[    1255] = 32'h0000059d;
    ram_cell[    1256] = 32'h000002b5;
    ram_cell[    1257] = 32'h0000063f;
    ram_cell[    1258] = 32'h000003f0;
    ram_cell[    1259] = 32'h000005f6;
    ram_cell[    1260] = 32'h000007e0;
    ram_cell[    1261] = 32'h00000662;
    ram_cell[    1262] = 32'h000003b1;
    ram_cell[    1263] = 32'h000006e8;
    ram_cell[    1264] = 32'h0000007c;
    ram_cell[    1265] = 32'h00000480;
    ram_cell[    1266] = 32'h0000023c;
    ram_cell[    1267] = 32'h00000105;
    ram_cell[    1268] = 32'h000004cf;
    ram_cell[    1269] = 32'h00000596;
    ram_cell[    1270] = 32'h00000269;
    ram_cell[    1271] = 32'h00000670;
    ram_cell[    1272] = 32'h00000336;
    ram_cell[    1273] = 32'h000000a5;
    ram_cell[    1274] = 32'h00000073;
    ram_cell[    1275] = 32'h00000698;
    ram_cell[    1276] = 32'h00000750;
    ram_cell[    1277] = 32'h0000043f;
    ram_cell[    1278] = 32'h0000076e;
    ram_cell[    1279] = 32'h0000002a;
    ram_cell[    1280] = 32'h00000602;
    ram_cell[    1281] = 32'h00000691;
    ram_cell[    1282] = 32'h00000789;
    ram_cell[    1283] = 32'h00000762;
    ram_cell[    1284] = 32'h0000046f;
    ram_cell[    1285] = 32'h00000761;
    ram_cell[    1286] = 32'h000005e2;
    ram_cell[    1287] = 32'h000004c0;
    ram_cell[    1288] = 32'h0000006f;
    ram_cell[    1289] = 32'h000003bc;
    ram_cell[    1290] = 32'h00000736;
    ram_cell[    1291] = 32'h0000026b;
    ram_cell[    1292] = 32'h000003a7;
    ram_cell[    1293] = 32'h000006f4;
    ram_cell[    1294] = 32'h000001da;
    ram_cell[    1295] = 32'h00000528;
    ram_cell[    1296] = 32'h00000730;
    ram_cell[    1297] = 32'h0000044c;
    ram_cell[    1298] = 32'h00000371;
    ram_cell[    1299] = 32'h00000655;
    ram_cell[    1300] = 32'h000005bf;
    ram_cell[    1301] = 32'h000001f5;
    ram_cell[    1302] = 32'h000001db;
    ram_cell[    1303] = 32'h0000026c;
    ram_cell[    1304] = 32'h000000cf;
    ram_cell[    1305] = 32'h000006fd;
    ram_cell[    1306] = 32'h0000047c;
    ram_cell[    1307] = 32'h00000680;
    ram_cell[    1308] = 32'h0000037d;
    ram_cell[    1309] = 32'h00000276;
    ram_cell[    1310] = 32'h0000067f;
    ram_cell[    1311] = 32'h0000014b;
    ram_cell[    1312] = 32'h00000075;
    ram_cell[    1313] = 32'h000003c2;
    ram_cell[    1314] = 32'h0000047b;
    ram_cell[    1315] = 32'h00000489;
    ram_cell[    1316] = 32'h00000460;
    ram_cell[    1317] = 32'h00000050;
    ram_cell[    1318] = 32'h000005e3;
    ram_cell[    1319] = 32'h0000000b;
    ram_cell[    1320] = 32'h000006dc;
    ram_cell[    1321] = 32'h00000737;
    ram_cell[    1322] = 32'h00000433;
    ram_cell[    1323] = 32'h00000732;
    ram_cell[    1324] = 32'h00000339;
    ram_cell[    1325] = 32'h0000073b;
    ram_cell[    1326] = 32'h000003a8;
    ram_cell[    1327] = 32'h00000470;
    ram_cell[    1328] = 32'h000007c0;
    ram_cell[    1329] = 32'h00000159;
    ram_cell[    1330] = 32'h00000785;
    ram_cell[    1331] = 32'h00000086;
    ram_cell[    1332] = 32'h00000141;
    ram_cell[    1333] = 32'h00000425;
    ram_cell[    1334] = 32'h0000018a;
    ram_cell[    1335] = 32'h00000472;
    ram_cell[    1336] = 32'h00000319;
    ram_cell[    1337] = 32'h000007ed;
    ram_cell[    1338] = 32'h000003d5;
    ram_cell[    1339] = 32'h000000fe;
    ram_cell[    1340] = 32'h0000047a;
    ram_cell[    1341] = 32'h00000639;
    ram_cell[    1342] = 32'h00000536;
    ram_cell[    1343] = 32'h00000385;
    ram_cell[    1344] = 32'h000005cb;
    ram_cell[    1345] = 32'h00000029;
    ram_cell[    1346] = 32'h00000236;
    ram_cell[    1347] = 32'h00000386;
    ram_cell[    1348] = 32'h00000441;
    ram_cell[    1349] = 32'h00000408;
    ram_cell[    1350] = 32'h00000716;
    ram_cell[    1351] = 32'h000004a8;
    ram_cell[    1352] = 32'h0000068b;
    ram_cell[    1353] = 32'h000004fe;
    ram_cell[    1354] = 32'h000004e8;
    ram_cell[    1355] = 32'h0000027f;
    ram_cell[    1356] = 32'h000001b5;
    ram_cell[    1357] = 32'h0000074f;
    ram_cell[    1358] = 32'h0000064f;
    ram_cell[    1359] = 32'h000005b3;
    ram_cell[    1360] = 32'h000003db;
    ram_cell[    1361] = 32'h00000060;
    ram_cell[    1362] = 32'h000005b2;
    ram_cell[    1363] = 32'h00000719;
    ram_cell[    1364] = 32'h00000078;
    ram_cell[    1365] = 32'h0000072c;
    ram_cell[    1366] = 32'h000005c5;
    ram_cell[    1367] = 32'h000005ae;
    ram_cell[    1368] = 32'h000004a5;
    ram_cell[    1369] = 32'h00000197;
    ram_cell[    1370] = 32'h00000367;
    ram_cell[    1371] = 32'h000004bf;
    ram_cell[    1372] = 32'h000000cb;
    ram_cell[    1373] = 32'h00000080;
    ram_cell[    1374] = 32'h00000465;
    ram_cell[    1375] = 32'h0000002f;
    ram_cell[    1376] = 32'h0000025c;
    ram_cell[    1377] = 32'h00000764;
    ram_cell[    1378] = 32'h0000069c;
    ram_cell[    1379] = 32'h00000556;
    ram_cell[    1380] = 32'h0000079e;
    ram_cell[    1381] = 32'h00000349;
    ram_cell[    1382] = 32'h000007be;
    ram_cell[    1383] = 32'h000007f1;
    ram_cell[    1384] = 32'h0000008d;
    ram_cell[    1385] = 32'h000002b3;
    ram_cell[    1386] = 32'h000005c0;
    ram_cell[    1387] = 32'h0000043d;
    ram_cell[    1388] = 32'h00000144;
    ram_cell[    1389] = 32'h00000101;
    ram_cell[    1390] = 32'h000006e7;
    ram_cell[    1391] = 32'h000004e5;
    ram_cell[    1392] = 32'h00000383;
    ram_cell[    1393] = 32'h000006b6;
    ram_cell[    1394] = 32'h000001c9;
    ram_cell[    1395] = 32'h00000604;
    ram_cell[    1396] = 32'h00000756;
    ram_cell[    1397] = 32'h0000075b;
    ram_cell[    1398] = 32'h000003ab;
    ram_cell[    1399] = 32'h00000388;
    ram_cell[    1400] = 32'h000000e7;
    ram_cell[    1401] = 32'h00000026;
    ram_cell[    1402] = 32'h0000041c;
    ram_cell[    1403] = 32'h00000064;
    ram_cell[    1404] = 32'h000000fc;
    ram_cell[    1405] = 32'h00000615;
    ram_cell[    1406] = 32'h000007ad;
    ram_cell[    1407] = 32'h00000121;
    ram_cell[    1408] = 32'h00000231;
    ram_cell[    1409] = 32'h000007c4;
    ram_cell[    1410] = 32'h000006c3;
    ram_cell[    1411] = 32'h00000377;
    ram_cell[    1412] = 32'h000006de;
    ram_cell[    1413] = 32'h00000218;
    ram_cell[    1414] = 32'h0000057c;
    ram_cell[    1415] = 32'h000002ed;
    ram_cell[    1416] = 32'h0000045a;
    ram_cell[    1417] = 32'h00000395;
    ram_cell[    1418] = 32'h0000052c;
    ram_cell[    1419] = 32'h00000479;
    ram_cell[    1420] = 32'h000002c0;
    ram_cell[    1421] = 32'h0000003e;
    ram_cell[    1422] = 32'h000001e1;
    ram_cell[    1423] = 32'h000003f2;
    ram_cell[    1424] = 32'h00000072;
    ram_cell[    1425] = 32'h000006ba;
    ram_cell[    1426] = 32'h000007a9;
    ram_cell[    1427] = 32'h00000384;
    ram_cell[    1428] = 32'h00000504;
    ram_cell[    1429] = 32'h000000eb;
    ram_cell[    1430] = 32'h000007c1;
    ram_cell[    1431] = 32'h000002fe;
    ram_cell[    1432] = 32'h00000162;
    ram_cell[    1433] = 32'h0000009d;
    ram_cell[    1434] = 32'h0000048c;
    ram_cell[    1435] = 32'h00000150;
    ram_cell[    1436] = 32'h0000077c;
    ram_cell[    1437] = 32'h000006a6;
    ram_cell[    1438] = 32'h00000363;
    ram_cell[    1439] = 32'h00000214;
    ram_cell[    1440] = 32'h000003e1;
    ram_cell[    1441] = 32'h00000332;
    ram_cell[    1442] = 32'h0000074e;
    ram_cell[    1443] = 32'h000006d6;
    ram_cell[    1444] = 32'h0000009a;
    ram_cell[    1445] = 32'h00000532;
    ram_cell[    1446] = 32'h000000d0;
    ram_cell[    1447] = 32'h0000053c;
    ram_cell[    1448] = 32'h00000463;
    ram_cell[    1449] = 32'h000006ee;
    ram_cell[    1450] = 32'h00000791;
    ram_cell[    1451] = 32'h0000015b;
    ram_cell[    1452] = 32'h000001f9;
    ram_cell[    1453] = 32'h000003c0;
    ram_cell[    1454] = 32'h00000563;
    ram_cell[    1455] = 32'h000001d3;
    ram_cell[    1456] = 32'h00000492;
    ram_cell[    1457] = 32'h00000635;
    ram_cell[    1458] = 32'h00000642;
    ram_cell[    1459] = 32'h00000138;
    ram_cell[    1460] = 32'h0000062d;
    ram_cell[    1461] = 32'h000007b2;
    ram_cell[    1462] = 32'h0000025e;
    ram_cell[    1463] = 32'h0000041b;
    ram_cell[    1464] = 32'h000007b7;
    ram_cell[    1465] = 32'h00000047;
    ram_cell[    1466] = 32'h00000038;
    ram_cell[    1467] = 32'h000001ec;
    ram_cell[    1468] = 32'h00000430;
    ram_cell[    1469] = 32'h00000679;
    ram_cell[    1470] = 32'h00000256;
    ram_cell[    1471] = 32'h00000132;
    ram_cell[    1472] = 32'h000003b0;
    ram_cell[    1473] = 32'h000001b4;
    ram_cell[    1474] = 32'h0000007f;
    ram_cell[    1475] = 32'h00000675;
    ram_cell[    1476] = 32'h000004f1;
    ram_cell[    1477] = 32'h00000129;
    ram_cell[    1478] = 32'h000002a0;
    ram_cell[    1479] = 32'h000004d0;
    ram_cell[    1480] = 32'h000004f3;
    ram_cell[    1481] = 32'h000002f8;
    ram_cell[    1482] = 32'h00000419;
    ram_cell[    1483] = 32'h00000244;
    ram_cell[    1484] = 32'h000002bd;
    ram_cell[    1485] = 32'h00000290;
    ram_cell[    1486] = 32'h0000021e;
    ram_cell[    1487] = 32'h00000672;
    ram_cell[    1488] = 32'h00000169;
    ram_cell[    1489] = 32'h00000069;
    ram_cell[    1490] = 32'h0000029d;
    ram_cell[    1491] = 32'h0000057d;
    ram_cell[    1492] = 32'h000000b8;
    ram_cell[    1493] = 32'h00000001;
    ram_cell[    1494] = 32'h0000030f;
    ram_cell[    1495] = 32'h00000530;
    ram_cell[    1496] = 32'h00000220;
    ram_cell[    1497] = 32'h000003f3;
    ram_cell[    1498] = 32'h00000020;
    ram_cell[    1499] = 32'h000002af;
    ram_cell[    1500] = 32'h0000060d;
    ram_cell[    1501] = 32'h000007b6;
    ram_cell[    1502] = 32'h000003da;
    ram_cell[    1503] = 32'h0000014d;
    ram_cell[    1504] = 32'h00000584;
    ram_cell[    1505] = 32'h000005a8;
    ram_cell[    1506] = 32'h00000694;
    ram_cell[    1507] = 32'h0000042d;
    ram_cell[    1508] = 32'h00000280;
    ram_cell[    1509] = 32'h000002ee;
    ram_cell[    1510] = 32'h000007ea;
    ram_cell[    1511] = 32'h000007aa;
    ram_cell[    1512] = 32'h000003a0;
    ram_cell[    1513] = 32'h000006aa;
    ram_cell[    1514] = 32'h00000021;
    ram_cell[    1515] = 32'h00000434;
    ram_cell[    1516] = 32'h0000065b;
    ram_cell[    1517] = 32'h00000781;
    ram_cell[    1518] = 32'h0000031e;
    ram_cell[    1519] = 32'h00000096;
    ram_cell[    1520] = 32'h000001ce;
    ram_cell[    1521] = 32'h000000de;
    ram_cell[    1522] = 32'h000001a1;
    ram_cell[    1523] = 32'h00000274;
    ram_cell[    1524] = 32'h00000428;
    ram_cell[    1525] = 32'h000001f1;
    ram_cell[    1526] = 32'h000005aa;
    ram_cell[    1527] = 32'h000004e3;
    ram_cell[    1528] = 32'h00000574;
    ram_cell[    1529] = 32'h00000669;
    ram_cell[    1530] = 32'h00000612;
    ram_cell[    1531] = 32'h00000076;
    ram_cell[    1532] = 32'h000005e0;
    ram_cell[    1533] = 32'h00000512;
    ram_cell[    1534] = 32'h000004dc;
    ram_cell[    1535] = 32'h00000366;
    ram_cell[    1536] = 32'h0000044a;
    ram_cell[    1537] = 32'h000002ef;
    ram_cell[    1538] = 32'h000003b9;
    ram_cell[    1539] = 32'h000005eb;
    ram_cell[    1540] = 32'h00000628;
    ram_cell[    1541] = 32'h000003c1;
    ram_cell[    1542] = 32'h0000022f;
    ram_cell[    1543] = 32'h00000797;
    ram_cell[    1544] = 32'h00000422;
    ram_cell[    1545] = 32'h00000589;
    ram_cell[    1546] = 32'h000001cb;
    ram_cell[    1547] = 32'h000004b0;
    ram_cell[    1548] = 32'h00000733;
    ram_cell[    1549] = 32'h00000217;
    ram_cell[    1550] = 32'h00000437;
    ram_cell[    1551] = 32'h0000020c;
    ram_cell[    1552] = 32'h00000436;
    ram_cell[    1553] = 32'h00000656;
    ram_cell[    1554] = 32'h000005e7;
    ram_cell[    1555] = 32'h00000540;
    ram_cell[    1556] = 32'h00000474;
    ram_cell[    1557] = 32'h00000250;
    ram_cell[    1558] = 32'h00000195;
    ram_cell[    1559] = 32'h00000058;
    ram_cell[    1560] = 32'h000002cc;
    ram_cell[    1561] = 32'h000000c2;
    ram_cell[    1562] = 32'h00000588;
    ram_cell[    1563] = 32'h0000058b;
    ram_cell[    1564] = 32'h00000713;
    ram_cell[    1565] = 32'h000004b9;
    ram_cell[    1566] = 32'h00000727;
    ram_cell[    1567] = 32'h0000013c;
    ram_cell[    1568] = 32'h0000069e;
    ram_cell[    1569] = 32'h00000577;
    ram_cell[    1570] = 32'h000003e3;
    ram_cell[    1571] = 32'h00000391;
    ram_cell[    1572] = 32'h000005f0;
    ram_cell[    1573] = 32'h00000594;
    ram_cell[    1574] = 32'h0000037e;
    ram_cell[    1575] = 32'h0000026d;
    ram_cell[    1576] = 32'h00000361;
    ram_cell[    1577] = 32'h0000022d;
    ram_cell[    1578] = 32'h00000104;
    ram_cell[    1579] = 32'h00000266;
    ram_cell[    1580] = 32'h0000074d;
    ram_cell[    1581] = 32'h0000054a;
    ram_cell[    1582] = 32'h000000af;
    ram_cell[    1583] = 32'h00000070;
    ram_cell[    1584] = 32'h0000061b;
    ram_cell[    1585] = 32'h000003d7;
    ram_cell[    1586] = 32'h000003d4;
    ram_cell[    1587] = 32'h00000005;
    ram_cell[    1588] = 32'h00000035;
    ram_cell[    1589] = 32'h00000097;
    ram_cell[    1590] = 32'h000005ee;
    ram_cell[    1591] = 32'h00000042;
    ram_cell[    1592] = 32'h000000be;
    ram_cell[    1593] = 32'h00000712;
    ram_cell[    1594] = 32'h000004e1;
    ram_cell[    1595] = 32'h00000208;
    ram_cell[    1596] = 32'h000006c5;
    ram_cell[    1597] = 32'h00000164;
    ram_cell[    1598] = 32'h00000711;
    ram_cell[    1599] = 32'h0000064a;
    ram_cell[    1600] = 32'h0000054f;
    ram_cell[    1601] = 32'h0000011b;
    ram_cell[    1602] = 32'h000000c0;
    ram_cell[    1603] = 32'h00000008;
    ram_cell[    1604] = 32'h000006ce;
    ram_cell[    1605] = 32'h000000b3;
    ram_cell[    1606] = 32'h0000044b;
    ram_cell[    1607] = 32'h0000074b;
    ram_cell[    1608] = 32'h000004ab;
    ram_cell[    1609] = 32'h00000115;
    ram_cell[    1610] = 32'h00000448;
    ram_cell[    1611] = 32'h00000766;
    ram_cell[    1612] = 32'h00000587;
    ram_cell[    1613] = 32'h00000475;
    ram_cell[    1614] = 32'h00000255;
    ram_cell[    1615] = 32'h0000062e;
    ram_cell[    1616] = 32'h000004d3;
    ram_cell[    1617] = 32'h00000285;
    ram_cell[    1618] = 32'h000004f7;
    ram_cell[    1619] = 32'h000003ba;
    ram_cell[    1620] = 32'h0000070a;
    ram_cell[    1621] = 32'h0000069d;
    ram_cell[    1622] = 32'h000000ee;
    ram_cell[    1623] = 32'h00000514;
    ram_cell[    1624] = 32'h0000074a;
    ram_cell[    1625] = 32'h00000375;
    ram_cell[    1626] = 32'h0000072f;
    ram_cell[    1627] = 32'h00000523;
    ram_cell[    1628] = 32'h000003cb;
    ram_cell[    1629] = 32'h000000e4;
    ram_cell[    1630] = 32'h0000004c;
    ram_cell[    1631] = 32'h00000610;
    ram_cell[    1632] = 32'h00000400;
    ram_cell[    1633] = 32'h00000406;
    ram_cell[    1634] = 32'h000004ea;
    ram_cell[    1635] = 32'h00000592;
    ram_cell[    1636] = 32'h00000799;
    ram_cell[    1637] = 32'h0000024c;
    ram_cell[    1638] = 32'h0000011a;
    ram_cell[    1639] = 32'h000002f9;
    ram_cell[    1640] = 32'h0000039f;
    ram_cell[    1641] = 32'h000002b6;
    ram_cell[    1642] = 32'h00000599;
    ram_cell[    1643] = 32'h00000623;
    ram_cell[    1644] = 32'h000004ef;
    ram_cell[    1645] = 32'h000007b0;
    ram_cell[    1646] = 32'h000007f2;
    ram_cell[    1647] = 32'h0000008a;
    ram_cell[    1648] = 32'h0000079d;
    ram_cell[    1649] = 32'h000002ca;
    ram_cell[    1650] = 32'h00000112;
    ram_cell[    1651] = 32'h00000160;
    ram_cell[    1652] = 32'h0000006a;
    ram_cell[    1653] = 32'h000000e8;
    ram_cell[    1654] = 32'h000002ff;
    ram_cell[    1655] = 32'h000002f0;
    ram_cell[    1656] = 32'h00000043;
    ram_cell[    1657] = 32'h00000033;
    ram_cell[    1658] = 32'h0000055a;
    ram_cell[    1659] = 32'h00000357;
    ram_cell[    1660] = 32'h000006d0;
    ram_cell[    1661] = 32'h0000057f;
    ram_cell[    1662] = 32'h00000091;
    ram_cell[    1663] = 32'h000007a6;
    ram_cell[    1664] = 32'h0000042b;
    ram_cell[    1665] = 32'h00000359;
    ram_cell[    1666] = 32'h000002c7;
    ram_cell[    1667] = 32'h00000511;
    ram_cell[    1668] = 32'h000003a6;
    ram_cell[    1669] = 32'h0000066f;
    ram_cell[    1670] = 32'h00000600;
    ram_cell[    1671] = 32'h000005e9;
    ram_cell[    1672] = 32'h0000067b;
    ram_cell[    1673] = 32'h00000179;
    ram_cell[    1674] = 32'h00000758;
    ram_cell[    1675] = 32'h000001a0;
    ram_cell[    1676] = 32'h0000003f;
    ram_cell[    1677] = 32'h00000649;
    ram_cell[    1678] = 32'h00000619;
    ram_cell[    1679] = 32'h00000109;
    ram_cell[    1680] = 32'h00000302;
    ram_cell[    1681] = 32'h000006e3;
    ram_cell[    1682] = 32'h00000583;
    ram_cell[    1683] = 32'h00000216;
    ram_cell[    1684] = 32'h0000019b;
    ram_cell[    1685] = 32'h000000b2;
    ram_cell[    1686] = 32'h0000038f;
    ram_cell[    1687] = 32'h00000779;
    ram_cell[    1688] = 32'h00000714;
    ram_cell[    1689] = 32'h00000753;
    ram_cell[    1690] = 32'h000001dd;
    ram_cell[    1691] = 32'h000003d3;
    ram_cell[    1692] = 32'h00000741;
    ram_cell[    1693] = 32'h000003a4;
    ram_cell[    1694] = 32'h000000e5;
    ram_cell[    1695] = 32'h00000455;
    ram_cell[    1696] = 32'h0000053e;
    ram_cell[    1697] = 32'h0000003a;
    ram_cell[    1698] = 32'h000000ff;
    ram_cell[    1699] = 32'h00000192;
    ram_cell[    1700] = 32'h000007c2;
    ram_cell[    1701] = 32'h000007a0;
    ram_cell[    1702] = 32'h00000093;
    ram_cell[    1703] = 32'h00000568;
    ram_cell[    1704] = 32'h00000149;
    ram_cell[    1705] = 32'h0000076b;
    ram_cell[    1706] = 32'h000002aa;
    ram_cell[    1707] = 32'h00000181;
    ram_cell[    1708] = 32'h00000152;
    ram_cell[    1709] = 32'h0000038e;
    ram_cell[    1710] = 32'h00000140;
    ram_cell[    1711] = 32'h000001e3;
    ram_cell[    1712] = 32'h000000dd;
    ram_cell[    1713] = 32'h00000340;
    ram_cell[    1714] = 32'h00000009;
    ram_cell[    1715] = 32'h000007cc;
    ram_cell[    1716] = 32'h00000543;
    ram_cell[    1717] = 32'h000005e4;
    ram_cell[    1718] = 32'h000003fe;
    ram_cell[    1719] = 32'h000001f4;
    ram_cell[    1720] = 32'h000003f4;
    ram_cell[    1721] = 32'h000002a4;
    ram_cell[    1722] = 32'h000003fa;
    ram_cell[    1723] = 32'h0000030d;
    ram_cell[    1724] = 32'h0000035a;
    ram_cell[    1725] = 32'h00000287;
    ram_cell[    1726] = 32'h000006ae;
    ram_cell[    1727] = 32'h00000180;
    ram_cell[    1728] = 32'h00000317;
    ram_cell[    1729] = 32'h000001eb;
    ram_cell[    1730] = 32'h00000134;
    ram_cell[    1731] = 32'h00000204;
    ram_cell[    1732] = 32'h00000617;
    ram_cell[    1733] = 32'h0000049d;
    ram_cell[    1734] = 32'h0000066a;
    ram_cell[    1735] = 32'h000007ff;
    ram_cell[    1736] = 32'h000006d9;
    ram_cell[    1737] = 32'h000005b5;
    ram_cell[    1738] = 32'h000006f3;
    ram_cell[    1739] = 32'h000002da;
    ram_cell[    1740] = 32'h00000777;
    ram_cell[    1741] = 32'h00000167;
    ram_cell[    1742] = 32'h000004bd;
    ram_cell[    1743] = 32'h000000c5;
    ram_cell[    1744] = 32'h00000019;
    ram_cell[    1745] = 32'h000002e9;
    ram_cell[    1746] = 32'h000003b3;
    ram_cell[    1747] = 32'h00000700;
    ram_cell[    1748] = 32'h000001fc;
    ram_cell[    1749] = 32'h000007b3;
    ram_cell[    1750] = 32'h00000488;
    ram_cell[    1751] = 32'h00000557;
    ram_cell[    1752] = 32'h000004e7;
    ram_cell[    1753] = 32'h000000cd;
    ram_cell[    1754] = 32'h000002b0;
    ram_cell[    1755] = 32'h0000059e;
    ram_cell[    1756] = 32'h000006c9;
    ram_cell[    1757] = 32'h0000044f;
    ram_cell[    1758] = 32'h00000697;
    ram_cell[    1759] = 32'h000004d7;
    ram_cell[    1760] = 32'h00000683;
    ram_cell[    1761] = 32'h00000633;
    ram_cell[    1762] = 32'h0000043e;
    ram_cell[    1763] = 32'h00000533;
    ram_cell[    1764] = 32'h0000061c;
    ram_cell[    1765] = 32'h00000110;
    ram_cell[    1766] = 32'h000003df;
    ram_cell[    1767] = 32'h000005a1;
    ram_cell[    1768] = 32'h000006da;
    ram_cell[    1769] = 32'h0000068d;
    ram_cell[    1770] = 32'h0000045b;
    ram_cell[    1771] = 32'h00000416;
    ram_cell[    1772] = 32'h000006d7;
    ram_cell[    1773] = 32'h00000307;
    ram_cell[    1774] = 32'h00000626;
    ram_cell[    1775] = 32'h000005d9;
    ram_cell[    1776] = 32'h00000145;
    ram_cell[    1777] = 32'h000001ff;
    ram_cell[    1778] = 32'h00000147;
    ram_cell[    1779] = 32'h00000555;
    ram_cell[    1780] = 32'h000001e0;
    ram_cell[    1781] = 32'h000002f2;
    ram_cell[    1782] = 32'h0000040a;
    ram_cell[    1783] = 32'h00000381;
    ram_cell[    1784] = 32'h000007e6;
    ram_cell[    1785] = 32'h00000327;
    ram_cell[    1786] = 32'h00000190;
    ram_cell[    1787] = 32'h000001b3;
    ram_cell[    1788] = 32'h000006eb;
    ram_cell[    1789] = 32'h0000055c;
    ram_cell[    1790] = 32'h000006f7;
    ram_cell[    1791] = 32'h00000687;
    ram_cell[    1792] = 32'h000003dd;
    ram_cell[    1793] = 32'h000004b3;
    ram_cell[    1794] = 32'h000007a1;
    ram_cell[    1795] = 32'h000006fb;
    ram_cell[    1796] = 32'h000007af;
    ram_cell[    1797] = 32'h000005e6;
    ram_cell[    1798] = 32'h00000759;
    ram_cell[    1799] = 32'h000002f5;
    ram_cell[    1800] = 32'h0000024a;
    ram_cell[    1801] = 32'h00000030;
    ram_cell[    1802] = 32'h0000017b;
    ram_cell[    1803] = 32'h000000b7;
    ram_cell[    1804] = 32'h000004be;
    ram_cell[    1805] = 32'h000006d2;
    ram_cell[    1806] = 32'h00000481;
    ram_cell[    1807] = 32'h000006bd;
    ram_cell[    1808] = 32'h000005bb;
    ram_cell[    1809] = 32'h00000742;
    ram_cell[    1810] = 32'h000003f6;
    ram_cell[    1811] = 32'h00000232;
    ram_cell[    1812] = 32'h00000579;
    ram_cell[    1813] = 32'h00000726;
    ram_cell[    1814] = 32'h000006cd;
    ram_cell[    1815] = 32'h00000341;
    ram_cell[    1816] = 32'h00000309;
    ram_cell[    1817] = 32'h0000005d;
    ram_cell[    1818] = 32'h000005f7;
    ram_cell[    1819] = 32'h000002e8;
    ram_cell[    1820] = 32'h000005c3;
    ram_cell[    1821] = 32'h00000310;
    ram_cell[    1822] = 32'h0000020e;
    ram_cell[    1823] = 32'h000004bb;
    ram_cell[    1824] = 32'h00000431;
    ram_cell[    1825] = 32'h000002f1;
    ram_cell[    1826] = 32'h00000067;
    ram_cell[    1827] = 32'h00000569;
    ram_cell[    1828] = 32'h000004fd;
    ram_cell[    1829] = 32'h0000000d;
    ram_cell[    1830] = 32'h00000443;
    ram_cell[    1831] = 32'h00000458;
    ram_cell[    1832] = 32'h00000497;
    ram_cell[    1833] = 32'h000004b2;
    ram_cell[    1834] = 32'h000007d5;
    ram_cell[    1835] = 32'h00000337;
    ram_cell[    1836] = 32'h0000048b;
    ram_cell[    1837] = 32'h00000382;
    ram_cell[    1838] = 32'h00000653;
    ram_cell[    1839] = 32'h00000240;
    ram_cell[    1840] = 32'h00000666;
    ram_cell[    1841] = 32'h00000325;
    ram_cell[    1842] = 32'h00000659;
    ram_cell[    1843] = 32'h000007df;
    ram_cell[    1844] = 32'h00000717;
    ram_cell[    1845] = 32'h00000439;
    ram_cell[    1846] = 32'h00000494;
    ram_cell[    1847] = 32'h000002d0;
    ram_cell[    1848] = 32'h00000183;
    ram_cell[    1849] = 32'h000004c4;
    ram_cell[    1850] = 32'h000000ca;
    ram_cell[    1851] = 32'h00000796;
    ram_cell[    1852] = 32'h00000295;
    ram_cell[    1853] = 32'h0000023b;
    ram_cell[    1854] = 32'h0000056f;
    ram_cell[    1855] = 32'h0000006b;
    ram_cell[    1856] = 32'h0000039c;
    ram_cell[    1857] = 32'h00000213;
    ram_cell[    1858] = 32'h000006ac;
    ram_cell[    1859] = 32'h00000718;
    ram_cell[    1860] = 32'h0000029e;
    ram_cell[    1861] = 32'h0000010d;
    ram_cell[    1862] = 32'h00000519;
    ram_cell[    1863] = 32'h0000052b;
    ram_cell[    1864] = 32'h00000211;
    ram_cell[    1865] = 32'h000003f8;
    ram_cell[    1866] = 32'h00000421;
    ram_cell[    1867] = 32'h0000077e;
    ram_cell[    1868] = 32'h000007dd;
    ram_cell[    1869] = 32'h000003e5;
    ram_cell[    1870] = 32'h00000292;
    ram_cell[    1871] = 32'h00000454;
    ram_cell[    1872] = 32'h00000165;
    ram_cell[    1873] = 32'h00000641;
    ram_cell[    1874] = 32'h000006a9;
    ram_cell[    1875] = 32'h000002c1;
    ram_cell[    1876] = 32'h000004f6;
    ram_cell[    1877] = 32'h00000024;
    ram_cell[    1878] = 32'h0000063b;
    ram_cell[    1879] = 32'h000004d4;
    ram_cell[    1880] = 32'h0000032c;
    ram_cell[    1881] = 32'h000001bd;
    ram_cell[    1882] = 32'h0000040c;
    ram_cell[    1883] = 32'h0000004b;
    ram_cell[    1884] = 32'h000000d9;
    ram_cell[    1885] = 32'h000000c8;
    ram_cell[    1886] = 32'h0000071f;
    ram_cell[    1887] = 32'h00000065;
    ram_cell[    1888] = 32'h0000009c;
    ram_cell[    1889] = 32'h00000551;
    ram_cell[    1890] = 32'h0000016d;
    ram_cell[    1891] = 32'h0000070c;
    ram_cell[    1892] = 32'h000001d7;
    ram_cell[    1893] = 32'h000003b2;
    ram_cell[    1894] = 32'h0000020d;
    ram_cell[    1895] = 32'h0000008f;
    ram_cell[    1896] = 32'h0000064d;
    ram_cell[    1897] = 32'h00000040;
    ram_cell[    1898] = 32'h0000078c;
    ram_cell[    1899] = 32'h00000477;
    ram_cell[    1900] = 32'h00000496;
    ram_cell[    1901] = 32'h000001b9;
    ram_cell[    1902] = 32'h0000073a;
    ram_cell[    1903] = 32'h00000404;
    ram_cell[    1904] = 32'h00000354;
    ram_cell[    1905] = 32'h000004e0;
    ram_cell[    1906] = 32'h0000028c;
    ram_cell[    1907] = 32'h0000009b;
    ram_cell[    1908] = 32'h00000262;
    ram_cell[    1909] = 32'h000003c5;
    ram_cell[    1910] = 32'h00000158;
    ram_cell[    1911] = 32'h00000000;
    ram_cell[    1912] = 32'h000007b4;
    ram_cell[    1913] = 32'h000005d4;
    ram_cell[    1914] = 32'h00000253;
    ram_cell[    1915] = 32'h00000350;
    ram_cell[    1916] = 32'h00000459;
    ram_cell[    1917] = 32'h00000664;
    ram_cell[    1918] = 32'h000002c8;
    ram_cell[    1919] = 32'h00000495;
    ram_cell[    1920] = 32'h000001a2;
    ram_cell[    1921] = 32'h000007bb;
    ram_cell[    1922] = 32'h0000047f;
    ram_cell[    1923] = 32'h000001e8;
    ram_cell[    1924] = 32'h00000752;
    ram_cell[    1925] = 32'h00000706;
    ram_cell[    1926] = 32'h00000345;
    ram_cell[    1927] = 32'h00000784;
    ram_cell[    1928] = 32'h00000674;
    ram_cell[    1929] = 32'h0000005a;
    ram_cell[    1930] = 32'h000007de;
    ram_cell[    1931] = 32'h000002a5;
    ram_cell[    1932] = 32'h0000028f;
    ram_cell[    1933] = 32'h0000015d;
    ram_cell[    1934] = 32'h0000008c;
    ram_cell[    1935] = 32'h0000067c;
    ram_cell[    1936] = 32'h00000261;
    ram_cell[    1937] = 32'h00000405;
    ram_cell[    1938] = 32'h000005d2;
    ram_cell[    1939] = 32'h000007fc;
    ram_cell[    1940] = 32'h0000077f;
    ram_cell[    1941] = 32'h000002b2;
    ram_cell[    1942] = 32'h000007d4;
    ram_cell[    1943] = 32'h0000039e;
    ram_cell[    1944] = 32'h0000022a;
    ram_cell[    1945] = 32'h000001bb;
    ram_cell[    1946] = 32'h0000034e;
    ram_cell[    1947] = 32'h0000060b;
    ram_cell[    1948] = 32'h00000738;
    ram_cell[    1949] = 32'h000006cc;
    ram_cell[    1950] = 32'h00000410;
    ram_cell[    1951] = 32'h00000521;
    ram_cell[    1952] = 32'h000004a6;
    ram_cell[    1953] = 32'h000007da;
    ram_cell[    1954] = 32'h0000036b;
    ram_cell[    1955] = 32'h000006f6;
    ram_cell[    1956] = 32'h00000660;
    ram_cell[    1957] = 32'h0000042e;
    ram_cell[    1958] = 32'h00000768;
    ram_cell[    1959] = 32'h00000194;
    ram_cell[    1960] = 32'h00000265;
    ram_cell[    1961] = 32'h00000170;
    ram_cell[    1962] = 32'h00000142;
    ram_cell[    1963] = 32'h000000bf;
    ram_cell[    1964] = 32'h00000355;
    ram_cell[    1965] = 32'h00000161;
    ram_cell[    1966] = 32'h0000043b;
    ram_cell[    1967] = 32'h0000075f;
    ram_cell[    1968] = 32'h000006a7;
    ram_cell[    1969] = 32'h00000423;
    ram_cell[    1970] = 32'h00000128;
    ram_cell[    1971] = 32'h00000701;
    ram_cell[    1972] = 32'h000006ec;
    ram_cell[    1973] = 32'h00000077;
    ram_cell[    1974] = 32'h000000b4;
    ram_cell[    1975] = 32'h00000277;
    ram_cell[    1976] = 32'h0000049e;
    ram_cell[    1977] = 32'h0000027a;
    ram_cell[    1978] = 32'h0000002e;
    ram_cell[    1979] = 32'h000000c1;
    ram_cell[    1980] = 32'h000005bd;
    ram_cell[    1981] = 32'h00000241;
    ram_cell[    1982] = 32'h000001ea;
    ram_cell[    1983] = 32'h000001dc;
    ram_cell[    1984] = 32'h00000071;
    ram_cell[    1985] = 32'h00000778;
    ram_cell[    1986] = 32'h000000d1;
    ram_cell[    1987] = 32'h000000bd;
    ram_cell[    1988] = 32'h00000535;
    ram_cell[    1989] = 32'h00000686;
    ram_cell[    1990] = 32'h000005b0;
    ram_cell[    1991] = 32'h000007bc;
    ram_cell[    1992] = 32'h000006fc;
    ram_cell[    1993] = 32'h000006ab;
    ram_cell[    1994] = 32'h000002b1;
    ram_cell[    1995] = 32'h0000050e;
    ram_cell[    1996] = 32'h00000390;
    ram_cell[    1997] = 32'h00000601;
    ram_cell[    1998] = 32'h00000725;
    ram_cell[    1999] = 32'h000007eb;
    ram_cell[    2000] = 32'h000004ae;
    ram_cell[    2001] = 32'h0000021a;
    ram_cell[    2002] = 32'h000002ad;
    ram_cell[    2003] = 32'h00000558;
    ram_cell[    2004] = 32'h000003be;
    ram_cell[    2005] = 32'h000001c6;
    ram_cell[    2006] = 32'h000001b7;
    ram_cell[    2007] = 32'h00000667;
    ram_cell[    2008] = 32'h0000015e;
    ram_cell[    2009] = 32'h00000565;
    ram_cell[    2010] = 32'h0000028a;
    ram_cell[    2011] = 32'h000006ea;
    ram_cell[    2012] = 32'h0000069b;
    ram_cell[    2013] = 32'h00000175;
    ram_cell[    2014] = 32'h00000450;
    ram_cell[    2015] = 32'h0000019c;
    ram_cell[    2016] = 32'h0000015a;
    ram_cell[    2017] = 32'h000000ab;
    ram_cell[    2018] = 32'h00000508;
    ram_cell[    2019] = 32'h000003e0;
    ram_cell[    2020] = 32'h000001e9;
    ram_cell[    2021] = 32'h0000031d;
    ram_cell[    2022] = 32'h000007a5;
    ram_cell[    2023] = 32'h000001e7;
    ram_cell[    2024] = 32'h00000209;
    ram_cell[    2025] = 32'h000005a4;
    ram_cell[    2026] = 32'h0000039b;
    ram_cell[    2027] = 32'h00000122;
    ram_cell[    2028] = 32'h00000629;
    ram_cell[    2029] = 32'h000007e3;
    ram_cell[    2030] = 32'h000005ad;
    ram_cell[    2031] = 32'h00000740;
    ram_cell[    2032] = 32'h00000765;
    ram_cell[    2033] = 32'h000003ed;
    ram_cell[    2034] = 32'h000003bd;
    ram_cell[    2035] = 32'h0000063e;
    ram_cell[    2036] = 32'h0000068a;
    ram_cell[    2037] = 32'h000003b6;
    ram_cell[    2038] = 32'h0000005e;
    ram_cell[    2039] = 32'h000002bb;
    ram_cell[    2040] = 32'h0000051a;
    ram_cell[    2041] = 32'h00000581;
    ram_cell[    2042] = 32'h0000037f;
    ram_cell[    2043] = 32'h000003a2;
    ram_cell[    2044] = 32'h000007ae;
    ram_cell[    2045] = 32'h00000620;
    ram_cell[    2046] = 32'h0000006d;
    ram_cell[    2047] = 32'h0000000c;
end

endmodule

