
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h13903f8a;
    ram_cell[       1] = 32'h0;  // 32'hb3362ab9;
    ram_cell[       2] = 32'h0;  // 32'hdfc4232c;
    ram_cell[       3] = 32'h0;  // 32'h8c84cdbc;
    ram_cell[       4] = 32'h0;  // 32'hd3bc0a15;
    ram_cell[       5] = 32'h0;  // 32'hc4f4ff03;
    ram_cell[       6] = 32'h0;  // 32'h3edeb501;
    ram_cell[       7] = 32'h0;  // 32'hf68a786e;
    ram_cell[       8] = 32'h0;  // 32'hb460706c;
    ram_cell[       9] = 32'h0;  // 32'hf883abd6;
    ram_cell[      10] = 32'h0;  // 32'h3bc63317;
    ram_cell[      11] = 32'h0;  // 32'h88d94cd8;
    ram_cell[      12] = 32'h0;  // 32'he3d6de7f;
    ram_cell[      13] = 32'h0;  // 32'h9d991d0c;
    ram_cell[      14] = 32'h0;  // 32'h1da2b2b5;
    ram_cell[      15] = 32'h0;  // 32'h82751f96;
    ram_cell[      16] = 32'h0;  // 32'h36ae4d93;
    ram_cell[      17] = 32'h0;  // 32'h8bd4f1d8;
    ram_cell[      18] = 32'h0;  // 32'h2cc11aa5;
    ram_cell[      19] = 32'h0;  // 32'h96b777af;
    ram_cell[      20] = 32'h0;  // 32'h222048db;
    ram_cell[      21] = 32'h0;  // 32'h37ce7efd;
    ram_cell[      22] = 32'h0;  // 32'hf64e32dd;
    ram_cell[      23] = 32'h0;  // 32'h890ca735;
    ram_cell[      24] = 32'h0;  // 32'h9faed061;
    ram_cell[      25] = 32'h0;  // 32'h46058b54;
    ram_cell[      26] = 32'h0;  // 32'hd1f76299;
    ram_cell[      27] = 32'h0;  // 32'h90c90852;
    ram_cell[      28] = 32'h0;  // 32'h0ae58c61;
    ram_cell[      29] = 32'h0;  // 32'he5364d10;
    ram_cell[      30] = 32'h0;  // 32'he0587ee7;
    ram_cell[      31] = 32'h0;  // 32'hda2bd3f8;
    ram_cell[      32] = 32'h0;  // 32'hcad982e6;
    ram_cell[      33] = 32'h0;  // 32'h772ae639;
    ram_cell[      34] = 32'h0;  // 32'h0e244c87;
    ram_cell[      35] = 32'h0;  // 32'hf330c9f6;
    ram_cell[      36] = 32'h0;  // 32'h7e32fa1e;
    ram_cell[      37] = 32'h0;  // 32'hfd799dd6;
    ram_cell[      38] = 32'h0;  // 32'h097b4f8e;
    ram_cell[      39] = 32'h0;  // 32'ha37310d4;
    ram_cell[      40] = 32'h0;  // 32'h6a34cb72;
    ram_cell[      41] = 32'h0;  // 32'hd06eb429;
    ram_cell[      42] = 32'h0;  // 32'hb954f8c9;
    ram_cell[      43] = 32'h0;  // 32'h3609231a;
    ram_cell[      44] = 32'h0;  // 32'h267339d6;
    ram_cell[      45] = 32'h0;  // 32'h92bec352;
    ram_cell[      46] = 32'h0;  // 32'h8140a46a;
    ram_cell[      47] = 32'h0;  // 32'h5bb12caa;
    ram_cell[      48] = 32'h0;  // 32'h663f8545;
    ram_cell[      49] = 32'h0;  // 32'hd3552b0b;
    ram_cell[      50] = 32'h0;  // 32'he97b93d1;
    ram_cell[      51] = 32'h0;  // 32'h455494fa;
    ram_cell[      52] = 32'h0;  // 32'h36c72389;
    ram_cell[      53] = 32'h0;  // 32'hc632a4b4;
    ram_cell[      54] = 32'h0;  // 32'hc3b4e2f0;
    ram_cell[      55] = 32'h0;  // 32'hb71c8bf2;
    ram_cell[      56] = 32'h0;  // 32'h3688a83e;
    ram_cell[      57] = 32'h0;  // 32'hc7df6b52;
    ram_cell[      58] = 32'h0;  // 32'h18cdb9d5;
    ram_cell[      59] = 32'h0;  // 32'h47a762f0;
    ram_cell[      60] = 32'h0;  // 32'hec7faf67;
    ram_cell[      61] = 32'h0;  // 32'h867e3a2a;
    ram_cell[      62] = 32'h0;  // 32'he36aeb8a;
    ram_cell[      63] = 32'h0;  // 32'h18220a54;
    ram_cell[      64] = 32'h0;  // 32'h4b3c158c;
    ram_cell[      65] = 32'h0;  // 32'ha3766d68;
    ram_cell[      66] = 32'h0;  // 32'h9d6dfc65;
    ram_cell[      67] = 32'h0;  // 32'heb0da816;
    ram_cell[      68] = 32'h0;  // 32'h34063062;
    ram_cell[      69] = 32'h0;  // 32'h68b37a49;
    ram_cell[      70] = 32'h0;  // 32'h0db577fb;
    ram_cell[      71] = 32'h0;  // 32'hc4c3d3b2;
    ram_cell[      72] = 32'h0;  // 32'h1f474d12;
    ram_cell[      73] = 32'h0;  // 32'h811f6592;
    ram_cell[      74] = 32'h0;  // 32'hba123769;
    ram_cell[      75] = 32'h0;  // 32'h4cba22b6;
    ram_cell[      76] = 32'h0;  // 32'h20ea8ebc;
    ram_cell[      77] = 32'h0;  // 32'ha243921c;
    ram_cell[      78] = 32'h0;  // 32'hcb8886f1;
    ram_cell[      79] = 32'h0;  // 32'hc4028d72;
    ram_cell[      80] = 32'h0;  // 32'he97b499b;
    ram_cell[      81] = 32'h0;  // 32'h5072fd56;
    ram_cell[      82] = 32'h0;  // 32'h247397cb;
    ram_cell[      83] = 32'h0;  // 32'h43b01f51;
    ram_cell[      84] = 32'h0;  // 32'h2b3940be;
    ram_cell[      85] = 32'h0;  // 32'h0fe26f84;
    ram_cell[      86] = 32'h0;  // 32'h345eaa5f;
    ram_cell[      87] = 32'h0;  // 32'hac5cdf00;
    ram_cell[      88] = 32'h0;  // 32'h853041d5;
    ram_cell[      89] = 32'h0;  // 32'h509e0077;
    ram_cell[      90] = 32'h0;  // 32'h54d6d4f4;
    ram_cell[      91] = 32'h0;  // 32'he96c61c8;
    ram_cell[      92] = 32'h0;  // 32'h46275211;
    ram_cell[      93] = 32'h0;  // 32'h9c95139a;
    ram_cell[      94] = 32'h0;  // 32'h437ed1af;
    ram_cell[      95] = 32'h0;  // 32'hf015ee63;
    ram_cell[      96] = 32'h0;  // 32'h8a4da902;
    ram_cell[      97] = 32'h0;  // 32'hcb8601e9;
    ram_cell[      98] = 32'h0;  // 32'h19098518;
    ram_cell[      99] = 32'h0;  // 32'h437c07bc;
    ram_cell[     100] = 32'h0;  // 32'h2dde82e4;
    ram_cell[     101] = 32'h0;  // 32'he0f1702d;
    ram_cell[     102] = 32'h0;  // 32'h78eca65c;
    ram_cell[     103] = 32'h0;  // 32'h377a1040;
    ram_cell[     104] = 32'h0;  // 32'hbd33cdf8;
    ram_cell[     105] = 32'h0;  // 32'hd2fcb6f9;
    ram_cell[     106] = 32'h0;  // 32'h2f434b09;
    ram_cell[     107] = 32'h0;  // 32'hab752abf;
    ram_cell[     108] = 32'h0;  // 32'hf11e95ae;
    ram_cell[     109] = 32'h0;  // 32'hc5cb6ce2;
    ram_cell[     110] = 32'h0;  // 32'hf5b1a143;
    ram_cell[     111] = 32'h0;  // 32'had459636;
    ram_cell[     112] = 32'h0;  // 32'h7988ae77;
    ram_cell[     113] = 32'h0;  // 32'h381cb6f3;
    ram_cell[     114] = 32'h0;  // 32'h0a692756;
    ram_cell[     115] = 32'h0;  // 32'h666fefe9;
    ram_cell[     116] = 32'h0;  // 32'hd2a6f96d;
    ram_cell[     117] = 32'h0;  // 32'hf1e665bc;
    ram_cell[     118] = 32'h0;  // 32'hb1e88e67;
    ram_cell[     119] = 32'h0;  // 32'he18bed27;
    ram_cell[     120] = 32'h0;  // 32'hb7ffec7d;
    ram_cell[     121] = 32'h0;  // 32'h845e2c44;
    ram_cell[     122] = 32'h0;  // 32'h553f2ed0;
    ram_cell[     123] = 32'h0;  // 32'hf9eb98ac;
    ram_cell[     124] = 32'h0;  // 32'he129d605;
    ram_cell[     125] = 32'h0;  // 32'h272fe068;
    ram_cell[     126] = 32'h0;  // 32'ha968bd65;
    ram_cell[     127] = 32'h0;  // 32'hd94c88e6;
    ram_cell[     128] = 32'h0;  // 32'h5900ec99;
    ram_cell[     129] = 32'h0;  // 32'h46d31544;
    ram_cell[     130] = 32'h0;  // 32'hca963eff;
    ram_cell[     131] = 32'h0;  // 32'h241fdecf;
    ram_cell[     132] = 32'h0;  // 32'hedba4dd7;
    ram_cell[     133] = 32'h0;  // 32'h9dffc104;
    ram_cell[     134] = 32'h0;  // 32'h4eec0c89;
    ram_cell[     135] = 32'h0;  // 32'h80fc3c8d;
    ram_cell[     136] = 32'h0;  // 32'h9c46b480;
    ram_cell[     137] = 32'h0;  // 32'h600e72ee;
    ram_cell[     138] = 32'h0;  // 32'h25445a60;
    ram_cell[     139] = 32'h0;  // 32'he9f4110d;
    ram_cell[     140] = 32'h0;  // 32'hb12ad61e;
    ram_cell[     141] = 32'h0;  // 32'h28c51563;
    ram_cell[     142] = 32'h0;  // 32'h8f0a15a7;
    ram_cell[     143] = 32'h0;  // 32'hf045855e;
    ram_cell[     144] = 32'h0;  // 32'h6c896f7d;
    ram_cell[     145] = 32'h0;  // 32'hbc8bc351;
    ram_cell[     146] = 32'h0;  // 32'hcbaeb545;
    ram_cell[     147] = 32'h0;  // 32'h1039b020;
    ram_cell[     148] = 32'h0;  // 32'he5e81a8a;
    ram_cell[     149] = 32'h0;  // 32'h3fde5bd0;
    ram_cell[     150] = 32'h0;  // 32'h9c3e1448;
    ram_cell[     151] = 32'h0;  // 32'hd816bd1d;
    ram_cell[     152] = 32'h0;  // 32'h08bc14b7;
    ram_cell[     153] = 32'h0;  // 32'hcfd59278;
    ram_cell[     154] = 32'h0;  // 32'hc7ecc080;
    ram_cell[     155] = 32'h0;  // 32'h901f611c;
    ram_cell[     156] = 32'h0;  // 32'hd3500c82;
    ram_cell[     157] = 32'h0;  // 32'h906fb23b;
    ram_cell[     158] = 32'h0;  // 32'h752d34a3;
    ram_cell[     159] = 32'h0;  // 32'ha6cfb1e3;
    ram_cell[     160] = 32'h0;  // 32'h634d5115;
    ram_cell[     161] = 32'h0;  // 32'h5e18d914;
    ram_cell[     162] = 32'h0;  // 32'ha9868eba;
    ram_cell[     163] = 32'h0;  // 32'h7832d3c6;
    ram_cell[     164] = 32'h0;  // 32'ha2a41233;
    ram_cell[     165] = 32'h0;  // 32'hdc89419c;
    ram_cell[     166] = 32'h0;  // 32'h203f9ca7;
    ram_cell[     167] = 32'h0;  // 32'hac5d2610;
    ram_cell[     168] = 32'h0;  // 32'haee58ca2;
    ram_cell[     169] = 32'h0;  // 32'h5d398498;
    ram_cell[     170] = 32'h0;  // 32'h40607688;
    ram_cell[     171] = 32'h0;  // 32'h9cbd552b;
    ram_cell[     172] = 32'h0;  // 32'h8b3b460e;
    ram_cell[     173] = 32'h0;  // 32'hed3c4617;
    ram_cell[     174] = 32'h0;  // 32'he4fa1e97;
    ram_cell[     175] = 32'h0;  // 32'hc155e316;
    ram_cell[     176] = 32'h0;  // 32'he8d18c2c;
    ram_cell[     177] = 32'h0;  // 32'h2c3e10fb;
    ram_cell[     178] = 32'h0;  // 32'h2cda63ff;
    ram_cell[     179] = 32'h0;  // 32'h10de725a;
    ram_cell[     180] = 32'h0;  // 32'h3e682f66;
    ram_cell[     181] = 32'h0;  // 32'h23cdef27;
    ram_cell[     182] = 32'h0;  // 32'h36d2deb8;
    ram_cell[     183] = 32'h0;  // 32'h1c4a435d;
    ram_cell[     184] = 32'h0;  // 32'hc8cac635;
    ram_cell[     185] = 32'h0;  // 32'h57e71557;
    ram_cell[     186] = 32'h0;  // 32'hdcaf8c69;
    ram_cell[     187] = 32'h0;  // 32'h9508bd3f;
    ram_cell[     188] = 32'h0;  // 32'h85b69186;
    ram_cell[     189] = 32'h0;  // 32'h5d6b1b47;
    ram_cell[     190] = 32'h0;  // 32'h7424edfe;
    ram_cell[     191] = 32'h0;  // 32'h49c43db1;
    ram_cell[     192] = 32'h0;  // 32'h2e1ee4c0;
    ram_cell[     193] = 32'h0;  // 32'h70d23c64;
    ram_cell[     194] = 32'h0;  // 32'hdab88ce5;
    ram_cell[     195] = 32'h0;  // 32'hab9087b6;
    ram_cell[     196] = 32'h0;  // 32'haa2b68f1;
    ram_cell[     197] = 32'h0;  // 32'h6a412d7c;
    ram_cell[     198] = 32'h0;  // 32'hb30972ff;
    ram_cell[     199] = 32'h0;  // 32'hbf1841ac;
    ram_cell[     200] = 32'h0;  // 32'he1abaa1b;
    ram_cell[     201] = 32'h0;  // 32'h897d6eac;
    ram_cell[     202] = 32'h0;  // 32'h2b571d68;
    ram_cell[     203] = 32'h0;  // 32'h8688ae60;
    ram_cell[     204] = 32'h0;  // 32'h20a22c44;
    ram_cell[     205] = 32'h0;  // 32'h06c0cdd4;
    ram_cell[     206] = 32'h0;  // 32'hba358472;
    ram_cell[     207] = 32'h0;  // 32'hd543c3ee;
    ram_cell[     208] = 32'h0;  // 32'hef568dff;
    ram_cell[     209] = 32'h0;  // 32'h6bfb06e5;
    ram_cell[     210] = 32'h0;  // 32'h463170dc;
    ram_cell[     211] = 32'h0;  // 32'hb1d6404c;
    ram_cell[     212] = 32'h0;  // 32'he08b3791;
    ram_cell[     213] = 32'h0;  // 32'hb5a40591;
    ram_cell[     214] = 32'h0;  // 32'h8a784158;
    ram_cell[     215] = 32'h0;  // 32'hf4c0221d;
    ram_cell[     216] = 32'h0;  // 32'h416dfb67;
    ram_cell[     217] = 32'h0;  // 32'h7f72cb1c;
    ram_cell[     218] = 32'h0;  // 32'hbbce2091;
    ram_cell[     219] = 32'h0;  // 32'h38782d32;
    ram_cell[     220] = 32'h0;  // 32'h3d9fa8fc;
    ram_cell[     221] = 32'h0;  // 32'h0afac61e;
    ram_cell[     222] = 32'h0;  // 32'h14f1859b;
    ram_cell[     223] = 32'h0;  // 32'h865e50a0;
    ram_cell[     224] = 32'h0;  // 32'h92012ef4;
    ram_cell[     225] = 32'h0;  // 32'h6b07475b;
    ram_cell[     226] = 32'h0;  // 32'hbdc50ecd;
    ram_cell[     227] = 32'h0;  // 32'hc4eaf022;
    ram_cell[     228] = 32'h0;  // 32'he1339cdf;
    ram_cell[     229] = 32'h0;  // 32'hfd44a3c2;
    ram_cell[     230] = 32'h0;  // 32'hf982ec43;
    ram_cell[     231] = 32'h0;  // 32'hafa1819a;
    ram_cell[     232] = 32'h0;  // 32'h3420cfb5;
    ram_cell[     233] = 32'h0;  // 32'ha10b8809;
    ram_cell[     234] = 32'h0;  // 32'hc741cfbb;
    ram_cell[     235] = 32'h0;  // 32'h0a2a2e00;
    ram_cell[     236] = 32'h0;  // 32'hddc9e138;
    ram_cell[     237] = 32'h0;  // 32'h01169329;
    ram_cell[     238] = 32'h0;  // 32'h5cfd6cba;
    ram_cell[     239] = 32'h0;  // 32'h961722be;
    ram_cell[     240] = 32'h0;  // 32'h2a1637a8;
    ram_cell[     241] = 32'h0;  // 32'h0a2d0d10;
    ram_cell[     242] = 32'h0;  // 32'hc69ba008;
    ram_cell[     243] = 32'h0;  // 32'h7fc8a085;
    ram_cell[     244] = 32'h0;  // 32'h6fce5c88;
    ram_cell[     245] = 32'h0;  // 32'h139f783b;
    ram_cell[     246] = 32'h0;  // 32'h2c920ef2;
    ram_cell[     247] = 32'h0;  // 32'h12f80c21;
    ram_cell[     248] = 32'h0;  // 32'hf7a951d4;
    ram_cell[     249] = 32'h0;  // 32'h3cbb950d;
    ram_cell[     250] = 32'h0;  // 32'hfd630dd0;
    ram_cell[     251] = 32'h0;  // 32'hcd371119;
    ram_cell[     252] = 32'h0;  // 32'hf3e61654;
    ram_cell[     253] = 32'h0;  // 32'h3549ee8d;
    ram_cell[     254] = 32'h0;  // 32'h5b9c8f00;
    ram_cell[     255] = 32'h0;  // 32'hba305bc2;
    ram_cell[     256] = 32'h0;  // 32'h78ffc057;
    ram_cell[     257] = 32'h0;  // 32'h52157990;
    ram_cell[     258] = 32'h0;  // 32'h3720db05;
    ram_cell[     259] = 32'h0;  // 32'h8c4ca512;
    ram_cell[     260] = 32'h0;  // 32'hd1c7fa9f;
    ram_cell[     261] = 32'h0;  // 32'h8eb00ea6;
    ram_cell[     262] = 32'h0;  // 32'hb8047aca;
    ram_cell[     263] = 32'h0;  // 32'h5a428b12;
    ram_cell[     264] = 32'h0;  // 32'h1a6616fd;
    ram_cell[     265] = 32'h0;  // 32'h4336f03d;
    ram_cell[     266] = 32'h0;  // 32'h316f51f2;
    ram_cell[     267] = 32'h0;  // 32'hd8fe388e;
    ram_cell[     268] = 32'h0;  // 32'h72ed098c;
    ram_cell[     269] = 32'h0;  // 32'hc5018cae;
    ram_cell[     270] = 32'h0;  // 32'h23612a22;
    ram_cell[     271] = 32'h0;  // 32'h41fffcf1;
    ram_cell[     272] = 32'h0;  // 32'hc8657752;
    ram_cell[     273] = 32'h0;  // 32'hd2a99fe7;
    ram_cell[     274] = 32'h0;  // 32'hbfab9632;
    ram_cell[     275] = 32'h0;  // 32'h06e045e0;
    ram_cell[     276] = 32'h0;  // 32'h33083d91;
    ram_cell[     277] = 32'h0;  // 32'heb87bf98;
    ram_cell[     278] = 32'h0;  // 32'h5cda9dad;
    ram_cell[     279] = 32'h0;  // 32'h217bd9bd;
    ram_cell[     280] = 32'h0;  // 32'heaa59e43;
    ram_cell[     281] = 32'h0;  // 32'h5c34b09f;
    ram_cell[     282] = 32'h0;  // 32'hc5656359;
    ram_cell[     283] = 32'h0;  // 32'h0dec6930;
    ram_cell[     284] = 32'h0;  // 32'h9084e52e;
    ram_cell[     285] = 32'h0;  // 32'hb1d564fc;
    ram_cell[     286] = 32'h0;  // 32'h0e41903f;
    ram_cell[     287] = 32'h0;  // 32'h3618cd3d;
    ram_cell[     288] = 32'h0;  // 32'h4ad9c325;
    ram_cell[     289] = 32'h0;  // 32'h59093419;
    ram_cell[     290] = 32'h0;  // 32'hc54cd6c8;
    ram_cell[     291] = 32'h0;  // 32'hc5ee244f;
    ram_cell[     292] = 32'h0;  // 32'h8398aa48;
    ram_cell[     293] = 32'h0;  // 32'hb0700f21;
    ram_cell[     294] = 32'h0;  // 32'hb36df84c;
    ram_cell[     295] = 32'h0;  // 32'h7a37d9ba;
    ram_cell[     296] = 32'h0;  // 32'h51130b38;
    ram_cell[     297] = 32'h0;  // 32'hcc6626e6;
    ram_cell[     298] = 32'h0;  // 32'h99c06c4a;
    ram_cell[     299] = 32'h0;  // 32'hbea7c917;
    ram_cell[     300] = 32'h0;  // 32'h206e9efc;
    ram_cell[     301] = 32'h0;  // 32'h5373e91e;
    ram_cell[     302] = 32'h0;  // 32'hda78b2bd;
    ram_cell[     303] = 32'h0;  // 32'h7c5e5c7a;
    ram_cell[     304] = 32'h0;  // 32'h882ecf29;
    ram_cell[     305] = 32'h0;  // 32'hd8192c23;
    ram_cell[     306] = 32'h0;  // 32'h3798a531;
    ram_cell[     307] = 32'h0;  // 32'hce2c7f40;
    ram_cell[     308] = 32'h0;  // 32'h5e48d1e0;
    ram_cell[     309] = 32'h0;  // 32'h710d5c2f;
    ram_cell[     310] = 32'h0;  // 32'hf10ec732;
    ram_cell[     311] = 32'h0;  // 32'hd12bdddc;
    ram_cell[     312] = 32'h0;  // 32'h04b218f2;
    ram_cell[     313] = 32'h0;  // 32'hd5efecc8;
    ram_cell[     314] = 32'h0;  // 32'hda186972;
    ram_cell[     315] = 32'h0;  // 32'hd5f1edb6;
    ram_cell[     316] = 32'h0;  // 32'haccb389c;
    ram_cell[     317] = 32'h0;  // 32'ha1e64991;
    ram_cell[     318] = 32'h0;  // 32'h475436b5;
    ram_cell[     319] = 32'h0;  // 32'h0ae24594;
    ram_cell[     320] = 32'h0;  // 32'h97aaea33;
    ram_cell[     321] = 32'h0;  // 32'hdb30e342;
    ram_cell[     322] = 32'h0;  // 32'h143d3046;
    ram_cell[     323] = 32'h0;  // 32'h3fbcd978;
    ram_cell[     324] = 32'h0;  // 32'hbd4ee99c;
    ram_cell[     325] = 32'h0;  // 32'hec5e15ad;
    ram_cell[     326] = 32'h0;  // 32'h830c0927;
    ram_cell[     327] = 32'h0;  // 32'h04fe87f1;
    ram_cell[     328] = 32'h0;  // 32'h51afb0ca;
    ram_cell[     329] = 32'h0;  // 32'hc37dc02e;
    ram_cell[     330] = 32'h0;  // 32'h7200b7c4;
    ram_cell[     331] = 32'h0;  // 32'hbfffa89d;
    ram_cell[     332] = 32'h0;  // 32'hf21ce264;
    ram_cell[     333] = 32'h0;  // 32'h9d8d2129;
    ram_cell[     334] = 32'h0;  // 32'h574afcac;
    ram_cell[     335] = 32'h0;  // 32'h54427880;
    ram_cell[     336] = 32'h0;  // 32'h8fd284bd;
    ram_cell[     337] = 32'h0;  // 32'h47afe4ff;
    ram_cell[     338] = 32'h0;  // 32'h147fbfb3;
    ram_cell[     339] = 32'h0;  // 32'ha9e463cf;
    ram_cell[     340] = 32'h0;  // 32'h4522b8ee;
    ram_cell[     341] = 32'h0;  // 32'h6aa5269f;
    ram_cell[     342] = 32'h0;  // 32'ha5d3565f;
    ram_cell[     343] = 32'h0;  // 32'h9eb0d2b3;
    ram_cell[     344] = 32'h0;  // 32'h09b98e74;
    ram_cell[     345] = 32'h0;  // 32'hc71b5c73;
    ram_cell[     346] = 32'h0;  // 32'hd1e15026;
    ram_cell[     347] = 32'h0;  // 32'h44a7c028;
    ram_cell[     348] = 32'h0;  // 32'h8ea849f9;
    ram_cell[     349] = 32'h0;  // 32'h4faac48f;
    ram_cell[     350] = 32'h0;  // 32'hd9a458fc;
    ram_cell[     351] = 32'h0;  // 32'h04cd948b;
    ram_cell[     352] = 32'h0;  // 32'h20447060;
    ram_cell[     353] = 32'h0;  // 32'h7f6672a3;
    ram_cell[     354] = 32'h0;  // 32'h017c852d;
    ram_cell[     355] = 32'h0;  // 32'he50003f0;
    ram_cell[     356] = 32'h0;  // 32'h711938ef;
    ram_cell[     357] = 32'h0;  // 32'h9bf142b0;
    ram_cell[     358] = 32'h0;  // 32'h37972e5c;
    ram_cell[     359] = 32'h0;  // 32'h87e4a635;
    ram_cell[     360] = 32'h0;  // 32'h68e04cbf;
    ram_cell[     361] = 32'h0;  // 32'hf32254b3;
    ram_cell[     362] = 32'h0;  // 32'ha893950f;
    ram_cell[     363] = 32'h0;  // 32'hc57e0587;
    ram_cell[     364] = 32'h0;  // 32'h4e65e2af;
    ram_cell[     365] = 32'h0;  // 32'h06dff286;
    ram_cell[     366] = 32'h0;  // 32'h3419108d;
    ram_cell[     367] = 32'h0;  // 32'hbbdfeedf;
    ram_cell[     368] = 32'h0;  // 32'h375e71e8;
    ram_cell[     369] = 32'h0;  // 32'hb92f383d;
    ram_cell[     370] = 32'h0;  // 32'hcf8f4eb0;
    ram_cell[     371] = 32'h0;  // 32'h413bda55;
    ram_cell[     372] = 32'h0;  // 32'hb3a72d2c;
    ram_cell[     373] = 32'h0;  // 32'he9d79da5;
    ram_cell[     374] = 32'h0;  // 32'h8b70f8cd;
    ram_cell[     375] = 32'h0;  // 32'hdbca5f72;
    ram_cell[     376] = 32'h0;  // 32'h8eb702fb;
    ram_cell[     377] = 32'h0;  // 32'h4ab29cf7;
    ram_cell[     378] = 32'h0;  // 32'h3d9ea919;
    ram_cell[     379] = 32'h0;  // 32'h1cff8c6c;
    ram_cell[     380] = 32'h0;  // 32'h1df189e4;
    ram_cell[     381] = 32'h0;  // 32'h1433157e;
    ram_cell[     382] = 32'h0;  // 32'ha2342625;
    ram_cell[     383] = 32'h0;  // 32'hb51ff798;
    ram_cell[     384] = 32'h0;  // 32'h24b8342d;
    ram_cell[     385] = 32'h0;  // 32'h28c411d7;
    ram_cell[     386] = 32'h0;  // 32'h7d9ec169;
    ram_cell[     387] = 32'h0;  // 32'h461441dd;
    ram_cell[     388] = 32'h0;  // 32'h4b35c3af;
    ram_cell[     389] = 32'h0;  // 32'h8c998026;
    ram_cell[     390] = 32'h0;  // 32'he37cb9f4;
    ram_cell[     391] = 32'h0;  // 32'h2d2ab05c;
    ram_cell[     392] = 32'h0;  // 32'hae627212;
    ram_cell[     393] = 32'h0;  // 32'hc81ef03c;
    ram_cell[     394] = 32'h0;  // 32'h88e097d0;
    ram_cell[     395] = 32'h0;  // 32'h58782bca;
    ram_cell[     396] = 32'h0;  // 32'h9b8e86a6;
    ram_cell[     397] = 32'h0;  // 32'h26890381;
    ram_cell[     398] = 32'h0;  // 32'hf976281c;
    ram_cell[     399] = 32'h0;  // 32'hb67ab27a;
    ram_cell[     400] = 32'h0;  // 32'hdfe7e77b;
    ram_cell[     401] = 32'h0;  // 32'h8e73863d;
    ram_cell[     402] = 32'h0;  // 32'h5f078fe1;
    ram_cell[     403] = 32'h0;  // 32'ha57ba379;
    ram_cell[     404] = 32'h0;  // 32'hc82bd14b;
    ram_cell[     405] = 32'h0;  // 32'hdc7341d7;
    ram_cell[     406] = 32'h0;  // 32'h6ccae4bf;
    ram_cell[     407] = 32'h0;  // 32'h58ee741c;
    ram_cell[     408] = 32'h0;  // 32'h9599a433;
    ram_cell[     409] = 32'h0;  // 32'hecf53f33;
    ram_cell[     410] = 32'h0;  // 32'h497d7d68;
    ram_cell[     411] = 32'h0;  // 32'he6b92c49;
    ram_cell[     412] = 32'h0;  // 32'h8d5877db;
    ram_cell[     413] = 32'h0;  // 32'h060b0c88;
    ram_cell[     414] = 32'h0;  // 32'h4fde709c;
    ram_cell[     415] = 32'h0;  // 32'h87523a32;
    ram_cell[     416] = 32'h0;  // 32'h8635c5e0;
    ram_cell[     417] = 32'h0;  // 32'h0f959b98;
    ram_cell[     418] = 32'h0;  // 32'h92820f0c;
    ram_cell[     419] = 32'h0;  // 32'hf90b4bf0;
    ram_cell[     420] = 32'h0;  // 32'ha03f71a8;
    ram_cell[     421] = 32'h0;  // 32'h3afa9c9f;
    ram_cell[     422] = 32'h0;  // 32'h394ee3e0;
    ram_cell[     423] = 32'h0;  // 32'h9fef7db2;
    ram_cell[     424] = 32'h0;  // 32'h1499b66e;
    ram_cell[     425] = 32'h0;  // 32'h950767c0;
    ram_cell[     426] = 32'h0;  // 32'hd957d959;
    ram_cell[     427] = 32'h0;  // 32'hf5968019;
    ram_cell[     428] = 32'h0;  // 32'h94ca81e8;
    ram_cell[     429] = 32'h0;  // 32'h985d0d42;
    ram_cell[     430] = 32'h0;  // 32'h8fc109b4;
    ram_cell[     431] = 32'h0;  // 32'hf750abb0;
    ram_cell[     432] = 32'h0;  // 32'h7ca68e0e;
    ram_cell[     433] = 32'h0;  // 32'h9413f051;
    ram_cell[     434] = 32'h0;  // 32'he7311577;
    ram_cell[     435] = 32'h0;  // 32'ha428036f;
    ram_cell[     436] = 32'h0;  // 32'habe5bf29;
    ram_cell[     437] = 32'h0;  // 32'he78eebd4;
    ram_cell[     438] = 32'h0;  // 32'hcd765cf5;
    ram_cell[     439] = 32'h0;  // 32'hf508517d;
    ram_cell[     440] = 32'h0;  // 32'h9a8e5b1d;
    ram_cell[     441] = 32'h0;  // 32'hc0031a53;
    ram_cell[     442] = 32'h0;  // 32'h2f2fc6f5;
    ram_cell[     443] = 32'h0;  // 32'h82822d98;
    ram_cell[     444] = 32'h0;  // 32'h32b8926d;
    ram_cell[     445] = 32'h0;  // 32'hd73da53d;
    ram_cell[     446] = 32'h0;  // 32'hc35ee584;
    ram_cell[     447] = 32'h0;  // 32'h80388862;
    ram_cell[     448] = 32'h0;  // 32'hde794744;
    ram_cell[     449] = 32'h0;  // 32'h7834b247;
    ram_cell[     450] = 32'h0;  // 32'h3bce0526;
    ram_cell[     451] = 32'h0;  // 32'h3eee7b91;
    ram_cell[     452] = 32'h0;  // 32'h7f943fcf;
    ram_cell[     453] = 32'h0;  // 32'ha87833c8;
    ram_cell[     454] = 32'h0;  // 32'hadd2ddf8;
    ram_cell[     455] = 32'h0;  // 32'h770daf96;
    ram_cell[     456] = 32'h0;  // 32'h30b5b182;
    ram_cell[     457] = 32'h0;  // 32'hf990b19d;
    ram_cell[     458] = 32'h0;  // 32'hd835aaa0;
    ram_cell[     459] = 32'h0;  // 32'h5f48749b;
    ram_cell[     460] = 32'h0;  // 32'hb7d68f9b;
    ram_cell[     461] = 32'h0;  // 32'hb32cc763;
    ram_cell[     462] = 32'h0;  // 32'h2ab1d4fb;
    ram_cell[     463] = 32'h0;  // 32'h7b084748;
    ram_cell[     464] = 32'h0;  // 32'h152e7c95;
    ram_cell[     465] = 32'h0;  // 32'h348782cd;
    ram_cell[     466] = 32'h0;  // 32'h74a8c274;
    ram_cell[     467] = 32'h0;  // 32'hd569efbc;
    ram_cell[     468] = 32'h0;  // 32'h304ff485;
    ram_cell[     469] = 32'h0;  // 32'hb950e783;
    ram_cell[     470] = 32'h0;  // 32'h9926aca9;
    ram_cell[     471] = 32'h0;  // 32'had767040;
    ram_cell[     472] = 32'h0;  // 32'h6f55981d;
    ram_cell[     473] = 32'h0;  // 32'hebc25da0;
    ram_cell[     474] = 32'h0;  // 32'h44986ddc;
    ram_cell[     475] = 32'h0;  // 32'ha58a4e3b;
    ram_cell[     476] = 32'h0;  // 32'h58c34b72;
    ram_cell[     477] = 32'h0;  // 32'h27ff209a;
    ram_cell[     478] = 32'h0;  // 32'h9eac2046;
    ram_cell[     479] = 32'h0;  // 32'hd4793e6b;
    ram_cell[     480] = 32'h0;  // 32'hf6174559;
    ram_cell[     481] = 32'h0;  // 32'hb415d4a9;
    ram_cell[     482] = 32'h0;  // 32'h3e736a77;
    ram_cell[     483] = 32'h0;  // 32'hc3c37a65;
    ram_cell[     484] = 32'h0;  // 32'h332cd02d;
    ram_cell[     485] = 32'h0;  // 32'h0d35c300;
    ram_cell[     486] = 32'h0;  // 32'ha5d52d44;
    ram_cell[     487] = 32'h0;  // 32'h80a7fd1c;
    ram_cell[     488] = 32'h0;  // 32'hee749fb7;
    ram_cell[     489] = 32'h0;  // 32'hab29ad1f;
    ram_cell[     490] = 32'h0;  // 32'h63866095;
    ram_cell[     491] = 32'h0;  // 32'he93bd52e;
    ram_cell[     492] = 32'h0;  // 32'h908a04b9;
    ram_cell[     493] = 32'h0;  // 32'h48d87d95;
    ram_cell[     494] = 32'h0;  // 32'haab94526;
    ram_cell[     495] = 32'h0;  // 32'h56ce7799;
    ram_cell[     496] = 32'h0;  // 32'h603d8419;
    ram_cell[     497] = 32'h0;  // 32'h54db84cc;
    ram_cell[     498] = 32'h0;  // 32'h77d5cd53;
    ram_cell[     499] = 32'h0;  // 32'hd9c8deb2;
    ram_cell[     500] = 32'h0;  // 32'h87f6bcd0;
    ram_cell[     501] = 32'h0;  // 32'he47c9f58;
    ram_cell[     502] = 32'h0;  // 32'h983f4d0b;
    ram_cell[     503] = 32'h0;  // 32'h17ee2c71;
    ram_cell[     504] = 32'h0;  // 32'h564ea279;
    ram_cell[     505] = 32'h0;  // 32'h7be19001;
    ram_cell[     506] = 32'h0;  // 32'h7c536831;
    ram_cell[     507] = 32'h0;  // 32'he58f517e;
    ram_cell[     508] = 32'h0;  // 32'hacbf7ea1;
    ram_cell[     509] = 32'h0;  // 32'h125347a3;
    ram_cell[     510] = 32'h0;  // 32'h3e7151f5;
    ram_cell[     511] = 32'h0;  // 32'h90b77298;
    ram_cell[     512] = 32'h0;  // 32'h396384e8;
    ram_cell[     513] = 32'h0;  // 32'h1c5e564d;
    ram_cell[     514] = 32'h0;  // 32'h57ecc870;
    ram_cell[     515] = 32'h0;  // 32'ha37eaf8f;
    ram_cell[     516] = 32'h0;  // 32'h83e8447a;
    ram_cell[     517] = 32'h0;  // 32'hcfaf3cca;
    ram_cell[     518] = 32'h0;  // 32'h80ec3f82;
    ram_cell[     519] = 32'h0;  // 32'h33a42d37;
    ram_cell[     520] = 32'h0;  // 32'h177bcd19;
    ram_cell[     521] = 32'h0;  // 32'h7ee1ecba;
    ram_cell[     522] = 32'h0;  // 32'h9696f9f9;
    ram_cell[     523] = 32'h0;  // 32'h74444988;
    ram_cell[     524] = 32'h0;  // 32'h6ce484e2;
    ram_cell[     525] = 32'h0;  // 32'h5609af52;
    ram_cell[     526] = 32'h0;  // 32'h7d92c182;
    ram_cell[     527] = 32'h0;  // 32'ha1402360;
    ram_cell[     528] = 32'h0;  // 32'h1b1ead71;
    ram_cell[     529] = 32'h0;  // 32'hbcbc823b;
    ram_cell[     530] = 32'h0;  // 32'h21a13279;
    ram_cell[     531] = 32'h0;  // 32'h9af12fcd;
    ram_cell[     532] = 32'h0;  // 32'h526fc522;
    ram_cell[     533] = 32'h0;  // 32'hec461642;
    ram_cell[     534] = 32'h0;  // 32'h29f5b428;
    ram_cell[     535] = 32'h0;  // 32'h8df1b6a4;
    ram_cell[     536] = 32'h0;  // 32'hc0cbed07;
    ram_cell[     537] = 32'h0;  // 32'heab16b85;
    ram_cell[     538] = 32'h0;  // 32'h7870870e;
    ram_cell[     539] = 32'h0;  // 32'hf09e9700;
    ram_cell[     540] = 32'h0;  // 32'h130768a9;
    ram_cell[     541] = 32'h0;  // 32'h51392da7;
    ram_cell[     542] = 32'h0;  // 32'h8e59cb63;
    ram_cell[     543] = 32'h0;  // 32'h0169b552;
    ram_cell[     544] = 32'h0;  // 32'h99340248;
    ram_cell[     545] = 32'h0;  // 32'h046c1c24;
    ram_cell[     546] = 32'h0;  // 32'h405d3342;
    ram_cell[     547] = 32'h0;  // 32'hf9ee7bc7;
    ram_cell[     548] = 32'h0;  // 32'h017cb6ea;
    ram_cell[     549] = 32'h0;  // 32'hfc87f0fa;
    ram_cell[     550] = 32'h0;  // 32'ha5e39b02;
    ram_cell[     551] = 32'h0;  // 32'h17ac0a8c;
    ram_cell[     552] = 32'h0;  // 32'h04b9ebf3;
    ram_cell[     553] = 32'h0;  // 32'h6679e00d;
    ram_cell[     554] = 32'h0;  // 32'hc1c92ae1;
    ram_cell[     555] = 32'h0;  // 32'h8e78234f;
    ram_cell[     556] = 32'h0;  // 32'h9806b6a1;
    ram_cell[     557] = 32'h0;  // 32'h6d31d76c;
    ram_cell[     558] = 32'h0;  // 32'h3b3ce753;
    ram_cell[     559] = 32'h0;  // 32'h7512c842;
    ram_cell[     560] = 32'h0;  // 32'h9e6e0be5;
    ram_cell[     561] = 32'h0;  // 32'h420d8879;
    ram_cell[     562] = 32'h0;  // 32'h5ff9ad95;
    ram_cell[     563] = 32'h0;  // 32'hf2c04dae;
    ram_cell[     564] = 32'h0;  // 32'hcf3b6e09;
    ram_cell[     565] = 32'h0;  // 32'he199c952;
    ram_cell[     566] = 32'h0;  // 32'h9c566022;
    ram_cell[     567] = 32'h0;  // 32'h4bc8fe70;
    ram_cell[     568] = 32'h0;  // 32'h04e3dd87;
    ram_cell[     569] = 32'h0;  // 32'h1acfe316;
    ram_cell[     570] = 32'h0;  // 32'h2fa2722b;
    ram_cell[     571] = 32'h0;  // 32'h1d951d54;
    ram_cell[     572] = 32'h0;  // 32'hc6d56cac;
    ram_cell[     573] = 32'h0;  // 32'h8996a647;
    ram_cell[     574] = 32'h0;  // 32'h7dfe2424;
    ram_cell[     575] = 32'h0;  // 32'h2634457a;
    ram_cell[     576] = 32'h0;  // 32'h30df62e7;
    ram_cell[     577] = 32'h0;  // 32'h73f3350e;
    ram_cell[     578] = 32'h0;  // 32'h4ac48e05;
    ram_cell[     579] = 32'h0;  // 32'h6a9bada8;
    ram_cell[     580] = 32'h0;  // 32'h4598ca86;
    ram_cell[     581] = 32'h0;  // 32'hc111fd63;
    ram_cell[     582] = 32'h0;  // 32'hc1bcc61b;
    ram_cell[     583] = 32'h0;  // 32'h031cfb1e;
    ram_cell[     584] = 32'h0;  // 32'hde28143b;
    ram_cell[     585] = 32'h0;  // 32'h06f722c4;
    ram_cell[     586] = 32'h0;  // 32'h8093ddf9;
    ram_cell[     587] = 32'h0;  // 32'h6653c39e;
    ram_cell[     588] = 32'h0;  // 32'h0ae77601;
    ram_cell[     589] = 32'h0;  // 32'h7c876014;
    ram_cell[     590] = 32'h0;  // 32'h1931de40;
    ram_cell[     591] = 32'h0;  // 32'hfe11d84b;
    ram_cell[     592] = 32'h0;  // 32'hefeb6041;
    ram_cell[     593] = 32'h0;  // 32'hfe843cb6;
    ram_cell[     594] = 32'h0;  // 32'hcf922dc1;
    ram_cell[     595] = 32'h0;  // 32'h65a9bb05;
    ram_cell[     596] = 32'h0;  // 32'ha87f48e8;
    ram_cell[     597] = 32'h0;  // 32'h906afbcf;
    ram_cell[     598] = 32'h0;  // 32'ha2d3c228;
    ram_cell[     599] = 32'h0;  // 32'hfdd66240;
    ram_cell[     600] = 32'h0;  // 32'hc3f9a149;
    ram_cell[     601] = 32'h0;  // 32'h3f671819;
    ram_cell[     602] = 32'h0;  // 32'h40fe419f;
    ram_cell[     603] = 32'h0;  // 32'ha9cd65d1;
    ram_cell[     604] = 32'h0;  // 32'h157eb61e;
    ram_cell[     605] = 32'h0;  // 32'h4d2d0fa8;
    ram_cell[     606] = 32'h0;  // 32'hb7b4a282;
    ram_cell[     607] = 32'h0;  // 32'hd0f5fdfe;
    ram_cell[     608] = 32'h0;  // 32'hb58615b2;
    ram_cell[     609] = 32'h0;  // 32'h34dae1c8;
    ram_cell[     610] = 32'h0;  // 32'hd53539b1;
    ram_cell[     611] = 32'h0;  // 32'h9251c830;
    ram_cell[     612] = 32'h0;  // 32'h444168b1;
    ram_cell[     613] = 32'h0;  // 32'he29e3ef1;
    ram_cell[     614] = 32'h0;  // 32'hd6305426;
    ram_cell[     615] = 32'h0;  // 32'h33a159cc;
    ram_cell[     616] = 32'h0;  // 32'h133e9ef9;
    ram_cell[     617] = 32'h0;  // 32'hcdd1fd86;
    ram_cell[     618] = 32'h0;  // 32'h2f89a4cd;
    ram_cell[     619] = 32'h0;  // 32'h1ec66c6b;
    ram_cell[     620] = 32'h0;  // 32'h0f8e1240;
    ram_cell[     621] = 32'h0;  // 32'hc0a0c9e4;
    ram_cell[     622] = 32'h0;  // 32'h3e30d5cc;
    ram_cell[     623] = 32'h0;  // 32'h6cea19b6;
    ram_cell[     624] = 32'h0;  // 32'hed790945;
    ram_cell[     625] = 32'h0;  // 32'h8b309af3;
    ram_cell[     626] = 32'h0;  // 32'h88a2a2d0;
    ram_cell[     627] = 32'h0;  // 32'h6a771332;
    ram_cell[     628] = 32'h0;  // 32'hbae0ac69;
    ram_cell[     629] = 32'h0;  // 32'h892adf51;
    ram_cell[     630] = 32'h0;  // 32'hafe2157d;
    ram_cell[     631] = 32'h0;  // 32'h968fd4e7;
    ram_cell[     632] = 32'h0;  // 32'hb436a5b8;
    ram_cell[     633] = 32'h0;  // 32'h8c73c1c4;
    ram_cell[     634] = 32'h0;  // 32'h44e504d4;
    ram_cell[     635] = 32'h0;  // 32'h819046ad;
    ram_cell[     636] = 32'h0;  // 32'h7defb92a;
    ram_cell[     637] = 32'h0;  // 32'h2339d525;
    ram_cell[     638] = 32'h0;  // 32'h66d6c3a5;
    ram_cell[     639] = 32'h0;  // 32'he4afc6c3;
    ram_cell[     640] = 32'h0;  // 32'hac9d5d17;
    ram_cell[     641] = 32'h0;  // 32'hc8095eda;
    ram_cell[     642] = 32'h0;  // 32'h05926025;
    ram_cell[     643] = 32'h0;  // 32'hc50993b2;
    ram_cell[     644] = 32'h0;  // 32'hfd097015;
    ram_cell[     645] = 32'h0;  // 32'he3d1f4cf;
    ram_cell[     646] = 32'h0;  // 32'hef47d148;
    ram_cell[     647] = 32'h0;  // 32'hd456713d;
    ram_cell[     648] = 32'h0;  // 32'h97311aed;
    ram_cell[     649] = 32'h0;  // 32'hc2c5ba65;
    ram_cell[     650] = 32'h0;  // 32'h6741ced0;
    ram_cell[     651] = 32'h0;  // 32'h2ba96930;
    ram_cell[     652] = 32'h0;  // 32'h474bfa96;
    ram_cell[     653] = 32'h0;  // 32'hd58a9868;
    ram_cell[     654] = 32'h0;  // 32'hbd1070aa;
    ram_cell[     655] = 32'h0;  // 32'h1e68e7b5;
    ram_cell[     656] = 32'h0;  // 32'hb4fcf396;
    ram_cell[     657] = 32'h0;  // 32'hdee6a776;
    ram_cell[     658] = 32'h0;  // 32'hd361c774;
    ram_cell[     659] = 32'h0;  // 32'he605e380;
    ram_cell[     660] = 32'h0;  // 32'hd5175230;
    ram_cell[     661] = 32'h0;  // 32'h59f9212c;
    ram_cell[     662] = 32'h0;  // 32'hb6bd7071;
    ram_cell[     663] = 32'h0;  // 32'h043c5a75;
    ram_cell[     664] = 32'h0;  // 32'h90c74fe9;
    ram_cell[     665] = 32'h0;  // 32'h8692f08f;
    ram_cell[     666] = 32'h0;  // 32'h24bc2234;
    ram_cell[     667] = 32'h0;  // 32'hea55df2c;
    ram_cell[     668] = 32'h0;  // 32'h04556d8b;
    ram_cell[     669] = 32'h0;  // 32'hca7003e9;
    ram_cell[     670] = 32'h0;  // 32'hd9f8c1a4;
    ram_cell[     671] = 32'h0;  // 32'hcc24775a;
    ram_cell[     672] = 32'h0;  // 32'h57b0ef10;
    ram_cell[     673] = 32'h0;  // 32'h24c969ff;
    ram_cell[     674] = 32'h0;  // 32'h7fb0171e;
    ram_cell[     675] = 32'h0;  // 32'hd7a71bb5;
    ram_cell[     676] = 32'h0;  // 32'h9127d488;
    ram_cell[     677] = 32'h0;  // 32'hd4154de0;
    ram_cell[     678] = 32'h0;  // 32'h78b16d85;
    ram_cell[     679] = 32'h0;  // 32'h74f86d5e;
    ram_cell[     680] = 32'h0;  // 32'h09f07409;
    ram_cell[     681] = 32'h0;  // 32'ha5e174ae;
    ram_cell[     682] = 32'h0;  // 32'hc25bf53d;
    ram_cell[     683] = 32'h0;  // 32'h5491af59;
    ram_cell[     684] = 32'h0;  // 32'h79589fad;
    ram_cell[     685] = 32'h0;  // 32'hb5f7d6fa;
    ram_cell[     686] = 32'h0;  // 32'h76c7ecbb;
    ram_cell[     687] = 32'h0;  // 32'hdd181479;
    ram_cell[     688] = 32'h0;  // 32'h894de597;
    ram_cell[     689] = 32'h0;  // 32'h94bf2397;
    ram_cell[     690] = 32'h0;  // 32'h9d5c2378;
    ram_cell[     691] = 32'h0;  // 32'hba779fd2;
    ram_cell[     692] = 32'h0;  // 32'hb259652f;
    ram_cell[     693] = 32'h0;  // 32'h82774290;
    ram_cell[     694] = 32'h0;  // 32'hf90cffa6;
    ram_cell[     695] = 32'h0;  // 32'h6db886ad;
    ram_cell[     696] = 32'h0;  // 32'hb4c6cdf3;
    ram_cell[     697] = 32'h0;  // 32'h615bfffb;
    ram_cell[     698] = 32'h0;  // 32'hbb022a63;
    ram_cell[     699] = 32'h0;  // 32'h47540c0c;
    ram_cell[     700] = 32'h0;  // 32'h697e0d13;
    ram_cell[     701] = 32'h0;  // 32'h007b6758;
    ram_cell[     702] = 32'h0;  // 32'h6d1329b5;
    ram_cell[     703] = 32'h0;  // 32'hf2c76715;
    ram_cell[     704] = 32'h0;  // 32'h3d9c253f;
    ram_cell[     705] = 32'h0;  // 32'h67b6da85;
    ram_cell[     706] = 32'h0;  // 32'h11650f78;
    ram_cell[     707] = 32'h0;  // 32'h5ad56b84;
    ram_cell[     708] = 32'h0;  // 32'ha64aa866;
    ram_cell[     709] = 32'h0;  // 32'h2bac812d;
    ram_cell[     710] = 32'h0;  // 32'h810665a0;
    ram_cell[     711] = 32'h0;  // 32'he990228e;
    ram_cell[     712] = 32'h0;  // 32'h11b582b8;
    ram_cell[     713] = 32'h0;  // 32'hb0fc7f90;
    ram_cell[     714] = 32'h0;  // 32'hb45cfa52;
    ram_cell[     715] = 32'h0;  // 32'he7ba39c9;
    ram_cell[     716] = 32'h0;  // 32'h70b83d8f;
    ram_cell[     717] = 32'h0;  // 32'hd0fdaf8a;
    ram_cell[     718] = 32'h0;  // 32'h3bc224c9;
    ram_cell[     719] = 32'h0;  // 32'h9bef8e59;
    ram_cell[     720] = 32'h0;  // 32'hff40abf5;
    ram_cell[     721] = 32'h0;  // 32'h3bcfaab4;
    ram_cell[     722] = 32'h0;  // 32'h0accb1ed;
    ram_cell[     723] = 32'h0;  // 32'he8e9d2ea;
    ram_cell[     724] = 32'h0;  // 32'h8e850498;
    ram_cell[     725] = 32'h0;  // 32'h9f9b42fc;
    ram_cell[     726] = 32'h0;  // 32'he45984cf;
    ram_cell[     727] = 32'h0;  // 32'h27573151;
    ram_cell[     728] = 32'h0;  // 32'h47723749;
    ram_cell[     729] = 32'h0;  // 32'h4835cb55;
    ram_cell[     730] = 32'h0;  // 32'hc7fc1800;
    ram_cell[     731] = 32'h0;  // 32'h01382d7f;
    ram_cell[     732] = 32'h0;  // 32'h05b4319a;
    ram_cell[     733] = 32'h0;  // 32'h19817ab4;
    ram_cell[     734] = 32'h0;  // 32'hc1927ccf;
    ram_cell[     735] = 32'h0;  // 32'hf781351d;
    ram_cell[     736] = 32'h0;  // 32'hfd46f033;
    ram_cell[     737] = 32'h0;  // 32'h6a1320e9;
    ram_cell[     738] = 32'h0;  // 32'h77d95837;
    ram_cell[     739] = 32'h0;  // 32'h90457af9;
    ram_cell[     740] = 32'h0;  // 32'h21a333b0;
    ram_cell[     741] = 32'h0;  // 32'h3c4b7c4b;
    ram_cell[     742] = 32'h0;  // 32'hf974ad79;
    ram_cell[     743] = 32'h0;  // 32'h94f27cc0;
    ram_cell[     744] = 32'h0;  // 32'h88daecd2;
    ram_cell[     745] = 32'h0;  // 32'h47dd9e45;
    ram_cell[     746] = 32'h0;  // 32'he30344b0;
    ram_cell[     747] = 32'h0;  // 32'ha08f36a0;
    ram_cell[     748] = 32'h0;  // 32'h0078a348;
    ram_cell[     749] = 32'h0;  // 32'h08675b9a;
    ram_cell[     750] = 32'h0;  // 32'ha4369925;
    ram_cell[     751] = 32'h0;  // 32'h7f62d93d;
    ram_cell[     752] = 32'h0;  // 32'h9448081b;
    ram_cell[     753] = 32'h0;  // 32'h6b5d44af;
    ram_cell[     754] = 32'h0;  // 32'hb5a33152;
    ram_cell[     755] = 32'h0;  // 32'hfbea6089;
    ram_cell[     756] = 32'h0;  // 32'h5e799192;
    ram_cell[     757] = 32'h0;  // 32'h8d026f04;
    ram_cell[     758] = 32'h0;  // 32'h766717d6;
    ram_cell[     759] = 32'h0;  // 32'h7276244b;
    ram_cell[     760] = 32'h0;  // 32'h2644ffb4;
    ram_cell[     761] = 32'h0;  // 32'h09a70430;
    ram_cell[     762] = 32'h0;  // 32'h6da8e30f;
    ram_cell[     763] = 32'h0;  // 32'hc784c1e6;
    ram_cell[     764] = 32'h0;  // 32'h0ce6ddce;
    ram_cell[     765] = 32'h0;  // 32'h167fb175;
    ram_cell[     766] = 32'h0;  // 32'h98ceb002;
    ram_cell[     767] = 32'h0;  // 32'heced95eb;
    ram_cell[     768] = 32'h0;  // 32'h19cfaf70;
    ram_cell[     769] = 32'h0;  // 32'h9ff0e0a3;
    ram_cell[     770] = 32'h0;  // 32'h9b619f36;
    ram_cell[     771] = 32'h0;  // 32'he36c3e71;
    ram_cell[     772] = 32'h0;  // 32'h44efd6e7;
    ram_cell[     773] = 32'h0;  // 32'he6c8b6ee;
    ram_cell[     774] = 32'h0;  // 32'h63cda373;
    ram_cell[     775] = 32'h0;  // 32'hef70277e;
    ram_cell[     776] = 32'h0;  // 32'h60f8702e;
    ram_cell[     777] = 32'h0;  // 32'h2347f351;
    ram_cell[     778] = 32'h0;  // 32'h50d4e3c1;
    ram_cell[     779] = 32'h0;  // 32'h3e1b9e04;
    ram_cell[     780] = 32'h0;  // 32'hc8d5cc03;
    ram_cell[     781] = 32'h0;  // 32'h52b1bb65;
    ram_cell[     782] = 32'h0;  // 32'h97277664;
    ram_cell[     783] = 32'h0;  // 32'h6f7e7c89;
    ram_cell[     784] = 32'h0;  // 32'h56ef3096;
    ram_cell[     785] = 32'h0;  // 32'h25862acf;
    ram_cell[     786] = 32'h0;  // 32'h1b2205a3;
    ram_cell[     787] = 32'h0;  // 32'heb454672;
    ram_cell[     788] = 32'h0;  // 32'ha367dc8b;
    ram_cell[     789] = 32'h0;  // 32'h62856fde;
    ram_cell[     790] = 32'h0;  // 32'h31efde08;
    ram_cell[     791] = 32'h0;  // 32'h05b7bacd;
    ram_cell[     792] = 32'h0;  // 32'h57277e1a;
    ram_cell[     793] = 32'h0;  // 32'h8294fed5;
    ram_cell[     794] = 32'h0;  // 32'h07e63b18;
    ram_cell[     795] = 32'h0;  // 32'hb744b430;
    ram_cell[     796] = 32'h0;  // 32'hdb8a6e27;
    ram_cell[     797] = 32'h0;  // 32'h48dd2e19;
    ram_cell[     798] = 32'h0;  // 32'h13a93d33;
    ram_cell[     799] = 32'h0;  // 32'h1b4669c7;
    ram_cell[     800] = 32'h0;  // 32'h937308cf;
    ram_cell[     801] = 32'h0;  // 32'ha421a9a8;
    ram_cell[     802] = 32'h0;  // 32'hb50d804b;
    ram_cell[     803] = 32'h0;  // 32'hbc1ae33d;
    ram_cell[     804] = 32'h0;  // 32'h0b6c9f79;
    ram_cell[     805] = 32'h0;  // 32'h01ff9d89;
    ram_cell[     806] = 32'h0;  // 32'ha4be9a37;
    ram_cell[     807] = 32'h0;  // 32'hff6f7c85;
    ram_cell[     808] = 32'h0;  // 32'h58b918a6;
    ram_cell[     809] = 32'h0;  // 32'h8bf486ce;
    ram_cell[     810] = 32'h0;  // 32'h28dbb2ff;
    ram_cell[     811] = 32'h0;  // 32'hfc1eabc5;
    ram_cell[     812] = 32'h0;  // 32'hba0164d0;
    ram_cell[     813] = 32'h0;  // 32'he7d75af4;
    ram_cell[     814] = 32'h0;  // 32'h99ac0886;
    ram_cell[     815] = 32'h0;  // 32'h84382aef;
    ram_cell[     816] = 32'h0;  // 32'h1a72aeb1;
    ram_cell[     817] = 32'h0;  // 32'hc3025690;
    ram_cell[     818] = 32'h0;  // 32'hec86c7ff;
    ram_cell[     819] = 32'h0;  // 32'h88eebc31;
    ram_cell[     820] = 32'h0;  // 32'h8d94ecf4;
    ram_cell[     821] = 32'h0;  // 32'h2b2dc464;
    ram_cell[     822] = 32'h0;  // 32'he1a64c4d;
    ram_cell[     823] = 32'h0;  // 32'hc4b38ed8;
    ram_cell[     824] = 32'h0;  // 32'h3f063ff5;
    ram_cell[     825] = 32'h0;  // 32'h14f0fa6e;
    ram_cell[     826] = 32'h0;  // 32'ha90b6448;
    ram_cell[     827] = 32'h0;  // 32'h59e2b73f;
    ram_cell[     828] = 32'h0;  // 32'h9d422321;
    ram_cell[     829] = 32'h0;  // 32'hf15da213;
    ram_cell[     830] = 32'h0;  // 32'h6129388c;
    ram_cell[     831] = 32'h0;  // 32'he65275f6;
    ram_cell[     832] = 32'h0;  // 32'h05a8f9f8;
    ram_cell[     833] = 32'h0;  // 32'h01b415c4;
    ram_cell[     834] = 32'h0;  // 32'hf66d7ef9;
    ram_cell[     835] = 32'h0;  // 32'hef90664c;
    ram_cell[     836] = 32'h0;  // 32'hc3655491;
    ram_cell[     837] = 32'h0;  // 32'h13a98f9e;
    ram_cell[     838] = 32'h0;  // 32'h5acab93b;
    ram_cell[     839] = 32'h0;  // 32'hc98eda96;
    ram_cell[     840] = 32'h0;  // 32'h65753b47;
    ram_cell[     841] = 32'h0;  // 32'hd73bfa11;
    ram_cell[     842] = 32'h0;  // 32'hc1ceb3e0;
    ram_cell[     843] = 32'h0;  // 32'hc41bd75f;
    ram_cell[     844] = 32'h0;  // 32'h29cabcee;
    ram_cell[     845] = 32'h0;  // 32'h0569eb07;
    ram_cell[     846] = 32'h0;  // 32'ha355e5a4;
    ram_cell[     847] = 32'h0;  // 32'hac68503a;
    ram_cell[     848] = 32'h0;  // 32'h40628111;
    ram_cell[     849] = 32'h0;  // 32'h5767f16a;
    ram_cell[     850] = 32'h0;  // 32'h78d5e437;
    ram_cell[     851] = 32'h0;  // 32'h7527b341;
    ram_cell[     852] = 32'h0;  // 32'hf4746647;
    ram_cell[     853] = 32'h0;  // 32'h7874c43a;
    ram_cell[     854] = 32'h0;  // 32'h33c6c0c7;
    ram_cell[     855] = 32'h0;  // 32'ha62edc0d;
    ram_cell[     856] = 32'h0;  // 32'h610c8764;
    ram_cell[     857] = 32'h0;  // 32'hbbc18266;
    ram_cell[     858] = 32'h0;  // 32'h5c8e0674;
    ram_cell[     859] = 32'h0;  // 32'hd92c5e25;
    ram_cell[     860] = 32'h0;  // 32'h9fbada59;
    ram_cell[     861] = 32'h0;  // 32'hf4c2497c;
    ram_cell[     862] = 32'h0;  // 32'hddccf9ba;
    ram_cell[     863] = 32'h0;  // 32'h70cde9c1;
    ram_cell[     864] = 32'h0;  // 32'h5c7dfb87;
    ram_cell[     865] = 32'h0;  // 32'hb767f5c1;
    ram_cell[     866] = 32'h0;  // 32'h7193b039;
    ram_cell[     867] = 32'h0;  // 32'hb8513ede;
    ram_cell[     868] = 32'h0;  // 32'h0a878e82;
    ram_cell[     869] = 32'h0;  // 32'hdee27dca;
    ram_cell[     870] = 32'h0;  // 32'hfa911b2f;
    ram_cell[     871] = 32'h0;  // 32'hadaf2437;
    ram_cell[     872] = 32'h0;  // 32'haf1228df;
    ram_cell[     873] = 32'h0;  // 32'hf13d67d2;
    ram_cell[     874] = 32'h0;  // 32'hc5bcfdfc;
    ram_cell[     875] = 32'h0;  // 32'hb6ee59d5;
    ram_cell[     876] = 32'h0;  // 32'h3113e703;
    ram_cell[     877] = 32'h0;  // 32'hbae8a7cc;
    ram_cell[     878] = 32'h0;  // 32'hd770c705;
    ram_cell[     879] = 32'h0;  // 32'ha47352aa;
    ram_cell[     880] = 32'h0;  // 32'hbdfbabc0;
    ram_cell[     881] = 32'h0;  // 32'hdbd7d757;
    ram_cell[     882] = 32'h0;  // 32'hd6680b48;
    ram_cell[     883] = 32'h0;  // 32'h546b527f;
    ram_cell[     884] = 32'h0;  // 32'hfcc61757;
    ram_cell[     885] = 32'h0;  // 32'h7bcc77c5;
    ram_cell[     886] = 32'h0;  // 32'hd1c82e7d;
    ram_cell[     887] = 32'h0;  // 32'h08ba92e5;
    ram_cell[     888] = 32'h0;  // 32'hdf6f2623;
    ram_cell[     889] = 32'h0;  // 32'h7191d400;
    ram_cell[     890] = 32'h0;  // 32'h5f855af1;
    ram_cell[     891] = 32'h0;  // 32'h9e5af64f;
    ram_cell[     892] = 32'h0;  // 32'h707e3908;
    ram_cell[     893] = 32'h0;  // 32'h5175e561;
    ram_cell[     894] = 32'h0;  // 32'h07f3c8c9;
    ram_cell[     895] = 32'h0;  // 32'h3c21dc45;
    ram_cell[     896] = 32'h0;  // 32'h9e8bfee0;
    ram_cell[     897] = 32'h0;  // 32'h89985e9b;
    ram_cell[     898] = 32'h0;  // 32'h10da453b;
    ram_cell[     899] = 32'h0;  // 32'h6d8bde53;
    ram_cell[     900] = 32'h0;  // 32'h3d15b443;
    ram_cell[     901] = 32'h0;  // 32'h6b819a6a;
    ram_cell[     902] = 32'h0;  // 32'he8c2a5fa;
    ram_cell[     903] = 32'h0;  // 32'h669a4f56;
    ram_cell[     904] = 32'h0;  // 32'hf4566d88;
    ram_cell[     905] = 32'h0;  // 32'hfe9680fb;
    ram_cell[     906] = 32'h0;  // 32'he1d6c1e9;
    ram_cell[     907] = 32'h0;  // 32'h584dc2b6;
    ram_cell[     908] = 32'h0;  // 32'h376ee917;
    ram_cell[     909] = 32'h0;  // 32'h3726d380;
    ram_cell[     910] = 32'h0;  // 32'h46b8997a;
    ram_cell[     911] = 32'h0;  // 32'h667b4d53;
    ram_cell[     912] = 32'h0;  // 32'hf30fba3a;
    ram_cell[     913] = 32'h0;  // 32'hf28e9bbd;
    ram_cell[     914] = 32'h0;  // 32'h95eceedb;
    ram_cell[     915] = 32'h0;  // 32'h9919533c;
    ram_cell[     916] = 32'h0;  // 32'h2667594f;
    ram_cell[     917] = 32'h0;  // 32'h9059aa08;
    ram_cell[     918] = 32'h0;  // 32'hf286d45f;
    ram_cell[     919] = 32'h0;  // 32'h21461e9a;
    ram_cell[     920] = 32'h0;  // 32'h58449a2c;
    ram_cell[     921] = 32'h0;  // 32'h772cf4dc;
    ram_cell[     922] = 32'h0;  // 32'hd699dea2;
    ram_cell[     923] = 32'h0;  // 32'h70d2c1e3;
    ram_cell[     924] = 32'h0;  // 32'h151c2ee0;
    ram_cell[     925] = 32'h0;  // 32'h9bf922f8;
    ram_cell[     926] = 32'h0;  // 32'h80009933;
    ram_cell[     927] = 32'h0;  // 32'h2cf44791;
    ram_cell[     928] = 32'h0;  // 32'hd15f1de2;
    ram_cell[     929] = 32'h0;  // 32'hecfb2514;
    ram_cell[     930] = 32'h0;  // 32'h05ca574b;
    ram_cell[     931] = 32'h0;  // 32'he8b85b39;
    ram_cell[     932] = 32'h0;  // 32'h44831bb1;
    ram_cell[     933] = 32'h0;  // 32'hf274ea73;
    ram_cell[     934] = 32'h0;  // 32'h11815770;
    ram_cell[     935] = 32'h0;  // 32'h725b2c56;
    ram_cell[     936] = 32'h0;  // 32'habf311f6;
    ram_cell[     937] = 32'h0;  // 32'h23da5f4d;
    ram_cell[     938] = 32'h0;  // 32'he2f48250;
    ram_cell[     939] = 32'h0;  // 32'h9e6d9824;
    ram_cell[     940] = 32'h0;  // 32'hcd0ad7cf;
    ram_cell[     941] = 32'h0;  // 32'hf5be6879;
    ram_cell[     942] = 32'h0;  // 32'h0dddaa2d;
    ram_cell[     943] = 32'h0;  // 32'h4d0f37be;
    ram_cell[     944] = 32'h0;  // 32'hcb7d99c9;
    ram_cell[     945] = 32'h0;  // 32'ha6bbf3e3;
    ram_cell[     946] = 32'h0;  // 32'h18571f5e;
    ram_cell[     947] = 32'h0;  // 32'ha5958ac4;
    ram_cell[     948] = 32'h0;  // 32'h6043bd25;
    ram_cell[     949] = 32'h0;  // 32'hbe8103af;
    ram_cell[     950] = 32'h0;  // 32'h7e6c13a6;
    ram_cell[     951] = 32'h0;  // 32'hfd1caa7e;
    ram_cell[     952] = 32'h0;  // 32'h42fc559e;
    ram_cell[     953] = 32'h0;  // 32'h76edc8fa;
    ram_cell[     954] = 32'h0;  // 32'hb63bd145;
    ram_cell[     955] = 32'h0;  // 32'h1e227c78;
    ram_cell[     956] = 32'h0;  // 32'h25e9ed3d;
    ram_cell[     957] = 32'h0;  // 32'h72dbabc5;
    ram_cell[     958] = 32'h0;  // 32'h210b9833;
    ram_cell[     959] = 32'h0;  // 32'h0d122b1b;
    ram_cell[     960] = 32'h0;  // 32'h126d8f7b;
    ram_cell[     961] = 32'h0;  // 32'ha3dcb1df;
    ram_cell[     962] = 32'h0;  // 32'h897fa936;
    ram_cell[     963] = 32'h0;  // 32'h944fcb42;
    ram_cell[     964] = 32'h0;  // 32'h3e645756;
    ram_cell[     965] = 32'h0;  // 32'hbce154bc;
    ram_cell[     966] = 32'h0;  // 32'h34f9a34d;
    ram_cell[     967] = 32'h0;  // 32'hdb59316c;
    ram_cell[     968] = 32'h0;  // 32'h56775f71;
    ram_cell[     969] = 32'h0;  // 32'hcea7503d;
    ram_cell[     970] = 32'h0;  // 32'ha7b09b67;
    ram_cell[     971] = 32'h0;  // 32'hfdd90b22;
    ram_cell[     972] = 32'h0;  // 32'h9cd5c2b5;
    ram_cell[     973] = 32'h0;  // 32'h08432dd3;
    ram_cell[     974] = 32'h0;  // 32'hf2ff4554;
    ram_cell[     975] = 32'h0;  // 32'h1a8f218c;
    ram_cell[     976] = 32'h0;  // 32'h74f3f7a8;
    ram_cell[     977] = 32'h0;  // 32'h13b2b4f4;
    ram_cell[     978] = 32'h0;  // 32'hff7efad0;
    ram_cell[     979] = 32'h0;  // 32'h5077ca02;
    ram_cell[     980] = 32'h0;  // 32'h93cd2c4d;
    ram_cell[     981] = 32'h0;  // 32'h47990589;
    ram_cell[     982] = 32'h0;  // 32'h53a40caa;
    ram_cell[     983] = 32'h0;  // 32'h4a703486;
    ram_cell[     984] = 32'h0;  // 32'hb25dc70a;
    ram_cell[     985] = 32'h0;  // 32'hff0db6ae;
    ram_cell[     986] = 32'h0;  // 32'h414ac351;
    ram_cell[     987] = 32'h0;  // 32'hb2c277b1;
    ram_cell[     988] = 32'h0;  // 32'h3801ce4e;
    ram_cell[     989] = 32'h0;  // 32'ha4abb19b;
    ram_cell[     990] = 32'h0;  // 32'h7b3b07df;
    ram_cell[     991] = 32'h0;  // 32'hc635e674;
    ram_cell[     992] = 32'h0;  // 32'ha0eca175;
    ram_cell[     993] = 32'h0;  // 32'h1486b36f;
    ram_cell[     994] = 32'h0;  // 32'h2360f826;
    ram_cell[     995] = 32'h0;  // 32'hb6b57293;
    ram_cell[     996] = 32'h0;  // 32'h8d1a901a;
    ram_cell[     997] = 32'h0;  // 32'h6be0333e;
    ram_cell[     998] = 32'h0;  // 32'h6ddb7457;
    ram_cell[     999] = 32'h0;  // 32'haea25c91;
    ram_cell[    1000] = 32'h0;  // 32'hf399d4ee;
    ram_cell[    1001] = 32'h0;  // 32'h0edfb9e2;
    ram_cell[    1002] = 32'h0;  // 32'h439778cd;
    ram_cell[    1003] = 32'h0;  // 32'h83138afb;
    ram_cell[    1004] = 32'h0;  // 32'h5ed2c0ca;
    ram_cell[    1005] = 32'h0;  // 32'h861ebfd1;
    ram_cell[    1006] = 32'h0;  // 32'h58fc28bf;
    ram_cell[    1007] = 32'h0;  // 32'h9734951b;
    ram_cell[    1008] = 32'h0;  // 32'h08c141b9;
    ram_cell[    1009] = 32'h0;  // 32'hcff444e7;
    ram_cell[    1010] = 32'h0;  // 32'h6cedca64;
    ram_cell[    1011] = 32'h0;  // 32'h95b88f3a;
    ram_cell[    1012] = 32'h0;  // 32'hf5d89fe1;
    ram_cell[    1013] = 32'h0;  // 32'hf10e3eeb;
    ram_cell[    1014] = 32'h0;  // 32'h28a104eb;
    ram_cell[    1015] = 32'h0;  // 32'h71368e34;
    ram_cell[    1016] = 32'h0;  // 32'h3ec20b5f;
    ram_cell[    1017] = 32'h0;  // 32'he6ac87c0;
    ram_cell[    1018] = 32'h0;  // 32'h3fa69436;
    ram_cell[    1019] = 32'h0;  // 32'hd06d3417;
    ram_cell[    1020] = 32'h0;  // 32'h586951da;
    ram_cell[    1021] = 32'h0;  // 32'h7df4aea3;
    ram_cell[    1022] = 32'h0;  // 32'hc611979f;
    ram_cell[    1023] = 32'h0;  // 32'h3e427e68;
    ram_cell[    1024] = 32'h0;  // 32'h62c30f63;
    ram_cell[    1025] = 32'h0;  // 32'hd922b076;
    ram_cell[    1026] = 32'h0;  // 32'heda6ff80;
    ram_cell[    1027] = 32'h0;  // 32'h882aebd9;
    ram_cell[    1028] = 32'h0;  // 32'h47660aee;
    ram_cell[    1029] = 32'h0;  // 32'h00e34672;
    ram_cell[    1030] = 32'h0;  // 32'h05339e0f;
    ram_cell[    1031] = 32'h0;  // 32'h1e44e5d9;
    ram_cell[    1032] = 32'h0;  // 32'hfbcc972d;
    ram_cell[    1033] = 32'h0;  // 32'h8d92d779;
    ram_cell[    1034] = 32'h0;  // 32'hab45880b;
    ram_cell[    1035] = 32'h0;  // 32'h457a6dd3;
    ram_cell[    1036] = 32'h0;  // 32'h27d05989;
    ram_cell[    1037] = 32'h0;  // 32'h0187b032;
    ram_cell[    1038] = 32'h0;  // 32'h4216baf9;
    ram_cell[    1039] = 32'h0;  // 32'hea82ff2f;
    ram_cell[    1040] = 32'h0;  // 32'h00bf78ea;
    ram_cell[    1041] = 32'h0;  // 32'hb736b57c;
    ram_cell[    1042] = 32'h0;  // 32'hf5a09ae7;
    ram_cell[    1043] = 32'h0;  // 32'hb5548f00;
    ram_cell[    1044] = 32'h0;  // 32'h44efe13f;
    ram_cell[    1045] = 32'h0;  // 32'h0f10c3cd;
    ram_cell[    1046] = 32'h0;  // 32'h3b9b3b1b;
    ram_cell[    1047] = 32'h0;  // 32'hdac9be44;
    ram_cell[    1048] = 32'h0;  // 32'h961e6ffa;
    ram_cell[    1049] = 32'h0;  // 32'hbc5e9bec;
    ram_cell[    1050] = 32'h0;  // 32'h9dddd846;
    ram_cell[    1051] = 32'h0;  // 32'hfba02262;
    ram_cell[    1052] = 32'h0;  // 32'h00f2b1ac;
    ram_cell[    1053] = 32'h0;  // 32'h177a17a0;
    ram_cell[    1054] = 32'h0;  // 32'hd8a1c4d6;
    ram_cell[    1055] = 32'h0;  // 32'h86a880c6;
    ram_cell[    1056] = 32'h0;  // 32'hcfcdfe8d;
    ram_cell[    1057] = 32'h0;  // 32'h6b27a782;
    ram_cell[    1058] = 32'h0;  // 32'h9edc9643;
    ram_cell[    1059] = 32'h0;  // 32'hf183ad12;
    ram_cell[    1060] = 32'h0;  // 32'h99900c67;
    ram_cell[    1061] = 32'h0;  // 32'he68d7277;
    ram_cell[    1062] = 32'h0;  // 32'h0d9e8d11;
    ram_cell[    1063] = 32'h0;  // 32'h26a82ab4;
    ram_cell[    1064] = 32'h0;  // 32'hd80bb7c7;
    ram_cell[    1065] = 32'h0;  // 32'h00fc66a1;
    ram_cell[    1066] = 32'h0;  // 32'h6a4b8ce1;
    ram_cell[    1067] = 32'h0;  // 32'hdc5079aa;
    ram_cell[    1068] = 32'h0;  // 32'h91fdfc6b;
    ram_cell[    1069] = 32'h0;  // 32'h6c72af97;
    ram_cell[    1070] = 32'h0;  // 32'h058bc936;
    ram_cell[    1071] = 32'h0;  // 32'hf38e490f;
    ram_cell[    1072] = 32'h0;  // 32'ha9bf973b;
    ram_cell[    1073] = 32'h0;  // 32'h45cdd392;
    ram_cell[    1074] = 32'h0;  // 32'hbd37238a;
    ram_cell[    1075] = 32'h0;  // 32'h78701d9a;
    ram_cell[    1076] = 32'h0;  // 32'hf9d67fb1;
    ram_cell[    1077] = 32'h0;  // 32'h4f850760;
    ram_cell[    1078] = 32'h0;  // 32'hc54ec1ee;
    ram_cell[    1079] = 32'h0;  // 32'hab5a91ab;
    ram_cell[    1080] = 32'h0;  // 32'ha3568257;
    ram_cell[    1081] = 32'h0;  // 32'he0d9fdb6;
    ram_cell[    1082] = 32'h0;  // 32'hf79512f2;
    ram_cell[    1083] = 32'h0;  // 32'hdec4f132;
    ram_cell[    1084] = 32'h0;  // 32'h32b380a4;
    ram_cell[    1085] = 32'h0;  // 32'h2b40a796;
    ram_cell[    1086] = 32'h0;  // 32'ha0c85ab6;
    ram_cell[    1087] = 32'h0;  // 32'h4e0f9e35;
    ram_cell[    1088] = 32'h0;  // 32'hd56696e5;
    ram_cell[    1089] = 32'h0;  // 32'h89967d0e;
    ram_cell[    1090] = 32'h0;  // 32'h05030d20;
    ram_cell[    1091] = 32'h0;  // 32'h20a71e60;
    ram_cell[    1092] = 32'h0;  // 32'haff84b70;
    ram_cell[    1093] = 32'h0;  // 32'h48ca36ee;
    ram_cell[    1094] = 32'h0;  // 32'hd6494bea;
    ram_cell[    1095] = 32'h0;  // 32'h1a3aed4a;
    ram_cell[    1096] = 32'h0;  // 32'hedd8dea4;
    ram_cell[    1097] = 32'h0;  // 32'hbfbb2b72;
    ram_cell[    1098] = 32'h0;  // 32'h12e42cad;
    ram_cell[    1099] = 32'h0;  // 32'h7a427e24;
    ram_cell[    1100] = 32'h0;  // 32'h7eb85482;
    ram_cell[    1101] = 32'h0;  // 32'h80101233;
    ram_cell[    1102] = 32'h0;  // 32'h3275bf72;
    ram_cell[    1103] = 32'h0;  // 32'h296d6d5d;
    ram_cell[    1104] = 32'h0;  // 32'hb829c213;
    ram_cell[    1105] = 32'h0;  // 32'hd2ce7da4;
    ram_cell[    1106] = 32'h0;  // 32'h9815e873;
    ram_cell[    1107] = 32'h0;  // 32'h67392747;
    ram_cell[    1108] = 32'h0;  // 32'h51327b75;
    ram_cell[    1109] = 32'h0;  // 32'hece530d2;
    ram_cell[    1110] = 32'h0;  // 32'h7acdbc76;
    ram_cell[    1111] = 32'h0;  // 32'h746ac487;
    ram_cell[    1112] = 32'h0;  // 32'hf029d045;
    ram_cell[    1113] = 32'h0;  // 32'h64be4346;
    ram_cell[    1114] = 32'h0;  // 32'h32d55cd5;
    ram_cell[    1115] = 32'h0;  // 32'h92c7e317;
    ram_cell[    1116] = 32'h0;  // 32'hd3be5a90;
    ram_cell[    1117] = 32'h0;  // 32'h633cf709;
    ram_cell[    1118] = 32'h0;  // 32'hdf3d52e6;
    ram_cell[    1119] = 32'h0;  // 32'h3890192b;
    ram_cell[    1120] = 32'h0;  // 32'hd793dfd8;
    ram_cell[    1121] = 32'h0;  // 32'h522fb61c;
    ram_cell[    1122] = 32'h0;  // 32'h7bd1361c;
    ram_cell[    1123] = 32'h0;  // 32'heb73e509;
    ram_cell[    1124] = 32'h0;  // 32'h7b0829b6;
    ram_cell[    1125] = 32'h0;  // 32'he1cba561;
    ram_cell[    1126] = 32'h0;  // 32'hc58117d0;
    ram_cell[    1127] = 32'h0;  // 32'h7ba2ea4f;
    ram_cell[    1128] = 32'h0;  // 32'he591d1ff;
    ram_cell[    1129] = 32'h0;  // 32'hc18fbc74;
    ram_cell[    1130] = 32'h0;  // 32'ha7738634;
    ram_cell[    1131] = 32'h0;  // 32'hc6eee2ee;
    ram_cell[    1132] = 32'h0;  // 32'h41cfb1b1;
    ram_cell[    1133] = 32'h0;  // 32'h53fbdf6d;
    ram_cell[    1134] = 32'h0;  // 32'hfbba4a62;
    ram_cell[    1135] = 32'h0;  // 32'h2f79e164;
    ram_cell[    1136] = 32'h0;  // 32'h492df19e;
    ram_cell[    1137] = 32'h0;  // 32'h7e43801b;
    ram_cell[    1138] = 32'h0;  // 32'h26bca0df;
    ram_cell[    1139] = 32'h0;  // 32'h29454c91;
    ram_cell[    1140] = 32'h0;  // 32'h91b43d18;
    ram_cell[    1141] = 32'h0;  // 32'h8746e722;
    ram_cell[    1142] = 32'h0;  // 32'h34c60762;
    ram_cell[    1143] = 32'h0;  // 32'h19b52b20;
    ram_cell[    1144] = 32'h0;  // 32'h5c941cb5;
    ram_cell[    1145] = 32'h0;  // 32'h7450a8b7;
    ram_cell[    1146] = 32'h0;  // 32'hc0fba47f;
    ram_cell[    1147] = 32'h0;  // 32'h89c272f7;
    ram_cell[    1148] = 32'h0;  // 32'h4db5be5e;
    ram_cell[    1149] = 32'h0;  // 32'h9a8d92f7;
    ram_cell[    1150] = 32'h0;  // 32'h752c7e06;
    ram_cell[    1151] = 32'h0;  // 32'h4ec1a720;
    ram_cell[    1152] = 32'h0;  // 32'hac2688f0;
    ram_cell[    1153] = 32'h0;  // 32'h3a438833;
    ram_cell[    1154] = 32'h0;  // 32'h81167a96;
    ram_cell[    1155] = 32'h0;  // 32'h5e026861;
    ram_cell[    1156] = 32'h0;  // 32'he8085c6a;
    ram_cell[    1157] = 32'h0;  // 32'h4d2d0f51;
    ram_cell[    1158] = 32'h0;  // 32'h6fa93783;
    ram_cell[    1159] = 32'h0;  // 32'hac338a17;
    ram_cell[    1160] = 32'h0;  // 32'he3773275;
    ram_cell[    1161] = 32'h0;  // 32'h496b5642;
    ram_cell[    1162] = 32'h0;  // 32'h0d3a070c;
    ram_cell[    1163] = 32'h0;  // 32'he9b512a3;
    ram_cell[    1164] = 32'h0;  // 32'h983ddd25;
    ram_cell[    1165] = 32'h0;  // 32'h400bae5c;
    ram_cell[    1166] = 32'h0;  // 32'h3761df0b;
    ram_cell[    1167] = 32'h0;  // 32'h81f24c0a;
    ram_cell[    1168] = 32'h0;  // 32'h1dd67839;
    ram_cell[    1169] = 32'h0;  // 32'hce3bd629;
    ram_cell[    1170] = 32'h0;  // 32'he4830cd0;
    ram_cell[    1171] = 32'h0;  // 32'h2776a2bb;
    ram_cell[    1172] = 32'h0;  // 32'h60f41a76;
    ram_cell[    1173] = 32'h0;  // 32'hebcbc46d;
    ram_cell[    1174] = 32'h0;  // 32'hef189bb9;
    ram_cell[    1175] = 32'h0;  // 32'hcef530be;
    ram_cell[    1176] = 32'h0;  // 32'hca06e200;
    ram_cell[    1177] = 32'h0;  // 32'h71adb1f9;
    ram_cell[    1178] = 32'h0;  // 32'h1159f05a;
    ram_cell[    1179] = 32'h0;  // 32'h21064ff5;
    ram_cell[    1180] = 32'h0;  // 32'h4b976e2a;
    ram_cell[    1181] = 32'h0;  // 32'h3b6856bc;
    ram_cell[    1182] = 32'h0;  // 32'h0d83958c;
    ram_cell[    1183] = 32'h0;  // 32'h242dbde8;
    ram_cell[    1184] = 32'h0;  // 32'h6a9275f3;
    ram_cell[    1185] = 32'h0;  // 32'h9cdffdfd;
    ram_cell[    1186] = 32'h0;  // 32'h6add3aff;
    ram_cell[    1187] = 32'h0;  // 32'h2b2b0435;
    ram_cell[    1188] = 32'h0;  // 32'heb896db2;
    ram_cell[    1189] = 32'h0;  // 32'h9f22b7e0;
    ram_cell[    1190] = 32'h0;  // 32'hcf4c60c4;
    ram_cell[    1191] = 32'h0;  // 32'hdd684c84;
    ram_cell[    1192] = 32'h0;  // 32'h1c79cfe0;
    ram_cell[    1193] = 32'h0;  // 32'h3769ec72;
    ram_cell[    1194] = 32'h0;  // 32'h71345bb8;
    ram_cell[    1195] = 32'h0;  // 32'h9de75d06;
    ram_cell[    1196] = 32'h0;  // 32'h3f1c1fce;
    ram_cell[    1197] = 32'h0;  // 32'h24f3b2c3;
    ram_cell[    1198] = 32'h0;  // 32'h5062d90c;
    ram_cell[    1199] = 32'h0;  // 32'hc416f1d4;
    ram_cell[    1200] = 32'h0;  // 32'h0a275756;
    ram_cell[    1201] = 32'h0;  // 32'h2cdc1733;
    ram_cell[    1202] = 32'h0;  // 32'hf80db7e0;
    ram_cell[    1203] = 32'h0;  // 32'he73ea4de;
    ram_cell[    1204] = 32'h0;  // 32'h80a78270;
    ram_cell[    1205] = 32'h0;  // 32'hc917b2ef;
    ram_cell[    1206] = 32'h0;  // 32'hb9a782b8;
    ram_cell[    1207] = 32'h0;  // 32'he819780c;
    ram_cell[    1208] = 32'h0;  // 32'hdb330064;
    ram_cell[    1209] = 32'h0;  // 32'hc0c9cbe9;
    ram_cell[    1210] = 32'h0;  // 32'h87e98065;
    ram_cell[    1211] = 32'h0;  // 32'h0dd2f156;
    ram_cell[    1212] = 32'h0;  // 32'h8ebbc107;
    ram_cell[    1213] = 32'h0;  // 32'h2a77c646;
    ram_cell[    1214] = 32'h0;  // 32'h98a1d74b;
    ram_cell[    1215] = 32'h0;  // 32'ha294f377;
    ram_cell[    1216] = 32'h0;  // 32'hc860f741;
    ram_cell[    1217] = 32'h0;  // 32'hdca17b3d;
    ram_cell[    1218] = 32'h0;  // 32'h18657bf1;
    ram_cell[    1219] = 32'h0;  // 32'h5ba766b7;
    ram_cell[    1220] = 32'h0;  // 32'h936cb5da;
    ram_cell[    1221] = 32'h0;  // 32'h428c78bc;
    ram_cell[    1222] = 32'h0;  // 32'h57065a24;
    ram_cell[    1223] = 32'h0;  // 32'h140dbded;
    ram_cell[    1224] = 32'h0;  // 32'h20b0b2df;
    ram_cell[    1225] = 32'h0;  // 32'h711fbb7a;
    ram_cell[    1226] = 32'h0;  // 32'h520f6825;
    ram_cell[    1227] = 32'h0;  // 32'h71e25790;
    ram_cell[    1228] = 32'h0;  // 32'hf9c39147;
    ram_cell[    1229] = 32'h0;  // 32'hd1e6330c;
    ram_cell[    1230] = 32'h0;  // 32'h19a60e92;
    ram_cell[    1231] = 32'h0;  // 32'h62c96cd0;
    ram_cell[    1232] = 32'h0;  // 32'h6abced54;
    ram_cell[    1233] = 32'h0;  // 32'hb6c16800;
    ram_cell[    1234] = 32'h0;  // 32'h01f2da08;
    ram_cell[    1235] = 32'h0;  // 32'h71cb1cb1;
    ram_cell[    1236] = 32'h0;  // 32'hf2317c7e;
    ram_cell[    1237] = 32'h0;  // 32'h5ecde094;
    ram_cell[    1238] = 32'h0;  // 32'ha443d201;
    ram_cell[    1239] = 32'h0;  // 32'hccf8e21a;
    ram_cell[    1240] = 32'h0;  // 32'ha9d991dc;
    ram_cell[    1241] = 32'h0;  // 32'hee21024b;
    ram_cell[    1242] = 32'h0;  // 32'hf2b53679;
    ram_cell[    1243] = 32'h0;  // 32'hec5050a9;
    ram_cell[    1244] = 32'h0;  // 32'h1d4640f7;
    ram_cell[    1245] = 32'h0;  // 32'h9fb79baf;
    ram_cell[    1246] = 32'h0;  // 32'hb0066449;
    ram_cell[    1247] = 32'h0;  // 32'h28de3050;
    ram_cell[    1248] = 32'h0;  // 32'h697642e3;
    ram_cell[    1249] = 32'h0;  // 32'h29fc2a75;
    ram_cell[    1250] = 32'h0;  // 32'ha9d5a574;
    ram_cell[    1251] = 32'h0;  // 32'h4286d565;
    ram_cell[    1252] = 32'h0;  // 32'hd8fe50ec;
    ram_cell[    1253] = 32'h0;  // 32'h6f6b2981;
    ram_cell[    1254] = 32'h0;  // 32'h452c554f;
    ram_cell[    1255] = 32'h0;  // 32'h1da354ce;
    ram_cell[    1256] = 32'h0;  // 32'h478f69ea;
    ram_cell[    1257] = 32'h0;  // 32'h7910d82c;
    ram_cell[    1258] = 32'h0;  // 32'h22cd4979;
    ram_cell[    1259] = 32'h0;  // 32'h9dc17d79;
    ram_cell[    1260] = 32'h0;  // 32'hda7ddc51;
    ram_cell[    1261] = 32'h0;  // 32'h3ae8b12d;
    ram_cell[    1262] = 32'h0;  // 32'h6dd03019;
    ram_cell[    1263] = 32'h0;  // 32'h5bb4e2a8;
    ram_cell[    1264] = 32'h0;  // 32'hbd1221f5;
    ram_cell[    1265] = 32'h0;  // 32'ha8e134c7;
    ram_cell[    1266] = 32'h0;  // 32'hd3b6610a;
    ram_cell[    1267] = 32'h0;  // 32'h3c6fec71;
    ram_cell[    1268] = 32'h0;  // 32'h3b5850fe;
    ram_cell[    1269] = 32'h0;  // 32'hcc3f3514;
    ram_cell[    1270] = 32'h0;  // 32'hb5e61bee;
    ram_cell[    1271] = 32'h0;  // 32'h5851b3c5;
    ram_cell[    1272] = 32'h0;  // 32'hddd62cce;
    ram_cell[    1273] = 32'h0;  // 32'h6494557c;
    ram_cell[    1274] = 32'h0;  // 32'h1df74335;
    ram_cell[    1275] = 32'h0;  // 32'h3a1bf446;
    ram_cell[    1276] = 32'h0;  // 32'h87f088c0;
    ram_cell[    1277] = 32'h0;  // 32'h54b8e12e;
    ram_cell[    1278] = 32'h0;  // 32'h2098a85e;
    ram_cell[    1279] = 32'h0;  // 32'h52dc1d31;
    ram_cell[    1280] = 32'h0;  // 32'h4c9c2acc;
    ram_cell[    1281] = 32'h0;  // 32'hc5c83414;
    ram_cell[    1282] = 32'h0;  // 32'h5a1108bb;
    ram_cell[    1283] = 32'h0;  // 32'h7345a8af;
    ram_cell[    1284] = 32'h0;  // 32'h984c12fb;
    ram_cell[    1285] = 32'h0;  // 32'hf6a53687;
    ram_cell[    1286] = 32'h0;  // 32'hb36bfb32;
    ram_cell[    1287] = 32'h0;  // 32'hc2d82452;
    ram_cell[    1288] = 32'h0;  // 32'h0447a452;
    ram_cell[    1289] = 32'h0;  // 32'h1fed4b64;
    ram_cell[    1290] = 32'h0;  // 32'h6da357e9;
    ram_cell[    1291] = 32'h0;  // 32'h579efcd2;
    ram_cell[    1292] = 32'h0;  // 32'h2fc992e6;
    ram_cell[    1293] = 32'h0;  // 32'hd83a6f54;
    ram_cell[    1294] = 32'h0;  // 32'h2fa90073;
    ram_cell[    1295] = 32'h0;  // 32'h355a1b55;
    ram_cell[    1296] = 32'h0;  // 32'h2ec8cb0c;
    ram_cell[    1297] = 32'h0;  // 32'h107fa111;
    ram_cell[    1298] = 32'h0;  // 32'h10945c2d;
    ram_cell[    1299] = 32'h0;  // 32'h7ca15e73;
    ram_cell[    1300] = 32'h0;  // 32'h555e37d2;
    ram_cell[    1301] = 32'h0;  // 32'h7f47bf72;
    ram_cell[    1302] = 32'h0;  // 32'h5347c967;
    ram_cell[    1303] = 32'h0;  // 32'hd935d8d3;
    ram_cell[    1304] = 32'h0;  // 32'hd312e747;
    ram_cell[    1305] = 32'h0;  // 32'hf19d96d1;
    ram_cell[    1306] = 32'h0;  // 32'h9ab59f4c;
    ram_cell[    1307] = 32'h0;  // 32'hd512b1c0;
    ram_cell[    1308] = 32'h0;  // 32'h1580c2bd;
    ram_cell[    1309] = 32'h0;  // 32'hb6244005;
    ram_cell[    1310] = 32'h0;  // 32'h2e2c859e;
    ram_cell[    1311] = 32'h0;  // 32'hdee4f8d2;
    ram_cell[    1312] = 32'h0;  // 32'ha4a4937b;
    ram_cell[    1313] = 32'h0;  // 32'h361a24d6;
    ram_cell[    1314] = 32'h0;  // 32'h7b827e07;
    ram_cell[    1315] = 32'h0;  // 32'h4000fc5b;
    ram_cell[    1316] = 32'h0;  // 32'h817f7339;
    ram_cell[    1317] = 32'h0;  // 32'hee71c693;
    ram_cell[    1318] = 32'h0;  // 32'hc65bc351;
    ram_cell[    1319] = 32'h0;  // 32'h249db596;
    ram_cell[    1320] = 32'h0;  // 32'hab378b40;
    ram_cell[    1321] = 32'h0;  // 32'h7eb8fb0e;
    ram_cell[    1322] = 32'h0;  // 32'h071bb679;
    ram_cell[    1323] = 32'h0;  // 32'h2ad671a4;
    ram_cell[    1324] = 32'h0;  // 32'h334594fc;
    ram_cell[    1325] = 32'h0;  // 32'hed91dec8;
    ram_cell[    1326] = 32'h0;  // 32'h3c000777;
    ram_cell[    1327] = 32'h0;  // 32'hd7f056d1;
    ram_cell[    1328] = 32'h0;  // 32'hff13b877;
    ram_cell[    1329] = 32'h0;  // 32'h2e187bbb;
    ram_cell[    1330] = 32'h0;  // 32'h40ef5945;
    ram_cell[    1331] = 32'h0;  // 32'h7b8f2418;
    ram_cell[    1332] = 32'h0;  // 32'h26dd7e2f;
    ram_cell[    1333] = 32'h0;  // 32'h5dfbe8aa;
    ram_cell[    1334] = 32'h0;  // 32'h232dc6ed;
    ram_cell[    1335] = 32'h0;  // 32'h429dbd5f;
    ram_cell[    1336] = 32'h0;  // 32'h3c9609b0;
    ram_cell[    1337] = 32'h0;  // 32'h3b5f236b;
    ram_cell[    1338] = 32'h0;  // 32'hfb71ab39;
    ram_cell[    1339] = 32'h0;  // 32'h4cc0fbb1;
    ram_cell[    1340] = 32'h0;  // 32'h9d433790;
    ram_cell[    1341] = 32'h0;  // 32'hcf9e047a;
    ram_cell[    1342] = 32'h0;  // 32'h856155a6;
    ram_cell[    1343] = 32'h0;  // 32'h1e02f5da;
    ram_cell[    1344] = 32'h0;  // 32'hbf5e360e;
    ram_cell[    1345] = 32'h0;  // 32'ha69771fc;
    ram_cell[    1346] = 32'h0;  // 32'hddf160ae;
    ram_cell[    1347] = 32'h0;  // 32'h05d33847;
    ram_cell[    1348] = 32'h0;  // 32'h3169f780;
    ram_cell[    1349] = 32'h0;  // 32'hb18ef269;
    ram_cell[    1350] = 32'h0;  // 32'hc7debc1a;
    ram_cell[    1351] = 32'h0;  // 32'h169ccb21;
    ram_cell[    1352] = 32'h0;  // 32'h4f8f9822;
    ram_cell[    1353] = 32'h0;  // 32'h4c87b0f4;
    ram_cell[    1354] = 32'h0;  // 32'h3740f26a;
    ram_cell[    1355] = 32'h0;  // 32'h252db84e;
    ram_cell[    1356] = 32'h0;  // 32'h7c966e00;
    ram_cell[    1357] = 32'h0;  // 32'ha5d6ce21;
    ram_cell[    1358] = 32'h0;  // 32'h4b4c3420;
    ram_cell[    1359] = 32'h0;  // 32'hff78d392;
    ram_cell[    1360] = 32'h0;  // 32'h7bd88560;
    ram_cell[    1361] = 32'h0;  // 32'h40f8b8d2;
    ram_cell[    1362] = 32'h0;  // 32'habc57002;
    ram_cell[    1363] = 32'h0;  // 32'h852afe45;
    ram_cell[    1364] = 32'h0;  // 32'hf8cdd255;
    ram_cell[    1365] = 32'h0;  // 32'hf9d2a945;
    ram_cell[    1366] = 32'h0;  // 32'h7b03c945;
    ram_cell[    1367] = 32'h0;  // 32'h8a142895;
    ram_cell[    1368] = 32'h0;  // 32'he7ff6630;
    ram_cell[    1369] = 32'h0;  // 32'hfe9af07b;
    ram_cell[    1370] = 32'h0;  // 32'h9ab13b4c;
    ram_cell[    1371] = 32'h0;  // 32'hf7aceda3;
    ram_cell[    1372] = 32'h0;  // 32'hc3432389;
    ram_cell[    1373] = 32'h0;  // 32'h83efd20c;
    ram_cell[    1374] = 32'h0;  // 32'h1233f082;
    ram_cell[    1375] = 32'h0;  // 32'hf2b4928d;
    ram_cell[    1376] = 32'h0;  // 32'h1c72b17c;
    ram_cell[    1377] = 32'h0;  // 32'h6ed7d98f;
    ram_cell[    1378] = 32'h0;  // 32'h4fa3952e;
    ram_cell[    1379] = 32'h0;  // 32'hfe4f536c;
    ram_cell[    1380] = 32'h0;  // 32'hff23b18f;
    ram_cell[    1381] = 32'h0;  // 32'he5fcc862;
    ram_cell[    1382] = 32'h0;  // 32'he79c510e;
    ram_cell[    1383] = 32'h0;  // 32'he7501778;
    ram_cell[    1384] = 32'h0;  // 32'h8276beae;
    ram_cell[    1385] = 32'h0;  // 32'h2adc0bef;
    ram_cell[    1386] = 32'h0;  // 32'hcc25ac3e;
    ram_cell[    1387] = 32'h0;  // 32'h26d31f53;
    ram_cell[    1388] = 32'h0;  // 32'h4842f48d;
    ram_cell[    1389] = 32'h0;  // 32'haaeebb99;
    ram_cell[    1390] = 32'h0;  // 32'haf8b1c30;
    ram_cell[    1391] = 32'h0;  // 32'h83bb5aaa;
    ram_cell[    1392] = 32'h0;  // 32'hbaafc29e;
    ram_cell[    1393] = 32'h0;  // 32'h7b4e2c24;
    ram_cell[    1394] = 32'h0;  // 32'h0155ce32;
    ram_cell[    1395] = 32'h0;  // 32'h9559b564;
    ram_cell[    1396] = 32'h0;  // 32'h57e9ed12;
    ram_cell[    1397] = 32'h0;  // 32'h7460be66;
    ram_cell[    1398] = 32'h0;  // 32'h245d04d3;
    ram_cell[    1399] = 32'h0;  // 32'h5c605a71;
    ram_cell[    1400] = 32'h0;  // 32'h4b51f70c;
    ram_cell[    1401] = 32'h0;  // 32'h097f0c21;
    ram_cell[    1402] = 32'h0;  // 32'h8cde46ea;
    ram_cell[    1403] = 32'h0;  // 32'h91c5a08b;
    ram_cell[    1404] = 32'h0;  // 32'h452842fd;
    ram_cell[    1405] = 32'h0;  // 32'h23ec963e;
    ram_cell[    1406] = 32'h0;  // 32'h57d612f8;
    ram_cell[    1407] = 32'h0;  // 32'h7c841bed;
    ram_cell[    1408] = 32'h0;  // 32'h91c57515;
    ram_cell[    1409] = 32'h0;  // 32'h9010e178;
    ram_cell[    1410] = 32'h0;  // 32'hdd5552cc;
    ram_cell[    1411] = 32'h0;  // 32'h1ac8c4d5;
    ram_cell[    1412] = 32'h0;  // 32'h1bf002ce;
    ram_cell[    1413] = 32'h0;  // 32'h6a697c33;
    ram_cell[    1414] = 32'h0;  // 32'h3c7d7f6b;
    ram_cell[    1415] = 32'h0;  // 32'hb227fc38;
    ram_cell[    1416] = 32'h0;  // 32'h8ed21b30;
    ram_cell[    1417] = 32'h0;  // 32'h077efb2d;
    ram_cell[    1418] = 32'h0;  // 32'h2920559f;
    ram_cell[    1419] = 32'h0;  // 32'hbbd583e1;
    ram_cell[    1420] = 32'h0;  // 32'h16923482;
    ram_cell[    1421] = 32'h0;  // 32'h81e7fd7e;
    ram_cell[    1422] = 32'h0;  // 32'h1bb9bf50;
    ram_cell[    1423] = 32'h0;  // 32'h1e93eb47;
    ram_cell[    1424] = 32'h0;  // 32'h4bfafe1d;
    ram_cell[    1425] = 32'h0;  // 32'hf64d3837;
    ram_cell[    1426] = 32'h0;  // 32'h26f70a02;
    ram_cell[    1427] = 32'h0;  // 32'h207e22f7;
    ram_cell[    1428] = 32'h0;  // 32'h7a58fdf2;
    ram_cell[    1429] = 32'h0;  // 32'h5d50eef5;
    ram_cell[    1430] = 32'h0;  // 32'had8f9a7e;
    ram_cell[    1431] = 32'h0;  // 32'he958d4dc;
    ram_cell[    1432] = 32'h0;  // 32'h31d89026;
    ram_cell[    1433] = 32'h0;  // 32'h0d9eddf6;
    ram_cell[    1434] = 32'h0;  // 32'h40f03091;
    ram_cell[    1435] = 32'h0;  // 32'h348d4eed;
    ram_cell[    1436] = 32'h0;  // 32'h44cd9eed;
    ram_cell[    1437] = 32'h0;  // 32'h5d01ddad;
    ram_cell[    1438] = 32'h0;  // 32'h6d0c580b;
    ram_cell[    1439] = 32'h0;  // 32'h8e4a7cb9;
    ram_cell[    1440] = 32'h0;  // 32'h42e99623;
    ram_cell[    1441] = 32'h0;  // 32'h729b491e;
    ram_cell[    1442] = 32'h0;  // 32'h4608981d;
    ram_cell[    1443] = 32'h0;  // 32'he023ea80;
    ram_cell[    1444] = 32'h0;  // 32'h642baf8f;
    ram_cell[    1445] = 32'h0;  // 32'h76acb5da;
    ram_cell[    1446] = 32'h0;  // 32'h91dd7f84;
    ram_cell[    1447] = 32'h0;  // 32'h49469d90;
    ram_cell[    1448] = 32'h0;  // 32'h20c4d448;
    ram_cell[    1449] = 32'h0;  // 32'h0c3e2ae1;
    ram_cell[    1450] = 32'h0;  // 32'he14efb2f;
    ram_cell[    1451] = 32'h0;  // 32'h34cb3a20;
    ram_cell[    1452] = 32'h0;  // 32'hc74d5216;
    ram_cell[    1453] = 32'h0;  // 32'he6208cfb;
    ram_cell[    1454] = 32'h0;  // 32'hc3503560;
    ram_cell[    1455] = 32'h0;  // 32'h63324c9f;
    ram_cell[    1456] = 32'h0;  // 32'h4441e38c;
    ram_cell[    1457] = 32'h0;  // 32'ha416b061;
    ram_cell[    1458] = 32'h0;  // 32'h15501c2c;
    ram_cell[    1459] = 32'h0;  // 32'h8797a505;
    ram_cell[    1460] = 32'h0;  // 32'h6f09772b;
    ram_cell[    1461] = 32'h0;  // 32'hc42eed6b;
    ram_cell[    1462] = 32'h0;  // 32'h62b5354e;
    ram_cell[    1463] = 32'h0;  // 32'h7e56a3de;
    ram_cell[    1464] = 32'h0;  // 32'h0fccd0f4;
    ram_cell[    1465] = 32'h0;  // 32'hda85726f;
    ram_cell[    1466] = 32'h0;  // 32'h9a8ef868;
    ram_cell[    1467] = 32'h0;  // 32'h4f33e75e;
    ram_cell[    1468] = 32'h0;  // 32'hdc6b5c36;
    ram_cell[    1469] = 32'h0;  // 32'h0ae37bff;
    ram_cell[    1470] = 32'h0;  // 32'hb8d3b0b9;
    ram_cell[    1471] = 32'h0;  // 32'h02204c9e;
    ram_cell[    1472] = 32'h0;  // 32'he0a5ed34;
    ram_cell[    1473] = 32'h0;  // 32'h0403222b;
    ram_cell[    1474] = 32'h0;  // 32'ha0bd89d9;
    ram_cell[    1475] = 32'h0;  // 32'h87fba828;
    ram_cell[    1476] = 32'h0;  // 32'hd48f19bf;
    ram_cell[    1477] = 32'h0;  // 32'h3abf457a;
    ram_cell[    1478] = 32'h0;  // 32'hb956b701;
    ram_cell[    1479] = 32'h0;  // 32'hcdd9bd2d;
    ram_cell[    1480] = 32'h0;  // 32'h2d4bd5cb;
    ram_cell[    1481] = 32'h0;  // 32'hf6c02865;
    ram_cell[    1482] = 32'h0;  // 32'h9f829fcf;
    ram_cell[    1483] = 32'h0;  // 32'h4f3c7d7e;
    ram_cell[    1484] = 32'h0;  // 32'hc4c7687f;
    ram_cell[    1485] = 32'h0;  // 32'h75c1cdfa;
    ram_cell[    1486] = 32'h0;  // 32'h22b81897;
    ram_cell[    1487] = 32'h0;  // 32'h4a949f36;
    ram_cell[    1488] = 32'h0;  // 32'hbc32c210;
    ram_cell[    1489] = 32'h0;  // 32'h58d5d57c;
    ram_cell[    1490] = 32'h0;  // 32'h0231e523;
    ram_cell[    1491] = 32'h0;  // 32'ha2b44685;
    ram_cell[    1492] = 32'h0;  // 32'h02e53c2b;
    ram_cell[    1493] = 32'h0;  // 32'ha69d0672;
    ram_cell[    1494] = 32'h0;  // 32'h26c67933;
    ram_cell[    1495] = 32'h0;  // 32'h91581ad2;
    ram_cell[    1496] = 32'h0;  // 32'hdd02d1e4;
    ram_cell[    1497] = 32'h0;  // 32'h62223551;
    ram_cell[    1498] = 32'h0;  // 32'hf77d5ce0;
    ram_cell[    1499] = 32'h0;  // 32'hf5d379ac;
    ram_cell[    1500] = 32'h0;  // 32'h5bffcd2a;
    ram_cell[    1501] = 32'h0;  // 32'h0721bfce;
    ram_cell[    1502] = 32'h0;  // 32'h83ebdf43;
    ram_cell[    1503] = 32'h0;  // 32'h40f47398;
    ram_cell[    1504] = 32'h0;  // 32'h7f311a58;
    ram_cell[    1505] = 32'h0;  // 32'hcc50c10d;
    ram_cell[    1506] = 32'h0;  // 32'ha1feb2e6;
    ram_cell[    1507] = 32'h0;  // 32'hf36357ff;
    ram_cell[    1508] = 32'h0;  // 32'he833eb7e;
    ram_cell[    1509] = 32'h0;  // 32'h8b57fdd8;
    ram_cell[    1510] = 32'h0;  // 32'h090d3925;
    ram_cell[    1511] = 32'h0;  // 32'hcbf16f5e;
    ram_cell[    1512] = 32'h0;  // 32'h1df226ed;
    ram_cell[    1513] = 32'h0;  // 32'ha82b5612;
    ram_cell[    1514] = 32'h0;  // 32'h1662ecc3;
    ram_cell[    1515] = 32'h0;  // 32'h7c1df5aa;
    ram_cell[    1516] = 32'h0;  // 32'hda35ac2c;
    ram_cell[    1517] = 32'h0;  // 32'h1b9171ee;
    ram_cell[    1518] = 32'h0;  // 32'h151da85a;
    ram_cell[    1519] = 32'h0;  // 32'h9aece32b;
    ram_cell[    1520] = 32'h0;  // 32'hc411de0a;
    ram_cell[    1521] = 32'h0;  // 32'hb5459bee;
    ram_cell[    1522] = 32'h0;  // 32'hfd775fac;
    ram_cell[    1523] = 32'h0;  // 32'h25567312;
    ram_cell[    1524] = 32'h0;  // 32'h8246b1b0;
    ram_cell[    1525] = 32'h0;  // 32'h72249794;
    ram_cell[    1526] = 32'h0;  // 32'h0f566947;
    ram_cell[    1527] = 32'h0;  // 32'h36e84fc9;
    ram_cell[    1528] = 32'h0;  // 32'h226799ff;
    ram_cell[    1529] = 32'h0;  // 32'h8eea4175;
    ram_cell[    1530] = 32'h0;  // 32'h87e3eb79;
    ram_cell[    1531] = 32'h0;  // 32'h8ecb1266;
    ram_cell[    1532] = 32'h0;  // 32'h0838f6ec;
    ram_cell[    1533] = 32'h0;  // 32'h7ce02225;
    ram_cell[    1534] = 32'h0;  // 32'h05be337e;
    ram_cell[    1535] = 32'h0;  // 32'h22e140d0;
    ram_cell[    1536] = 32'h0;  // 32'h72561958;
    ram_cell[    1537] = 32'h0;  // 32'h90b3fcf7;
    ram_cell[    1538] = 32'h0;  // 32'h2026d1cc;
    ram_cell[    1539] = 32'h0;  // 32'h6ca8e401;
    ram_cell[    1540] = 32'h0;  // 32'had45b4c0;
    ram_cell[    1541] = 32'h0;  // 32'he0f810f0;
    ram_cell[    1542] = 32'h0;  // 32'h9f310802;
    ram_cell[    1543] = 32'h0;  // 32'h526479c4;
    ram_cell[    1544] = 32'h0;  // 32'h97381437;
    ram_cell[    1545] = 32'h0;  // 32'hba4a56c6;
    ram_cell[    1546] = 32'h0;  // 32'h5a680d40;
    ram_cell[    1547] = 32'h0;  // 32'h074c7bbb;
    ram_cell[    1548] = 32'h0;  // 32'h0d0a94ce;
    ram_cell[    1549] = 32'h0;  // 32'hbe04560d;
    ram_cell[    1550] = 32'h0;  // 32'h49b140cb;
    ram_cell[    1551] = 32'h0;  // 32'h584eb687;
    ram_cell[    1552] = 32'h0;  // 32'h9a8510e4;
    ram_cell[    1553] = 32'h0;  // 32'heb3719b1;
    ram_cell[    1554] = 32'h0;  // 32'h020359d4;
    ram_cell[    1555] = 32'h0;  // 32'h15f766e9;
    ram_cell[    1556] = 32'h0;  // 32'h773505ec;
    ram_cell[    1557] = 32'h0;  // 32'h3a9b927e;
    ram_cell[    1558] = 32'h0;  // 32'h97482710;
    ram_cell[    1559] = 32'h0;  // 32'h40a02ce6;
    ram_cell[    1560] = 32'h0;  // 32'h422e3f0c;
    ram_cell[    1561] = 32'h0;  // 32'h26fa96de;
    ram_cell[    1562] = 32'h0;  // 32'h1570556f;
    ram_cell[    1563] = 32'h0;  // 32'h36d0093b;
    ram_cell[    1564] = 32'h0;  // 32'h97c848c6;
    ram_cell[    1565] = 32'h0;  // 32'h2a15987e;
    ram_cell[    1566] = 32'h0;  // 32'h80512e69;
    ram_cell[    1567] = 32'h0;  // 32'hd9ac7490;
    ram_cell[    1568] = 32'h0;  // 32'h8f782268;
    ram_cell[    1569] = 32'h0;  // 32'h8bcef1be;
    ram_cell[    1570] = 32'h0;  // 32'h359dd991;
    ram_cell[    1571] = 32'h0;  // 32'h7d2d247c;
    ram_cell[    1572] = 32'h0;  // 32'h924d133a;
    ram_cell[    1573] = 32'h0;  // 32'h95d1dd6f;
    ram_cell[    1574] = 32'h0;  // 32'h2531a1ff;
    ram_cell[    1575] = 32'h0;  // 32'h838276f6;
    ram_cell[    1576] = 32'h0;  // 32'h6a7e7f27;
    ram_cell[    1577] = 32'h0;  // 32'h32714ffa;
    ram_cell[    1578] = 32'h0;  // 32'hbab36dae;
    ram_cell[    1579] = 32'h0;  // 32'h9dc1242c;
    ram_cell[    1580] = 32'h0;  // 32'h33a0d6f7;
    ram_cell[    1581] = 32'h0;  // 32'hd21a7a2d;
    ram_cell[    1582] = 32'h0;  // 32'hd8c06010;
    ram_cell[    1583] = 32'h0;  // 32'h0fa772cc;
    ram_cell[    1584] = 32'h0;  // 32'h757a9a91;
    ram_cell[    1585] = 32'h0;  // 32'h24fd88fa;
    ram_cell[    1586] = 32'h0;  // 32'h462a5783;
    ram_cell[    1587] = 32'h0;  // 32'h462d25ac;
    ram_cell[    1588] = 32'h0;  // 32'he6b05168;
    ram_cell[    1589] = 32'h0;  // 32'h00092943;
    ram_cell[    1590] = 32'h0;  // 32'hd181e5af;
    ram_cell[    1591] = 32'h0;  // 32'h3e195061;
    ram_cell[    1592] = 32'h0;  // 32'h3b254adf;
    ram_cell[    1593] = 32'h0;  // 32'h59faedf8;
    ram_cell[    1594] = 32'h0;  // 32'h1aa26e45;
    ram_cell[    1595] = 32'h0;  // 32'h36730fc3;
    ram_cell[    1596] = 32'h0;  // 32'h99791a44;
    ram_cell[    1597] = 32'h0;  // 32'he005692d;
    ram_cell[    1598] = 32'h0;  // 32'hd35e0f0e;
    ram_cell[    1599] = 32'h0;  // 32'h76974c01;
    ram_cell[    1600] = 32'h0;  // 32'h5b23e598;
    ram_cell[    1601] = 32'h0;  // 32'h10219110;
    ram_cell[    1602] = 32'h0;  // 32'h8b8d7283;
    ram_cell[    1603] = 32'h0;  // 32'h2b089631;
    ram_cell[    1604] = 32'h0;  // 32'hdecec111;
    ram_cell[    1605] = 32'h0;  // 32'h8f7b62a9;
    ram_cell[    1606] = 32'h0;  // 32'hba6aa587;
    ram_cell[    1607] = 32'h0;  // 32'h4497ff9a;
    ram_cell[    1608] = 32'h0;  // 32'h63303d8a;
    ram_cell[    1609] = 32'h0;  // 32'he25e3d90;
    ram_cell[    1610] = 32'h0;  // 32'hcbe6e380;
    ram_cell[    1611] = 32'h0;  // 32'hd95a9e90;
    ram_cell[    1612] = 32'h0;  // 32'hafc0818d;
    ram_cell[    1613] = 32'h0;  // 32'hbaa45b19;
    ram_cell[    1614] = 32'h0;  // 32'h12498205;
    ram_cell[    1615] = 32'h0;  // 32'hebefda61;
    ram_cell[    1616] = 32'h0;  // 32'h645dd994;
    ram_cell[    1617] = 32'h0;  // 32'hb303c705;
    ram_cell[    1618] = 32'h0;  // 32'h985df127;
    ram_cell[    1619] = 32'h0;  // 32'h888ea35a;
    ram_cell[    1620] = 32'h0;  // 32'h74f71e65;
    ram_cell[    1621] = 32'h0;  // 32'ha460878f;
    ram_cell[    1622] = 32'h0;  // 32'h2335a883;
    ram_cell[    1623] = 32'h0;  // 32'h80f05bc6;
    ram_cell[    1624] = 32'h0;  // 32'hbf672365;
    ram_cell[    1625] = 32'h0;  // 32'h8cec63c3;
    ram_cell[    1626] = 32'h0;  // 32'h21b13f22;
    ram_cell[    1627] = 32'h0;  // 32'hc3c6d3e0;
    ram_cell[    1628] = 32'h0;  // 32'hccc36315;
    ram_cell[    1629] = 32'h0;  // 32'h065ff6c2;
    ram_cell[    1630] = 32'h0;  // 32'he8ef9ede;
    ram_cell[    1631] = 32'h0;  // 32'ha1fe7b6c;
    ram_cell[    1632] = 32'h0;  // 32'he2456b98;
    ram_cell[    1633] = 32'h0;  // 32'h8c8d6558;
    ram_cell[    1634] = 32'h0;  // 32'h0778b3ea;
    ram_cell[    1635] = 32'h0;  // 32'h2153fb3c;
    ram_cell[    1636] = 32'h0;  // 32'hc9743775;
    ram_cell[    1637] = 32'h0;  // 32'hdf798122;
    ram_cell[    1638] = 32'h0;  // 32'h416af10f;
    ram_cell[    1639] = 32'h0;  // 32'h025f17c5;
    ram_cell[    1640] = 32'h0;  // 32'hf79029e1;
    ram_cell[    1641] = 32'h0;  // 32'h943ba43d;
    ram_cell[    1642] = 32'h0;  // 32'h98b695f1;
    ram_cell[    1643] = 32'h0;  // 32'haac23776;
    ram_cell[    1644] = 32'h0;  // 32'hec83ac52;
    ram_cell[    1645] = 32'h0;  // 32'haf99d15b;
    ram_cell[    1646] = 32'h0;  // 32'hd71df0bc;
    ram_cell[    1647] = 32'h0;  // 32'hb8c81b33;
    ram_cell[    1648] = 32'h0;  // 32'h2d46ff43;
    ram_cell[    1649] = 32'h0;  // 32'ha1c9dbe7;
    ram_cell[    1650] = 32'h0;  // 32'h639d81f5;
    ram_cell[    1651] = 32'h0;  // 32'h0820dcee;
    ram_cell[    1652] = 32'h0;  // 32'h68df2890;
    ram_cell[    1653] = 32'h0;  // 32'ha67c683c;
    ram_cell[    1654] = 32'h0;  // 32'hd00411a7;
    ram_cell[    1655] = 32'h0;  // 32'h7c99cd60;
    ram_cell[    1656] = 32'h0;  // 32'h9093c0cb;
    ram_cell[    1657] = 32'h0;  // 32'haeba69c4;
    ram_cell[    1658] = 32'h0;  // 32'h423168ad;
    ram_cell[    1659] = 32'h0;  // 32'h817d7d62;
    ram_cell[    1660] = 32'h0;  // 32'hda52ebf9;
    ram_cell[    1661] = 32'h0;  // 32'h9b169583;
    ram_cell[    1662] = 32'h0;  // 32'hee0a25f0;
    ram_cell[    1663] = 32'h0;  // 32'hce0b7136;
    ram_cell[    1664] = 32'h0;  // 32'h22a2a5cc;
    ram_cell[    1665] = 32'h0;  // 32'ha291375c;
    ram_cell[    1666] = 32'h0;  // 32'hb1d283cf;
    ram_cell[    1667] = 32'h0;  // 32'hb4826339;
    ram_cell[    1668] = 32'h0;  // 32'h85e25ddc;
    ram_cell[    1669] = 32'h0;  // 32'h30a428eb;
    ram_cell[    1670] = 32'h0;  // 32'hc21ff14a;
    ram_cell[    1671] = 32'h0;  // 32'hf302d51c;
    ram_cell[    1672] = 32'h0;  // 32'h84135e57;
    ram_cell[    1673] = 32'h0;  // 32'h682c5f4a;
    ram_cell[    1674] = 32'h0;  // 32'h44def31a;
    ram_cell[    1675] = 32'h0;  // 32'h402b2183;
    ram_cell[    1676] = 32'h0;  // 32'he13cc092;
    ram_cell[    1677] = 32'h0;  // 32'h94a9831c;
    ram_cell[    1678] = 32'h0;  // 32'hea634532;
    ram_cell[    1679] = 32'h0;  // 32'hf6d66f38;
    ram_cell[    1680] = 32'h0;  // 32'h2fe36084;
    ram_cell[    1681] = 32'h0;  // 32'hb6dbef15;
    ram_cell[    1682] = 32'h0;  // 32'h629bd02d;
    ram_cell[    1683] = 32'h0;  // 32'hcaab8a08;
    ram_cell[    1684] = 32'h0;  // 32'hdfd3a9ba;
    ram_cell[    1685] = 32'h0;  // 32'hb1cbf646;
    ram_cell[    1686] = 32'h0;  // 32'hd7741871;
    ram_cell[    1687] = 32'h0;  // 32'h58e6ef14;
    ram_cell[    1688] = 32'h0;  // 32'hb52f8761;
    ram_cell[    1689] = 32'h0;  // 32'h2bfb8cb2;
    ram_cell[    1690] = 32'h0;  // 32'h285a8982;
    ram_cell[    1691] = 32'h0;  // 32'h3d733f09;
    ram_cell[    1692] = 32'h0;  // 32'ha79c471c;
    ram_cell[    1693] = 32'h0;  // 32'hc645e1b7;
    ram_cell[    1694] = 32'h0;  // 32'h6ca3517d;
    ram_cell[    1695] = 32'h0;  // 32'h0647bc04;
    ram_cell[    1696] = 32'h0;  // 32'h3c1d1684;
    ram_cell[    1697] = 32'h0;  // 32'hd7e831f2;
    ram_cell[    1698] = 32'h0;  // 32'h8d379a02;
    ram_cell[    1699] = 32'h0;  // 32'hc9ee7751;
    ram_cell[    1700] = 32'h0;  // 32'hdd4a6989;
    ram_cell[    1701] = 32'h0;  // 32'hc26382e1;
    ram_cell[    1702] = 32'h0;  // 32'h5d127bcc;
    ram_cell[    1703] = 32'h0;  // 32'hfb783d63;
    ram_cell[    1704] = 32'h0;  // 32'hf572c781;
    ram_cell[    1705] = 32'h0;  // 32'h814bbe38;
    ram_cell[    1706] = 32'h0;  // 32'h55f73d06;
    ram_cell[    1707] = 32'h0;  // 32'h4d88ef96;
    ram_cell[    1708] = 32'h0;  // 32'h6629d57d;
    ram_cell[    1709] = 32'h0;  // 32'h284270d2;
    ram_cell[    1710] = 32'h0;  // 32'h22acb847;
    ram_cell[    1711] = 32'h0;  // 32'hb0ee50be;
    ram_cell[    1712] = 32'h0;  // 32'hb4502372;
    ram_cell[    1713] = 32'h0;  // 32'h36093889;
    ram_cell[    1714] = 32'h0;  // 32'h5adb9c44;
    ram_cell[    1715] = 32'h0;  // 32'hf31709d8;
    ram_cell[    1716] = 32'h0;  // 32'had0d9d52;
    ram_cell[    1717] = 32'h0;  // 32'h471874e7;
    ram_cell[    1718] = 32'h0;  // 32'h29fb238e;
    ram_cell[    1719] = 32'h0;  // 32'ha56cf322;
    ram_cell[    1720] = 32'h0;  // 32'hf8ed5e0a;
    ram_cell[    1721] = 32'h0;  // 32'h96d877b3;
    ram_cell[    1722] = 32'h0;  // 32'h93767d0f;
    ram_cell[    1723] = 32'h0;  // 32'h198edadc;
    ram_cell[    1724] = 32'h0;  // 32'h61980f64;
    ram_cell[    1725] = 32'h0;  // 32'h4b51fb08;
    ram_cell[    1726] = 32'h0;  // 32'h2b16c0fe;
    ram_cell[    1727] = 32'h0;  // 32'h4b1548be;
    ram_cell[    1728] = 32'h0;  // 32'hb42d06dd;
    ram_cell[    1729] = 32'h0;  // 32'hcde72ad3;
    ram_cell[    1730] = 32'h0;  // 32'h3bc579e4;
    ram_cell[    1731] = 32'h0;  // 32'h7992fd71;
    ram_cell[    1732] = 32'h0;  // 32'h69056f60;
    ram_cell[    1733] = 32'h0;  // 32'h59bd53d5;
    ram_cell[    1734] = 32'h0;  // 32'hbf8ad96d;
    ram_cell[    1735] = 32'h0;  // 32'h4d7f022a;
    ram_cell[    1736] = 32'h0;  // 32'h166338be;
    ram_cell[    1737] = 32'h0;  // 32'h24043878;
    ram_cell[    1738] = 32'h0;  // 32'h25a99d07;
    ram_cell[    1739] = 32'h0;  // 32'hbc882eb1;
    ram_cell[    1740] = 32'h0;  // 32'h4c5d7e25;
    ram_cell[    1741] = 32'h0;  // 32'ha9b0fe27;
    ram_cell[    1742] = 32'h0;  // 32'h95bfaa72;
    ram_cell[    1743] = 32'h0;  // 32'h071c9b42;
    ram_cell[    1744] = 32'h0;  // 32'h2a7f2a16;
    ram_cell[    1745] = 32'h0;  // 32'h34a35d91;
    ram_cell[    1746] = 32'h0;  // 32'hd2641649;
    ram_cell[    1747] = 32'h0;  // 32'h33d925d3;
    ram_cell[    1748] = 32'h0;  // 32'h8fe6a7b7;
    ram_cell[    1749] = 32'h0;  // 32'h83f1f442;
    ram_cell[    1750] = 32'h0;  // 32'h79675eb3;
    ram_cell[    1751] = 32'h0;  // 32'h28e2332d;
    ram_cell[    1752] = 32'h0;  // 32'h56e2321d;
    ram_cell[    1753] = 32'h0;  // 32'he9ddbf93;
    ram_cell[    1754] = 32'h0;  // 32'h36f74260;
    ram_cell[    1755] = 32'h0;  // 32'h4b5e9716;
    ram_cell[    1756] = 32'h0;  // 32'h664b3817;
    ram_cell[    1757] = 32'h0;  // 32'hda88a930;
    ram_cell[    1758] = 32'h0;  // 32'h6d362dea;
    ram_cell[    1759] = 32'h0;  // 32'h6a90ac4f;
    ram_cell[    1760] = 32'h0;  // 32'h7ded075e;
    ram_cell[    1761] = 32'h0;  // 32'h354961c3;
    ram_cell[    1762] = 32'h0;  // 32'h63ee9d50;
    ram_cell[    1763] = 32'h0;  // 32'h0522af4f;
    ram_cell[    1764] = 32'h0;  // 32'hb33bc090;
    ram_cell[    1765] = 32'h0;  // 32'h956efbe0;
    ram_cell[    1766] = 32'h0;  // 32'h3d63d6af;
    ram_cell[    1767] = 32'h0;  // 32'ha4fcb540;
    ram_cell[    1768] = 32'h0;  // 32'h86e79b07;
    ram_cell[    1769] = 32'h0;  // 32'h1d5a6401;
    ram_cell[    1770] = 32'h0;  // 32'h9cefcf18;
    ram_cell[    1771] = 32'h0;  // 32'h9e4e6123;
    ram_cell[    1772] = 32'h0;  // 32'h7be0a4d2;
    ram_cell[    1773] = 32'h0;  // 32'h2ceaedca;
    ram_cell[    1774] = 32'h0;  // 32'h7781ab08;
    ram_cell[    1775] = 32'h0;  // 32'hadf2dc17;
    ram_cell[    1776] = 32'h0;  // 32'h333c3971;
    ram_cell[    1777] = 32'h0;  // 32'hd86cf3c5;
    ram_cell[    1778] = 32'h0;  // 32'hef547531;
    ram_cell[    1779] = 32'h0;  // 32'hfd71c65d;
    ram_cell[    1780] = 32'h0;  // 32'haafdeba2;
    ram_cell[    1781] = 32'h0;  // 32'h8fcffeb4;
    ram_cell[    1782] = 32'h0;  // 32'h535b8c07;
    ram_cell[    1783] = 32'h0;  // 32'h64e9d377;
    ram_cell[    1784] = 32'h0;  // 32'h312d732d;
    ram_cell[    1785] = 32'h0;  // 32'hb0bd592a;
    ram_cell[    1786] = 32'h0;  // 32'haa763bef;
    ram_cell[    1787] = 32'h0;  // 32'h6e870c65;
    ram_cell[    1788] = 32'h0;  // 32'h893eecb7;
    ram_cell[    1789] = 32'h0;  // 32'h055d4ff1;
    ram_cell[    1790] = 32'h0;  // 32'h53359e05;
    ram_cell[    1791] = 32'h0;  // 32'habdd1b9c;
    ram_cell[    1792] = 32'h0;  // 32'hd059151b;
    ram_cell[    1793] = 32'h0;  // 32'hedb26b3f;
    ram_cell[    1794] = 32'h0;  // 32'hd7e5ea45;
    ram_cell[    1795] = 32'h0;  // 32'h90558814;
    ram_cell[    1796] = 32'h0;  // 32'h2fab1803;
    ram_cell[    1797] = 32'h0;  // 32'h05a7f0fb;
    ram_cell[    1798] = 32'h0;  // 32'h53da006b;
    ram_cell[    1799] = 32'h0;  // 32'h11d3260f;
    ram_cell[    1800] = 32'h0;  // 32'ha49c5b0a;
    ram_cell[    1801] = 32'h0;  // 32'h8d9d3177;
    ram_cell[    1802] = 32'h0;  // 32'h53aa8cfb;
    ram_cell[    1803] = 32'h0;  // 32'h21b771f3;
    ram_cell[    1804] = 32'h0;  // 32'h0d0d7c40;
    ram_cell[    1805] = 32'h0;  // 32'h6ef76eda;
    ram_cell[    1806] = 32'h0;  // 32'h3e3b103b;
    ram_cell[    1807] = 32'h0;  // 32'h3e600465;
    ram_cell[    1808] = 32'h0;  // 32'h7a3a161d;
    ram_cell[    1809] = 32'h0;  // 32'hbaa13814;
    ram_cell[    1810] = 32'h0;  // 32'h9e05c79c;
    ram_cell[    1811] = 32'h0;  // 32'h12cf7d39;
    ram_cell[    1812] = 32'h0;  // 32'h2546aff2;
    ram_cell[    1813] = 32'h0;  // 32'h23555ae8;
    ram_cell[    1814] = 32'h0;  // 32'h5f6ee0bc;
    ram_cell[    1815] = 32'h0;  // 32'h0f153d4b;
    ram_cell[    1816] = 32'h0;  // 32'h2109b3d2;
    ram_cell[    1817] = 32'h0;  // 32'h51d160f4;
    ram_cell[    1818] = 32'h0;  // 32'h07e69168;
    ram_cell[    1819] = 32'h0;  // 32'hed52bdea;
    ram_cell[    1820] = 32'h0;  // 32'h60ab4681;
    ram_cell[    1821] = 32'h0;  // 32'h08a5e69f;
    ram_cell[    1822] = 32'h0;  // 32'h58c404e7;
    ram_cell[    1823] = 32'h0;  // 32'h9fc7c87d;
    ram_cell[    1824] = 32'h0;  // 32'hf88f4edc;
    ram_cell[    1825] = 32'h0;  // 32'h7b3bbd49;
    ram_cell[    1826] = 32'h0;  // 32'h963a6981;
    ram_cell[    1827] = 32'h0;  // 32'h27a19427;
    ram_cell[    1828] = 32'h0;  // 32'he812f01f;
    ram_cell[    1829] = 32'h0;  // 32'h97a51335;
    ram_cell[    1830] = 32'h0;  // 32'h29100aba;
    ram_cell[    1831] = 32'h0;  // 32'hb48e2c4a;
    ram_cell[    1832] = 32'h0;  // 32'h77e23952;
    ram_cell[    1833] = 32'h0;  // 32'h5593d4c1;
    ram_cell[    1834] = 32'h0;  // 32'h66701678;
    ram_cell[    1835] = 32'h0;  // 32'hb729ab10;
    ram_cell[    1836] = 32'h0;  // 32'ha8869bd0;
    ram_cell[    1837] = 32'h0;  // 32'hc9b920c1;
    ram_cell[    1838] = 32'h0;  // 32'h2b6ab906;
    ram_cell[    1839] = 32'h0;  // 32'h5104ca41;
    ram_cell[    1840] = 32'h0;  // 32'hccd5f335;
    ram_cell[    1841] = 32'h0;  // 32'h693961d6;
    ram_cell[    1842] = 32'h0;  // 32'h720ae9b6;
    ram_cell[    1843] = 32'h0;  // 32'h49858505;
    ram_cell[    1844] = 32'h0;  // 32'h2aea8aed;
    ram_cell[    1845] = 32'h0;  // 32'h356210f6;
    ram_cell[    1846] = 32'h0;  // 32'h148f1252;
    ram_cell[    1847] = 32'h0;  // 32'h5244866c;
    ram_cell[    1848] = 32'h0;  // 32'h7c7934f6;
    ram_cell[    1849] = 32'h0;  // 32'hc55e77ea;
    ram_cell[    1850] = 32'h0;  // 32'h17a0d0bf;
    ram_cell[    1851] = 32'h0;  // 32'h2e8c058a;
    ram_cell[    1852] = 32'h0;  // 32'h6b4f52f4;
    ram_cell[    1853] = 32'h0;  // 32'h28a54156;
    ram_cell[    1854] = 32'h0;  // 32'ha1e69131;
    ram_cell[    1855] = 32'h0;  // 32'h3e3e11c0;
    ram_cell[    1856] = 32'h0;  // 32'h4eeeab58;
    ram_cell[    1857] = 32'h0;  // 32'h28ad3c2a;
    ram_cell[    1858] = 32'h0;  // 32'hcb30e5ca;
    ram_cell[    1859] = 32'h0;  // 32'h59d53913;
    ram_cell[    1860] = 32'h0;  // 32'hc3f71ef1;
    ram_cell[    1861] = 32'h0;  // 32'h660d44e8;
    ram_cell[    1862] = 32'h0;  // 32'h584bd25e;
    ram_cell[    1863] = 32'h0;  // 32'ha95d0415;
    ram_cell[    1864] = 32'h0;  // 32'hf5855381;
    ram_cell[    1865] = 32'h0;  // 32'h5d390832;
    ram_cell[    1866] = 32'h0;  // 32'h32b66e63;
    ram_cell[    1867] = 32'h0;  // 32'hc997d92d;
    ram_cell[    1868] = 32'h0;  // 32'h142ce4b3;
    ram_cell[    1869] = 32'h0;  // 32'h6e0051c8;
    ram_cell[    1870] = 32'h0;  // 32'he22f9eeb;
    ram_cell[    1871] = 32'h0;  // 32'h36aa0a1b;
    ram_cell[    1872] = 32'h0;  // 32'h65d7a54a;
    ram_cell[    1873] = 32'h0;  // 32'ha0c4caf6;
    ram_cell[    1874] = 32'h0;  // 32'hf0fd1a8a;
    ram_cell[    1875] = 32'h0;  // 32'hef335191;
    ram_cell[    1876] = 32'h0;  // 32'hb4159e65;
    ram_cell[    1877] = 32'h0;  // 32'h7c852cb1;
    ram_cell[    1878] = 32'h0;  // 32'h28106444;
    ram_cell[    1879] = 32'h0;  // 32'hdb5b6881;
    ram_cell[    1880] = 32'h0;  // 32'h461ff9bf;
    ram_cell[    1881] = 32'h0;  // 32'h3feb01ea;
    ram_cell[    1882] = 32'h0;  // 32'h44cd97ea;
    ram_cell[    1883] = 32'h0;  // 32'h631f43f6;
    ram_cell[    1884] = 32'h0;  // 32'h38cde948;
    ram_cell[    1885] = 32'h0;  // 32'h4e9ab97a;
    ram_cell[    1886] = 32'h0;  // 32'h86a204be;
    ram_cell[    1887] = 32'h0;  // 32'h9fd4f56a;
    ram_cell[    1888] = 32'h0;  // 32'h488da0d7;
    ram_cell[    1889] = 32'h0;  // 32'hc65d6669;
    ram_cell[    1890] = 32'h0;  // 32'h52bd1eac;
    ram_cell[    1891] = 32'h0;  // 32'h518ae018;
    ram_cell[    1892] = 32'h0;  // 32'h0af39838;
    ram_cell[    1893] = 32'h0;  // 32'hac14f6d4;
    ram_cell[    1894] = 32'h0;  // 32'h3ad0261a;
    ram_cell[    1895] = 32'h0;  // 32'hca82e066;
    ram_cell[    1896] = 32'h0;  // 32'ha6654700;
    ram_cell[    1897] = 32'h0;  // 32'h71c2415a;
    ram_cell[    1898] = 32'h0;  // 32'he86f3a58;
    ram_cell[    1899] = 32'h0;  // 32'he824fabe;
    ram_cell[    1900] = 32'h0;  // 32'h31b11d5a;
    ram_cell[    1901] = 32'h0;  // 32'h46f7b5ca;
    ram_cell[    1902] = 32'h0;  // 32'h0bc86472;
    ram_cell[    1903] = 32'h0;  // 32'h4f7df0c8;
    ram_cell[    1904] = 32'h0;  // 32'h38113c4e;
    ram_cell[    1905] = 32'h0;  // 32'h6c4ea5d6;
    ram_cell[    1906] = 32'h0;  // 32'hb5431116;
    ram_cell[    1907] = 32'h0;  // 32'h6eb9cc3a;
    ram_cell[    1908] = 32'h0;  // 32'h78f18ae3;
    ram_cell[    1909] = 32'h0;  // 32'hf7d42762;
    ram_cell[    1910] = 32'h0;  // 32'hb2cbb991;
    ram_cell[    1911] = 32'h0;  // 32'h3ca56a4a;
    ram_cell[    1912] = 32'h0;  // 32'h39d6df4e;
    ram_cell[    1913] = 32'h0;  // 32'h56899a62;
    ram_cell[    1914] = 32'h0;  // 32'h3d831c56;
    ram_cell[    1915] = 32'h0;  // 32'h5cf8de19;
    ram_cell[    1916] = 32'h0;  // 32'h4e38b06c;
    ram_cell[    1917] = 32'h0;  // 32'h7a6360b4;
    ram_cell[    1918] = 32'h0;  // 32'h1f6d7132;
    ram_cell[    1919] = 32'h0;  // 32'hf9c871fc;
    ram_cell[    1920] = 32'h0;  // 32'h4ab02aaf;
    ram_cell[    1921] = 32'h0;  // 32'h1cf24e1b;
    ram_cell[    1922] = 32'h0;  // 32'hbf072e36;
    ram_cell[    1923] = 32'h0;  // 32'h5aef77f7;
    ram_cell[    1924] = 32'h0;  // 32'h658be380;
    ram_cell[    1925] = 32'h0;  // 32'h96627b69;
    ram_cell[    1926] = 32'h0;  // 32'he88f8381;
    ram_cell[    1927] = 32'h0;  // 32'h735c759f;
    ram_cell[    1928] = 32'h0;  // 32'h3394a8c2;
    ram_cell[    1929] = 32'h0;  // 32'hd8cc1c8a;
    ram_cell[    1930] = 32'h0;  // 32'h603dcf59;
    ram_cell[    1931] = 32'h0;  // 32'h8b21c1e6;
    ram_cell[    1932] = 32'h0;  // 32'h8fdb97cb;
    ram_cell[    1933] = 32'h0;  // 32'h7bd73303;
    ram_cell[    1934] = 32'h0;  // 32'h4078c3dc;
    ram_cell[    1935] = 32'h0;  // 32'h893125df;
    ram_cell[    1936] = 32'h0;  // 32'h6d13b053;
    ram_cell[    1937] = 32'h0;  // 32'hf8b07be2;
    ram_cell[    1938] = 32'h0;  // 32'h1c734cfa;
    ram_cell[    1939] = 32'h0;  // 32'he7506f4c;
    ram_cell[    1940] = 32'h0;  // 32'hcbd54faf;
    ram_cell[    1941] = 32'h0;  // 32'h61dd0ad8;
    ram_cell[    1942] = 32'h0;  // 32'he284e7da;
    ram_cell[    1943] = 32'h0;  // 32'h245eb719;
    ram_cell[    1944] = 32'h0;  // 32'h61e8ef36;
    ram_cell[    1945] = 32'h0;  // 32'h1985f4ef;
    ram_cell[    1946] = 32'h0;  // 32'h3b047956;
    ram_cell[    1947] = 32'h0;  // 32'h12f9513f;
    ram_cell[    1948] = 32'h0;  // 32'h610c113b;
    ram_cell[    1949] = 32'h0;  // 32'he7654d83;
    ram_cell[    1950] = 32'h0;  // 32'ha53fc188;
    ram_cell[    1951] = 32'h0;  // 32'ha044826c;
    ram_cell[    1952] = 32'h0;  // 32'he23f91e2;
    ram_cell[    1953] = 32'h0;  // 32'hd4052b81;
    ram_cell[    1954] = 32'h0;  // 32'hebeef22c;
    ram_cell[    1955] = 32'h0;  // 32'hca116a99;
    ram_cell[    1956] = 32'h0;  // 32'hdf05e9a6;
    ram_cell[    1957] = 32'h0;  // 32'ha18eb86a;
    ram_cell[    1958] = 32'h0;  // 32'h4c7dafd0;
    ram_cell[    1959] = 32'h0;  // 32'h26ed1c27;
    ram_cell[    1960] = 32'h0;  // 32'h552deb9f;
    ram_cell[    1961] = 32'h0;  // 32'h007c089b;
    ram_cell[    1962] = 32'h0;  // 32'hb2b30e67;
    ram_cell[    1963] = 32'h0;  // 32'h08c7f730;
    ram_cell[    1964] = 32'h0;  // 32'hcf5c5ca8;
    ram_cell[    1965] = 32'h0;  // 32'hd20d9721;
    ram_cell[    1966] = 32'h0;  // 32'hef6a1d51;
    ram_cell[    1967] = 32'h0;  // 32'he460ccbd;
    ram_cell[    1968] = 32'h0;  // 32'h3095c3ef;
    ram_cell[    1969] = 32'h0;  // 32'h2b8f88a9;
    ram_cell[    1970] = 32'h0;  // 32'h8df6181e;
    ram_cell[    1971] = 32'h0;  // 32'hda08e6b1;
    ram_cell[    1972] = 32'h0;  // 32'hbee241a3;
    ram_cell[    1973] = 32'h0;  // 32'ha63ecacb;
    ram_cell[    1974] = 32'h0;  // 32'hf5c8bb5d;
    ram_cell[    1975] = 32'h0;  // 32'hdaf550ca;
    ram_cell[    1976] = 32'h0;  // 32'h84776256;
    ram_cell[    1977] = 32'h0;  // 32'h391c0cd8;
    ram_cell[    1978] = 32'h0;  // 32'h89a8b35e;
    ram_cell[    1979] = 32'h0;  // 32'h698fab8f;
    ram_cell[    1980] = 32'h0;  // 32'h242a49ae;
    ram_cell[    1981] = 32'h0;  // 32'haab95d6f;
    ram_cell[    1982] = 32'h0;  // 32'ha8f20c89;
    ram_cell[    1983] = 32'h0;  // 32'h7174e462;
    ram_cell[    1984] = 32'h0;  // 32'haf64bdfc;
    ram_cell[    1985] = 32'h0;  // 32'h4d544d21;
    ram_cell[    1986] = 32'h0;  // 32'h05747f2f;
    ram_cell[    1987] = 32'h0;  // 32'h138b1408;
    ram_cell[    1988] = 32'h0;  // 32'h7fedfd25;
    ram_cell[    1989] = 32'h0;  // 32'h48757906;
    ram_cell[    1990] = 32'h0;  // 32'hd852d110;
    ram_cell[    1991] = 32'h0;  // 32'hf8475c52;
    ram_cell[    1992] = 32'h0;  // 32'h6a59706f;
    ram_cell[    1993] = 32'h0;  // 32'ha661fcdc;
    ram_cell[    1994] = 32'h0;  // 32'h755b0c91;
    ram_cell[    1995] = 32'h0;  // 32'he6720c8a;
    ram_cell[    1996] = 32'h0;  // 32'h3d9f5943;
    ram_cell[    1997] = 32'h0;  // 32'h26416642;
    ram_cell[    1998] = 32'h0;  // 32'ha08663ba;
    ram_cell[    1999] = 32'h0;  // 32'h0129dba0;
    ram_cell[    2000] = 32'h0;  // 32'h30df9c09;
    ram_cell[    2001] = 32'h0;  // 32'h576af07b;
    ram_cell[    2002] = 32'h0;  // 32'h93062b80;
    ram_cell[    2003] = 32'h0;  // 32'h3d1d1f75;
    ram_cell[    2004] = 32'h0;  // 32'h5507587c;
    ram_cell[    2005] = 32'h0;  // 32'hf744e149;
    ram_cell[    2006] = 32'h0;  // 32'h336e02a9;
    ram_cell[    2007] = 32'h0;  // 32'h96f93998;
    ram_cell[    2008] = 32'h0;  // 32'he60914ae;
    ram_cell[    2009] = 32'h0;  // 32'h232b1484;
    ram_cell[    2010] = 32'h0;  // 32'h97077d90;
    ram_cell[    2011] = 32'h0;  // 32'hcae2e9f5;
    ram_cell[    2012] = 32'h0;  // 32'h4aa70119;
    ram_cell[    2013] = 32'h0;  // 32'h2ad04d8c;
    ram_cell[    2014] = 32'h0;  // 32'h6ad5059d;
    ram_cell[    2015] = 32'h0;  // 32'h4d637bfb;
    ram_cell[    2016] = 32'h0;  // 32'hcb4dd87c;
    ram_cell[    2017] = 32'h0;  // 32'hf723f3a2;
    ram_cell[    2018] = 32'h0;  // 32'h152c5f7f;
    ram_cell[    2019] = 32'h0;  // 32'h805e7c45;
    ram_cell[    2020] = 32'h0;  // 32'h37bd1ed8;
    ram_cell[    2021] = 32'h0;  // 32'hd360e935;
    ram_cell[    2022] = 32'h0;  // 32'h0675bffe;
    ram_cell[    2023] = 32'h0;  // 32'h80778280;
    ram_cell[    2024] = 32'h0;  // 32'h43535a08;
    ram_cell[    2025] = 32'h0;  // 32'h75ac5619;
    ram_cell[    2026] = 32'h0;  // 32'ha4bdec11;
    ram_cell[    2027] = 32'h0;  // 32'he99ce9ed;
    ram_cell[    2028] = 32'h0;  // 32'h3ad0be88;
    ram_cell[    2029] = 32'h0;  // 32'hae660d4f;
    ram_cell[    2030] = 32'h0;  // 32'hcc8783b1;
    ram_cell[    2031] = 32'h0;  // 32'h0d089ef4;
    ram_cell[    2032] = 32'h0;  // 32'hadf1e591;
    ram_cell[    2033] = 32'h0;  // 32'h99e5f5f6;
    ram_cell[    2034] = 32'h0;  // 32'h03d685eb;
    ram_cell[    2035] = 32'h0;  // 32'h3fa74318;
    ram_cell[    2036] = 32'h0;  // 32'h37924906;
    ram_cell[    2037] = 32'h0;  // 32'hdc1d548f;
    ram_cell[    2038] = 32'h0;  // 32'h0365fadf;
    ram_cell[    2039] = 32'h0;  // 32'hfed31001;
    ram_cell[    2040] = 32'h0;  // 32'h2a3f9bd4;
    ram_cell[    2041] = 32'h0;  // 32'hf78843f7;
    ram_cell[    2042] = 32'h0;  // 32'hd9c9b81b;
    ram_cell[    2043] = 32'h0;  // 32'h772e4dd0;
    ram_cell[    2044] = 32'h0;  // 32'h318dcc9d;
    ram_cell[    2045] = 32'h0;  // 32'h9e5d3dff;
    ram_cell[    2046] = 32'h0;  // 32'h2af6fbae;
    ram_cell[    2047] = 32'h0;  // 32'h268ff1ea;
    ram_cell[    2048] = 32'h0;  // 32'h65d20e56;
    ram_cell[    2049] = 32'h0;  // 32'hc7f34bd6;
    ram_cell[    2050] = 32'h0;  // 32'h20b350af;
    ram_cell[    2051] = 32'h0;  // 32'h2bb7ccb1;
    ram_cell[    2052] = 32'h0;  // 32'hca5dddbc;
    ram_cell[    2053] = 32'h0;  // 32'ha581adc2;
    ram_cell[    2054] = 32'h0;  // 32'h5d419eea;
    ram_cell[    2055] = 32'h0;  // 32'hf6d4570d;
    ram_cell[    2056] = 32'h0;  // 32'h9b508fec;
    ram_cell[    2057] = 32'h0;  // 32'hcf5d14a1;
    ram_cell[    2058] = 32'h0;  // 32'hb3c1e7bf;
    ram_cell[    2059] = 32'h0;  // 32'hf0bdedf3;
    ram_cell[    2060] = 32'h0;  // 32'h6bac317a;
    ram_cell[    2061] = 32'h0;  // 32'h270e61ed;
    ram_cell[    2062] = 32'h0;  // 32'h2c08fb08;
    ram_cell[    2063] = 32'h0;  // 32'h9060e1a5;
    ram_cell[    2064] = 32'h0;  // 32'h55fd8f06;
    ram_cell[    2065] = 32'h0;  // 32'h233ebf2c;
    ram_cell[    2066] = 32'h0;  // 32'h63a97ccf;
    ram_cell[    2067] = 32'h0;  // 32'h7ea9f58d;
    ram_cell[    2068] = 32'h0;  // 32'h17303c03;
    ram_cell[    2069] = 32'h0;  // 32'hf639147f;
    ram_cell[    2070] = 32'h0;  // 32'h43957edb;
    ram_cell[    2071] = 32'h0;  // 32'h5f47a41a;
    ram_cell[    2072] = 32'h0;  // 32'hec319ebd;
    ram_cell[    2073] = 32'h0;  // 32'h06a47855;
    ram_cell[    2074] = 32'h0;  // 32'ha34b7090;
    ram_cell[    2075] = 32'h0;  // 32'hd2477da4;
    ram_cell[    2076] = 32'h0;  // 32'hdc0e01da;
    ram_cell[    2077] = 32'h0;  // 32'h973832e2;
    ram_cell[    2078] = 32'h0;  // 32'he6f7c508;
    ram_cell[    2079] = 32'h0;  // 32'hd979e666;
    ram_cell[    2080] = 32'h0;  // 32'h453a0250;
    ram_cell[    2081] = 32'h0;  // 32'h97ce8c1b;
    ram_cell[    2082] = 32'h0;  // 32'hbda367e5;
    ram_cell[    2083] = 32'h0;  // 32'hda7d14bf;
    ram_cell[    2084] = 32'h0;  // 32'he2f7bc3a;
    ram_cell[    2085] = 32'h0;  // 32'h67ef62f1;
    ram_cell[    2086] = 32'h0;  // 32'h71c51d82;
    ram_cell[    2087] = 32'h0;  // 32'he57d41b2;
    ram_cell[    2088] = 32'h0;  // 32'hd06411f0;
    ram_cell[    2089] = 32'h0;  // 32'h084cd489;
    ram_cell[    2090] = 32'h0;  // 32'h18465a69;
    ram_cell[    2091] = 32'h0;  // 32'h5d10f57a;
    ram_cell[    2092] = 32'h0;  // 32'h4e350d55;
    ram_cell[    2093] = 32'h0;  // 32'hb20d6076;
    ram_cell[    2094] = 32'h0;  // 32'h20ad4c62;
    ram_cell[    2095] = 32'h0;  // 32'h1c406bb3;
    ram_cell[    2096] = 32'h0;  // 32'h6c318074;
    ram_cell[    2097] = 32'h0;  // 32'h8cfa152a;
    ram_cell[    2098] = 32'h0;  // 32'ha897bcb4;
    ram_cell[    2099] = 32'h0;  // 32'h2e40025e;
    ram_cell[    2100] = 32'h0;  // 32'hc42e20ee;
    ram_cell[    2101] = 32'h0;  // 32'h2c2fce26;
    ram_cell[    2102] = 32'h0;  // 32'h5bd800ac;
    ram_cell[    2103] = 32'h0;  // 32'h4526c463;
    ram_cell[    2104] = 32'h0;  // 32'h502c574a;
    ram_cell[    2105] = 32'h0;  // 32'h3f618b8b;
    ram_cell[    2106] = 32'h0;  // 32'h17e76277;
    ram_cell[    2107] = 32'h0;  // 32'h4fd2ec83;
    ram_cell[    2108] = 32'h0;  // 32'h5672dd57;
    ram_cell[    2109] = 32'h0;  // 32'h99866479;
    ram_cell[    2110] = 32'h0;  // 32'h834d90b7;
    ram_cell[    2111] = 32'h0;  // 32'h10bbd6b5;
    ram_cell[    2112] = 32'h0;  // 32'h114086d5;
    ram_cell[    2113] = 32'h0;  // 32'h993f483e;
    ram_cell[    2114] = 32'h0;  // 32'h3bb43eb2;
    ram_cell[    2115] = 32'h0;  // 32'h93adff2f;
    ram_cell[    2116] = 32'h0;  // 32'ha337d9c7;
    ram_cell[    2117] = 32'h0;  // 32'h8164ef78;
    ram_cell[    2118] = 32'h0;  // 32'h51fe5dc8;
    ram_cell[    2119] = 32'h0;  // 32'h1c248498;
    ram_cell[    2120] = 32'h0;  // 32'h65d3ee6f;
    ram_cell[    2121] = 32'h0;  // 32'h6e4535ff;
    ram_cell[    2122] = 32'h0;  // 32'he9eb05dc;
    ram_cell[    2123] = 32'h0;  // 32'h6ef80ede;
    ram_cell[    2124] = 32'h0;  // 32'h27f90bce;
    ram_cell[    2125] = 32'h0;  // 32'h1ab35437;
    ram_cell[    2126] = 32'h0;  // 32'hc58a8588;
    ram_cell[    2127] = 32'h0;  // 32'h17b7e52d;
    ram_cell[    2128] = 32'h0;  // 32'hfcd14170;
    ram_cell[    2129] = 32'h0;  // 32'he46e1bb0;
    ram_cell[    2130] = 32'h0;  // 32'h61987b47;
    ram_cell[    2131] = 32'h0;  // 32'hbdf12d2e;
    ram_cell[    2132] = 32'h0;  // 32'h36a59990;
    ram_cell[    2133] = 32'h0;  // 32'h72f8bdf1;
    ram_cell[    2134] = 32'h0;  // 32'h0859bdd1;
    ram_cell[    2135] = 32'h0;  // 32'hc7f86758;
    ram_cell[    2136] = 32'h0;  // 32'hea4423ef;
    ram_cell[    2137] = 32'h0;  // 32'hd4b96f1a;
    ram_cell[    2138] = 32'h0;  // 32'h4fecdacf;
    ram_cell[    2139] = 32'h0;  // 32'h15a392c0;
    ram_cell[    2140] = 32'h0;  // 32'ha028fd92;
    ram_cell[    2141] = 32'h0;  // 32'h96749d86;
    ram_cell[    2142] = 32'h0;  // 32'he9053e32;
    ram_cell[    2143] = 32'h0;  // 32'h8942cd3b;
    ram_cell[    2144] = 32'h0;  // 32'hebd89fcb;
    ram_cell[    2145] = 32'h0;  // 32'h5325f862;
    ram_cell[    2146] = 32'h0;  // 32'hb97fcbb5;
    ram_cell[    2147] = 32'h0;  // 32'h2e0e99a0;
    ram_cell[    2148] = 32'h0;  // 32'ha259148e;
    ram_cell[    2149] = 32'h0;  // 32'h2e2a63ba;
    ram_cell[    2150] = 32'h0;  // 32'h811a8a17;
    ram_cell[    2151] = 32'h0;  // 32'hafe84807;
    ram_cell[    2152] = 32'h0;  // 32'h99a19399;
    ram_cell[    2153] = 32'h0;  // 32'h536bf003;
    ram_cell[    2154] = 32'h0;  // 32'hbddf116e;
    ram_cell[    2155] = 32'h0;  // 32'h335c84e7;
    ram_cell[    2156] = 32'h0;  // 32'h436e7988;
    ram_cell[    2157] = 32'h0;  // 32'h598d8e22;
    ram_cell[    2158] = 32'h0;  // 32'hd07e91bd;
    ram_cell[    2159] = 32'h0;  // 32'h7768129c;
    ram_cell[    2160] = 32'h0;  // 32'hd528d6a7;
    ram_cell[    2161] = 32'h0;  // 32'hccfd630d;
    ram_cell[    2162] = 32'h0;  // 32'h79f88bc4;
    ram_cell[    2163] = 32'h0;  // 32'h1e1a7bb8;
    ram_cell[    2164] = 32'h0;  // 32'h9fdd1d23;
    ram_cell[    2165] = 32'h0;  // 32'h115f229d;
    ram_cell[    2166] = 32'h0;  // 32'h7ce13e0b;
    ram_cell[    2167] = 32'h0;  // 32'haf8ab5f1;
    ram_cell[    2168] = 32'h0;  // 32'heeb07886;
    ram_cell[    2169] = 32'h0;  // 32'hdb504303;
    ram_cell[    2170] = 32'h0;  // 32'h8fab83ce;
    ram_cell[    2171] = 32'h0;  // 32'h171d88a0;
    ram_cell[    2172] = 32'h0;  // 32'h6c1327b2;
    ram_cell[    2173] = 32'h0;  // 32'h87b3fff6;
    ram_cell[    2174] = 32'h0;  // 32'h82b076b9;
    ram_cell[    2175] = 32'h0;  // 32'h18f9e591;
    ram_cell[    2176] = 32'h0;  // 32'h92a3990d;
    ram_cell[    2177] = 32'h0;  // 32'h11931c4d;
    ram_cell[    2178] = 32'h0;  // 32'h394dfb7e;
    ram_cell[    2179] = 32'h0;  // 32'hb68a1428;
    ram_cell[    2180] = 32'h0;  // 32'h7a7e719b;
    ram_cell[    2181] = 32'h0;  // 32'h3cf7b873;
    ram_cell[    2182] = 32'h0;  // 32'hda5c7fc9;
    ram_cell[    2183] = 32'h0;  // 32'h2c3f886a;
    ram_cell[    2184] = 32'h0;  // 32'hdf30ce8c;
    ram_cell[    2185] = 32'h0;  // 32'hd813e2ff;
    ram_cell[    2186] = 32'h0;  // 32'h16cf502e;
    ram_cell[    2187] = 32'h0;  // 32'h1f6090a4;
    ram_cell[    2188] = 32'h0;  // 32'h482ae693;
    ram_cell[    2189] = 32'h0;  // 32'hafc8ae35;
    ram_cell[    2190] = 32'h0;  // 32'h27a1d777;
    ram_cell[    2191] = 32'h0;  // 32'h10af1811;
    ram_cell[    2192] = 32'h0;  // 32'h88a4c2c5;
    ram_cell[    2193] = 32'h0;  // 32'h50289cc6;
    ram_cell[    2194] = 32'h0;  // 32'h96c8a22f;
    ram_cell[    2195] = 32'h0;  // 32'hbe15316e;
    ram_cell[    2196] = 32'h0;  // 32'hd02dacc3;
    ram_cell[    2197] = 32'h0;  // 32'hc0dc70a6;
    ram_cell[    2198] = 32'h0;  // 32'hbce63c2e;
    ram_cell[    2199] = 32'h0;  // 32'h049662da;
    ram_cell[    2200] = 32'h0;  // 32'hbd73bc04;
    ram_cell[    2201] = 32'h0;  // 32'h28856a9d;
    ram_cell[    2202] = 32'h0;  // 32'hd87f15a0;
    ram_cell[    2203] = 32'h0;  // 32'h37e7e8c9;
    ram_cell[    2204] = 32'h0;  // 32'h0e34d74c;
    ram_cell[    2205] = 32'h0;  // 32'h23745087;
    ram_cell[    2206] = 32'h0;  // 32'h1c5bcf59;
    ram_cell[    2207] = 32'h0;  // 32'he3f0c379;
    ram_cell[    2208] = 32'h0;  // 32'hc66c795b;
    ram_cell[    2209] = 32'h0;  // 32'ha6388ab6;
    ram_cell[    2210] = 32'h0;  // 32'h57ededde;
    ram_cell[    2211] = 32'h0;  // 32'hd5619c99;
    ram_cell[    2212] = 32'h0;  // 32'h009b1fce;
    ram_cell[    2213] = 32'h0;  // 32'h2a3f4683;
    ram_cell[    2214] = 32'h0;  // 32'hbaf414d5;
    ram_cell[    2215] = 32'h0;  // 32'haf6e0ac7;
    ram_cell[    2216] = 32'h0;  // 32'h128e25d9;
    ram_cell[    2217] = 32'h0;  // 32'hbcf0ff6e;
    ram_cell[    2218] = 32'h0;  // 32'h2a3fb802;
    ram_cell[    2219] = 32'h0;  // 32'h6b07a7d9;
    ram_cell[    2220] = 32'h0;  // 32'hba038630;
    ram_cell[    2221] = 32'h0;  // 32'h7da1fdcf;
    ram_cell[    2222] = 32'h0;  // 32'h3a9ed689;
    ram_cell[    2223] = 32'h0;  // 32'h9df7aeee;
    ram_cell[    2224] = 32'h0;  // 32'h93331c22;
    ram_cell[    2225] = 32'h0;  // 32'hcbb7a36c;
    ram_cell[    2226] = 32'h0;  // 32'h55cf94e9;
    ram_cell[    2227] = 32'h0;  // 32'ha97d9666;
    ram_cell[    2228] = 32'h0;  // 32'hb59bef6a;
    ram_cell[    2229] = 32'h0;  // 32'hc680a4f3;
    ram_cell[    2230] = 32'h0;  // 32'h3de56835;
    ram_cell[    2231] = 32'h0;  // 32'h22b3f13b;
    ram_cell[    2232] = 32'h0;  // 32'h7ec4984a;
    ram_cell[    2233] = 32'h0;  // 32'h3c49a6a1;
    ram_cell[    2234] = 32'h0;  // 32'h09d5a130;
    ram_cell[    2235] = 32'h0;  // 32'hd3ca908a;
    ram_cell[    2236] = 32'h0;  // 32'h9d7f5a31;
    ram_cell[    2237] = 32'h0;  // 32'hccc3f027;
    ram_cell[    2238] = 32'h0;  // 32'hc58418c5;
    ram_cell[    2239] = 32'h0;  // 32'hcb7c14dd;
    ram_cell[    2240] = 32'h0;  // 32'h5ed371c2;
    ram_cell[    2241] = 32'h0;  // 32'h43c346b8;
    ram_cell[    2242] = 32'h0;  // 32'hadad4c81;
    ram_cell[    2243] = 32'h0;  // 32'h4e599be7;
    ram_cell[    2244] = 32'h0;  // 32'hd432e078;
    ram_cell[    2245] = 32'h0;  // 32'h9a36d816;
    ram_cell[    2246] = 32'h0;  // 32'hec4c394b;
    ram_cell[    2247] = 32'h0;  // 32'hfaba1cdf;
    ram_cell[    2248] = 32'h0;  // 32'h79105e53;
    ram_cell[    2249] = 32'h0;  // 32'h5e3953a7;
    ram_cell[    2250] = 32'h0;  // 32'ha6df47e7;
    ram_cell[    2251] = 32'h0;  // 32'hab436a96;
    ram_cell[    2252] = 32'h0;  // 32'hd1f318ee;
    ram_cell[    2253] = 32'h0;  // 32'h219cb5e0;
    ram_cell[    2254] = 32'h0;  // 32'hc864bc8c;
    ram_cell[    2255] = 32'h0;  // 32'hed543b39;
    ram_cell[    2256] = 32'h0;  // 32'h8cbe1333;
    ram_cell[    2257] = 32'h0;  // 32'h0d306f3c;
    ram_cell[    2258] = 32'h0;  // 32'h489af48c;
    ram_cell[    2259] = 32'h0;  // 32'h398506f4;
    ram_cell[    2260] = 32'h0;  // 32'h8256aceb;
    ram_cell[    2261] = 32'h0;  // 32'h78fde63f;
    ram_cell[    2262] = 32'h0;  // 32'ha2330a08;
    ram_cell[    2263] = 32'h0;  // 32'h45d0f071;
    ram_cell[    2264] = 32'h0;  // 32'hc916944f;
    ram_cell[    2265] = 32'h0;  // 32'h97a4c100;
    ram_cell[    2266] = 32'h0;  // 32'h375e789b;
    ram_cell[    2267] = 32'h0;  // 32'he2f4080c;
    ram_cell[    2268] = 32'h0;  // 32'h5b8f1a56;
    ram_cell[    2269] = 32'h0;  // 32'hcf8cfe75;
    ram_cell[    2270] = 32'h0;  // 32'h7ec8b1be;
    ram_cell[    2271] = 32'h0;  // 32'h020f6ee8;
    ram_cell[    2272] = 32'h0;  // 32'hc5fcdc93;
    ram_cell[    2273] = 32'h0;  // 32'h0077a02b;
    ram_cell[    2274] = 32'h0;  // 32'h53ec55b5;
    ram_cell[    2275] = 32'h0;  // 32'h06c532ac;
    ram_cell[    2276] = 32'h0;  // 32'hfb16d2c7;
    ram_cell[    2277] = 32'h0;  // 32'h5c8e15d5;
    ram_cell[    2278] = 32'h0;  // 32'h25635b83;
    ram_cell[    2279] = 32'h0;  // 32'h48f48d47;
    ram_cell[    2280] = 32'h0;  // 32'hca231305;
    ram_cell[    2281] = 32'h0;  // 32'h06120290;
    ram_cell[    2282] = 32'h0;  // 32'h2c838e13;
    ram_cell[    2283] = 32'h0;  // 32'h78e06a3f;
    ram_cell[    2284] = 32'h0;  // 32'h85aed490;
    ram_cell[    2285] = 32'h0;  // 32'h698da53b;
    ram_cell[    2286] = 32'h0;  // 32'h62cdfe0f;
    ram_cell[    2287] = 32'h0;  // 32'h8ad87ac2;
    ram_cell[    2288] = 32'h0;  // 32'h7ccc10f9;
    ram_cell[    2289] = 32'h0;  // 32'h06f8f7c4;
    ram_cell[    2290] = 32'h0;  // 32'hf2beaa0a;
    ram_cell[    2291] = 32'h0;  // 32'hfbcaa99e;
    ram_cell[    2292] = 32'h0;  // 32'hb090b2c4;
    ram_cell[    2293] = 32'h0;  // 32'h459703b6;
    ram_cell[    2294] = 32'h0;  // 32'hd7cb27fb;
    ram_cell[    2295] = 32'h0;  // 32'h9983ba32;
    ram_cell[    2296] = 32'h0;  // 32'hb775c749;
    ram_cell[    2297] = 32'h0;  // 32'h8562ebd2;
    ram_cell[    2298] = 32'h0;  // 32'h0e0d43a7;
    ram_cell[    2299] = 32'h0;  // 32'h56e93a63;
    ram_cell[    2300] = 32'h0;  // 32'h0cdb9fbb;
    ram_cell[    2301] = 32'h0;  // 32'ha03791c4;
    ram_cell[    2302] = 32'h0;  // 32'ha2796ea7;
    ram_cell[    2303] = 32'h0;  // 32'h1a994add;
    ram_cell[    2304] = 32'h0;  // 32'h53a6abaf;
    ram_cell[    2305] = 32'h0;  // 32'hc5736bf3;
    ram_cell[    2306] = 32'h0;  // 32'h33c687a0;
    ram_cell[    2307] = 32'h0;  // 32'hba680cd5;
    ram_cell[    2308] = 32'h0;  // 32'h6b521a84;
    ram_cell[    2309] = 32'h0;  // 32'h2ca3a540;
    ram_cell[    2310] = 32'h0;  // 32'h0d94babb;
    ram_cell[    2311] = 32'h0;  // 32'hdc5b8e70;
    ram_cell[    2312] = 32'h0;  // 32'h879119bc;
    ram_cell[    2313] = 32'h0;  // 32'h78f89cc9;
    ram_cell[    2314] = 32'h0;  // 32'h2cdb9693;
    ram_cell[    2315] = 32'h0;  // 32'h9642574d;
    ram_cell[    2316] = 32'h0;  // 32'h87901122;
    ram_cell[    2317] = 32'h0;  // 32'h29a8cdf1;
    ram_cell[    2318] = 32'h0;  // 32'h6e1236e9;
    ram_cell[    2319] = 32'h0;  // 32'h18d717c9;
    ram_cell[    2320] = 32'h0;  // 32'hd1d5a026;
    ram_cell[    2321] = 32'h0;  // 32'hba713437;
    ram_cell[    2322] = 32'h0;  // 32'h94d9e3bc;
    ram_cell[    2323] = 32'h0;  // 32'h31450d83;
    ram_cell[    2324] = 32'h0;  // 32'he8ffd47e;
    ram_cell[    2325] = 32'h0;  // 32'hd1f1e4ae;
    ram_cell[    2326] = 32'h0;  // 32'h66e856ea;
    ram_cell[    2327] = 32'h0;  // 32'hf8a738ff;
    ram_cell[    2328] = 32'h0;  // 32'h4c97fe6d;
    ram_cell[    2329] = 32'h0;  // 32'haa113cc3;
    ram_cell[    2330] = 32'h0;  // 32'h153f734c;
    ram_cell[    2331] = 32'h0;  // 32'h38b05c78;
    ram_cell[    2332] = 32'h0;  // 32'h32ab660b;
    ram_cell[    2333] = 32'h0;  // 32'hb776625c;
    ram_cell[    2334] = 32'h0;  // 32'h8b1361ab;
    ram_cell[    2335] = 32'h0;  // 32'hbf399b93;
    ram_cell[    2336] = 32'h0;  // 32'hc538ddaa;
    ram_cell[    2337] = 32'h0;  // 32'hec72ddf1;
    ram_cell[    2338] = 32'h0;  // 32'hfdee0f17;
    ram_cell[    2339] = 32'h0;  // 32'h892bcc46;
    ram_cell[    2340] = 32'h0;  // 32'h3e0014bd;
    ram_cell[    2341] = 32'h0;  // 32'ha95227c7;
    ram_cell[    2342] = 32'h0;  // 32'h278f8ef4;
    ram_cell[    2343] = 32'h0;  // 32'h315cb6f8;
    ram_cell[    2344] = 32'h0;  // 32'h44e186ab;
    ram_cell[    2345] = 32'h0;  // 32'hcc832d64;
    ram_cell[    2346] = 32'h0;  // 32'haae79bc6;
    ram_cell[    2347] = 32'h0;  // 32'h75c175b0;
    ram_cell[    2348] = 32'h0;  // 32'h03e45ac2;
    ram_cell[    2349] = 32'h0;  // 32'h74417f16;
    ram_cell[    2350] = 32'h0;  // 32'h41df1b44;
    ram_cell[    2351] = 32'h0;  // 32'ha02ef34f;
    ram_cell[    2352] = 32'h0;  // 32'hd12a1d15;
    ram_cell[    2353] = 32'h0;  // 32'hbf6e0eac;
    ram_cell[    2354] = 32'h0;  // 32'hcedb0d60;
    ram_cell[    2355] = 32'h0;  // 32'h0c11b9ab;
    ram_cell[    2356] = 32'h0;  // 32'hedfbdf0b;
    ram_cell[    2357] = 32'h0;  // 32'h3737a555;
    ram_cell[    2358] = 32'h0;  // 32'h6246a0d9;
    ram_cell[    2359] = 32'h0;  // 32'h4d96737a;
    ram_cell[    2360] = 32'h0;  // 32'h6696dd15;
    ram_cell[    2361] = 32'h0;  // 32'h18c1a9a7;
    ram_cell[    2362] = 32'h0;  // 32'h0287e01d;
    ram_cell[    2363] = 32'h0;  // 32'h95b5ff97;
    ram_cell[    2364] = 32'h0;  // 32'hcbd715d5;
    ram_cell[    2365] = 32'h0;  // 32'h9242da37;
    ram_cell[    2366] = 32'h0;  // 32'he88993c9;
    ram_cell[    2367] = 32'h0;  // 32'hec07fab5;
    ram_cell[    2368] = 32'h0;  // 32'h27ce3604;
    ram_cell[    2369] = 32'h0;  // 32'hf5f679c5;
    ram_cell[    2370] = 32'h0;  // 32'hc7f4ee95;
    ram_cell[    2371] = 32'h0;  // 32'h0b890d7f;
    ram_cell[    2372] = 32'h0;  // 32'h3e277cb1;
    ram_cell[    2373] = 32'h0;  // 32'hb8aac4dc;
    ram_cell[    2374] = 32'h0;  // 32'h76227d37;
    ram_cell[    2375] = 32'h0;  // 32'h4d3e7127;
    ram_cell[    2376] = 32'h0;  // 32'h1e574682;
    ram_cell[    2377] = 32'h0;  // 32'hdae004a4;
    ram_cell[    2378] = 32'h0;  // 32'h8584abf8;
    ram_cell[    2379] = 32'h0;  // 32'h378a7bbb;
    ram_cell[    2380] = 32'h0;  // 32'h696f8f1d;
    ram_cell[    2381] = 32'h0;  // 32'h4562b9ed;
    ram_cell[    2382] = 32'h0;  // 32'he86ba293;
    ram_cell[    2383] = 32'h0;  // 32'hffe4af82;
    ram_cell[    2384] = 32'h0;  // 32'h8df603f7;
    ram_cell[    2385] = 32'h0;  // 32'h57b764b7;
    ram_cell[    2386] = 32'h0;  // 32'hcaa22ab1;
    ram_cell[    2387] = 32'h0;  // 32'h2c1b0a0a;
    ram_cell[    2388] = 32'h0;  // 32'h9a007e9f;
    ram_cell[    2389] = 32'h0;  // 32'h54e57d5b;
    ram_cell[    2390] = 32'h0;  // 32'h4a01b707;
    ram_cell[    2391] = 32'h0;  // 32'ha436c37b;
    ram_cell[    2392] = 32'h0;  // 32'h1d4ed4af;
    ram_cell[    2393] = 32'h0;  // 32'h41241c2f;
    ram_cell[    2394] = 32'h0;  // 32'h2908f3d1;
    ram_cell[    2395] = 32'h0;  // 32'h6e437445;
    ram_cell[    2396] = 32'h0;  // 32'h0a6c28aa;
    ram_cell[    2397] = 32'h0;  // 32'h1bdb7117;
    ram_cell[    2398] = 32'h0;  // 32'h80edc493;
    ram_cell[    2399] = 32'h0;  // 32'h4b112722;
    ram_cell[    2400] = 32'h0;  // 32'h9a32a9ee;
    ram_cell[    2401] = 32'h0;  // 32'h2dc22059;
    ram_cell[    2402] = 32'h0;  // 32'h8af959b4;
    ram_cell[    2403] = 32'h0;  // 32'h4d9a1c22;
    ram_cell[    2404] = 32'h0;  // 32'h7f3e04ae;
    ram_cell[    2405] = 32'h0;  // 32'h7201d350;
    ram_cell[    2406] = 32'h0;  // 32'h1d53068b;
    ram_cell[    2407] = 32'h0;  // 32'hb9748988;
    ram_cell[    2408] = 32'h0;  // 32'h0262616f;
    ram_cell[    2409] = 32'h0;  // 32'he91039f7;
    ram_cell[    2410] = 32'h0;  // 32'h8ba99f14;
    ram_cell[    2411] = 32'h0;  // 32'h242971eb;
    ram_cell[    2412] = 32'h0;  // 32'h40a883fb;
    ram_cell[    2413] = 32'h0;  // 32'h3aff0bbc;
    ram_cell[    2414] = 32'h0;  // 32'hc09532ab;
    ram_cell[    2415] = 32'h0;  // 32'hdbdb2e26;
    ram_cell[    2416] = 32'h0;  // 32'hce33e262;
    ram_cell[    2417] = 32'h0;  // 32'hd0b37ea0;
    ram_cell[    2418] = 32'h0;  // 32'ha9b45875;
    ram_cell[    2419] = 32'h0;  // 32'hc8b555ab;
    ram_cell[    2420] = 32'h0;  // 32'hfafec4db;
    ram_cell[    2421] = 32'h0;  // 32'h1012489d;
    ram_cell[    2422] = 32'h0;  // 32'he5c75d7a;
    ram_cell[    2423] = 32'h0;  // 32'h608313fe;
    ram_cell[    2424] = 32'h0;  // 32'h73cb26d5;
    ram_cell[    2425] = 32'h0;  // 32'h9cb64106;
    ram_cell[    2426] = 32'h0;  // 32'hb0e6d734;
    ram_cell[    2427] = 32'h0;  // 32'he15b410c;
    ram_cell[    2428] = 32'h0;  // 32'h5bda8634;
    ram_cell[    2429] = 32'h0;  // 32'he0d808c9;
    ram_cell[    2430] = 32'h0;  // 32'heb994385;
    ram_cell[    2431] = 32'h0;  // 32'hf8713e29;
    ram_cell[    2432] = 32'h0;  // 32'h2e4b5350;
    ram_cell[    2433] = 32'h0;  // 32'hf1c37671;
    ram_cell[    2434] = 32'h0;  // 32'hb22e1254;
    ram_cell[    2435] = 32'h0;  // 32'h0f15a6e5;
    ram_cell[    2436] = 32'h0;  // 32'h2cd7b579;
    ram_cell[    2437] = 32'h0;  // 32'h6400c14a;
    ram_cell[    2438] = 32'h0;  // 32'h485d2b66;
    ram_cell[    2439] = 32'h0;  // 32'h571e81be;
    ram_cell[    2440] = 32'h0;  // 32'he9e1631e;
    ram_cell[    2441] = 32'h0;  // 32'h13ec5d05;
    ram_cell[    2442] = 32'h0;  // 32'heb10e286;
    ram_cell[    2443] = 32'h0;  // 32'h004f60f8;
    ram_cell[    2444] = 32'h0;  // 32'hec989702;
    ram_cell[    2445] = 32'h0;  // 32'h15a61440;
    ram_cell[    2446] = 32'h0;  // 32'h5fd53781;
    ram_cell[    2447] = 32'h0;  // 32'h52a04267;
    ram_cell[    2448] = 32'h0;  // 32'h7cb5811b;
    ram_cell[    2449] = 32'h0;  // 32'h7d41a39b;
    ram_cell[    2450] = 32'h0;  // 32'h55d5367e;
    ram_cell[    2451] = 32'h0;  // 32'h2ebd6faf;
    ram_cell[    2452] = 32'h0;  // 32'h79f7c225;
    ram_cell[    2453] = 32'h0;  // 32'h69abca53;
    ram_cell[    2454] = 32'h0;  // 32'h82784c8e;
    ram_cell[    2455] = 32'h0;  // 32'hff49eedb;
    ram_cell[    2456] = 32'h0;  // 32'hd6d9aaed;
    ram_cell[    2457] = 32'h0;  // 32'h1f963f0e;
    ram_cell[    2458] = 32'h0;  // 32'ha91b5f1e;
    ram_cell[    2459] = 32'h0;  // 32'h2cee8013;
    ram_cell[    2460] = 32'h0;  // 32'hcfc6cc43;
    ram_cell[    2461] = 32'h0;  // 32'h5954c3af;
    ram_cell[    2462] = 32'h0;  // 32'h41c8a860;
    ram_cell[    2463] = 32'h0;  // 32'ha053b5c4;
    ram_cell[    2464] = 32'h0;  // 32'h388dcd36;
    ram_cell[    2465] = 32'h0;  // 32'h764c0081;
    ram_cell[    2466] = 32'h0;  // 32'h706e1f48;
    ram_cell[    2467] = 32'h0;  // 32'h9d72d07c;
    ram_cell[    2468] = 32'h0;  // 32'h68b9588e;
    ram_cell[    2469] = 32'h0;  // 32'hfadfb4f2;
    ram_cell[    2470] = 32'h0;  // 32'h78346a13;
    ram_cell[    2471] = 32'h0;  // 32'hf002593f;
    ram_cell[    2472] = 32'h0;  // 32'h2a6d5b43;
    ram_cell[    2473] = 32'h0;  // 32'h3825d0f3;
    ram_cell[    2474] = 32'h0;  // 32'ha501bd5b;
    ram_cell[    2475] = 32'h0;  // 32'h8a1ea4fa;
    ram_cell[    2476] = 32'h0;  // 32'h0b29724d;
    ram_cell[    2477] = 32'h0;  // 32'h3f136474;
    ram_cell[    2478] = 32'h0;  // 32'h8ba0be2c;
    ram_cell[    2479] = 32'h0;  // 32'h73f7954f;
    ram_cell[    2480] = 32'h0;  // 32'h7d3c9eea;
    ram_cell[    2481] = 32'h0;  // 32'h3157104a;
    ram_cell[    2482] = 32'h0;  // 32'h4d433dc8;
    ram_cell[    2483] = 32'h0;  // 32'ha3843c4a;
    ram_cell[    2484] = 32'h0;  // 32'h81181321;
    ram_cell[    2485] = 32'h0;  // 32'h4a852bb1;
    ram_cell[    2486] = 32'h0;  // 32'h0ef7ead5;
    ram_cell[    2487] = 32'h0;  // 32'h5765b993;
    ram_cell[    2488] = 32'h0;  // 32'h7775cd89;
    ram_cell[    2489] = 32'h0;  // 32'hf333f8bb;
    ram_cell[    2490] = 32'h0;  // 32'hf6068799;
    ram_cell[    2491] = 32'h0;  // 32'h330b0dbf;
    ram_cell[    2492] = 32'h0;  // 32'he045e100;
    ram_cell[    2493] = 32'h0;  // 32'h3ff372bb;
    ram_cell[    2494] = 32'h0;  // 32'h0ac7d21f;
    ram_cell[    2495] = 32'h0;  // 32'hceae1c8a;
    ram_cell[    2496] = 32'h0;  // 32'h9f76c465;
    ram_cell[    2497] = 32'h0;  // 32'hdd9368e4;
    ram_cell[    2498] = 32'h0;  // 32'h8b04d3e2;
    ram_cell[    2499] = 32'h0;  // 32'hd33cf93d;
    ram_cell[    2500] = 32'h0;  // 32'h0caca5f8;
    ram_cell[    2501] = 32'h0;  // 32'ha5a0ccdf;
    ram_cell[    2502] = 32'h0;  // 32'hae1642ed;
    ram_cell[    2503] = 32'h0;  // 32'hbe33bc6a;
    ram_cell[    2504] = 32'h0;  // 32'hd8d07d86;
    ram_cell[    2505] = 32'h0;  // 32'h52fd8b8b;
    ram_cell[    2506] = 32'h0;  // 32'h4031c4f3;
    ram_cell[    2507] = 32'h0;  // 32'h64c5e0d7;
    ram_cell[    2508] = 32'h0;  // 32'h8034ee26;
    ram_cell[    2509] = 32'h0;  // 32'h3fffa628;
    ram_cell[    2510] = 32'h0;  // 32'h6d17da7b;
    ram_cell[    2511] = 32'h0;  // 32'hd7c9a866;
    ram_cell[    2512] = 32'h0;  // 32'h83066cc9;
    ram_cell[    2513] = 32'h0;  // 32'h2ee56038;
    ram_cell[    2514] = 32'h0;  // 32'haf04485b;
    ram_cell[    2515] = 32'h0;  // 32'ha45898b4;
    ram_cell[    2516] = 32'h0;  // 32'h816ed133;
    ram_cell[    2517] = 32'h0;  // 32'h69fb4eab;
    ram_cell[    2518] = 32'h0;  // 32'h9ffec63b;
    ram_cell[    2519] = 32'h0;  // 32'he20d8b98;
    ram_cell[    2520] = 32'h0;  // 32'h8c1aca86;
    ram_cell[    2521] = 32'h0;  // 32'h669a9500;
    ram_cell[    2522] = 32'h0;  // 32'hdfc38b0c;
    ram_cell[    2523] = 32'h0;  // 32'h862ac2f1;
    ram_cell[    2524] = 32'h0;  // 32'h8fdd61a6;
    ram_cell[    2525] = 32'h0;  // 32'h53e148fc;
    ram_cell[    2526] = 32'h0;  // 32'he0ec465a;
    ram_cell[    2527] = 32'h0;  // 32'he67c8070;
    ram_cell[    2528] = 32'h0;  // 32'h84a0455e;
    ram_cell[    2529] = 32'h0;  // 32'hdab4dcc6;
    ram_cell[    2530] = 32'h0;  // 32'h6a56adf8;
    ram_cell[    2531] = 32'h0;  // 32'h17a07045;
    ram_cell[    2532] = 32'h0;  // 32'hce2625f1;
    ram_cell[    2533] = 32'h0;  // 32'hd7f193f2;
    ram_cell[    2534] = 32'h0;  // 32'h414dc064;
    ram_cell[    2535] = 32'h0;  // 32'h79764edb;
    ram_cell[    2536] = 32'h0;  // 32'h040fc545;
    ram_cell[    2537] = 32'h0;  // 32'h787e56dd;
    ram_cell[    2538] = 32'h0;  // 32'h61391907;
    ram_cell[    2539] = 32'h0;  // 32'hb18988c8;
    ram_cell[    2540] = 32'h0;  // 32'hdde8ca26;
    ram_cell[    2541] = 32'h0;  // 32'h661e9cbc;
    ram_cell[    2542] = 32'h0;  // 32'hb1cac3ac;
    ram_cell[    2543] = 32'h0;  // 32'h4a4b4f11;
    ram_cell[    2544] = 32'h0;  // 32'h237f333f;
    ram_cell[    2545] = 32'h0;  // 32'h561c3e5b;
    ram_cell[    2546] = 32'h0;  // 32'hd66b9b48;
    ram_cell[    2547] = 32'h0;  // 32'h97b8cb72;
    ram_cell[    2548] = 32'h0;  // 32'hc3d5f55c;
    ram_cell[    2549] = 32'h0;  // 32'h5485365d;
    ram_cell[    2550] = 32'h0;  // 32'he416a6ed;
    ram_cell[    2551] = 32'h0;  // 32'hbde6a053;
    ram_cell[    2552] = 32'h0;  // 32'ha11a7ac6;
    ram_cell[    2553] = 32'h0;  // 32'h7a55bc7d;
    ram_cell[    2554] = 32'h0;  // 32'h30fb95ef;
    ram_cell[    2555] = 32'h0;  // 32'hf6ef4195;
    ram_cell[    2556] = 32'h0;  // 32'h34aec710;
    ram_cell[    2557] = 32'h0;  // 32'hb2045c98;
    ram_cell[    2558] = 32'h0;  // 32'h2c4be3e3;
    ram_cell[    2559] = 32'h0;  // 32'h6951c2f2;
    ram_cell[    2560] = 32'h0;  // 32'h629ee994;
    ram_cell[    2561] = 32'h0;  // 32'hddfd5f21;
    ram_cell[    2562] = 32'h0;  // 32'hed3691d4;
    ram_cell[    2563] = 32'h0;  // 32'hade53da4;
    ram_cell[    2564] = 32'h0;  // 32'h4b610f94;
    ram_cell[    2565] = 32'h0;  // 32'h4112875b;
    ram_cell[    2566] = 32'h0;  // 32'hd595af96;
    ram_cell[    2567] = 32'h0;  // 32'he4ed076d;
    ram_cell[    2568] = 32'h0;  // 32'h24fc66bc;
    ram_cell[    2569] = 32'h0;  // 32'h4b936e9f;
    ram_cell[    2570] = 32'h0;  // 32'h230a5d1e;
    ram_cell[    2571] = 32'h0;  // 32'h90f915d9;
    ram_cell[    2572] = 32'h0;  // 32'hef790810;
    ram_cell[    2573] = 32'h0;  // 32'h38f716d8;
    ram_cell[    2574] = 32'h0;  // 32'h2e4def42;
    ram_cell[    2575] = 32'h0;  // 32'h7635285e;
    ram_cell[    2576] = 32'h0;  // 32'hb9cfa386;
    ram_cell[    2577] = 32'h0;  // 32'hc45ec5af;
    ram_cell[    2578] = 32'h0;  // 32'h4c9e8526;
    ram_cell[    2579] = 32'h0;  // 32'hb7c24fd6;
    ram_cell[    2580] = 32'h0;  // 32'h0fd1a3d6;
    ram_cell[    2581] = 32'h0;  // 32'h0d9a1ac7;
    ram_cell[    2582] = 32'h0;  // 32'h77b00164;
    ram_cell[    2583] = 32'h0;  // 32'ha208c554;
    ram_cell[    2584] = 32'h0;  // 32'hd5030569;
    ram_cell[    2585] = 32'h0;  // 32'he78b8ea5;
    ram_cell[    2586] = 32'h0;  // 32'hcc5fdffe;
    ram_cell[    2587] = 32'h0;  // 32'h0d9866a7;
    ram_cell[    2588] = 32'h0;  // 32'h7699de77;
    ram_cell[    2589] = 32'h0;  // 32'hf3c380cc;
    ram_cell[    2590] = 32'h0;  // 32'he436ce94;
    ram_cell[    2591] = 32'h0;  // 32'h3c607dd3;
    ram_cell[    2592] = 32'h0;  // 32'hf02119d4;
    ram_cell[    2593] = 32'h0;  // 32'h1c2d81e6;
    ram_cell[    2594] = 32'h0;  // 32'h075377af;
    ram_cell[    2595] = 32'h0;  // 32'h92b051cb;
    ram_cell[    2596] = 32'h0;  // 32'hc8d78f27;
    ram_cell[    2597] = 32'h0;  // 32'ha22b5dd3;
    ram_cell[    2598] = 32'h0;  // 32'ha7c35a66;
    ram_cell[    2599] = 32'h0;  // 32'h564d3bc1;
    ram_cell[    2600] = 32'h0;  // 32'h0105e75a;
    ram_cell[    2601] = 32'h0;  // 32'hbc33e665;
    ram_cell[    2602] = 32'h0;  // 32'h69459a7b;
    ram_cell[    2603] = 32'h0;  // 32'h9271f18f;
    ram_cell[    2604] = 32'h0;  // 32'h84f4d113;
    ram_cell[    2605] = 32'h0;  // 32'h1dce9675;
    ram_cell[    2606] = 32'h0;  // 32'heb543cfe;
    ram_cell[    2607] = 32'h0;  // 32'h59c3fa9d;
    ram_cell[    2608] = 32'h0;  // 32'h7caa853b;
    ram_cell[    2609] = 32'h0;  // 32'hec8a87df;
    ram_cell[    2610] = 32'h0;  // 32'hee556d4c;
    ram_cell[    2611] = 32'h0;  // 32'h02ef7b13;
    ram_cell[    2612] = 32'h0;  // 32'h66bba118;
    ram_cell[    2613] = 32'h0;  // 32'h85e529f3;
    ram_cell[    2614] = 32'h0;  // 32'h7f7eec08;
    ram_cell[    2615] = 32'h0;  // 32'h68ccd15a;
    ram_cell[    2616] = 32'h0;  // 32'h25588f43;
    ram_cell[    2617] = 32'h0;  // 32'hb95d795e;
    ram_cell[    2618] = 32'h0;  // 32'hbc22df29;
    ram_cell[    2619] = 32'h0;  // 32'h59821d54;
    ram_cell[    2620] = 32'h0;  // 32'haa5e1ff8;
    ram_cell[    2621] = 32'h0;  // 32'h4c546549;
    ram_cell[    2622] = 32'h0;  // 32'h90a3c82d;
    ram_cell[    2623] = 32'h0;  // 32'hea8b875c;
    ram_cell[    2624] = 32'h0;  // 32'h1545ec3f;
    ram_cell[    2625] = 32'h0;  // 32'h89f87c67;
    ram_cell[    2626] = 32'h0;  // 32'h81b0e474;
    ram_cell[    2627] = 32'h0;  // 32'h81711262;
    ram_cell[    2628] = 32'h0;  // 32'hb9e67c05;
    ram_cell[    2629] = 32'h0;  // 32'h80572599;
    ram_cell[    2630] = 32'h0;  // 32'h1370e42e;
    ram_cell[    2631] = 32'h0;  // 32'h05f7c381;
    ram_cell[    2632] = 32'h0;  // 32'h9eea2041;
    ram_cell[    2633] = 32'h0;  // 32'h4207fc0d;
    ram_cell[    2634] = 32'h0;  // 32'hb7b90f34;
    ram_cell[    2635] = 32'h0;  // 32'h3ef353ca;
    ram_cell[    2636] = 32'h0;  // 32'ha5c4a89e;
    ram_cell[    2637] = 32'h0;  // 32'h1e87dc67;
    ram_cell[    2638] = 32'h0;  // 32'h8c79141c;
    ram_cell[    2639] = 32'h0;  // 32'hf3577299;
    ram_cell[    2640] = 32'h0;  // 32'he789483a;
    ram_cell[    2641] = 32'h0;  // 32'h2bab9671;
    ram_cell[    2642] = 32'h0;  // 32'hc0d77829;
    ram_cell[    2643] = 32'h0;  // 32'h7da93a68;
    ram_cell[    2644] = 32'h0;  // 32'h05229dc8;
    ram_cell[    2645] = 32'h0;  // 32'h7a0afb7d;
    ram_cell[    2646] = 32'h0;  // 32'h06783f78;
    ram_cell[    2647] = 32'h0;  // 32'hf0d5f720;
    ram_cell[    2648] = 32'h0;  // 32'h71dc480f;
    ram_cell[    2649] = 32'h0;  // 32'h7cd67f7b;
    ram_cell[    2650] = 32'h0;  // 32'h68cefa77;
    ram_cell[    2651] = 32'h0;  // 32'h03d8aeb2;
    ram_cell[    2652] = 32'h0;  // 32'h59f96a30;
    ram_cell[    2653] = 32'h0;  // 32'hec2774d6;
    ram_cell[    2654] = 32'h0;  // 32'hfcab7ea2;
    ram_cell[    2655] = 32'h0;  // 32'h4ecdd20b;
    ram_cell[    2656] = 32'h0;  // 32'h6b25af0b;
    ram_cell[    2657] = 32'h0;  // 32'hbac0d753;
    ram_cell[    2658] = 32'h0;  // 32'h6de070f9;
    ram_cell[    2659] = 32'h0;  // 32'hc8b5896b;
    ram_cell[    2660] = 32'h0;  // 32'hcc170ff7;
    ram_cell[    2661] = 32'h0;  // 32'h8cb05618;
    ram_cell[    2662] = 32'h0;  // 32'hada6b51e;
    ram_cell[    2663] = 32'h0;  // 32'h6b67f52f;
    ram_cell[    2664] = 32'h0;  // 32'h291b8e72;
    ram_cell[    2665] = 32'h0;  // 32'hf9c023c1;
    ram_cell[    2666] = 32'h0;  // 32'h92f77a24;
    ram_cell[    2667] = 32'h0;  // 32'h1a6d974b;
    ram_cell[    2668] = 32'h0;  // 32'h2b37b3a9;
    ram_cell[    2669] = 32'h0;  // 32'h142f9036;
    ram_cell[    2670] = 32'h0;  // 32'he5f3cf1e;
    ram_cell[    2671] = 32'h0;  // 32'h0bc39023;
    ram_cell[    2672] = 32'h0;  // 32'h8b725c7b;
    ram_cell[    2673] = 32'h0;  // 32'h81595aae;
    ram_cell[    2674] = 32'h0;  // 32'h60a6a018;
    ram_cell[    2675] = 32'h0;  // 32'h18ea2564;
    ram_cell[    2676] = 32'h0;  // 32'hb8de1a87;
    ram_cell[    2677] = 32'h0;  // 32'h1469af1b;
    ram_cell[    2678] = 32'h0;  // 32'h2c637e78;
    ram_cell[    2679] = 32'h0;  // 32'h869e8698;
    ram_cell[    2680] = 32'h0;  // 32'hc7ecd7f4;
    ram_cell[    2681] = 32'h0;  // 32'hb99ea219;
    ram_cell[    2682] = 32'h0;  // 32'h66b7f9ec;
    ram_cell[    2683] = 32'h0;  // 32'h2a2156ff;
    ram_cell[    2684] = 32'h0;  // 32'h0cb5dbe8;
    ram_cell[    2685] = 32'h0;  // 32'hec47d7dc;
    ram_cell[    2686] = 32'h0;  // 32'hcf37b872;
    ram_cell[    2687] = 32'h0;  // 32'hc9b53c59;
    ram_cell[    2688] = 32'h0;  // 32'hcafeadc3;
    ram_cell[    2689] = 32'h0;  // 32'h1ab2f376;
    ram_cell[    2690] = 32'h0;  // 32'hb8f7c2ff;
    ram_cell[    2691] = 32'h0;  // 32'hf45db526;
    ram_cell[    2692] = 32'h0;  // 32'he81af193;
    ram_cell[    2693] = 32'h0;  // 32'h1c032679;
    ram_cell[    2694] = 32'h0;  // 32'hf6705979;
    ram_cell[    2695] = 32'h0;  // 32'hf7fa5e8e;
    ram_cell[    2696] = 32'h0;  // 32'h5db04a1a;
    ram_cell[    2697] = 32'h0;  // 32'ha24db3ee;
    ram_cell[    2698] = 32'h0;  // 32'h00dce58d;
    ram_cell[    2699] = 32'h0;  // 32'hd3b8939b;
    ram_cell[    2700] = 32'h0;  // 32'h2916477f;
    ram_cell[    2701] = 32'h0;  // 32'h6c951dab;
    ram_cell[    2702] = 32'h0;  // 32'heee86c78;
    ram_cell[    2703] = 32'h0;  // 32'h0472e126;
    ram_cell[    2704] = 32'h0;  // 32'h17e9d9ec;
    ram_cell[    2705] = 32'h0;  // 32'h2f981c1c;
    ram_cell[    2706] = 32'h0;  // 32'h4f9dec93;
    ram_cell[    2707] = 32'h0;  // 32'h4c0f179f;
    ram_cell[    2708] = 32'h0;  // 32'h77554887;
    ram_cell[    2709] = 32'h0;  // 32'hf547b254;
    ram_cell[    2710] = 32'h0;  // 32'hbb3ebe7f;
    ram_cell[    2711] = 32'h0;  // 32'hf91dce19;
    ram_cell[    2712] = 32'h0;  // 32'hbd87212a;
    ram_cell[    2713] = 32'h0;  // 32'hf39feae3;
    ram_cell[    2714] = 32'h0;  // 32'hcff01393;
    ram_cell[    2715] = 32'h0;  // 32'h611f262b;
    ram_cell[    2716] = 32'h0;  // 32'h0b6519de;
    ram_cell[    2717] = 32'h0;  // 32'hb366ff04;
    ram_cell[    2718] = 32'h0;  // 32'he92c169c;
    ram_cell[    2719] = 32'h0;  // 32'h285e9b5e;
    ram_cell[    2720] = 32'h0;  // 32'h81c65536;
    ram_cell[    2721] = 32'h0;  // 32'h11769f94;
    ram_cell[    2722] = 32'h0;  // 32'h0e09fa91;
    ram_cell[    2723] = 32'h0;  // 32'h0f72384b;
    ram_cell[    2724] = 32'h0;  // 32'h56f0c9d1;
    ram_cell[    2725] = 32'h0;  // 32'hf47fb239;
    ram_cell[    2726] = 32'h0;  // 32'hf85d3512;
    ram_cell[    2727] = 32'h0;  // 32'h9e2f0d02;
    ram_cell[    2728] = 32'h0;  // 32'h8d709452;
    ram_cell[    2729] = 32'h0;  // 32'hb9d53fe2;
    ram_cell[    2730] = 32'h0;  // 32'he148e451;
    ram_cell[    2731] = 32'h0;  // 32'h2d9ef0f1;
    ram_cell[    2732] = 32'h0;  // 32'hda0ec204;
    ram_cell[    2733] = 32'h0;  // 32'h6f2f1e47;
    ram_cell[    2734] = 32'h0;  // 32'h5e129cd0;
    ram_cell[    2735] = 32'h0;  // 32'hdf4013d1;
    ram_cell[    2736] = 32'h0;  // 32'hc502059a;
    ram_cell[    2737] = 32'h0;  // 32'h8d26860d;
    ram_cell[    2738] = 32'h0;  // 32'h15addaa3;
    ram_cell[    2739] = 32'h0;  // 32'hd5ea3957;
    ram_cell[    2740] = 32'h0;  // 32'h5f1b1b55;
    ram_cell[    2741] = 32'h0;  // 32'h7e3fdc83;
    ram_cell[    2742] = 32'h0;  // 32'h5f5d83b2;
    ram_cell[    2743] = 32'h0;  // 32'h763f33d4;
    ram_cell[    2744] = 32'h0;  // 32'hfe9089b6;
    ram_cell[    2745] = 32'h0;  // 32'hf32b4f08;
    ram_cell[    2746] = 32'h0;  // 32'hef4241e0;
    ram_cell[    2747] = 32'h0;  // 32'h02d6a570;
    ram_cell[    2748] = 32'h0;  // 32'h482d0aae;
    ram_cell[    2749] = 32'h0;  // 32'h03f47402;
    ram_cell[    2750] = 32'h0;  // 32'hb7d3e8e2;
    ram_cell[    2751] = 32'h0;  // 32'h6893a684;
    ram_cell[    2752] = 32'h0;  // 32'h79c39d1c;
    ram_cell[    2753] = 32'h0;  // 32'hf713a78e;
    ram_cell[    2754] = 32'h0;  // 32'h462fc6a2;
    ram_cell[    2755] = 32'h0;  // 32'ha3079ace;
    ram_cell[    2756] = 32'h0;  // 32'hf179ed89;
    ram_cell[    2757] = 32'h0;  // 32'h82f0a1a2;
    ram_cell[    2758] = 32'h0;  // 32'hcda36ddc;
    ram_cell[    2759] = 32'h0;  // 32'h973172a4;
    ram_cell[    2760] = 32'h0;  // 32'hfc55828f;
    ram_cell[    2761] = 32'h0;  // 32'h486930a4;
    ram_cell[    2762] = 32'h0;  // 32'hd6e19046;
    ram_cell[    2763] = 32'h0;  // 32'h9c90021a;
    ram_cell[    2764] = 32'h0;  // 32'h2a7cf83f;
    ram_cell[    2765] = 32'h0;  // 32'hdffe243d;
    ram_cell[    2766] = 32'h0;  // 32'h9dfdb907;
    ram_cell[    2767] = 32'h0;  // 32'h34bb141a;
    ram_cell[    2768] = 32'h0;  // 32'h80ce2f9c;
    ram_cell[    2769] = 32'h0;  // 32'hef9f32c9;
    ram_cell[    2770] = 32'h0;  // 32'hbf42c4f9;
    ram_cell[    2771] = 32'h0;  // 32'hdfe6345f;
    ram_cell[    2772] = 32'h0;  // 32'hce9e5cfa;
    ram_cell[    2773] = 32'h0;  // 32'h50330324;
    ram_cell[    2774] = 32'h0;  // 32'h84d31a9a;
    ram_cell[    2775] = 32'h0;  // 32'heffc06a9;
    ram_cell[    2776] = 32'h0;  // 32'hb5b498d4;
    ram_cell[    2777] = 32'h0;  // 32'h3e0ec93a;
    ram_cell[    2778] = 32'h0;  // 32'h87cbac92;
    ram_cell[    2779] = 32'h0;  // 32'h9121b137;
    ram_cell[    2780] = 32'h0;  // 32'hd65c838a;
    ram_cell[    2781] = 32'h0;  // 32'h66cbda11;
    ram_cell[    2782] = 32'h0;  // 32'h130c4469;
    ram_cell[    2783] = 32'h0;  // 32'h79f8af01;
    ram_cell[    2784] = 32'h0;  // 32'hadbddfa8;
    ram_cell[    2785] = 32'h0;  // 32'h03d7989e;
    ram_cell[    2786] = 32'h0;  // 32'he6f3b2bd;
    ram_cell[    2787] = 32'h0;  // 32'h6c158eb9;
    ram_cell[    2788] = 32'h0;  // 32'h85ee9d41;
    ram_cell[    2789] = 32'h0;  // 32'h9e60c2ad;
    ram_cell[    2790] = 32'h0;  // 32'h2a1c8910;
    ram_cell[    2791] = 32'h0;  // 32'hfa2fab73;
    ram_cell[    2792] = 32'h0;  // 32'h8e719f7a;
    ram_cell[    2793] = 32'h0;  // 32'ha65e8f04;
    ram_cell[    2794] = 32'h0;  // 32'h7cd65679;
    ram_cell[    2795] = 32'h0;  // 32'h8c367989;
    ram_cell[    2796] = 32'h0;  // 32'h223b96e7;
    ram_cell[    2797] = 32'h0;  // 32'hc555e536;
    ram_cell[    2798] = 32'h0;  // 32'h22888f2f;
    ram_cell[    2799] = 32'h0;  // 32'h9d574353;
    ram_cell[    2800] = 32'h0;  // 32'h8c4375e1;
    ram_cell[    2801] = 32'h0;  // 32'h186691aa;
    ram_cell[    2802] = 32'h0;  // 32'haf9decaa;
    ram_cell[    2803] = 32'h0;  // 32'h132c5103;
    ram_cell[    2804] = 32'h0;  // 32'h7dd7109f;
    ram_cell[    2805] = 32'h0;  // 32'h6754be4b;
    ram_cell[    2806] = 32'h0;  // 32'hb41d89ed;
    ram_cell[    2807] = 32'h0;  // 32'h7f4855e7;
    ram_cell[    2808] = 32'h0;  // 32'ha7055017;
    ram_cell[    2809] = 32'h0;  // 32'h54020744;
    ram_cell[    2810] = 32'h0;  // 32'hc20ded05;
    ram_cell[    2811] = 32'h0;  // 32'h881f26a5;
    ram_cell[    2812] = 32'h0;  // 32'hecb89169;
    ram_cell[    2813] = 32'h0;  // 32'ha97954df;
    ram_cell[    2814] = 32'h0;  // 32'ha4f2ef49;
    ram_cell[    2815] = 32'h0;  // 32'h425baf31;
    ram_cell[    2816] = 32'h0;  // 32'h61af350b;
    ram_cell[    2817] = 32'h0;  // 32'h726b88b0;
    ram_cell[    2818] = 32'h0;  // 32'hee60a7d9;
    ram_cell[    2819] = 32'h0;  // 32'hc235e905;
    ram_cell[    2820] = 32'h0;  // 32'h1cffbc3b;
    ram_cell[    2821] = 32'h0;  // 32'h7d46ec41;
    ram_cell[    2822] = 32'h0;  // 32'h6f13049c;
    ram_cell[    2823] = 32'h0;  // 32'hcb385c5a;
    ram_cell[    2824] = 32'h0;  // 32'h133bad84;
    ram_cell[    2825] = 32'h0;  // 32'he92cd8a3;
    ram_cell[    2826] = 32'h0;  // 32'h3f363a55;
    ram_cell[    2827] = 32'h0;  // 32'hfa32d2a4;
    ram_cell[    2828] = 32'h0;  // 32'h899acc8b;
    ram_cell[    2829] = 32'h0;  // 32'h1783be59;
    ram_cell[    2830] = 32'h0;  // 32'hb7178bc1;
    ram_cell[    2831] = 32'h0;  // 32'h1ec2fbb8;
    ram_cell[    2832] = 32'h0;  // 32'h7705635f;
    ram_cell[    2833] = 32'h0;  // 32'h54bf9917;
    ram_cell[    2834] = 32'h0;  // 32'h383e75a2;
    ram_cell[    2835] = 32'h0;  // 32'h7a641638;
    ram_cell[    2836] = 32'h0;  // 32'h6e622390;
    ram_cell[    2837] = 32'h0;  // 32'h125e41bb;
    ram_cell[    2838] = 32'h0;  // 32'h42d1bef0;
    ram_cell[    2839] = 32'h0;  // 32'hf2b6494a;
    ram_cell[    2840] = 32'h0;  // 32'hc03a2338;
    ram_cell[    2841] = 32'h0;  // 32'hb9f31e8e;
    ram_cell[    2842] = 32'h0;  // 32'h2446760e;
    ram_cell[    2843] = 32'h0;  // 32'hd290b1e5;
    ram_cell[    2844] = 32'h0;  // 32'hb51d6016;
    ram_cell[    2845] = 32'h0;  // 32'ha7917163;
    ram_cell[    2846] = 32'h0;  // 32'hd26f268c;
    ram_cell[    2847] = 32'h0;  // 32'h2d8b43c8;
    ram_cell[    2848] = 32'h0;  // 32'h11e2b078;
    ram_cell[    2849] = 32'h0;  // 32'hee93c890;
    ram_cell[    2850] = 32'h0;  // 32'h6c39ef30;
    ram_cell[    2851] = 32'h0;  // 32'hac3663e2;
    ram_cell[    2852] = 32'h0;  // 32'h1a96fb38;
    ram_cell[    2853] = 32'h0;  // 32'hc1c334c4;
    ram_cell[    2854] = 32'h0;  // 32'h7215a97a;
    ram_cell[    2855] = 32'h0;  // 32'h9f952320;
    ram_cell[    2856] = 32'h0;  // 32'h48e1aa54;
    ram_cell[    2857] = 32'h0;  // 32'h82e37e7c;
    ram_cell[    2858] = 32'h0;  // 32'h17a5c237;
    ram_cell[    2859] = 32'h0;  // 32'h31338013;
    ram_cell[    2860] = 32'h0;  // 32'h8d56c7c2;
    ram_cell[    2861] = 32'h0;  // 32'hef002915;
    ram_cell[    2862] = 32'h0;  // 32'hed6c412e;
    ram_cell[    2863] = 32'h0;  // 32'h953f5c82;
    ram_cell[    2864] = 32'h0;  // 32'h0014b897;
    ram_cell[    2865] = 32'h0;  // 32'h6161a05b;
    ram_cell[    2866] = 32'h0;  // 32'h29a431cc;
    ram_cell[    2867] = 32'h0;  // 32'h86cbd843;
    ram_cell[    2868] = 32'h0;  // 32'h3be155b0;
    ram_cell[    2869] = 32'h0;  // 32'h6fcb9cc0;
    ram_cell[    2870] = 32'h0;  // 32'h9fdb14e4;
    ram_cell[    2871] = 32'h0;  // 32'h20717174;
    ram_cell[    2872] = 32'h0;  // 32'h7ac1f25a;
    ram_cell[    2873] = 32'h0;  // 32'hbaae0c94;
    ram_cell[    2874] = 32'h0;  // 32'h1deff51f;
    ram_cell[    2875] = 32'h0;  // 32'h10709962;
    ram_cell[    2876] = 32'h0;  // 32'h35d1f959;
    ram_cell[    2877] = 32'h0;  // 32'hd1ea2771;
    ram_cell[    2878] = 32'h0;  // 32'ha052a4e9;
    ram_cell[    2879] = 32'h0;  // 32'h21188e8d;
    ram_cell[    2880] = 32'h0;  // 32'haa9127b3;
    ram_cell[    2881] = 32'h0;  // 32'h7a6d6ea1;
    ram_cell[    2882] = 32'h0;  // 32'h0edad89d;
    ram_cell[    2883] = 32'h0;  // 32'h5b6f0ebd;
    ram_cell[    2884] = 32'h0;  // 32'h29ad611f;
    ram_cell[    2885] = 32'h0;  // 32'h604bc6be;
    ram_cell[    2886] = 32'h0;  // 32'h0a4331c4;
    ram_cell[    2887] = 32'h0;  // 32'h3ca1a7df;
    ram_cell[    2888] = 32'h0;  // 32'h827147c1;
    ram_cell[    2889] = 32'h0;  // 32'hfb7918c6;
    ram_cell[    2890] = 32'h0;  // 32'ha9f7230f;
    ram_cell[    2891] = 32'h0;  // 32'hd4176601;
    ram_cell[    2892] = 32'h0;  // 32'h9ca906f6;
    ram_cell[    2893] = 32'h0;  // 32'h264e2be4;
    ram_cell[    2894] = 32'h0;  // 32'hb50d1ce9;
    ram_cell[    2895] = 32'h0;  // 32'h9c58aaad;
    ram_cell[    2896] = 32'h0;  // 32'h0066cc4e;
    ram_cell[    2897] = 32'h0;  // 32'h7bb555ab;
    ram_cell[    2898] = 32'h0;  // 32'hdec940c4;
    ram_cell[    2899] = 32'h0;  // 32'hff271bcf;
    ram_cell[    2900] = 32'h0;  // 32'h09b86214;
    ram_cell[    2901] = 32'h0;  // 32'hd69414e2;
    ram_cell[    2902] = 32'h0;  // 32'h376c7473;
    ram_cell[    2903] = 32'h0;  // 32'h0e8030e2;
    ram_cell[    2904] = 32'h0;  // 32'h9ea521ea;
    ram_cell[    2905] = 32'h0;  // 32'h015d6123;
    ram_cell[    2906] = 32'h0;  // 32'h4dd519c7;
    ram_cell[    2907] = 32'h0;  // 32'h05e39b8c;
    ram_cell[    2908] = 32'h0;  // 32'hd202fc53;
    ram_cell[    2909] = 32'h0;  // 32'hc8238a2b;
    ram_cell[    2910] = 32'h0;  // 32'h23285871;
    ram_cell[    2911] = 32'h0;  // 32'h420ded9f;
    ram_cell[    2912] = 32'h0;  // 32'hb949cb4d;
    ram_cell[    2913] = 32'h0;  // 32'hf9db3201;
    ram_cell[    2914] = 32'h0;  // 32'h1a22946f;
    ram_cell[    2915] = 32'h0;  // 32'h362aeb21;
    ram_cell[    2916] = 32'h0;  // 32'h7b6b418d;
    ram_cell[    2917] = 32'h0;  // 32'hdafbf875;
    ram_cell[    2918] = 32'h0;  // 32'h3c46fe69;
    ram_cell[    2919] = 32'h0;  // 32'hc0a877d6;
    ram_cell[    2920] = 32'h0;  // 32'hbe54c414;
    ram_cell[    2921] = 32'h0;  // 32'h7f15fe2d;
    ram_cell[    2922] = 32'h0;  // 32'h064232fd;
    ram_cell[    2923] = 32'h0;  // 32'h9ba5baae;
    ram_cell[    2924] = 32'h0;  // 32'hdc1cfa7b;
    ram_cell[    2925] = 32'h0;  // 32'h2088e6e2;
    ram_cell[    2926] = 32'h0;  // 32'h10a8b85c;
    ram_cell[    2927] = 32'h0;  // 32'h6fd35c01;
    ram_cell[    2928] = 32'h0;  // 32'hc6c46fdc;
    ram_cell[    2929] = 32'h0;  // 32'hfa8c73b8;
    ram_cell[    2930] = 32'h0;  // 32'hccaad090;
    ram_cell[    2931] = 32'h0;  // 32'hd455fdf3;
    ram_cell[    2932] = 32'h0;  // 32'h5ffee396;
    ram_cell[    2933] = 32'h0;  // 32'h3c595175;
    ram_cell[    2934] = 32'h0;  // 32'hf36ce3ce;
    ram_cell[    2935] = 32'h0;  // 32'h2701caf0;
    ram_cell[    2936] = 32'h0;  // 32'h728def41;
    ram_cell[    2937] = 32'h0;  // 32'hec3a7902;
    ram_cell[    2938] = 32'h0;  // 32'h56d83dff;
    ram_cell[    2939] = 32'h0;  // 32'hd2287ad4;
    ram_cell[    2940] = 32'h0;  // 32'h6cf37e79;
    ram_cell[    2941] = 32'h0;  // 32'haf72ae5d;
    ram_cell[    2942] = 32'h0;  // 32'h9c65ca5b;
    ram_cell[    2943] = 32'h0;  // 32'he084a710;
    ram_cell[    2944] = 32'h0;  // 32'h4cf0288b;
    ram_cell[    2945] = 32'h0;  // 32'ha389e177;
    ram_cell[    2946] = 32'h0;  // 32'h94612ea8;
    ram_cell[    2947] = 32'h0;  // 32'h3f327e19;
    ram_cell[    2948] = 32'h0;  // 32'h3e83f22d;
    ram_cell[    2949] = 32'h0;  // 32'h0688372c;
    ram_cell[    2950] = 32'h0;  // 32'h3bc65b2e;
    ram_cell[    2951] = 32'h0;  // 32'he11b809e;
    ram_cell[    2952] = 32'h0;  // 32'hc58d5df2;
    ram_cell[    2953] = 32'h0;  // 32'h766d8ac5;
    ram_cell[    2954] = 32'h0;  // 32'h5d3d5863;
    ram_cell[    2955] = 32'h0;  // 32'h460f75bb;
    ram_cell[    2956] = 32'h0;  // 32'hcadff64f;
    ram_cell[    2957] = 32'h0;  // 32'h333b8ed4;
    ram_cell[    2958] = 32'h0;  // 32'h6c483a51;
    ram_cell[    2959] = 32'h0;  // 32'h66e743a3;
    ram_cell[    2960] = 32'h0;  // 32'hb78704f5;
    ram_cell[    2961] = 32'h0;  // 32'h6d6c80df;
    ram_cell[    2962] = 32'h0;  // 32'hdb2f56d2;
    ram_cell[    2963] = 32'h0;  // 32'h86267408;
    ram_cell[    2964] = 32'h0;  // 32'h3bfdb622;
    ram_cell[    2965] = 32'h0;  // 32'hbef2ceaf;
    ram_cell[    2966] = 32'h0;  // 32'h112ac2f2;
    ram_cell[    2967] = 32'h0;  // 32'h1d11b2fc;
    ram_cell[    2968] = 32'h0;  // 32'h059dab9a;
    ram_cell[    2969] = 32'h0;  // 32'h70877168;
    ram_cell[    2970] = 32'h0;  // 32'h47f95a30;
    ram_cell[    2971] = 32'h0;  // 32'h94adf1a5;
    ram_cell[    2972] = 32'h0;  // 32'h0500dbb1;
    ram_cell[    2973] = 32'h0;  // 32'hfebf2092;
    ram_cell[    2974] = 32'h0;  // 32'ha2b6dd41;
    ram_cell[    2975] = 32'h0;  // 32'h673aa1d6;
    ram_cell[    2976] = 32'h0;  // 32'h33e1f538;
    ram_cell[    2977] = 32'h0;  // 32'hf72af03e;
    ram_cell[    2978] = 32'h0;  // 32'hf5dcf0c8;
    ram_cell[    2979] = 32'h0;  // 32'ha653a2aa;
    ram_cell[    2980] = 32'h0;  // 32'h4c8f3353;
    ram_cell[    2981] = 32'h0;  // 32'h3a9cfa51;
    ram_cell[    2982] = 32'h0;  // 32'h2ccb0bd4;
    ram_cell[    2983] = 32'h0;  // 32'ha12456e0;
    ram_cell[    2984] = 32'h0;  // 32'h5d83268c;
    ram_cell[    2985] = 32'h0;  // 32'h5ad2aa53;
    ram_cell[    2986] = 32'h0;  // 32'h035ea02c;
    ram_cell[    2987] = 32'h0;  // 32'h3d440906;
    ram_cell[    2988] = 32'h0;  // 32'hb4c6a15b;
    ram_cell[    2989] = 32'h0;  // 32'h592b9101;
    ram_cell[    2990] = 32'h0;  // 32'hb1544896;
    ram_cell[    2991] = 32'h0;  // 32'h2cef07ac;
    ram_cell[    2992] = 32'h0;  // 32'h489aba33;
    ram_cell[    2993] = 32'h0;  // 32'hd37938da;
    ram_cell[    2994] = 32'h0;  // 32'h8887e946;
    ram_cell[    2995] = 32'h0;  // 32'hfd333856;
    ram_cell[    2996] = 32'h0;  // 32'h1a326abf;
    ram_cell[    2997] = 32'h0;  // 32'h5365288a;
    ram_cell[    2998] = 32'h0;  // 32'he1d723c0;
    ram_cell[    2999] = 32'h0;  // 32'hfc5575da;
    ram_cell[    3000] = 32'h0;  // 32'h48f08b77;
    ram_cell[    3001] = 32'h0;  // 32'h665b35dd;
    ram_cell[    3002] = 32'h0;  // 32'h2fb94629;
    ram_cell[    3003] = 32'h0;  // 32'h0aaed971;
    ram_cell[    3004] = 32'h0;  // 32'hfe3b4f61;
    ram_cell[    3005] = 32'h0;  // 32'h48dbf39a;
    ram_cell[    3006] = 32'h0;  // 32'hca1c41b9;
    ram_cell[    3007] = 32'h0;  // 32'h53644673;
    ram_cell[    3008] = 32'h0;  // 32'hed06122f;
    ram_cell[    3009] = 32'h0;  // 32'h14137055;
    ram_cell[    3010] = 32'h0;  // 32'h6fe22d64;
    ram_cell[    3011] = 32'h0;  // 32'hfb03ae5d;
    ram_cell[    3012] = 32'h0;  // 32'h18e47f7a;
    ram_cell[    3013] = 32'h0;  // 32'h7442f7e1;
    ram_cell[    3014] = 32'h0;  // 32'hd4be745d;
    ram_cell[    3015] = 32'h0;  // 32'h32fd391d;
    ram_cell[    3016] = 32'h0;  // 32'h4e8849c9;
    ram_cell[    3017] = 32'h0;  // 32'h7648ce5e;
    ram_cell[    3018] = 32'h0;  // 32'ha07e16ff;
    ram_cell[    3019] = 32'h0;  // 32'he4ace4d9;
    ram_cell[    3020] = 32'h0;  // 32'hcc935f3e;
    ram_cell[    3021] = 32'h0;  // 32'hb2579ffd;
    ram_cell[    3022] = 32'h0;  // 32'he977d281;
    ram_cell[    3023] = 32'h0;  // 32'hd9dd5fc2;
    ram_cell[    3024] = 32'h0;  // 32'ha6696b35;
    ram_cell[    3025] = 32'h0;  // 32'hfd9b702f;
    ram_cell[    3026] = 32'h0;  // 32'h5b9d8da4;
    ram_cell[    3027] = 32'h0;  // 32'h3108c2ed;
    ram_cell[    3028] = 32'h0;  // 32'hca9df364;
    ram_cell[    3029] = 32'h0;  // 32'h8fc440ed;
    ram_cell[    3030] = 32'h0;  // 32'h1fe50e5e;
    ram_cell[    3031] = 32'h0;  // 32'h9b769001;
    ram_cell[    3032] = 32'h0;  // 32'h6adc32a0;
    ram_cell[    3033] = 32'h0;  // 32'hab6672a2;
    ram_cell[    3034] = 32'h0;  // 32'h803b0cf4;
    ram_cell[    3035] = 32'h0;  // 32'hbb434376;
    ram_cell[    3036] = 32'h0;  // 32'h84ec9bba;
    ram_cell[    3037] = 32'h0;  // 32'h3da01c72;
    ram_cell[    3038] = 32'h0;  // 32'h3d8e3a58;
    ram_cell[    3039] = 32'h0;  // 32'hc242f71f;
    ram_cell[    3040] = 32'h0;  // 32'h3c5da12f;
    ram_cell[    3041] = 32'h0;  // 32'hf62b6930;
    ram_cell[    3042] = 32'h0;  // 32'hbe05e793;
    ram_cell[    3043] = 32'h0;  // 32'hb2a6c78a;
    ram_cell[    3044] = 32'h0;  // 32'hfc5bdeab;
    ram_cell[    3045] = 32'h0;  // 32'he71c67d8;
    ram_cell[    3046] = 32'h0;  // 32'heafad8cf;
    ram_cell[    3047] = 32'h0;  // 32'h9c9afa58;
    ram_cell[    3048] = 32'h0;  // 32'hfef917e0;
    ram_cell[    3049] = 32'h0;  // 32'h443add17;
    ram_cell[    3050] = 32'h0;  // 32'h2a11e94d;
    ram_cell[    3051] = 32'h0;  // 32'hd10eeb98;
    ram_cell[    3052] = 32'h0;  // 32'heb5ae179;
    ram_cell[    3053] = 32'h0;  // 32'hd77b7942;
    ram_cell[    3054] = 32'h0;  // 32'h51c6d851;
    ram_cell[    3055] = 32'h0;  // 32'h2fa99fa6;
    ram_cell[    3056] = 32'h0;  // 32'h3b1fb95a;
    ram_cell[    3057] = 32'h0;  // 32'hd83a5283;
    ram_cell[    3058] = 32'h0;  // 32'h771949a2;
    ram_cell[    3059] = 32'h0;  // 32'hef1a025c;
    ram_cell[    3060] = 32'h0;  // 32'h63fc38f1;
    ram_cell[    3061] = 32'h0;  // 32'hf4fede0a;
    ram_cell[    3062] = 32'h0;  // 32'h735f45db;
    ram_cell[    3063] = 32'h0;  // 32'hb34caee4;
    ram_cell[    3064] = 32'h0;  // 32'haf205da6;
    ram_cell[    3065] = 32'h0;  // 32'hac136cb1;
    ram_cell[    3066] = 32'h0;  // 32'h680dd254;
    ram_cell[    3067] = 32'h0;  // 32'h22e2417e;
    ram_cell[    3068] = 32'h0;  // 32'hbced93ab;
    ram_cell[    3069] = 32'h0;  // 32'h3a882612;
    ram_cell[    3070] = 32'h0;  // 32'h7bf58651;
    ram_cell[    3071] = 32'h0;  // 32'hbca75ad0;
    ram_cell[    3072] = 32'h0;  // 32'hfb0d082a;
    ram_cell[    3073] = 32'h0;  // 32'heffc68f6;
    ram_cell[    3074] = 32'h0;  // 32'hdd742674;
    ram_cell[    3075] = 32'h0;  // 32'h47efe1d2;
    ram_cell[    3076] = 32'h0;  // 32'hb46ff446;
    ram_cell[    3077] = 32'h0;  // 32'h5dad6896;
    ram_cell[    3078] = 32'h0;  // 32'h56e05fef;
    ram_cell[    3079] = 32'h0;  // 32'h4c1081e0;
    ram_cell[    3080] = 32'h0;  // 32'he47187d4;
    ram_cell[    3081] = 32'h0;  // 32'h42d92190;
    ram_cell[    3082] = 32'h0;  // 32'h6d76f0ad;
    ram_cell[    3083] = 32'h0;  // 32'h637adc9c;
    ram_cell[    3084] = 32'h0;  // 32'h572cbba4;
    ram_cell[    3085] = 32'h0;  // 32'hcb8de18b;
    ram_cell[    3086] = 32'h0;  // 32'ha854ebd7;
    ram_cell[    3087] = 32'h0;  // 32'h0cf322df;
    ram_cell[    3088] = 32'h0;  // 32'he879453a;
    ram_cell[    3089] = 32'h0;  // 32'hf53ad3b1;
    ram_cell[    3090] = 32'h0;  // 32'h6d550d2b;
    ram_cell[    3091] = 32'h0;  // 32'h4b359807;
    ram_cell[    3092] = 32'h0;  // 32'h7fdc9f41;
    ram_cell[    3093] = 32'h0;  // 32'h331e3702;
    ram_cell[    3094] = 32'h0;  // 32'h6f91d170;
    ram_cell[    3095] = 32'h0;  // 32'hd63af841;
    ram_cell[    3096] = 32'h0;  // 32'h0867edf7;
    ram_cell[    3097] = 32'h0;  // 32'hb66f7618;
    ram_cell[    3098] = 32'h0;  // 32'hc4c3c861;
    ram_cell[    3099] = 32'h0;  // 32'h76a0c802;
    ram_cell[    3100] = 32'h0;  // 32'h48313c62;
    ram_cell[    3101] = 32'h0;  // 32'hcbe3c832;
    ram_cell[    3102] = 32'h0;  // 32'h1e8312cc;
    ram_cell[    3103] = 32'h0;  // 32'h464363b7;
    ram_cell[    3104] = 32'h0;  // 32'h3ddb5387;
    ram_cell[    3105] = 32'h0;  // 32'haeca632a;
    ram_cell[    3106] = 32'h0;  // 32'h5943ddfa;
    ram_cell[    3107] = 32'h0;  // 32'h99d47336;
    ram_cell[    3108] = 32'h0;  // 32'hbd94a7a6;
    ram_cell[    3109] = 32'h0;  // 32'he8226d8a;
    ram_cell[    3110] = 32'h0;  // 32'hbad33402;
    ram_cell[    3111] = 32'h0;  // 32'h1205d940;
    ram_cell[    3112] = 32'h0;  // 32'h14e9a705;
    ram_cell[    3113] = 32'h0;  // 32'hda2a35b2;
    ram_cell[    3114] = 32'h0;  // 32'h19c22740;
    ram_cell[    3115] = 32'h0;  // 32'h7be6f4a4;
    ram_cell[    3116] = 32'h0;  // 32'h83c027e2;
    ram_cell[    3117] = 32'h0;  // 32'h3fb41a6d;
    ram_cell[    3118] = 32'h0;  // 32'h7dace408;
    ram_cell[    3119] = 32'h0;  // 32'h901320bf;
    ram_cell[    3120] = 32'h0;  // 32'h0ef447e3;
    ram_cell[    3121] = 32'h0;  // 32'he69ba8f8;
    ram_cell[    3122] = 32'h0;  // 32'hc81c4e45;
    ram_cell[    3123] = 32'h0;  // 32'hd35185bd;
    ram_cell[    3124] = 32'h0;  // 32'h9d91017c;
    ram_cell[    3125] = 32'h0;  // 32'h92077340;
    ram_cell[    3126] = 32'h0;  // 32'h9b334ec9;
    ram_cell[    3127] = 32'h0;  // 32'h5c0360f3;
    ram_cell[    3128] = 32'h0;  // 32'hdb6f9e97;
    ram_cell[    3129] = 32'h0;  // 32'h8ad0d94a;
    ram_cell[    3130] = 32'h0;  // 32'hcef7030f;
    ram_cell[    3131] = 32'h0;  // 32'h1c8fc97c;
    ram_cell[    3132] = 32'h0;  // 32'hb8ad13e3;
    ram_cell[    3133] = 32'h0;  // 32'hb56f4cc9;
    ram_cell[    3134] = 32'h0;  // 32'h296d6674;
    ram_cell[    3135] = 32'h0;  // 32'hfc5bc2ee;
    ram_cell[    3136] = 32'h0;  // 32'h54a3d086;
    ram_cell[    3137] = 32'h0;  // 32'hebed33e6;
    ram_cell[    3138] = 32'h0;  // 32'hb3155c34;
    ram_cell[    3139] = 32'h0;  // 32'hc3fedd49;
    ram_cell[    3140] = 32'h0;  // 32'hae36d864;
    ram_cell[    3141] = 32'h0;  // 32'heba5503c;
    ram_cell[    3142] = 32'h0;  // 32'h20b05b19;
    ram_cell[    3143] = 32'h0;  // 32'ha96e6dfe;
    ram_cell[    3144] = 32'h0;  // 32'hadc40bb3;
    ram_cell[    3145] = 32'h0;  // 32'he8462b33;
    ram_cell[    3146] = 32'h0;  // 32'h5f59db3a;
    ram_cell[    3147] = 32'h0;  // 32'h9b9067ed;
    ram_cell[    3148] = 32'h0;  // 32'h0b7394ab;
    ram_cell[    3149] = 32'h0;  // 32'h496efbb9;
    ram_cell[    3150] = 32'h0;  // 32'haf8bfbe2;
    ram_cell[    3151] = 32'h0;  // 32'h383d36da;
    ram_cell[    3152] = 32'h0;  // 32'hd9d98781;
    ram_cell[    3153] = 32'h0;  // 32'h7ea0dcf1;
    ram_cell[    3154] = 32'h0;  // 32'h2a2bbed3;
    ram_cell[    3155] = 32'h0;  // 32'he85564da;
    ram_cell[    3156] = 32'h0;  // 32'ha1289106;
    ram_cell[    3157] = 32'h0;  // 32'hb1d9d1d2;
    ram_cell[    3158] = 32'h0;  // 32'h441c3a98;
    ram_cell[    3159] = 32'h0;  // 32'ha7e4756f;
    ram_cell[    3160] = 32'h0;  // 32'h004feede;
    ram_cell[    3161] = 32'h0;  // 32'h3577ff1d;
    ram_cell[    3162] = 32'h0;  // 32'ha3a3b986;
    ram_cell[    3163] = 32'h0;  // 32'h1ddbac66;
    ram_cell[    3164] = 32'h0;  // 32'h9b05456b;
    ram_cell[    3165] = 32'h0;  // 32'hfb03e2e1;
    ram_cell[    3166] = 32'h0;  // 32'h11fdd411;
    ram_cell[    3167] = 32'h0;  // 32'ha9080f80;
    ram_cell[    3168] = 32'h0;  // 32'h1bfe6f02;
    ram_cell[    3169] = 32'h0;  // 32'h34a78fb3;
    ram_cell[    3170] = 32'h0;  // 32'h64799c1b;
    ram_cell[    3171] = 32'h0;  // 32'h799239f8;
    ram_cell[    3172] = 32'h0;  // 32'h9dbafa18;
    ram_cell[    3173] = 32'h0;  // 32'hd42fc91a;
    ram_cell[    3174] = 32'h0;  // 32'hb31e6492;
    ram_cell[    3175] = 32'h0;  // 32'h6c35716b;
    ram_cell[    3176] = 32'h0;  // 32'h6873989c;
    ram_cell[    3177] = 32'h0;  // 32'h776ab452;
    ram_cell[    3178] = 32'h0;  // 32'h0125a964;
    ram_cell[    3179] = 32'h0;  // 32'h369457f9;
    ram_cell[    3180] = 32'h0;  // 32'h13f63daf;
    ram_cell[    3181] = 32'h0;  // 32'hd57fbc2e;
    ram_cell[    3182] = 32'h0;  // 32'hec9a4e18;
    ram_cell[    3183] = 32'h0;  // 32'hf0c06146;
    ram_cell[    3184] = 32'h0;  // 32'h79d9d95d;
    ram_cell[    3185] = 32'h0;  // 32'h40a3edcf;
    ram_cell[    3186] = 32'h0;  // 32'h3f9b2500;
    ram_cell[    3187] = 32'h0;  // 32'hfe70fe1c;
    ram_cell[    3188] = 32'h0;  // 32'hd7a27de3;
    ram_cell[    3189] = 32'h0;  // 32'h2f325e52;
    ram_cell[    3190] = 32'h0;  // 32'h2698cdf2;
    ram_cell[    3191] = 32'h0;  // 32'h341b37d9;
    ram_cell[    3192] = 32'h0;  // 32'h9d9c3a21;
    ram_cell[    3193] = 32'h0;  // 32'h2e177aff;
    ram_cell[    3194] = 32'h0;  // 32'h4b608f19;
    ram_cell[    3195] = 32'h0;  // 32'h56ec1503;
    ram_cell[    3196] = 32'h0;  // 32'h77070298;
    ram_cell[    3197] = 32'h0;  // 32'hf9574a2b;
    ram_cell[    3198] = 32'h0;  // 32'h349bdcae;
    ram_cell[    3199] = 32'h0;  // 32'h751a790a;
    ram_cell[    3200] = 32'h0;  // 32'h34c0e032;
    ram_cell[    3201] = 32'h0;  // 32'h14ba8157;
    ram_cell[    3202] = 32'h0;  // 32'h76ce00da;
    ram_cell[    3203] = 32'h0;  // 32'h697435c9;
    ram_cell[    3204] = 32'h0;  // 32'h4d147b2a;
    ram_cell[    3205] = 32'h0;  // 32'h11abd739;
    ram_cell[    3206] = 32'h0;  // 32'h7d66cc75;
    ram_cell[    3207] = 32'h0;  // 32'h0c87ce8b;
    ram_cell[    3208] = 32'h0;  // 32'hef11381d;
    ram_cell[    3209] = 32'h0;  // 32'h135d9d1a;
    ram_cell[    3210] = 32'h0;  // 32'h99342cac;
    ram_cell[    3211] = 32'h0;  // 32'h08f9217c;
    ram_cell[    3212] = 32'h0;  // 32'h08cca187;
    ram_cell[    3213] = 32'h0;  // 32'hc566fb39;
    ram_cell[    3214] = 32'h0;  // 32'h467c0fae;
    ram_cell[    3215] = 32'h0;  // 32'hfcd7c81e;
    ram_cell[    3216] = 32'h0;  // 32'h77865248;
    ram_cell[    3217] = 32'h0;  // 32'ha61c87a0;
    ram_cell[    3218] = 32'h0;  // 32'h78752969;
    ram_cell[    3219] = 32'h0;  // 32'hca1bd02a;
    ram_cell[    3220] = 32'h0;  // 32'hd63d0069;
    ram_cell[    3221] = 32'h0;  // 32'h85d628a2;
    ram_cell[    3222] = 32'h0;  // 32'hc7c0b03c;
    ram_cell[    3223] = 32'h0;  // 32'hdc603ba9;
    ram_cell[    3224] = 32'h0;  // 32'ha147a1ad;
    ram_cell[    3225] = 32'h0;  // 32'ha542d26f;
    ram_cell[    3226] = 32'h0;  // 32'ha248ddfb;
    ram_cell[    3227] = 32'h0;  // 32'hcc9e13b4;
    ram_cell[    3228] = 32'h0;  // 32'hc3c9e9e4;
    ram_cell[    3229] = 32'h0;  // 32'hf2771a40;
    ram_cell[    3230] = 32'h0;  // 32'hfd0c877a;
    ram_cell[    3231] = 32'h0;  // 32'h439ccdc6;
    ram_cell[    3232] = 32'h0;  // 32'he7f846b0;
    ram_cell[    3233] = 32'h0;  // 32'hb8e7aeae;
    ram_cell[    3234] = 32'h0;  // 32'h38aba4c1;
    ram_cell[    3235] = 32'h0;  // 32'hc4b160f0;
    ram_cell[    3236] = 32'h0;  // 32'h817d0f22;
    ram_cell[    3237] = 32'h0;  // 32'h7711768f;
    ram_cell[    3238] = 32'h0;  // 32'hb60677d2;
    ram_cell[    3239] = 32'h0;  // 32'h9c79075f;
    ram_cell[    3240] = 32'h0;  // 32'h62b8353f;
    ram_cell[    3241] = 32'h0;  // 32'h12709b67;
    ram_cell[    3242] = 32'h0;  // 32'h05f1ce4b;
    ram_cell[    3243] = 32'h0;  // 32'h2fa0afc9;
    ram_cell[    3244] = 32'h0;  // 32'hf8fa35e3;
    ram_cell[    3245] = 32'h0;  // 32'h7dbedb22;
    ram_cell[    3246] = 32'h0;  // 32'hc3e1c5f1;
    ram_cell[    3247] = 32'h0;  // 32'h3cc4225f;
    ram_cell[    3248] = 32'h0;  // 32'he9e7d304;
    ram_cell[    3249] = 32'h0;  // 32'heb79e137;
    ram_cell[    3250] = 32'h0;  // 32'hb549dcf5;
    ram_cell[    3251] = 32'h0;  // 32'he7fdfbf7;
    ram_cell[    3252] = 32'h0;  // 32'h751213d0;
    ram_cell[    3253] = 32'h0;  // 32'hf1571c5b;
    ram_cell[    3254] = 32'h0;  // 32'h678c5442;
    ram_cell[    3255] = 32'h0;  // 32'h5be39122;
    ram_cell[    3256] = 32'h0;  // 32'hc6e945da;
    ram_cell[    3257] = 32'h0;  // 32'hadfe7031;
    ram_cell[    3258] = 32'h0;  // 32'hfb20c81b;
    ram_cell[    3259] = 32'h0;  // 32'h89051e70;
    ram_cell[    3260] = 32'h0;  // 32'hc8a4c0b0;
    ram_cell[    3261] = 32'h0;  // 32'ha14a1857;
    ram_cell[    3262] = 32'h0;  // 32'haaf887d4;
    ram_cell[    3263] = 32'h0;  // 32'h035c234c;
    ram_cell[    3264] = 32'h0;  // 32'h6702a85a;
    ram_cell[    3265] = 32'h0;  // 32'h5e7b25bd;
    ram_cell[    3266] = 32'h0;  // 32'h6143564e;
    ram_cell[    3267] = 32'h0;  // 32'h746b5778;
    ram_cell[    3268] = 32'h0;  // 32'h779175d7;
    ram_cell[    3269] = 32'h0;  // 32'hbe2f230d;
    ram_cell[    3270] = 32'h0;  // 32'hf4bce7cd;
    ram_cell[    3271] = 32'h0;  // 32'h7af6d2c8;
    ram_cell[    3272] = 32'h0;  // 32'hb9086f67;
    ram_cell[    3273] = 32'h0;  // 32'hd353842e;
    ram_cell[    3274] = 32'h0;  // 32'h786a2485;
    ram_cell[    3275] = 32'h0;  // 32'he79a33ef;
    ram_cell[    3276] = 32'h0;  // 32'hc93f219b;
    ram_cell[    3277] = 32'h0;  // 32'he400522b;
    ram_cell[    3278] = 32'h0;  // 32'h3d427c5e;
    ram_cell[    3279] = 32'h0;  // 32'hfd8ce6ac;
    ram_cell[    3280] = 32'h0;  // 32'h45797936;
    ram_cell[    3281] = 32'h0;  // 32'h7e7985fa;
    ram_cell[    3282] = 32'h0;  // 32'h13ad6f02;
    ram_cell[    3283] = 32'h0;  // 32'h4e7614c7;
    ram_cell[    3284] = 32'h0;  // 32'h06d5163c;
    ram_cell[    3285] = 32'h0;  // 32'hbe1305f9;
    ram_cell[    3286] = 32'h0;  // 32'hf856b468;
    ram_cell[    3287] = 32'h0;  // 32'h81e093ab;
    ram_cell[    3288] = 32'h0;  // 32'hdf76defb;
    ram_cell[    3289] = 32'h0;  // 32'h13c331be;
    ram_cell[    3290] = 32'h0;  // 32'h5779b5af;
    ram_cell[    3291] = 32'h0;  // 32'hb6eae942;
    ram_cell[    3292] = 32'h0;  // 32'hab69ee1c;
    ram_cell[    3293] = 32'h0;  // 32'ha7b77dc9;
    ram_cell[    3294] = 32'h0;  // 32'h260a04a2;
    ram_cell[    3295] = 32'h0;  // 32'hf9cf928c;
    ram_cell[    3296] = 32'h0;  // 32'h57f18465;
    ram_cell[    3297] = 32'h0;  // 32'hcea3375f;
    ram_cell[    3298] = 32'h0;  // 32'hee89cf0b;
    ram_cell[    3299] = 32'h0;  // 32'he0bdb3cc;
    ram_cell[    3300] = 32'h0;  // 32'hac190896;
    ram_cell[    3301] = 32'h0;  // 32'h84330b5f;
    ram_cell[    3302] = 32'h0;  // 32'ha10adb5e;
    ram_cell[    3303] = 32'h0;  // 32'h4e70faca;
    ram_cell[    3304] = 32'h0;  // 32'h49734a2b;
    ram_cell[    3305] = 32'h0;  // 32'h5537a193;
    ram_cell[    3306] = 32'h0;  // 32'h573079ae;
    ram_cell[    3307] = 32'h0;  // 32'hfe8547ae;
    ram_cell[    3308] = 32'h0;  // 32'had171be9;
    ram_cell[    3309] = 32'h0;  // 32'h769d7309;
    ram_cell[    3310] = 32'h0;  // 32'h28a95d00;
    ram_cell[    3311] = 32'h0;  // 32'hdaeb5d58;
    ram_cell[    3312] = 32'h0;  // 32'h5c00ec79;
    ram_cell[    3313] = 32'h0;  // 32'h2e2a4a44;
    ram_cell[    3314] = 32'h0;  // 32'h7214d2ee;
    ram_cell[    3315] = 32'h0;  // 32'h9a833421;
    ram_cell[    3316] = 32'h0;  // 32'h2cbc67c3;
    ram_cell[    3317] = 32'h0;  // 32'h99c5e411;
    ram_cell[    3318] = 32'h0;  // 32'h639c14a3;
    ram_cell[    3319] = 32'h0;  // 32'hfbf767b4;
    ram_cell[    3320] = 32'h0;  // 32'ha29b8d76;
    ram_cell[    3321] = 32'h0;  // 32'h95f48305;
    ram_cell[    3322] = 32'h0;  // 32'h3f10196a;
    ram_cell[    3323] = 32'h0;  // 32'h59187bda;
    ram_cell[    3324] = 32'h0;  // 32'haca232de;
    ram_cell[    3325] = 32'h0;  // 32'h46854c1b;
    ram_cell[    3326] = 32'h0;  // 32'hc05b605d;
    ram_cell[    3327] = 32'h0;  // 32'hfa339b75;
    ram_cell[    3328] = 32'h0;  // 32'h0f08e8d6;
    ram_cell[    3329] = 32'h0;  // 32'he5a408e2;
    ram_cell[    3330] = 32'h0;  // 32'h75a9f2f2;
    ram_cell[    3331] = 32'h0;  // 32'h146ce4fa;
    ram_cell[    3332] = 32'h0;  // 32'h3ae5dc52;
    ram_cell[    3333] = 32'h0;  // 32'hc4ced1a9;
    ram_cell[    3334] = 32'h0;  // 32'h1439df00;
    ram_cell[    3335] = 32'h0;  // 32'h7a5e498b;
    ram_cell[    3336] = 32'h0;  // 32'h85d12f90;
    ram_cell[    3337] = 32'h0;  // 32'h68130eb2;
    ram_cell[    3338] = 32'h0;  // 32'h7544c102;
    ram_cell[    3339] = 32'h0;  // 32'h9cca1d4a;
    ram_cell[    3340] = 32'h0;  // 32'h5535f9cc;
    ram_cell[    3341] = 32'h0;  // 32'h19e205f3;
    ram_cell[    3342] = 32'h0;  // 32'h798135d0;
    ram_cell[    3343] = 32'h0;  // 32'h66abd4c5;
    ram_cell[    3344] = 32'h0;  // 32'hb0aa0d2a;
    ram_cell[    3345] = 32'h0;  // 32'h0b1ee7f7;
    ram_cell[    3346] = 32'h0;  // 32'h994f4614;
    ram_cell[    3347] = 32'h0;  // 32'h59520c10;
    ram_cell[    3348] = 32'h0;  // 32'h924e1f08;
    ram_cell[    3349] = 32'h0;  // 32'had65de26;
    ram_cell[    3350] = 32'h0;  // 32'he5dc8bb7;
    ram_cell[    3351] = 32'h0;  // 32'hf66f1521;
    ram_cell[    3352] = 32'h0;  // 32'hb54a3bfe;
    ram_cell[    3353] = 32'h0;  // 32'h787c9b74;
    ram_cell[    3354] = 32'h0;  // 32'h4eb6c318;
    ram_cell[    3355] = 32'h0;  // 32'hc558bb00;
    ram_cell[    3356] = 32'h0;  // 32'h9c9b4262;
    ram_cell[    3357] = 32'h0;  // 32'h74c3ce5f;
    ram_cell[    3358] = 32'h0;  // 32'hf80d146c;
    ram_cell[    3359] = 32'h0;  // 32'h517e7fec;
    ram_cell[    3360] = 32'h0;  // 32'hc1797fd1;
    ram_cell[    3361] = 32'h0;  // 32'h4a1b06f8;
    ram_cell[    3362] = 32'h0;  // 32'h1abfa9f5;
    ram_cell[    3363] = 32'h0;  // 32'hfcbc86e9;
    ram_cell[    3364] = 32'h0;  // 32'h7a5b9fe8;
    ram_cell[    3365] = 32'h0;  // 32'h94c6aaa2;
    ram_cell[    3366] = 32'h0;  // 32'h19df5cf6;
    ram_cell[    3367] = 32'h0;  // 32'hfef5833b;
    ram_cell[    3368] = 32'h0;  // 32'h310799c5;
    ram_cell[    3369] = 32'h0;  // 32'hacc551d0;
    ram_cell[    3370] = 32'h0;  // 32'hf4872a99;
    ram_cell[    3371] = 32'h0;  // 32'h50e6d247;
    ram_cell[    3372] = 32'h0;  // 32'ha6f95a49;
    ram_cell[    3373] = 32'h0;  // 32'h2ace7ba5;
    ram_cell[    3374] = 32'h0;  // 32'h6718eb37;
    ram_cell[    3375] = 32'h0;  // 32'h2b47e77a;
    ram_cell[    3376] = 32'h0;  // 32'h6f268c53;
    ram_cell[    3377] = 32'h0;  // 32'h50a38c2d;
    ram_cell[    3378] = 32'h0;  // 32'h0bcb1aca;
    ram_cell[    3379] = 32'h0;  // 32'h2f8825fb;
    ram_cell[    3380] = 32'h0;  // 32'ha2d59d39;
    ram_cell[    3381] = 32'h0;  // 32'h94e8a5a6;
    ram_cell[    3382] = 32'h0;  // 32'h5130165b;
    ram_cell[    3383] = 32'h0;  // 32'h21301925;
    ram_cell[    3384] = 32'h0;  // 32'h97df2b0a;
    ram_cell[    3385] = 32'h0;  // 32'h74e172d4;
    ram_cell[    3386] = 32'h0;  // 32'h77774f4c;
    ram_cell[    3387] = 32'h0;  // 32'hb6879a04;
    ram_cell[    3388] = 32'h0;  // 32'h70b722d6;
    ram_cell[    3389] = 32'h0;  // 32'h8435a5a3;
    ram_cell[    3390] = 32'h0;  // 32'h73e215cf;
    ram_cell[    3391] = 32'h0;  // 32'ha88494dd;
    ram_cell[    3392] = 32'h0;  // 32'h2e2e8e64;
    ram_cell[    3393] = 32'h0;  // 32'h82f5b239;
    ram_cell[    3394] = 32'h0;  // 32'h043d314e;
    ram_cell[    3395] = 32'h0;  // 32'h4e5987ca;
    ram_cell[    3396] = 32'h0;  // 32'h51289f42;
    ram_cell[    3397] = 32'h0;  // 32'h5c52f14f;
    ram_cell[    3398] = 32'h0;  // 32'he7006137;
    ram_cell[    3399] = 32'h0;  // 32'h44401772;
    ram_cell[    3400] = 32'h0;  // 32'h50be70fb;
    ram_cell[    3401] = 32'h0;  // 32'hdba455b8;
    ram_cell[    3402] = 32'h0;  // 32'hbd3af496;
    ram_cell[    3403] = 32'h0;  // 32'h6f3d7952;
    ram_cell[    3404] = 32'h0;  // 32'h959b0ad6;
    ram_cell[    3405] = 32'h0;  // 32'he84355be;
    ram_cell[    3406] = 32'h0;  // 32'hd5f938d8;
    ram_cell[    3407] = 32'h0;  // 32'h0d24ebbd;
    ram_cell[    3408] = 32'h0;  // 32'he44a34e5;
    ram_cell[    3409] = 32'h0;  // 32'h9ce4ac5c;
    ram_cell[    3410] = 32'h0;  // 32'h24fab819;
    ram_cell[    3411] = 32'h0;  // 32'h60a21aa1;
    ram_cell[    3412] = 32'h0;  // 32'hc2b00d5a;
    ram_cell[    3413] = 32'h0;  // 32'h787eee59;
    ram_cell[    3414] = 32'h0;  // 32'hdd9ac00c;
    ram_cell[    3415] = 32'h0;  // 32'h2e81c33d;
    ram_cell[    3416] = 32'h0;  // 32'hef5d00a8;
    ram_cell[    3417] = 32'h0;  // 32'h43a9f6d4;
    ram_cell[    3418] = 32'h0;  // 32'heee5066c;
    ram_cell[    3419] = 32'h0;  // 32'h00d1096d;
    ram_cell[    3420] = 32'h0;  // 32'h2a4e0f32;
    ram_cell[    3421] = 32'h0;  // 32'h84fe1cee;
    ram_cell[    3422] = 32'h0;  // 32'h18c4912a;
    ram_cell[    3423] = 32'h0;  // 32'h2cc43b43;
    ram_cell[    3424] = 32'h0;  // 32'h5ace8922;
    ram_cell[    3425] = 32'h0;  // 32'hed1b53ca;
    ram_cell[    3426] = 32'h0;  // 32'h36647bd6;
    ram_cell[    3427] = 32'h0;  // 32'h3db24a91;
    ram_cell[    3428] = 32'h0;  // 32'h807bb21b;
    ram_cell[    3429] = 32'h0;  // 32'h69e02900;
    ram_cell[    3430] = 32'h0;  // 32'hd7865625;
    ram_cell[    3431] = 32'h0;  // 32'h79833daa;
    ram_cell[    3432] = 32'h0;  // 32'h7361d0e1;
    ram_cell[    3433] = 32'h0;  // 32'hd5091b31;
    ram_cell[    3434] = 32'h0;  // 32'h9ecb41b9;
    ram_cell[    3435] = 32'h0;  // 32'h8a51e695;
    ram_cell[    3436] = 32'h0;  // 32'h95eb8871;
    ram_cell[    3437] = 32'h0;  // 32'h3defd4db;
    ram_cell[    3438] = 32'h0;  // 32'heee4a2b2;
    ram_cell[    3439] = 32'h0;  // 32'h6182ce96;
    ram_cell[    3440] = 32'h0;  // 32'hba3ed6e2;
    ram_cell[    3441] = 32'h0;  // 32'h00941e76;
    ram_cell[    3442] = 32'h0;  // 32'h3099d962;
    ram_cell[    3443] = 32'h0;  // 32'h4a27289a;
    ram_cell[    3444] = 32'h0;  // 32'h490bde9a;
    ram_cell[    3445] = 32'h0;  // 32'hac249b78;
    ram_cell[    3446] = 32'h0;  // 32'hb1b0a885;
    ram_cell[    3447] = 32'h0;  // 32'hbec1d40f;
    ram_cell[    3448] = 32'h0;  // 32'h926a8b7a;
    ram_cell[    3449] = 32'h0;  // 32'h2ab0da8e;
    ram_cell[    3450] = 32'h0;  // 32'haa7ee8e0;
    ram_cell[    3451] = 32'h0;  // 32'h78cd140a;
    ram_cell[    3452] = 32'h0;  // 32'h938b7e8c;
    ram_cell[    3453] = 32'h0;  // 32'h07b5dfc6;
    ram_cell[    3454] = 32'h0;  // 32'h2a9c9000;
    ram_cell[    3455] = 32'h0;  // 32'h865fa394;
    ram_cell[    3456] = 32'h0;  // 32'he16a142d;
    ram_cell[    3457] = 32'h0;  // 32'h3b9594fd;
    ram_cell[    3458] = 32'h0;  // 32'hab647366;
    ram_cell[    3459] = 32'h0;  // 32'h4492d160;
    ram_cell[    3460] = 32'h0;  // 32'h324b3391;
    ram_cell[    3461] = 32'h0;  // 32'h1437041e;
    ram_cell[    3462] = 32'h0;  // 32'h9f94a1fa;
    ram_cell[    3463] = 32'h0;  // 32'hb9b7c9ee;
    ram_cell[    3464] = 32'h0;  // 32'h2b8a5314;
    ram_cell[    3465] = 32'h0;  // 32'hab059162;
    ram_cell[    3466] = 32'h0;  // 32'hc30a40e8;
    ram_cell[    3467] = 32'h0;  // 32'h0fda4556;
    ram_cell[    3468] = 32'h0;  // 32'h5c4233a1;
    ram_cell[    3469] = 32'h0;  // 32'h312b5027;
    ram_cell[    3470] = 32'h0;  // 32'h7236c5fd;
    ram_cell[    3471] = 32'h0;  // 32'h3be2f526;
    ram_cell[    3472] = 32'h0;  // 32'h6b5e16ad;
    ram_cell[    3473] = 32'h0;  // 32'hab0e9f46;
    ram_cell[    3474] = 32'h0;  // 32'h4f1bc13d;
    ram_cell[    3475] = 32'h0;  // 32'ha266f178;
    ram_cell[    3476] = 32'h0;  // 32'hc7f8fb0e;
    ram_cell[    3477] = 32'h0;  // 32'h6a4791f5;
    ram_cell[    3478] = 32'h0;  // 32'hf934bf53;
    ram_cell[    3479] = 32'h0;  // 32'h7c809789;
    ram_cell[    3480] = 32'h0;  // 32'h4ddfef41;
    ram_cell[    3481] = 32'h0;  // 32'h9de3cbc2;
    ram_cell[    3482] = 32'h0;  // 32'h7f86b3ee;
    ram_cell[    3483] = 32'h0;  // 32'h01998d17;
    ram_cell[    3484] = 32'h0;  // 32'h38cd36ad;
    ram_cell[    3485] = 32'h0;  // 32'hc30bb043;
    ram_cell[    3486] = 32'h0;  // 32'h6ff36f1d;
    ram_cell[    3487] = 32'h0;  // 32'h90b47f57;
    ram_cell[    3488] = 32'h0;  // 32'h1e146f2c;
    ram_cell[    3489] = 32'h0;  // 32'h34676038;
    ram_cell[    3490] = 32'h0;  // 32'hf8489780;
    ram_cell[    3491] = 32'h0;  // 32'hc3bcd6ad;
    ram_cell[    3492] = 32'h0;  // 32'h602f1c84;
    ram_cell[    3493] = 32'h0;  // 32'h0054d59d;
    ram_cell[    3494] = 32'h0;  // 32'hec2e1a1d;
    ram_cell[    3495] = 32'h0;  // 32'h1dd8552f;
    ram_cell[    3496] = 32'h0;  // 32'hc01df45e;
    ram_cell[    3497] = 32'h0;  // 32'h96d8af36;
    ram_cell[    3498] = 32'h0;  // 32'h1152aa9e;
    ram_cell[    3499] = 32'h0;  // 32'h8736a125;
    ram_cell[    3500] = 32'h0;  // 32'hf00a148b;
    ram_cell[    3501] = 32'h0;  // 32'hc673efe3;
    ram_cell[    3502] = 32'h0;  // 32'hc708c4de;
    ram_cell[    3503] = 32'h0;  // 32'h38be2d09;
    ram_cell[    3504] = 32'h0;  // 32'hf682791d;
    ram_cell[    3505] = 32'h0;  // 32'h9b277242;
    ram_cell[    3506] = 32'h0;  // 32'hf9aebf0f;
    ram_cell[    3507] = 32'h0;  // 32'h84b16180;
    ram_cell[    3508] = 32'h0;  // 32'hb37d7a7e;
    ram_cell[    3509] = 32'h0;  // 32'h59747e21;
    ram_cell[    3510] = 32'h0;  // 32'h43105001;
    ram_cell[    3511] = 32'h0;  // 32'h7b297f7d;
    ram_cell[    3512] = 32'h0;  // 32'hfe29982f;
    ram_cell[    3513] = 32'h0;  // 32'h651e1377;
    ram_cell[    3514] = 32'h0;  // 32'heae0f52d;
    ram_cell[    3515] = 32'h0;  // 32'h583b5143;
    ram_cell[    3516] = 32'h0;  // 32'hb3689161;
    ram_cell[    3517] = 32'h0;  // 32'h6dbac6a1;
    ram_cell[    3518] = 32'h0;  // 32'hed1f80b9;
    ram_cell[    3519] = 32'h0;  // 32'h46ef536c;
    ram_cell[    3520] = 32'h0;  // 32'h9dd04fae;
    ram_cell[    3521] = 32'h0;  // 32'h4d7851e2;
    ram_cell[    3522] = 32'h0;  // 32'h7165be92;
    ram_cell[    3523] = 32'h0;  // 32'h725da9c9;
    ram_cell[    3524] = 32'h0;  // 32'h800d4bf8;
    ram_cell[    3525] = 32'h0;  // 32'h7e532a9b;
    ram_cell[    3526] = 32'h0;  // 32'hedc3fffc;
    ram_cell[    3527] = 32'h0;  // 32'h4f7781de;
    ram_cell[    3528] = 32'h0;  // 32'he6dc4e69;
    ram_cell[    3529] = 32'h0;  // 32'h2dc237f9;
    ram_cell[    3530] = 32'h0;  // 32'h10000518;
    ram_cell[    3531] = 32'h0;  // 32'hf50cea77;
    ram_cell[    3532] = 32'h0;  // 32'h2c05d927;
    ram_cell[    3533] = 32'h0;  // 32'h10396ace;
    ram_cell[    3534] = 32'h0;  // 32'hdf119550;
    ram_cell[    3535] = 32'h0;  // 32'hf3a2d0aa;
    ram_cell[    3536] = 32'h0;  // 32'h1f40204e;
    ram_cell[    3537] = 32'h0;  // 32'h88f3916b;
    ram_cell[    3538] = 32'h0;  // 32'h608346c3;
    ram_cell[    3539] = 32'h0;  // 32'h2808e124;
    ram_cell[    3540] = 32'h0;  // 32'heca55cf6;
    ram_cell[    3541] = 32'h0;  // 32'he6f42fa0;
    ram_cell[    3542] = 32'h0;  // 32'h3ee2ee7d;
    ram_cell[    3543] = 32'h0;  // 32'h20a8e7c3;
    ram_cell[    3544] = 32'h0;  // 32'h6b0f5e8e;
    ram_cell[    3545] = 32'h0;  // 32'h25b40807;
    ram_cell[    3546] = 32'h0;  // 32'h37ece0bd;
    ram_cell[    3547] = 32'h0;  // 32'h7f95449d;
    ram_cell[    3548] = 32'h0;  // 32'hf440087e;
    ram_cell[    3549] = 32'h0;  // 32'hf7be3f22;
    ram_cell[    3550] = 32'h0;  // 32'he40ef317;
    ram_cell[    3551] = 32'h0;  // 32'h0d4fb0af;
    ram_cell[    3552] = 32'h0;  // 32'h35d452ed;
    ram_cell[    3553] = 32'h0;  // 32'h61daa056;
    ram_cell[    3554] = 32'h0;  // 32'h9aca330e;
    ram_cell[    3555] = 32'h0;  // 32'h1bdb57e3;
    ram_cell[    3556] = 32'h0;  // 32'hb8a598db;
    ram_cell[    3557] = 32'h0;  // 32'h4fe48704;
    ram_cell[    3558] = 32'h0;  // 32'hf15f3ff0;
    ram_cell[    3559] = 32'h0;  // 32'haf58af56;
    ram_cell[    3560] = 32'h0;  // 32'hbfb76a52;
    ram_cell[    3561] = 32'h0;  // 32'hd37b2cea;
    ram_cell[    3562] = 32'h0;  // 32'hea1b6831;
    ram_cell[    3563] = 32'h0;  // 32'h3b2f2046;
    ram_cell[    3564] = 32'h0;  // 32'h54bb434c;
    ram_cell[    3565] = 32'h0;  // 32'hc4d6baab;
    ram_cell[    3566] = 32'h0;  // 32'hb0301be8;
    ram_cell[    3567] = 32'h0;  // 32'h03d0c91e;
    ram_cell[    3568] = 32'h0;  // 32'h4d0eee63;
    ram_cell[    3569] = 32'h0;  // 32'hee87dae9;
    ram_cell[    3570] = 32'h0;  // 32'ha4c8ae37;
    ram_cell[    3571] = 32'h0;  // 32'h1e8dee93;
    ram_cell[    3572] = 32'h0;  // 32'h979be43f;
    ram_cell[    3573] = 32'h0;  // 32'h8cc7fceb;
    ram_cell[    3574] = 32'h0;  // 32'h78239d9c;
    ram_cell[    3575] = 32'h0;  // 32'h5a2f4a2e;
    ram_cell[    3576] = 32'h0;  // 32'hb90c4b77;
    ram_cell[    3577] = 32'h0;  // 32'hdb9eb78b;
    ram_cell[    3578] = 32'h0;  // 32'h733e9206;
    ram_cell[    3579] = 32'h0;  // 32'heb24355f;
    ram_cell[    3580] = 32'h0;  // 32'h2aee1750;
    ram_cell[    3581] = 32'h0;  // 32'ha006e4b9;
    ram_cell[    3582] = 32'h0;  // 32'h29caaf28;
    ram_cell[    3583] = 32'h0;  // 32'h38a413fb;
    ram_cell[    3584] = 32'h0;  // 32'h16beb31d;
    ram_cell[    3585] = 32'h0;  // 32'hf8fd5be3;
    ram_cell[    3586] = 32'h0;  // 32'h97186f01;
    ram_cell[    3587] = 32'h0;  // 32'h953d7ffb;
    ram_cell[    3588] = 32'h0;  // 32'hc56742a1;
    ram_cell[    3589] = 32'h0;  // 32'h868fc63c;
    ram_cell[    3590] = 32'h0;  // 32'h0f707a17;
    ram_cell[    3591] = 32'h0;  // 32'h3aa359c8;
    ram_cell[    3592] = 32'h0;  // 32'h754172fc;
    ram_cell[    3593] = 32'h0;  // 32'ha77fe6b3;
    ram_cell[    3594] = 32'h0;  // 32'hdb0d9a77;
    ram_cell[    3595] = 32'h0;  // 32'hf5de675d;
    ram_cell[    3596] = 32'h0;  // 32'hd1113730;
    ram_cell[    3597] = 32'h0;  // 32'h6d0aae41;
    ram_cell[    3598] = 32'h0;  // 32'h4250d5d1;
    ram_cell[    3599] = 32'h0;  // 32'h8678a27f;
    ram_cell[    3600] = 32'h0;  // 32'h973e663c;
    ram_cell[    3601] = 32'h0;  // 32'h820c9383;
    ram_cell[    3602] = 32'h0;  // 32'hbaaa6cc4;
    ram_cell[    3603] = 32'h0;  // 32'hc4f3f512;
    ram_cell[    3604] = 32'h0;  // 32'h797a5ef6;
    ram_cell[    3605] = 32'h0;  // 32'h89a9638b;
    ram_cell[    3606] = 32'h0;  // 32'h8c1866e2;
    ram_cell[    3607] = 32'h0;  // 32'h7303b920;
    ram_cell[    3608] = 32'h0;  // 32'h79872940;
    ram_cell[    3609] = 32'h0;  // 32'h09f7c314;
    ram_cell[    3610] = 32'h0;  // 32'h1314bd8d;
    ram_cell[    3611] = 32'h0;  // 32'hd13aa1ee;
    ram_cell[    3612] = 32'h0;  // 32'hd49db33f;
    ram_cell[    3613] = 32'h0;  // 32'h3e69ea03;
    ram_cell[    3614] = 32'h0;  // 32'hf90699c2;
    ram_cell[    3615] = 32'h0;  // 32'h32fa787c;
    ram_cell[    3616] = 32'h0;  // 32'h98a6f4f3;
    ram_cell[    3617] = 32'h0;  // 32'h31a5e14f;
    ram_cell[    3618] = 32'h0;  // 32'h8f1b4ed5;
    ram_cell[    3619] = 32'h0;  // 32'h625fe8af;
    ram_cell[    3620] = 32'h0;  // 32'hf05ac579;
    ram_cell[    3621] = 32'h0;  // 32'h763f503d;
    ram_cell[    3622] = 32'h0;  // 32'hc423d143;
    ram_cell[    3623] = 32'h0;  // 32'hb526810f;
    ram_cell[    3624] = 32'h0;  // 32'he14fe3b5;
    ram_cell[    3625] = 32'h0;  // 32'h5fc1849b;
    ram_cell[    3626] = 32'h0;  // 32'hcbe4556c;
    ram_cell[    3627] = 32'h0;  // 32'hf04d9f81;
    ram_cell[    3628] = 32'h0;  // 32'h9564ea38;
    ram_cell[    3629] = 32'h0;  // 32'h814882b2;
    ram_cell[    3630] = 32'h0;  // 32'h524bb11d;
    ram_cell[    3631] = 32'h0;  // 32'h9feef0f6;
    ram_cell[    3632] = 32'h0;  // 32'h70660f0a;
    ram_cell[    3633] = 32'h0;  // 32'h02788395;
    ram_cell[    3634] = 32'h0;  // 32'h1a348972;
    ram_cell[    3635] = 32'h0;  // 32'habd94b9a;
    ram_cell[    3636] = 32'h0;  // 32'hcc4771d5;
    ram_cell[    3637] = 32'h0;  // 32'h00d0f3f6;
    ram_cell[    3638] = 32'h0;  // 32'h64d55001;
    ram_cell[    3639] = 32'h0;  // 32'h6ec0cf9f;
    ram_cell[    3640] = 32'h0;  // 32'h61aaebe7;
    ram_cell[    3641] = 32'h0;  // 32'hbcf2261b;
    ram_cell[    3642] = 32'h0;  // 32'hd44d16b1;
    ram_cell[    3643] = 32'h0;  // 32'heee11d1f;
    ram_cell[    3644] = 32'h0;  // 32'h559a23bf;
    ram_cell[    3645] = 32'h0;  // 32'h8dc7ea9b;
    ram_cell[    3646] = 32'h0;  // 32'h6f96436f;
    ram_cell[    3647] = 32'h0;  // 32'h21cd11fa;
    ram_cell[    3648] = 32'h0;  // 32'h5ec350a6;
    ram_cell[    3649] = 32'h0;  // 32'hfdc444a1;
    ram_cell[    3650] = 32'h0;  // 32'h520c684c;
    ram_cell[    3651] = 32'h0;  // 32'h494f9168;
    ram_cell[    3652] = 32'h0;  // 32'h714abb17;
    ram_cell[    3653] = 32'h0;  // 32'hd971efe5;
    ram_cell[    3654] = 32'h0;  // 32'h3e8ce752;
    ram_cell[    3655] = 32'h0;  // 32'hded63318;
    ram_cell[    3656] = 32'h0;  // 32'h752bd77a;
    ram_cell[    3657] = 32'h0;  // 32'hd169496d;
    ram_cell[    3658] = 32'h0;  // 32'h7b9fe8f9;
    ram_cell[    3659] = 32'h0;  // 32'ha42d81be;
    ram_cell[    3660] = 32'h0;  // 32'h06bc2357;
    ram_cell[    3661] = 32'h0;  // 32'haf372d4d;
    ram_cell[    3662] = 32'h0;  // 32'hfb785549;
    ram_cell[    3663] = 32'h0;  // 32'h20420485;
    ram_cell[    3664] = 32'h0;  // 32'hf82e6f46;
    ram_cell[    3665] = 32'h0;  // 32'h6fd91b88;
    ram_cell[    3666] = 32'h0;  // 32'hbd5d9ec3;
    ram_cell[    3667] = 32'h0;  // 32'ha6f73608;
    ram_cell[    3668] = 32'h0;  // 32'h03f28b92;
    ram_cell[    3669] = 32'h0;  // 32'h3d0ac6d4;
    ram_cell[    3670] = 32'h0;  // 32'h6aee5983;
    ram_cell[    3671] = 32'h0;  // 32'h191047eb;
    ram_cell[    3672] = 32'h0;  // 32'h64e121b7;
    ram_cell[    3673] = 32'h0;  // 32'h9c52cc24;
    ram_cell[    3674] = 32'h0;  // 32'h602213a6;
    ram_cell[    3675] = 32'h0;  // 32'he5e19f9a;
    ram_cell[    3676] = 32'h0;  // 32'h80ceb3e2;
    ram_cell[    3677] = 32'h0;  // 32'h19b2cf90;
    ram_cell[    3678] = 32'h0;  // 32'h5d58c417;
    ram_cell[    3679] = 32'h0;  // 32'hc86339f0;
    ram_cell[    3680] = 32'h0;  // 32'h0f421122;
    ram_cell[    3681] = 32'h0;  // 32'h8c0f74f0;
    ram_cell[    3682] = 32'h0;  // 32'h341b1b09;
    ram_cell[    3683] = 32'h0;  // 32'h08da9802;
    ram_cell[    3684] = 32'h0;  // 32'h13e5c7f2;
    ram_cell[    3685] = 32'h0;  // 32'hecf69782;
    ram_cell[    3686] = 32'h0;  // 32'hf929b5fb;
    ram_cell[    3687] = 32'h0;  // 32'h21e39a04;
    ram_cell[    3688] = 32'h0;  // 32'h64be7c70;
    ram_cell[    3689] = 32'h0;  // 32'hc4381927;
    ram_cell[    3690] = 32'h0;  // 32'h4aa95590;
    ram_cell[    3691] = 32'h0;  // 32'h66145f8d;
    ram_cell[    3692] = 32'h0;  // 32'h57264c8f;
    ram_cell[    3693] = 32'h0;  // 32'hfd1909ba;
    ram_cell[    3694] = 32'h0;  // 32'he3157de7;
    ram_cell[    3695] = 32'h0;  // 32'heb605b6f;
    ram_cell[    3696] = 32'h0;  // 32'h27dd172b;
    ram_cell[    3697] = 32'h0;  // 32'hed1c079c;
    ram_cell[    3698] = 32'h0;  // 32'h203fcf15;
    ram_cell[    3699] = 32'h0;  // 32'h4f8b5f12;
    ram_cell[    3700] = 32'h0;  // 32'hd72ed678;
    ram_cell[    3701] = 32'h0;  // 32'h7ceefe1d;
    ram_cell[    3702] = 32'h0;  // 32'h7965c164;
    ram_cell[    3703] = 32'h0;  // 32'h84374940;
    ram_cell[    3704] = 32'h0;  // 32'h4a1c039e;
    ram_cell[    3705] = 32'h0;  // 32'h1df72664;
    ram_cell[    3706] = 32'h0;  // 32'h12ca8b41;
    ram_cell[    3707] = 32'h0;  // 32'hb0e7cec0;
    ram_cell[    3708] = 32'h0;  // 32'ha6801d8f;
    ram_cell[    3709] = 32'h0;  // 32'h4c21eb8d;
    ram_cell[    3710] = 32'h0;  // 32'hbfdb059b;
    ram_cell[    3711] = 32'h0;  // 32'h81891729;
    ram_cell[    3712] = 32'h0;  // 32'hf96be5c9;
    ram_cell[    3713] = 32'h0;  // 32'h3ca96b7a;
    ram_cell[    3714] = 32'h0;  // 32'h12be1823;
    ram_cell[    3715] = 32'h0;  // 32'h0bc8bfde;
    ram_cell[    3716] = 32'h0;  // 32'h654cc430;
    ram_cell[    3717] = 32'h0;  // 32'heb4e60e0;
    ram_cell[    3718] = 32'h0;  // 32'h140087a0;
    ram_cell[    3719] = 32'h0;  // 32'hd447f65a;
    ram_cell[    3720] = 32'h0;  // 32'h4263a33c;
    ram_cell[    3721] = 32'h0;  // 32'h5d794b16;
    ram_cell[    3722] = 32'h0;  // 32'he8910196;
    ram_cell[    3723] = 32'h0;  // 32'h94dbd388;
    ram_cell[    3724] = 32'h0;  // 32'he49a6f80;
    ram_cell[    3725] = 32'h0;  // 32'hf7cb2177;
    ram_cell[    3726] = 32'h0;  // 32'h0b9efbe3;
    ram_cell[    3727] = 32'h0;  // 32'hb5fb39cc;
    ram_cell[    3728] = 32'h0;  // 32'h1c35f303;
    ram_cell[    3729] = 32'h0;  // 32'hb7f2fec3;
    ram_cell[    3730] = 32'h0;  // 32'hfa7fae0c;
    ram_cell[    3731] = 32'h0;  // 32'h7eef82b1;
    ram_cell[    3732] = 32'h0;  // 32'h555ef38d;
    ram_cell[    3733] = 32'h0;  // 32'hac62b3be;
    ram_cell[    3734] = 32'h0;  // 32'hc4f2db02;
    ram_cell[    3735] = 32'h0;  // 32'h55ad7874;
    ram_cell[    3736] = 32'h0;  // 32'h5c86e610;
    ram_cell[    3737] = 32'h0;  // 32'h30c95790;
    ram_cell[    3738] = 32'h0;  // 32'h9a02152e;
    ram_cell[    3739] = 32'h0;  // 32'h86555149;
    ram_cell[    3740] = 32'h0;  // 32'hf335da6f;
    ram_cell[    3741] = 32'h0;  // 32'hf071ed18;
    ram_cell[    3742] = 32'h0;  // 32'h496663b2;
    ram_cell[    3743] = 32'h0;  // 32'h933f1f96;
    ram_cell[    3744] = 32'h0;  // 32'h614972f9;
    ram_cell[    3745] = 32'h0;  // 32'hb0ab4256;
    ram_cell[    3746] = 32'h0;  // 32'h6c76799c;
    ram_cell[    3747] = 32'h0;  // 32'h06d3669c;
    ram_cell[    3748] = 32'h0;  // 32'h23cc77f6;
    ram_cell[    3749] = 32'h0;  // 32'hd51d9086;
    ram_cell[    3750] = 32'h0;  // 32'hf0f6959f;
    ram_cell[    3751] = 32'h0;  // 32'h44b0a04c;
    ram_cell[    3752] = 32'h0;  // 32'h75bcfe6b;
    ram_cell[    3753] = 32'h0;  // 32'heb09cdb8;
    ram_cell[    3754] = 32'h0;  // 32'h5c153bf7;
    ram_cell[    3755] = 32'h0;  // 32'h98c027bb;
    ram_cell[    3756] = 32'h0;  // 32'h0e4317eb;
    ram_cell[    3757] = 32'h0;  // 32'h7c99884c;
    ram_cell[    3758] = 32'h0;  // 32'heeadf4eb;
    ram_cell[    3759] = 32'h0;  // 32'h06700299;
    ram_cell[    3760] = 32'h0;  // 32'h55cfd17d;
    ram_cell[    3761] = 32'h0;  // 32'h88d31036;
    ram_cell[    3762] = 32'h0;  // 32'h0128e9d6;
    ram_cell[    3763] = 32'h0;  // 32'h3f388368;
    ram_cell[    3764] = 32'h0;  // 32'h7d09edcd;
    ram_cell[    3765] = 32'h0;  // 32'h03ccdb1c;
    ram_cell[    3766] = 32'h0;  // 32'h6fc0b2d8;
    ram_cell[    3767] = 32'h0;  // 32'h78e74c4e;
    ram_cell[    3768] = 32'h0;  // 32'hecf3217a;
    ram_cell[    3769] = 32'h0;  // 32'he07d189a;
    ram_cell[    3770] = 32'h0;  // 32'h78cad052;
    ram_cell[    3771] = 32'h0;  // 32'h8b2550da;
    ram_cell[    3772] = 32'h0;  // 32'h758b24de;
    ram_cell[    3773] = 32'h0;  // 32'h39243c04;
    ram_cell[    3774] = 32'h0;  // 32'h1335a278;
    ram_cell[    3775] = 32'h0;  // 32'h2a5dde93;
    ram_cell[    3776] = 32'h0;  // 32'h3931d047;
    ram_cell[    3777] = 32'h0;  // 32'h04d15a71;
    ram_cell[    3778] = 32'h0;  // 32'h03102279;
    ram_cell[    3779] = 32'h0;  // 32'h59fd279f;
    ram_cell[    3780] = 32'h0;  // 32'h4f3d41ff;
    ram_cell[    3781] = 32'h0;  // 32'h78b7444a;
    ram_cell[    3782] = 32'h0;  // 32'h6ec37031;
    ram_cell[    3783] = 32'h0;  // 32'h5da6983a;
    ram_cell[    3784] = 32'h0;  // 32'h086ad4dd;
    ram_cell[    3785] = 32'h0;  // 32'h1d335d5a;
    ram_cell[    3786] = 32'h0;  // 32'ha960e04b;
    ram_cell[    3787] = 32'h0;  // 32'h755be199;
    ram_cell[    3788] = 32'h0;  // 32'hccddee6f;
    ram_cell[    3789] = 32'h0;  // 32'h5f848a39;
    ram_cell[    3790] = 32'h0;  // 32'hac4d3e9f;
    ram_cell[    3791] = 32'h0;  // 32'h716e4a30;
    ram_cell[    3792] = 32'h0;  // 32'h5affb3a7;
    ram_cell[    3793] = 32'h0;  // 32'hc3ef0819;
    ram_cell[    3794] = 32'h0;  // 32'hae7bba4d;
    ram_cell[    3795] = 32'h0;  // 32'h4177d5c8;
    ram_cell[    3796] = 32'h0;  // 32'hdaf4e1c5;
    ram_cell[    3797] = 32'h0;  // 32'hcc19e183;
    ram_cell[    3798] = 32'h0;  // 32'hacaa9543;
    ram_cell[    3799] = 32'h0;  // 32'he0efcb8c;
    ram_cell[    3800] = 32'h0;  // 32'ha746fb42;
    ram_cell[    3801] = 32'h0;  // 32'h4c506158;
    ram_cell[    3802] = 32'h0;  // 32'ha1353b1b;
    ram_cell[    3803] = 32'h0;  // 32'h949137a1;
    ram_cell[    3804] = 32'h0;  // 32'h1db686e5;
    ram_cell[    3805] = 32'h0;  // 32'h05fe2cb1;
    ram_cell[    3806] = 32'h0;  // 32'h5bf3f495;
    ram_cell[    3807] = 32'h0;  // 32'h3757c756;
    ram_cell[    3808] = 32'h0;  // 32'h66308a95;
    ram_cell[    3809] = 32'h0;  // 32'ha3d0297b;
    ram_cell[    3810] = 32'h0;  // 32'h174dcdbb;
    ram_cell[    3811] = 32'h0;  // 32'h96d88081;
    ram_cell[    3812] = 32'h0;  // 32'h0e3fb73a;
    ram_cell[    3813] = 32'h0;  // 32'h7d028a3c;
    ram_cell[    3814] = 32'h0;  // 32'h985e1426;
    ram_cell[    3815] = 32'h0;  // 32'hd05c19af;
    ram_cell[    3816] = 32'h0;  // 32'ha1c28e52;
    ram_cell[    3817] = 32'h0;  // 32'h4510d215;
    ram_cell[    3818] = 32'h0;  // 32'h1bb2adae;
    ram_cell[    3819] = 32'h0;  // 32'ha40c5394;
    ram_cell[    3820] = 32'h0;  // 32'h30c5b70a;
    ram_cell[    3821] = 32'h0;  // 32'h950dc16e;
    ram_cell[    3822] = 32'h0;  // 32'hb0c95b08;
    ram_cell[    3823] = 32'h0;  // 32'h7876d2fd;
    ram_cell[    3824] = 32'h0;  // 32'h8ccaee39;
    ram_cell[    3825] = 32'h0;  // 32'ha3d64f45;
    ram_cell[    3826] = 32'h0;  // 32'ha3cad2b0;
    ram_cell[    3827] = 32'h0;  // 32'h1dcea258;
    ram_cell[    3828] = 32'h0;  // 32'h4af3e318;
    ram_cell[    3829] = 32'h0;  // 32'ha36f13e9;
    ram_cell[    3830] = 32'h0;  // 32'hf01d2d7a;
    ram_cell[    3831] = 32'h0;  // 32'hc4e0b4e0;
    ram_cell[    3832] = 32'h0;  // 32'h04822304;
    ram_cell[    3833] = 32'h0;  // 32'h5eb6d6c1;
    ram_cell[    3834] = 32'h0;  // 32'h02cc2d2c;
    ram_cell[    3835] = 32'h0;  // 32'hf605f40b;
    ram_cell[    3836] = 32'h0;  // 32'h3fed6664;
    ram_cell[    3837] = 32'h0;  // 32'hc9633c73;
    ram_cell[    3838] = 32'h0;  // 32'h8af1de1c;
    ram_cell[    3839] = 32'h0;  // 32'hec1324b9;
    ram_cell[    3840] = 32'h0;  // 32'h948df5fb;
    ram_cell[    3841] = 32'h0;  // 32'h97d2dff0;
    ram_cell[    3842] = 32'h0;  // 32'hf4384e2b;
    ram_cell[    3843] = 32'h0;  // 32'hde903226;
    ram_cell[    3844] = 32'h0;  // 32'he294f744;
    ram_cell[    3845] = 32'h0;  // 32'h6429f154;
    ram_cell[    3846] = 32'h0;  // 32'he47d65ca;
    ram_cell[    3847] = 32'h0;  // 32'h6da048c9;
    ram_cell[    3848] = 32'h0;  // 32'h4723ed8b;
    ram_cell[    3849] = 32'h0;  // 32'hbe6a2cae;
    ram_cell[    3850] = 32'h0;  // 32'h6ebbbca1;
    ram_cell[    3851] = 32'h0;  // 32'h79a0307a;
    ram_cell[    3852] = 32'h0;  // 32'h22642392;
    ram_cell[    3853] = 32'h0;  // 32'h07832a06;
    ram_cell[    3854] = 32'h0;  // 32'hb40765cc;
    ram_cell[    3855] = 32'h0;  // 32'hda9ab92a;
    ram_cell[    3856] = 32'h0;  // 32'h18109600;
    ram_cell[    3857] = 32'h0;  // 32'h7c6aad16;
    ram_cell[    3858] = 32'h0;  // 32'h76002dcc;
    ram_cell[    3859] = 32'h0;  // 32'h4142d32b;
    ram_cell[    3860] = 32'h0;  // 32'h8a39f1ca;
    ram_cell[    3861] = 32'h0;  // 32'h8b465301;
    ram_cell[    3862] = 32'h0;  // 32'h91548080;
    ram_cell[    3863] = 32'h0;  // 32'he46698eb;
    ram_cell[    3864] = 32'h0;  // 32'h68b58e5d;
    ram_cell[    3865] = 32'h0;  // 32'h9407dd8a;
    ram_cell[    3866] = 32'h0;  // 32'h77b613f5;
    ram_cell[    3867] = 32'h0;  // 32'h46b87cf4;
    ram_cell[    3868] = 32'h0;  // 32'h26dbcf41;
    ram_cell[    3869] = 32'h0;  // 32'h4cfde0a4;
    ram_cell[    3870] = 32'h0;  // 32'h06c1d14d;
    ram_cell[    3871] = 32'h0;  // 32'hb8246eef;
    ram_cell[    3872] = 32'h0;  // 32'h02c863bd;
    ram_cell[    3873] = 32'h0;  // 32'he5bb25a8;
    ram_cell[    3874] = 32'h0;  // 32'h7c2c5461;
    ram_cell[    3875] = 32'h0;  // 32'h918940b1;
    ram_cell[    3876] = 32'h0;  // 32'hb867819c;
    ram_cell[    3877] = 32'h0;  // 32'hcde41a93;
    ram_cell[    3878] = 32'h0;  // 32'h331d2cbf;
    ram_cell[    3879] = 32'h0;  // 32'hf45d1895;
    ram_cell[    3880] = 32'h0;  // 32'h519a4ee1;
    ram_cell[    3881] = 32'h0;  // 32'h985ecc02;
    ram_cell[    3882] = 32'h0;  // 32'h76756378;
    ram_cell[    3883] = 32'h0;  // 32'h2c23fe89;
    ram_cell[    3884] = 32'h0;  // 32'ha0f257e3;
    ram_cell[    3885] = 32'h0;  // 32'h18881e61;
    ram_cell[    3886] = 32'h0;  // 32'hec011ae7;
    ram_cell[    3887] = 32'h0;  // 32'h71278e31;
    ram_cell[    3888] = 32'h0;  // 32'hdd183250;
    ram_cell[    3889] = 32'h0;  // 32'ha3e570e9;
    ram_cell[    3890] = 32'h0;  // 32'hebf78895;
    ram_cell[    3891] = 32'h0;  // 32'ha7ed4d4e;
    ram_cell[    3892] = 32'h0;  // 32'ha30fdce8;
    ram_cell[    3893] = 32'h0;  // 32'h0f219e00;
    ram_cell[    3894] = 32'h0;  // 32'h7f9d24b5;
    ram_cell[    3895] = 32'h0;  // 32'h89caaec4;
    ram_cell[    3896] = 32'h0;  // 32'h08132d9a;
    ram_cell[    3897] = 32'h0;  // 32'hc3ce701b;
    ram_cell[    3898] = 32'h0;  // 32'h4c69a18d;
    ram_cell[    3899] = 32'h0;  // 32'h16ab7766;
    ram_cell[    3900] = 32'h0;  // 32'h86051b72;
    ram_cell[    3901] = 32'h0;  // 32'hd0b2e4a3;
    ram_cell[    3902] = 32'h0;  // 32'h5736f3f6;
    ram_cell[    3903] = 32'h0;  // 32'hf22e8440;
    ram_cell[    3904] = 32'h0;  // 32'hf618d8e5;
    ram_cell[    3905] = 32'h0;  // 32'h70228dc0;
    ram_cell[    3906] = 32'h0;  // 32'h70dcf4f5;
    ram_cell[    3907] = 32'h0;  // 32'h0433740f;
    ram_cell[    3908] = 32'h0;  // 32'he310ebfa;
    ram_cell[    3909] = 32'h0;  // 32'ha7e4f907;
    ram_cell[    3910] = 32'h0;  // 32'h88956e73;
    ram_cell[    3911] = 32'h0;  // 32'hf2d2c23f;
    ram_cell[    3912] = 32'h0;  // 32'ha332ff20;
    ram_cell[    3913] = 32'h0;  // 32'h1fc25d7b;
    ram_cell[    3914] = 32'h0;  // 32'hae9f2cca;
    ram_cell[    3915] = 32'h0;  // 32'hc6096c62;
    ram_cell[    3916] = 32'h0;  // 32'hce3528f6;
    ram_cell[    3917] = 32'h0;  // 32'h9e280483;
    ram_cell[    3918] = 32'h0;  // 32'hbcb66f12;
    ram_cell[    3919] = 32'h0;  // 32'h9430ee27;
    ram_cell[    3920] = 32'h0;  // 32'h38214d8e;
    ram_cell[    3921] = 32'h0;  // 32'h479d3ff8;
    ram_cell[    3922] = 32'h0;  // 32'h5fd1de41;
    ram_cell[    3923] = 32'h0;  // 32'hdf082f45;
    ram_cell[    3924] = 32'h0;  // 32'h4a37306d;
    ram_cell[    3925] = 32'h0;  // 32'h2b38ac07;
    ram_cell[    3926] = 32'h0;  // 32'h2fc3a66d;
    ram_cell[    3927] = 32'h0;  // 32'ha10b347f;
    ram_cell[    3928] = 32'h0;  // 32'hb488ea4e;
    ram_cell[    3929] = 32'h0;  // 32'h8713153d;
    ram_cell[    3930] = 32'h0;  // 32'hf3dcfffc;
    ram_cell[    3931] = 32'h0;  // 32'ha17d5908;
    ram_cell[    3932] = 32'h0;  // 32'h6ce4b83a;
    ram_cell[    3933] = 32'h0;  // 32'h245a09ee;
    ram_cell[    3934] = 32'h0;  // 32'haebedcf1;
    ram_cell[    3935] = 32'h0;  // 32'h1a9fd38d;
    ram_cell[    3936] = 32'h0;  // 32'h348d2795;
    ram_cell[    3937] = 32'h0;  // 32'h5e9b87a8;
    ram_cell[    3938] = 32'h0;  // 32'hf00aa1d9;
    ram_cell[    3939] = 32'h0;  // 32'h7818e6dd;
    ram_cell[    3940] = 32'h0;  // 32'h275bba9a;
    ram_cell[    3941] = 32'h0;  // 32'ha51d5999;
    ram_cell[    3942] = 32'h0;  // 32'hdceb57b3;
    ram_cell[    3943] = 32'h0;  // 32'he6166562;
    ram_cell[    3944] = 32'h0;  // 32'h1dec2bed;
    ram_cell[    3945] = 32'h0;  // 32'he3bfc0f4;
    ram_cell[    3946] = 32'h0;  // 32'h97a5e99b;
    ram_cell[    3947] = 32'h0;  // 32'h4326797b;
    ram_cell[    3948] = 32'h0;  // 32'h2d8b444f;
    ram_cell[    3949] = 32'h0;  // 32'h20064913;
    ram_cell[    3950] = 32'h0;  // 32'hba1fbca6;
    ram_cell[    3951] = 32'h0;  // 32'hb36a8385;
    ram_cell[    3952] = 32'h0;  // 32'ha82a0d99;
    ram_cell[    3953] = 32'h0;  // 32'h369d8bd1;
    ram_cell[    3954] = 32'h0;  // 32'hea4175cf;
    ram_cell[    3955] = 32'h0;  // 32'ha2dfbd16;
    ram_cell[    3956] = 32'h0;  // 32'h1132ca94;
    ram_cell[    3957] = 32'h0;  // 32'h86830404;
    ram_cell[    3958] = 32'h0;  // 32'hfa6eb68f;
    ram_cell[    3959] = 32'h0;  // 32'he0339150;
    ram_cell[    3960] = 32'h0;  // 32'h529d3afe;
    ram_cell[    3961] = 32'h0;  // 32'hea784326;
    ram_cell[    3962] = 32'h0;  // 32'h80c01d4b;
    ram_cell[    3963] = 32'h0;  // 32'hdbbd0047;
    ram_cell[    3964] = 32'h0;  // 32'hbc903682;
    ram_cell[    3965] = 32'h0;  // 32'h501dd4b1;
    ram_cell[    3966] = 32'h0;  // 32'h6a562087;
    ram_cell[    3967] = 32'h0;  // 32'hfcf13545;
    ram_cell[    3968] = 32'h0;  // 32'hf35aec3c;
    ram_cell[    3969] = 32'h0;  // 32'h7a1b7226;
    ram_cell[    3970] = 32'h0;  // 32'h6f1048a0;
    ram_cell[    3971] = 32'h0;  // 32'h22e346b2;
    ram_cell[    3972] = 32'h0;  // 32'hef665b2b;
    ram_cell[    3973] = 32'h0;  // 32'h51f15614;
    ram_cell[    3974] = 32'h0;  // 32'ha37be50b;
    ram_cell[    3975] = 32'h0;  // 32'hecfaa532;
    ram_cell[    3976] = 32'h0;  // 32'h6b90a275;
    ram_cell[    3977] = 32'h0;  // 32'hb85c837a;
    ram_cell[    3978] = 32'h0;  // 32'h2b81c23e;
    ram_cell[    3979] = 32'h0;  // 32'h384ae32b;
    ram_cell[    3980] = 32'h0;  // 32'h3f46acc5;
    ram_cell[    3981] = 32'h0;  // 32'h769d5c27;
    ram_cell[    3982] = 32'h0;  // 32'ha2dce98a;
    ram_cell[    3983] = 32'h0;  // 32'h55b49fb0;
    ram_cell[    3984] = 32'h0;  // 32'hab763c46;
    ram_cell[    3985] = 32'h0;  // 32'h6b8f4d11;
    ram_cell[    3986] = 32'h0;  // 32'hed50c986;
    ram_cell[    3987] = 32'h0;  // 32'h5cc19f87;
    ram_cell[    3988] = 32'h0;  // 32'hea871468;
    ram_cell[    3989] = 32'h0;  // 32'hf427827c;
    ram_cell[    3990] = 32'h0;  // 32'h18512f53;
    ram_cell[    3991] = 32'h0;  // 32'h6973aeb7;
    ram_cell[    3992] = 32'h0;  // 32'hd1c2324f;
    ram_cell[    3993] = 32'h0;  // 32'ha2d14bb6;
    ram_cell[    3994] = 32'h0;  // 32'h6b1b0e88;
    ram_cell[    3995] = 32'h0;  // 32'h0be5ed09;
    ram_cell[    3996] = 32'h0;  // 32'hb8031ba7;
    ram_cell[    3997] = 32'h0;  // 32'hb6f5722d;
    ram_cell[    3998] = 32'h0;  // 32'hb9706f75;
    ram_cell[    3999] = 32'h0;  // 32'h47a5c6b1;
    ram_cell[    4000] = 32'h0;  // 32'h49fc5bf4;
    ram_cell[    4001] = 32'h0;  // 32'h6619e299;
    ram_cell[    4002] = 32'h0;  // 32'h1ce86504;
    ram_cell[    4003] = 32'h0;  // 32'h4f0ef4b6;
    ram_cell[    4004] = 32'h0;  // 32'h000d12de;
    ram_cell[    4005] = 32'h0;  // 32'h249d5fa4;
    ram_cell[    4006] = 32'h0;  // 32'h5e8dc896;
    ram_cell[    4007] = 32'h0;  // 32'h3fb74588;
    ram_cell[    4008] = 32'h0;  // 32'hbffdcdcd;
    ram_cell[    4009] = 32'h0;  // 32'h050a83d2;
    ram_cell[    4010] = 32'h0;  // 32'h42b9dab7;
    ram_cell[    4011] = 32'h0;  // 32'h89bc59fb;
    ram_cell[    4012] = 32'h0;  // 32'hded50717;
    ram_cell[    4013] = 32'h0;  // 32'h5e24c0d7;
    ram_cell[    4014] = 32'h0;  // 32'hedcd2263;
    ram_cell[    4015] = 32'h0;  // 32'hbf6d2918;
    ram_cell[    4016] = 32'h0;  // 32'h52453ee1;
    ram_cell[    4017] = 32'h0;  // 32'ha3657558;
    ram_cell[    4018] = 32'h0;  // 32'h9a53a0a6;
    ram_cell[    4019] = 32'h0;  // 32'hb1cc3bda;
    ram_cell[    4020] = 32'h0;  // 32'hfd2f9450;
    ram_cell[    4021] = 32'h0;  // 32'hc0eb18e2;
    ram_cell[    4022] = 32'h0;  // 32'h53707d83;
    ram_cell[    4023] = 32'h0;  // 32'he13ab64f;
    ram_cell[    4024] = 32'h0;  // 32'h25c57974;
    ram_cell[    4025] = 32'h0;  // 32'h1fcade55;
    ram_cell[    4026] = 32'h0;  // 32'h01257b1f;
    ram_cell[    4027] = 32'h0;  // 32'hb596c797;
    ram_cell[    4028] = 32'h0;  // 32'ha415a32e;
    ram_cell[    4029] = 32'h0;  // 32'h1946d50b;
    ram_cell[    4030] = 32'h0;  // 32'h0709554a;
    ram_cell[    4031] = 32'h0;  // 32'h240cdb30;
    ram_cell[    4032] = 32'h0;  // 32'he4f986f2;
    ram_cell[    4033] = 32'h0;  // 32'ha93e71b0;
    ram_cell[    4034] = 32'h0;  // 32'h17e90305;
    ram_cell[    4035] = 32'h0;  // 32'h918e6b39;
    ram_cell[    4036] = 32'h0;  // 32'h6459d63e;
    ram_cell[    4037] = 32'h0;  // 32'h8f3035bc;
    ram_cell[    4038] = 32'h0;  // 32'h2da056f2;
    ram_cell[    4039] = 32'h0;  // 32'h82616dc3;
    ram_cell[    4040] = 32'h0;  // 32'h7bac8588;
    ram_cell[    4041] = 32'h0;  // 32'h2e995b0e;
    ram_cell[    4042] = 32'h0;  // 32'h72537f1a;
    ram_cell[    4043] = 32'h0;  // 32'h20a06bc5;
    ram_cell[    4044] = 32'h0;  // 32'h18e58ea0;
    ram_cell[    4045] = 32'h0;  // 32'h7cf05197;
    ram_cell[    4046] = 32'h0;  // 32'h1f72a605;
    ram_cell[    4047] = 32'h0;  // 32'h674e06db;
    ram_cell[    4048] = 32'h0;  // 32'hedaa6053;
    ram_cell[    4049] = 32'h0;  // 32'h5595d690;
    ram_cell[    4050] = 32'h0;  // 32'hd10d18ab;
    ram_cell[    4051] = 32'h0;  // 32'h294ec038;
    ram_cell[    4052] = 32'h0;  // 32'hb699c53b;
    ram_cell[    4053] = 32'h0;  // 32'h10c8ebe2;
    ram_cell[    4054] = 32'h0;  // 32'h18093da6;
    ram_cell[    4055] = 32'h0;  // 32'hc01a1873;
    ram_cell[    4056] = 32'h0;  // 32'h479395ac;
    ram_cell[    4057] = 32'h0;  // 32'h484c3228;
    ram_cell[    4058] = 32'h0;  // 32'hd0f5b55f;
    ram_cell[    4059] = 32'h0;  // 32'h0acbf7e0;
    ram_cell[    4060] = 32'h0;  // 32'h0dfb6613;
    ram_cell[    4061] = 32'h0;  // 32'h6898f41e;
    ram_cell[    4062] = 32'h0;  // 32'ha43e0562;
    ram_cell[    4063] = 32'h0;  // 32'he6be3dbf;
    ram_cell[    4064] = 32'h0;  // 32'h313e35c3;
    ram_cell[    4065] = 32'h0;  // 32'h282f60db;
    ram_cell[    4066] = 32'h0;  // 32'hc2104445;
    ram_cell[    4067] = 32'h0;  // 32'hd644cf86;
    ram_cell[    4068] = 32'h0;  // 32'had94f574;
    ram_cell[    4069] = 32'h0;  // 32'hf50aa5c6;
    ram_cell[    4070] = 32'h0;  // 32'h94d1e811;
    ram_cell[    4071] = 32'h0;  // 32'h04b8bf77;
    ram_cell[    4072] = 32'h0;  // 32'ha0b6f399;
    ram_cell[    4073] = 32'h0;  // 32'h90270eea;
    ram_cell[    4074] = 32'h0;  // 32'hdc670f78;
    ram_cell[    4075] = 32'h0;  // 32'h20e8dac6;
    ram_cell[    4076] = 32'h0;  // 32'h89fe0b8d;
    ram_cell[    4077] = 32'h0;  // 32'ha8968c2a;
    ram_cell[    4078] = 32'h0;  // 32'h254ddfe7;
    ram_cell[    4079] = 32'h0;  // 32'h117c3954;
    ram_cell[    4080] = 32'h0;  // 32'h8ea41118;
    ram_cell[    4081] = 32'h0;  // 32'hdec83751;
    ram_cell[    4082] = 32'h0;  // 32'heb23b8d7;
    ram_cell[    4083] = 32'h0;  // 32'h231e91ae;
    ram_cell[    4084] = 32'h0;  // 32'h72647d54;
    ram_cell[    4085] = 32'h0;  // 32'h24cbd514;
    ram_cell[    4086] = 32'h0;  // 32'hc761085a;
    ram_cell[    4087] = 32'h0;  // 32'he45c7909;
    ram_cell[    4088] = 32'h0;  // 32'ha4faa151;
    ram_cell[    4089] = 32'h0;  // 32'hfbcc6c06;
    ram_cell[    4090] = 32'h0;  // 32'hb9a359d8;
    ram_cell[    4091] = 32'h0;  // 32'h4ef8737d;
    ram_cell[    4092] = 32'h0;  // 32'h06ec51b9;
    ram_cell[    4093] = 32'h0;  // 32'h0043efbe;
    ram_cell[    4094] = 32'h0;  // 32'ha25069de;
    ram_cell[    4095] = 32'h0;  // 32'h4f4c8c9f;
    ram_cell[    4096] = 32'h0;  // 32'hf16c6305;
    ram_cell[    4097] = 32'h0;  // 32'h43164f8e;
    ram_cell[    4098] = 32'h0;  // 32'hf4f8e449;
    ram_cell[    4099] = 32'h0;  // 32'h58f599c9;
    ram_cell[    4100] = 32'h0;  // 32'h202d5fa0;
    ram_cell[    4101] = 32'h0;  // 32'h284c044e;
    ram_cell[    4102] = 32'h0;  // 32'hc9fba34e;
    ram_cell[    4103] = 32'h0;  // 32'hcb457fa3;
    ram_cell[    4104] = 32'h0;  // 32'h3be75f61;
    ram_cell[    4105] = 32'h0;  // 32'hc84240a1;
    ram_cell[    4106] = 32'h0;  // 32'h62c4b997;
    ram_cell[    4107] = 32'h0;  // 32'h930007c9;
    ram_cell[    4108] = 32'h0;  // 32'hcdfdf309;
    ram_cell[    4109] = 32'h0;  // 32'h963b1357;
    ram_cell[    4110] = 32'h0;  // 32'h6b835ee8;
    ram_cell[    4111] = 32'h0;  // 32'hb4df378c;
    ram_cell[    4112] = 32'h0;  // 32'h69d0c5aa;
    ram_cell[    4113] = 32'h0;  // 32'hcd436fba;
    ram_cell[    4114] = 32'h0;  // 32'h99d63e92;
    ram_cell[    4115] = 32'h0;  // 32'h7e2a38ad;
    ram_cell[    4116] = 32'h0;  // 32'h19b48ba2;
    ram_cell[    4117] = 32'h0;  // 32'hd0b9df86;
    ram_cell[    4118] = 32'h0;  // 32'ha6948efb;
    ram_cell[    4119] = 32'h0;  // 32'h491fd3e5;
    ram_cell[    4120] = 32'h0;  // 32'hf1fc445b;
    ram_cell[    4121] = 32'h0;  // 32'hd2cd2a28;
    ram_cell[    4122] = 32'h0;  // 32'h3341e4dd;
    ram_cell[    4123] = 32'h0;  // 32'h3181df5d;
    ram_cell[    4124] = 32'h0;  // 32'h1efece65;
    ram_cell[    4125] = 32'h0;  // 32'h2e64a506;
    ram_cell[    4126] = 32'h0;  // 32'hd093af12;
    ram_cell[    4127] = 32'h0;  // 32'h3e1a0085;
    ram_cell[    4128] = 32'h0;  // 32'h6b1b781c;
    ram_cell[    4129] = 32'h0;  // 32'ha198c2f8;
    ram_cell[    4130] = 32'h0;  // 32'h73e82428;
    ram_cell[    4131] = 32'h0;  // 32'hc0213419;
    ram_cell[    4132] = 32'h0;  // 32'h20a5bc0d;
    ram_cell[    4133] = 32'h0;  // 32'h9acc06cc;
    ram_cell[    4134] = 32'h0;  // 32'h402d3a8c;
    ram_cell[    4135] = 32'h0;  // 32'hf99a9b00;
    ram_cell[    4136] = 32'h0;  // 32'h86d23250;
    ram_cell[    4137] = 32'h0;  // 32'h8cd7dbec;
    ram_cell[    4138] = 32'h0;  // 32'h41f7113f;
    ram_cell[    4139] = 32'h0;  // 32'h69cb7a5b;
    ram_cell[    4140] = 32'h0;  // 32'hbde9f39f;
    ram_cell[    4141] = 32'h0;  // 32'hdf52159a;
    ram_cell[    4142] = 32'h0;  // 32'hbe4c43f7;
    ram_cell[    4143] = 32'h0;  // 32'h97a5b34e;
    ram_cell[    4144] = 32'h0;  // 32'he5bba0b4;
    ram_cell[    4145] = 32'h0;  // 32'hb5128be8;
    ram_cell[    4146] = 32'h0;  // 32'h9207c1bb;
    ram_cell[    4147] = 32'h0;  // 32'h5608afcd;
    ram_cell[    4148] = 32'h0;  // 32'h05da1d58;
    ram_cell[    4149] = 32'h0;  // 32'h9b0d753f;
    ram_cell[    4150] = 32'h0;  // 32'hbbe83ffd;
    ram_cell[    4151] = 32'h0;  // 32'hde6d1d43;
    ram_cell[    4152] = 32'h0;  // 32'hb095b738;
    ram_cell[    4153] = 32'h0;  // 32'hecfb658f;
    ram_cell[    4154] = 32'h0;  // 32'hfe9cb37a;
    ram_cell[    4155] = 32'h0;  // 32'h38bfc533;
    ram_cell[    4156] = 32'h0;  // 32'h50b6d2b1;
    ram_cell[    4157] = 32'h0;  // 32'h6831adb3;
    ram_cell[    4158] = 32'h0;  // 32'h746e03b1;
    ram_cell[    4159] = 32'h0;  // 32'h300ac901;
    ram_cell[    4160] = 32'h0;  // 32'h2bbd9352;
    ram_cell[    4161] = 32'h0;  // 32'h0598d768;
    ram_cell[    4162] = 32'h0;  // 32'hc8ce1031;
    ram_cell[    4163] = 32'h0;  // 32'hff7b8b72;
    ram_cell[    4164] = 32'h0;  // 32'h1465af6f;
    ram_cell[    4165] = 32'h0;  // 32'h08cedebf;
    ram_cell[    4166] = 32'h0;  // 32'h5a6e48a0;
    ram_cell[    4167] = 32'h0;  // 32'hf2b0d945;
    ram_cell[    4168] = 32'h0;  // 32'ha3cdb847;
    ram_cell[    4169] = 32'h0;  // 32'hd3082b22;
    ram_cell[    4170] = 32'h0;  // 32'h88364a44;
    ram_cell[    4171] = 32'h0;  // 32'h4415de1d;
    ram_cell[    4172] = 32'h0;  // 32'h67df84ea;
    ram_cell[    4173] = 32'h0;  // 32'h32abe333;
    ram_cell[    4174] = 32'h0;  // 32'hfc5b03b7;
    ram_cell[    4175] = 32'h0;  // 32'hbae537ae;
    ram_cell[    4176] = 32'h0;  // 32'he00847bd;
    ram_cell[    4177] = 32'h0;  // 32'h115c129b;
    ram_cell[    4178] = 32'h0;  // 32'hf83c9e85;
    ram_cell[    4179] = 32'h0;  // 32'h720fa092;
    ram_cell[    4180] = 32'h0;  // 32'h8ae01719;
    ram_cell[    4181] = 32'h0;  // 32'hff235e23;
    ram_cell[    4182] = 32'h0;  // 32'h4bd2f789;
    ram_cell[    4183] = 32'h0;  // 32'h93959086;
    ram_cell[    4184] = 32'h0;  // 32'hb8fef4b8;
    ram_cell[    4185] = 32'h0;  // 32'h0f87f77c;
    ram_cell[    4186] = 32'h0;  // 32'h85456fc7;
    ram_cell[    4187] = 32'h0;  // 32'h4ea1057d;
    ram_cell[    4188] = 32'h0;  // 32'h25cf98cc;
    ram_cell[    4189] = 32'h0;  // 32'h499c3d15;
    ram_cell[    4190] = 32'h0;  // 32'h6ee1250a;
    ram_cell[    4191] = 32'h0;  // 32'h6a06de49;
    ram_cell[    4192] = 32'h0;  // 32'he40fc197;
    ram_cell[    4193] = 32'h0;  // 32'he94f30b1;
    ram_cell[    4194] = 32'h0;  // 32'h6eed30ca;
    ram_cell[    4195] = 32'h0;  // 32'h8385d3a9;
    ram_cell[    4196] = 32'h0;  // 32'ha8ee8694;
    ram_cell[    4197] = 32'h0;  // 32'h6539bc42;
    ram_cell[    4198] = 32'h0;  // 32'h66d4495c;
    ram_cell[    4199] = 32'h0;  // 32'ha0ffc614;
    ram_cell[    4200] = 32'h0;  // 32'hbe9fe0df;
    ram_cell[    4201] = 32'h0;  // 32'hdcde9e82;
    ram_cell[    4202] = 32'h0;  // 32'h934acd07;
    ram_cell[    4203] = 32'h0;  // 32'h9c11471c;
    ram_cell[    4204] = 32'h0;  // 32'hef0bf5b6;
    ram_cell[    4205] = 32'h0;  // 32'hc7eb7446;
    ram_cell[    4206] = 32'h0;  // 32'h62a275ff;
    ram_cell[    4207] = 32'h0;  // 32'h52550fe1;
    ram_cell[    4208] = 32'h0;  // 32'h644d0512;
    ram_cell[    4209] = 32'h0;  // 32'h192e3fff;
    ram_cell[    4210] = 32'h0;  // 32'h6f94408c;
    ram_cell[    4211] = 32'h0;  // 32'h96c0ac24;
    ram_cell[    4212] = 32'h0;  // 32'hf8b129f1;
    ram_cell[    4213] = 32'h0;  // 32'h8e253b19;
    ram_cell[    4214] = 32'h0;  // 32'he4011f7a;
    ram_cell[    4215] = 32'h0;  // 32'hfbeccbf5;
    ram_cell[    4216] = 32'h0;  // 32'h6369048a;
    ram_cell[    4217] = 32'h0;  // 32'hcdb1db35;
    ram_cell[    4218] = 32'h0;  // 32'h4ef4aad7;
    ram_cell[    4219] = 32'h0;  // 32'h3611007e;
    ram_cell[    4220] = 32'h0;  // 32'h3703ca30;
    ram_cell[    4221] = 32'h0;  // 32'h5c5c49f1;
    ram_cell[    4222] = 32'h0;  // 32'h6e376476;
    ram_cell[    4223] = 32'h0;  // 32'hb0988c80;
    ram_cell[    4224] = 32'h0;  // 32'hcdde5873;
    ram_cell[    4225] = 32'h0;  // 32'hbf0b95b5;
    ram_cell[    4226] = 32'h0;  // 32'h899e04d0;
    ram_cell[    4227] = 32'h0;  // 32'hd7199628;
    ram_cell[    4228] = 32'h0;  // 32'h7a2d2494;
    ram_cell[    4229] = 32'h0;  // 32'h7b4f096e;
    ram_cell[    4230] = 32'h0;  // 32'h2dba5a44;
    ram_cell[    4231] = 32'h0;  // 32'hcf3e2179;
    ram_cell[    4232] = 32'h0;  // 32'h7babcc8c;
    ram_cell[    4233] = 32'h0;  // 32'h874c38a7;
    ram_cell[    4234] = 32'h0;  // 32'h98a99590;
    ram_cell[    4235] = 32'h0;  // 32'hb883f299;
    ram_cell[    4236] = 32'h0;  // 32'h6694173b;
    ram_cell[    4237] = 32'h0;  // 32'he382891d;
    ram_cell[    4238] = 32'h0;  // 32'h7a88c191;
    ram_cell[    4239] = 32'h0;  // 32'hef657a6a;
    ram_cell[    4240] = 32'h0;  // 32'h31bded6c;
    ram_cell[    4241] = 32'h0;  // 32'heb987919;
    ram_cell[    4242] = 32'h0;  // 32'h064dc628;
    ram_cell[    4243] = 32'h0;  // 32'h038733b5;
    ram_cell[    4244] = 32'h0;  // 32'h768e8dd4;
    ram_cell[    4245] = 32'h0;  // 32'h2687a26d;
    ram_cell[    4246] = 32'h0;  // 32'h0c1b50ce;
    ram_cell[    4247] = 32'h0;  // 32'hf056ba18;
    ram_cell[    4248] = 32'h0;  // 32'hed73da17;
    ram_cell[    4249] = 32'h0;  // 32'h0ef92794;
    ram_cell[    4250] = 32'h0;  // 32'h665ba81d;
    ram_cell[    4251] = 32'h0;  // 32'hd2b69bd1;
    ram_cell[    4252] = 32'h0;  // 32'h0bed2f24;
    ram_cell[    4253] = 32'h0;  // 32'hb5678f4f;
    ram_cell[    4254] = 32'h0;  // 32'h7af87636;
    ram_cell[    4255] = 32'h0;  // 32'h508a3025;
    ram_cell[    4256] = 32'h0;  // 32'hbfdd91fc;
    ram_cell[    4257] = 32'h0;  // 32'hb7d965ad;
    ram_cell[    4258] = 32'h0;  // 32'hc42f100b;
    ram_cell[    4259] = 32'h0;  // 32'h7fbc2e0d;
    ram_cell[    4260] = 32'h0;  // 32'hcc970dc3;
    ram_cell[    4261] = 32'h0;  // 32'h73b020bc;
    ram_cell[    4262] = 32'h0;  // 32'ha1ab0c2b;
    ram_cell[    4263] = 32'h0;  // 32'h110025a7;
    ram_cell[    4264] = 32'h0;  // 32'h26363420;
    ram_cell[    4265] = 32'h0;  // 32'h9e5848bb;
    ram_cell[    4266] = 32'h0;  // 32'hafa20807;
    ram_cell[    4267] = 32'h0;  // 32'h56f56f12;
    ram_cell[    4268] = 32'h0;  // 32'hbec85927;
    ram_cell[    4269] = 32'h0;  // 32'h79c5d966;
    ram_cell[    4270] = 32'h0;  // 32'h940f7fac;
    ram_cell[    4271] = 32'h0;  // 32'h64222bd7;
    ram_cell[    4272] = 32'h0;  // 32'h39775296;
    ram_cell[    4273] = 32'h0;  // 32'hd8e036eb;
    ram_cell[    4274] = 32'h0;  // 32'h76ef48a9;
    ram_cell[    4275] = 32'h0;  // 32'h9e403ce5;
    ram_cell[    4276] = 32'h0;  // 32'h7f0a3330;
    ram_cell[    4277] = 32'h0;  // 32'hf93fdd29;
    ram_cell[    4278] = 32'h0;  // 32'h2a88eee3;
    ram_cell[    4279] = 32'h0;  // 32'h049216cc;
    ram_cell[    4280] = 32'h0;  // 32'hd865f4d7;
    ram_cell[    4281] = 32'h0;  // 32'hf93c4177;
    ram_cell[    4282] = 32'h0;  // 32'h9364b256;
    ram_cell[    4283] = 32'h0;  // 32'h317f765d;
    ram_cell[    4284] = 32'h0;  // 32'hbb0e55a4;
    ram_cell[    4285] = 32'h0;  // 32'h76d583fe;
    ram_cell[    4286] = 32'h0;  // 32'h9372a218;
    ram_cell[    4287] = 32'h0;  // 32'h32206c05;
    ram_cell[    4288] = 32'h0;  // 32'hc56b85e4;
    ram_cell[    4289] = 32'h0;  // 32'h77845c45;
    ram_cell[    4290] = 32'h0;  // 32'hf0008350;
    ram_cell[    4291] = 32'h0;  // 32'h4467e528;
    ram_cell[    4292] = 32'h0;  // 32'h5ce3b273;
    ram_cell[    4293] = 32'h0;  // 32'h0ccbb4ca;
    ram_cell[    4294] = 32'h0;  // 32'h8d40dcd8;
    ram_cell[    4295] = 32'h0;  // 32'h9224743e;
    ram_cell[    4296] = 32'h0;  // 32'h300df73a;
    ram_cell[    4297] = 32'h0;  // 32'h79d37bbe;
    ram_cell[    4298] = 32'h0;  // 32'ha18b711c;
    ram_cell[    4299] = 32'h0;  // 32'h570a3fb3;
    ram_cell[    4300] = 32'h0;  // 32'hdee35738;
    ram_cell[    4301] = 32'h0;  // 32'hc7098583;
    ram_cell[    4302] = 32'h0;  // 32'hf33abef1;
    ram_cell[    4303] = 32'h0;  // 32'h4b772314;
    ram_cell[    4304] = 32'h0;  // 32'h01013bdb;
    ram_cell[    4305] = 32'h0;  // 32'h0712e6f6;
    ram_cell[    4306] = 32'h0;  // 32'h6ba47dbc;
    ram_cell[    4307] = 32'h0;  // 32'h47120281;
    ram_cell[    4308] = 32'h0;  // 32'h0547eae3;
    ram_cell[    4309] = 32'h0;  // 32'h61d374e2;
    ram_cell[    4310] = 32'h0;  // 32'hae24cc81;
    ram_cell[    4311] = 32'h0;  // 32'h8a6773ba;
    ram_cell[    4312] = 32'h0;  // 32'hb86037bc;
    ram_cell[    4313] = 32'h0;  // 32'had01b231;
    ram_cell[    4314] = 32'h0;  // 32'h1f10c229;
    ram_cell[    4315] = 32'h0;  // 32'h7bb37ebf;
    ram_cell[    4316] = 32'h0;  // 32'h373ad6a1;
    ram_cell[    4317] = 32'h0;  // 32'h6ec1a8cd;
    ram_cell[    4318] = 32'h0;  // 32'h3bbae38f;
    ram_cell[    4319] = 32'h0;  // 32'h2da8649a;
    ram_cell[    4320] = 32'h0;  // 32'h11699385;
    ram_cell[    4321] = 32'h0;  // 32'hc010f9c7;
    ram_cell[    4322] = 32'h0;  // 32'hbbf706c4;
    ram_cell[    4323] = 32'h0;  // 32'h230e4cd1;
    ram_cell[    4324] = 32'h0;  // 32'ha2b666ff;
    ram_cell[    4325] = 32'h0;  // 32'hcd71774f;
    ram_cell[    4326] = 32'h0;  // 32'h5d6971e1;
    ram_cell[    4327] = 32'h0;  // 32'h6e8a9d8d;
    ram_cell[    4328] = 32'h0;  // 32'h4303d64c;
    ram_cell[    4329] = 32'h0;  // 32'h187e7f66;
    ram_cell[    4330] = 32'h0;  // 32'h4a68ee0e;
    ram_cell[    4331] = 32'h0;  // 32'hd38296df;
    ram_cell[    4332] = 32'h0;  // 32'h3465e54e;
    ram_cell[    4333] = 32'h0;  // 32'h402a4fcf;
    ram_cell[    4334] = 32'h0;  // 32'h1d717362;
    ram_cell[    4335] = 32'h0;  // 32'h5aec176f;
    ram_cell[    4336] = 32'h0;  // 32'hca6c0c05;
    ram_cell[    4337] = 32'h0;  // 32'hb519a9bb;
    ram_cell[    4338] = 32'h0;  // 32'h824d55f1;
    ram_cell[    4339] = 32'h0;  // 32'h29c96a38;
    ram_cell[    4340] = 32'h0;  // 32'hc44d21f1;
    ram_cell[    4341] = 32'h0;  // 32'hc015a2e4;
    ram_cell[    4342] = 32'h0;  // 32'hb86d1d71;
    ram_cell[    4343] = 32'h0;  // 32'h63de4bab;
    ram_cell[    4344] = 32'h0;  // 32'h21eef753;
    ram_cell[    4345] = 32'h0;  // 32'ha20e31ac;
    ram_cell[    4346] = 32'h0;  // 32'hf9dd04d9;
    ram_cell[    4347] = 32'h0;  // 32'h7ce18dac;
    ram_cell[    4348] = 32'h0;  // 32'hb2a21c06;
    ram_cell[    4349] = 32'h0;  // 32'h635b0533;
    ram_cell[    4350] = 32'h0;  // 32'ha879c035;
    ram_cell[    4351] = 32'h0;  // 32'h6e4a1cf1;
    ram_cell[    4352] = 32'h0;  // 32'h57cccca2;
    ram_cell[    4353] = 32'h0;  // 32'h21f17744;
    ram_cell[    4354] = 32'h0;  // 32'hd6997060;
    ram_cell[    4355] = 32'h0;  // 32'he21a9c6e;
    ram_cell[    4356] = 32'h0;  // 32'hcc35f748;
    ram_cell[    4357] = 32'h0;  // 32'hfcd92b1e;
    ram_cell[    4358] = 32'h0;  // 32'heb1ff16d;
    ram_cell[    4359] = 32'h0;  // 32'heccbebc2;
    ram_cell[    4360] = 32'h0;  // 32'hbbbc963b;
    ram_cell[    4361] = 32'h0;  // 32'h4a98e1b8;
    ram_cell[    4362] = 32'h0;  // 32'he62fc624;
    ram_cell[    4363] = 32'h0;  // 32'hb7fd1dc7;
    ram_cell[    4364] = 32'h0;  // 32'h4a3369b9;
    ram_cell[    4365] = 32'h0;  // 32'h5eed89b0;
    ram_cell[    4366] = 32'h0;  // 32'hcaa7def4;
    ram_cell[    4367] = 32'h0;  // 32'h370b1492;
    ram_cell[    4368] = 32'h0;  // 32'h32c916c6;
    ram_cell[    4369] = 32'h0;  // 32'h83664238;
    ram_cell[    4370] = 32'h0;  // 32'h3cbdc9c6;
    ram_cell[    4371] = 32'h0;  // 32'h6c53aff0;
    ram_cell[    4372] = 32'h0;  // 32'h0e9180fd;
    ram_cell[    4373] = 32'h0;  // 32'h8938dda6;
    ram_cell[    4374] = 32'h0;  // 32'h5786dc57;
    ram_cell[    4375] = 32'h0;  // 32'h6422c81c;
    ram_cell[    4376] = 32'h0;  // 32'hd14976ad;
    ram_cell[    4377] = 32'h0;  // 32'h2589769f;
    ram_cell[    4378] = 32'h0;  // 32'h6d2f40e9;
    ram_cell[    4379] = 32'h0;  // 32'h9b228a03;
    ram_cell[    4380] = 32'h0;  // 32'h2a5c4d5e;
    ram_cell[    4381] = 32'h0;  // 32'ha0e87276;
    ram_cell[    4382] = 32'h0;  // 32'he1ed4a31;
    ram_cell[    4383] = 32'h0;  // 32'hbd0de437;
    ram_cell[    4384] = 32'h0;  // 32'heb628fa0;
    ram_cell[    4385] = 32'h0;  // 32'h66397ba0;
    ram_cell[    4386] = 32'h0;  // 32'h883df170;
    ram_cell[    4387] = 32'h0;  // 32'h794bf560;
    ram_cell[    4388] = 32'h0;  // 32'h07e7b092;
    ram_cell[    4389] = 32'h0;  // 32'h7178c9dd;
    ram_cell[    4390] = 32'h0;  // 32'h7b406daf;
    ram_cell[    4391] = 32'h0;  // 32'h96804971;
    ram_cell[    4392] = 32'h0;  // 32'h9e355bc0;
    ram_cell[    4393] = 32'h0;  // 32'haacfa4aa;
    ram_cell[    4394] = 32'h0;  // 32'hc370b8f9;
    ram_cell[    4395] = 32'h0;  // 32'h690a796a;
    ram_cell[    4396] = 32'h0;  // 32'hb4f8dddd;
    ram_cell[    4397] = 32'h0;  // 32'hc185b55f;
    ram_cell[    4398] = 32'h0;  // 32'h94072a49;
    ram_cell[    4399] = 32'h0;  // 32'h89a184b3;
    ram_cell[    4400] = 32'h0;  // 32'hc5c3617e;
    ram_cell[    4401] = 32'h0;  // 32'h2fd7b519;
    ram_cell[    4402] = 32'h0;  // 32'h0f0d248a;
    ram_cell[    4403] = 32'h0;  // 32'hecf4075d;
    ram_cell[    4404] = 32'h0;  // 32'h013d0393;
    ram_cell[    4405] = 32'h0;  // 32'hd44f3502;
    ram_cell[    4406] = 32'h0;  // 32'haeb535ae;
    ram_cell[    4407] = 32'h0;  // 32'h3d341fac;
    ram_cell[    4408] = 32'h0;  // 32'ha4308956;
    ram_cell[    4409] = 32'h0;  // 32'h4bd41434;
    ram_cell[    4410] = 32'h0;  // 32'hc416678a;
    ram_cell[    4411] = 32'h0;  // 32'h2ebda68f;
    ram_cell[    4412] = 32'h0;  // 32'h2bbf9bef;
    ram_cell[    4413] = 32'h0;  // 32'hdc974119;
    ram_cell[    4414] = 32'h0;  // 32'h41e4899f;
    ram_cell[    4415] = 32'h0;  // 32'h2032311c;
    ram_cell[    4416] = 32'h0;  // 32'h332dbcd8;
    ram_cell[    4417] = 32'h0;  // 32'h8448b393;
    ram_cell[    4418] = 32'h0;  // 32'hd93f11ef;
    ram_cell[    4419] = 32'h0;  // 32'hcb09751a;
    ram_cell[    4420] = 32'h0;  // 32'h1f582ea5;
    ram_cell[    4421] = 32'h0;  // 32'haa3524a5;
    ram_cell[    4422] = 32'h0;  // 32'h134c61cc;
    ram_cell[    4423] = 32'h0;  // 32'h49081166;
    ram_cell[    4424] = 32'h0;  // 32'hb521255d;
    ram_cell[    4425] = 32'h0;  // 32'h59e7f67c;
    ram_cell[    4426] = 32'h0;  // 32'h2f127ec3;
    ram_cell[    4427] = 32'h0;  // 32'h72040577;
    ram_cell[    4428] = 32'h0;  // 32'h75c0dea0;
    ram_cell[    4429] = 32'h0;  // 32'h5c3a8934;
    ram_cell[    4430] = 32'h0;  // 32'h59a57f25;
    ram_cell[    4431] = 32'h0;  // 32'hb5a8b48d;
    ram_cell[    4432] = 32'h0;  // 32'h751f2181;
    ram_cell[    4433] = 32'h0;  // 32'h1e5a0610;
    ram_cell[    4434] = 32'h0;  // 32'hf9010595;
    ram_cell[    4435] = 32'h0;  // 32'h3777138d;
    ram_cell[    4436] = 32'h0;  // 32'h85b19ce7;
    ram_cell[    4437] = 32'h0;  // 32'h311e617f;
    ram_cell[    4438] = 32'h0;  // 32'hfbb96f77;
    ram_cell[    4439] = 32'h0;  // 32'h6342ce0e;
    ram_cell[    4440] = 32'h0;  // 32'h986ce0cc;
    ram_cell[    4441] = 32'h0;  // 32'h1ff71fbf;
    ram_cell[    4442] = 32'h0;  // 32'h5a84385a;
    ram_cell[    4443] = 32'h0;  // 32'h44946009;
    ram_cell[    4444] = 32'h0;  // 32'hbd4a5e47;
    ram_cell[    4445] = 32'h0;  // 32'hc633f302;
    ram_cell[    4446] = 32'h0;  // 32'h1f228354;
    ram_cell[    4447] = 32'h0;  // 32'h9c2da7e2;
    ram_cell[    4448] = 32'h0;  // 32'h9f4e2beb;
    ram_cell[    4449] = 32'h0;  // 32'h9b7a6fb3;
    ram_cell[    4450] = 32'h0;  // 32'h3294683c;
    ram_cell[    4451] = 32'h0;  // 32'h2e5a3447;
    ram_cell[    4452] = 32'h0;  // 32'h58f6307d;
    ram_cell[    4453] = 32'h0;  // 32'hbe8cbe79;
    ram_cell[    4454] = 32'h0;  // 32'h89b65971;
    ram_cell[    4455] = 32'h0;  // 32'ha421616a;
    ram_cell[    4456] = 32'h0;  // 32'hcaff689c;
    ram_cell[    4457] = 32'h0;  // 32'h2ec667e2;
    ram_cell[    4458] = 32'h0;  // 32'hc538a5d6;
    ram_cell[    4459] = 32'h0;  // 32'hc8483a60;
    ram_cell[    4460] = 32'h0;  // 32'h9486e58f;
    ram_cell[    4461] = 32'h0;  // 32'h72539d88;
    ram_cell[    4462] = 32'h0;  // 32'h6f76b9ac;
    ram_cell[    4463] = 32'h0;  // 32'h57654e7a;
    ram_cell[    4464] = 32'h0;  // 32'hb7a1edd4;
    ram_cell[    4465] = 32'h0;  // 32'h311d3d6b;
    ram_cell[    4466] = 32'h0;  // 32'h92e7b610;
    ram_cell[    4467] = 32'h0;  // 32'ha6fca518;
    ram_cell[    4468] = 32'h0;  // 32'h0f6c929c;
    ram_cell[    4469] = 32'h0;  // 32'h394f4a75;
    ram_cell[    4470] = 32'h0;  // 32'h9f406625;
    ram_cell[    4471] = 32'h0;  // 32'h2ac634cb;
    ram_cell[    4472] = 32'h0;  // 32'h7dd08993;
    ram_cell[    4473] = 32'h0;  // 32'h838f0ebb;
    ram_cell[    4474] = 32'h0;  // 32'h9e4e4fa7;
    ram_cell[    4475] = 32'h0;  // 32'h89561ab0;
    ram_cell[    4476] = 32'h0;  // 32'ha6b4006a;
    ram_cell[    4477] = 32'h0;  // 32'he1d68f1b;
    ram_cell[    4478] = 32'h0;  // 32'hb19e758e;
    ram_cell[    4479] = 32'h0;  // 32'ha2d62f5c;
    ram_cell[    4480] = 32'h0;  // 32'hf980d861;
    ram_cell[    4481] = 32'h0;  // 32'h941175f1;
    ram_cell[    4482] = 32'h0;  // 32'h57902399;
    ram_cell[    4483] = 32'h0;  // 32'h385a4d7b;
    ram_cell[    4484] = 32'h0;  // 32'h307af5e9;
    ram_cell[    4485] = 32'h0;  // 32'h41dee637;
    ram_cell[    4486] = 32'h0;  // 32'hc3c53bab;
    ram_cell[    4487] = 32'h0;  // 32'h33213e60;
    ram_cell[    4488] = 32'h0;  // 32'h16294da0;
    ram_cell[    4489] = 32'h0;  // 32'hb87066a0;
    ram_cell[    4490] = 32'h0;  // 32'h7ac3e44c;
    ram_cell[    4491] = 32'h0;  // 32'h82cc056e;
    ram_cell[    4492] = 32'h0;  // 32'hdccaafeb;
    ram_cell[    4493] = 32'h0;  // 32'hfcd2d7f7;
    ram_cell[    4494] = 32'h0;  // 32'h6648d908;
    ram_cell[    4495] = 32'h0;  // 32'hf5506296;
    ram_cell[    4496] = 32'h0;  // 32'h2ab6a478;
    ram_cell[    4497] = 32'h0;  // 32'h2c5c4fe2;
    ram_cell[    4498] = 32'h0;  // 32'h23167f47;
    ram_cell[    4499] = 32'h0;  // 32'hfdd2535a;
    ram_cell[    4500] = 32'h0;  // 32'h389def87;
    ram_cell[    4501] = 32'h0;  // 32'h288ef338;
    ram_cell[    4502] = 32'h0;  // 32'h8253d00c;
    ram_cell[    4503] = 32'h0;  // 32'h6d49b8ca;
    ram_cell[    4504] = 32'h0;  // 32'ha6e2e58a;
    ram_cell[    4505] = 32'h0;  // 32'hac4a3302;
    ram_cell[    4506] = 32'h0;  // 32'h009d20b2;
    ram_cell[    4507] = 32'h0;  // 32'h48455955;
    ram_cell[    4508] = 32'h0;  // 32'he1696f3e;
    ram_cell[    4509] = 32'h0;  // 32'hb765c364;
    ram_cell[    4510] = 32'h0;  // 32'h96d0de75;
    ram_cell[    4511] = 32'h0;  // 32'h53bc7f01;
    ram_cell[    4512] = 32'h0;  // 32'hf7757a67;
    ram_cell[    4513] = 32'h0;  // 32'h95751ab8;
    ram_cell[    4514] = 32'h0;  // 32'h86992a7d;
    ram_cell[    4515] = 32'h0;  // 32'h84d13756;
    ram_cell[    4516] = 32'h0;  // 32'haa50c3a5;
    ram_cell[    4517] = 32'h0;  // 32'hae4a8c67;
    ram_cell[    4518] = 32'h0;  // 32'h14dd6718;
    ram_cell[    4519] = 32'h0;  // 32'hf8fd046c;
    ram_cell[    4520] = 32'h0;  // 32'h55d8122f;
    ram_cell[    4521] = 32'h0;  // 32'h87a396fd;
    ram_cell[    4522] = 32'h0;  // 32'hb2823ffd;
    ram_cell[    4523] = 32'h0;  // 32'h0692755b;
    ram_cell[    4524] = 32'h0;  // 32'hcf0d659a;
    ram_cell[    4525] = 32'h0;  // 32'ha078bbf2;
    ram_cell[    4526] = 32'h0;  // 32'h3d7b4165;
    ram_cell[    4527] = 32'h0;  // 32'h8a4d9b5c;
    ram_cell[    4528] = 32'h0;  // 32'h35a2467d;
    ram_cell[    4529] = 32'h0;  // 32'hc14a66e7;
    ram_cell[    4530] = 32'h0;  // 32'hf9e47d0a;
    ram_cell[    4531] = 32'h0;  // 32'h5f7cffc9;
    ram_cell[    4532] = 32'h0;  // 32'h2163bdf1;
    ram_cell[    4533] = 32'h0;  // 32'h1a29a257;
    ram_cell[    4534] = 32'h0;  // 32'hd2ec8904;
    ram_cell[    4535] = 32'h0;  // 32'hee864a8b;
    ram_cell[    4536] = 32'h0;  // 32'hc0024031;
    ram_cell[    4537] = 32'h0;  // 32'h3e00effc;
    ram_cell[    4538] = 32'h0;  // 32'h2539a540;
    ram_cell[    4539] = 32'h0;  // 32'h9a3091a9;
    ram_cell[    4540] = 32'h0;  // 32'hf6ac914e;
    ram_cell[    4541] = 32'h0;  // 32'hd687c056;
    ram_cell[    4542] = 32'h0;  // 32'h67070906;
    ram_cell[    4543] = 32'h0;  // 32'hd6bcbbb8;
    ram_cell[    4544] = 32'h0;  // 32'h4578c56a;
    ram_cell[    4545] = 32'h0;  // 32'h250878b8;
    ram_cell[    4546] = 32'h0;  // 32'h5283fbb6;
    ram_cell[    4547] = 32'h0;  // 32'h13623472;
    ram_cell[    4548] = 32'h0;  // 32'h188e2df2;
    ram_cell[    4549] = 32'h0;  // 32'h08dcd26b;
    ram_cell[    4550] = 32'h0;  // 32'h66e02bbb;
    ram_cell[    4551] = 32'h0;  // 32'hf61cefe5;
    ram_cell[    4552] = 32'h0;  // 32'hfd7597ef;
    ram_cell[    4553] = 32'h0;  // 32'h96215417;
    ram_cell[    4554] = 32'h0;  // 32'hc7cd3637;
    ram_cell[    4555] = 32'h0;  // 32'hda10de4d;
    ram_cell[    4556] = 32'h0;  // 32'hbe79ea87;
    ram_cell[    4557] = 32'h0;  // 32'he89c0444;
    ram_cell[    4558] = 32'h0;  // 32'he48d5746;
    ram_cell[    4559] = 32'h0;  // 32'hfcaeccd3;
    ram_cell[    4560] = 32'h0;  // 32'h617e5c39;
    ram_cell[    4561] = 32'h0;  // 32'hc6133e88;
    ram_cell[    4562] = 32'h0;  // 32'h862eeb08;
    ram_cell[    4563] = 32'h0;  // 32'hd7999095;
    ram_cell[    4564] = 32'h0;  // 32'h11653665;
    ram_cell[    4565] = 32'h0;  // 32'hf7788c68;
    ram_cell[    4566] = 32'h0;  // 32'h945055de;
    ram_cell[    4567] = 32'h0;  // 32'h8bb65289;
    ram_cell[    4568] = 32'h0;  // 32'h081c65de;
    ram_cell[    4569] = 32'h0;  // 32'hfbbf231d;
    ram_cell[    4570] = 32'h0;  // 32'h1c24bae8;
    ram_cell[    4571] = 32'h0;  // 32'hf4cbdbde;
    ram_cell[    4572] = 32'h0;  // 32'h95e49526;
    ram_cell[    4573] = 32'h0;  // 32'hec131e06;
    ram_cell[    4574] = 32'h0;  // 32'h796bef00;
    ram_cell[    4575] = 32'h0;  // 32'h38685bac;
    ram_cell[    4576] = 32'h0;  // 32'h1601f0b7;
    ram_cell[    4577] = 32'h0;  // 32'h1b020491;
    ram_cell[    4578] = 32'h0;  // 32'h79529d1f;
    ram_cell[    4579] = 32'h0;  // 32'h8dbeda4c;
    ram_cell[    4580] = 32'h0;  // 32'h7e513f48;
    ram_cell[    4581] = 32'h0;  // 32'h42e33071;
    ram_cell[    4582] = 32'h0;  // 32'h8415e85d;
    ram_cell[    4583] = 32'h0;  // 32'h818dbe9d;
    ram_cell[    4584] = 32'h0;  // 32'h4b208955;
    ram_cell[    4585] = 32'h0;  // 32'h04d38ea2;
    ram_cell[    4586] = 32'h0;  // 32'hd62418e4;
    ram_cell[    4587] = 32'h0;  // 32'hc05a74d4;
    ram_cell[    4588] = 32'h0;  // 32'hb9f9bd8c;
    ram_cell[    4589] = 32'h0;  // 32'h5a742d56;
    ram_cell[    4590] = 32'h0;  // 32'h9bd78dc9;
    ram_cell[    4591] = 32'h0;  // 32'h58b984ae;
    ram_cell[    4592] = 32'h0;  // 32'ha4f6996c;
    ram_cell[    4593] = 32'h0;  // 32'h519188ac;
    ram_cell[    4594] = 32'h0;  // 32'h6944d8f7;
    ram_cell[    4595] = 32'h0;  // 32'h59886bd9;
    ram_cell[    4596] = 32'h0;  // 32'h1e97c4c4;
    ram_cell[    4597] = 32'h0;  // 32'h0f485728;
    ram_cell[    4598] = 32'h0;  // 32'h73c7d65f;
    ram_cell[    4599] = 32'h0;  // 32'h103bea06;
    ram_cell[    4600] = 32'h0;  // 32'hc4701cea;
    ram_cell[    4601] = 32'h0;  // 32'hb179affc;
    ram_cell[    4602] = 32'h0;  // 32'h0bd1fcc9;
    ram_cell[    4603] = 32'h0;  // 32'hcc3112cd;
    ram_cell[    4604] = 32'h0;  // 32'hdce4eab1;
    ram_cell[    4605] = 32'h0;  // 32'h7024dca2;
    ram_cell[    4606] = 32'h0;  // 32'h0558ed37;
    ram_cell[    4607] = 32'h0;  // 32'hc27e29b8;
    ram_cell[    4608] = 32'h0;  // 32'h9dceb892;
    ram_cell[    4609] = 32'h0;  // 32'h91748553;
    ram_cell[    4610] = 32'h0;  // 32'h13ad576d;
    ram_cell[    4611] = 32'h0;  // 32'hef067d80;
    ram_cell[    4612] = 32'h0;  // 32'h18a18230;
    ram_cell[    4613] = 32'h0;  // 32'hbbe6052a;
    ram_cell[    4614] = 32'h0;  // 32'h9a63594e;
    ram_cell[    4615] = 32'h0;  // 32'h6bf46a3e;
    ram_cell[    4616] = 32'h0;  // 32'h74c0807d;
    ram_cell[    4617] = 32'h0;  // 32'hf73b643e;
    ram_cell[    4618] = 32'h0;  // 32'h63d20b48;
    ram_cell[    4619] = 32'h0;  // 32'h2138eb14;
    ram_cell[    4620] = 32'h0;  // 32'h311d84ee;
    ram_cell[    4621] = 32'h0;  // 32'hf5a0fe2a;
    ram_cell[    4622] = 32'h0;  // 32'h9f3c6882;
    ram_cell[    4623] = 32'h0;  // 32'hb61479f4;
    ram_cell[    4624] = 32'h0;  // 32'h7c6eda77;
    ram_cell[    4625] = 32'h0;  // 32'h33c8c7b3;
    ram_cell[    4626] = 32'h0;  // 32'h7f3ff326;
    ram_cell[    4627] = 32'h0;  // 32'h697c1c64;
    ram_cell[    4628] = 32'h0;  // 32'h85504416;
    ram_cell[    4629] = 32'h0;  // 32'h82a0b399;
    ram_cell[    4630] = 32'h0;  // 32'hef371f1f;
    ram_cell[    4631] = 32'h0;  // 32'hd7e25802;
    ram_cell[    4632] = 32'h0;  // 32'h865e87d1;
    ram_cell[    4633] = 32'h0;  // 32'h95987485;
    ram_cell[    4634] = 32'h0;  // 32'haf370e53;
    ram_cell[    4635] = 32'h0;  // 32'h7d55df2e;
    ram_cell[    4636] = 32'h0;  // 32'hfbcb5e85;
    ram_cell[    4637] = 32'h0;  // 32'h92d48bf3;
    ram_cell[    4638] = 32'h0;  // 32'hefaebabe;
    ram_cell[    4639] = 32'h0;  // 32'h13ec7b6a;
    ram_cell[    4640] = 32'h0;  // 32'hd0eb2c2a;
    ram_cell[    4641] = 32'h0;  // 32'hd6fe026a;
    ram_cell[    4642] = 32'h0;  // 32'h60dd4e1f;
    ram_cell[    4643] = 32'h0;  // 32'h4907a3e8;
    ram_cell[    4644] = 32'h0;  // 32'h273ef324;
    ram_cell[    4645] = 32'h0;  // 32'hf5d17e86;
    ram_cell[    4646] = 32'h0;  // 32'h8d197592;
    ram_cell[    4647] = 32'h0;  // 32'h5e9f16da;
    ram_cell[    4648] = 32'h0;  // 32'hcca1c37b;
    ram_cell[    4649] = 32'h0;  // 32'hc3cfd397;
    ram_cell[    4650] = 32'h0;  // 32'he96ff691;
    ram_cell[    4651] = 32'h0;  // 32'hfb2b0590;
    ram_cell[    4652] = 32'h0;  // 32'h5bdf3c83;
    ram_cell[    4653] = 32'h0;  // 32'ha090562b;
    ram_cell[    4654] = 32'h0;  // 32'h8fb2caa4;
    ram_cell[    4655] = 32'h0;  // 32'h0d38aeb7;
    ram_cell[    4656] = 32'h0;  // 32'h0c819783;
    ram_cell[    4657] = 32'h0;  // 32'h914ad3a0;
    ram_cell[    4658] = 32'h0;  // 32'h67fc80cf;
    ram_cell[    4659] = 32'h0;  // 32'h786585a5;
    ram_cell[    4660] = 32'h0;  // 32'hd0611c65;
    ram_cell[    4661] = 32'h0;  // 32'h47d9758c;
    ram_cell[    4662] = 32'h0;  // 32'hab42a85e;
    ram_cell[    4663] = 32'h0;  // 32'h51dc56e3;
    ram_cell[    4664] = 32'h0;  // 32'hf0533896;
    ram_cell[    4665] = 32'h0;  // 32'h508be4b3;
    ram_cell[    4666] = 32'h0;  // 32'h7220f88f;
    ram_cell[    4667] = 32'h0;  // 32'hf43d1f24;
    ram_cell[    4668] = 32'h0;  // 32'h162eba45;
    ram_cell[    4669] = 32'h0;  // 32'h08f0dfe7;
    ram_cell[    4670] = 32'h0;  // 32'h032269aa;
    ram_cell[    4671] = 32'h0;  // 32'h1b5e1109;
    ram_cell[    4672] = 32'h0;  // 32'hc08bedc4;
    ram_cell[    4673] = 32'h0;  // 32'h796e33d4;
    ram_cell[    4674] = 32'h0;  // 32'hd3caccb2;
    ram_cell[    4675] = 32'h0;  // 32'h4eecf65c;
    ram_cell[    4676] = 32'h0;  // 32'h175259a8;
    ram_cell[    4677] = 32'h0;  // 32'hf909d1c9;
    ram_cell[    4678] = 32'h0;  // 32'h54448972;
    ram_cell[    4679] = 32'h0;  // 32'h272a99d0;
    ram_cell[    4680] = 32'h0;  // 32'h26a3fd48;
    ram_cell[    4681] = 32'h0;  // 32'hf4b68362;
    ram_cell[    4682] = 32'h0;  // 32'h673a7477;
    ram_cell[    4683] = 32'h0;  // 32'hc280141c;
    ram_cell[    4684] = 32'h0;  // 32'h405c1fde;
    ram_cell[    4685] = 32'h0;  // 32'h31a23f7d;
    ram_cell[    4686] = 32'h0;  // 32'hd22c3009;
    ram_cell[    4687] = 32'h0;  // 32'h2fca2ec7;
    ram_cell[    4688] = 32'h0;  // 32'hc6fbc07b;
    ram_cell[    4689] = 32'h0;  // 32'h4ef62d85;
    ram_cell[    4690] = 32'h0;  // 32'he4168baf;
    ram_cell[    4691] = 32'h0;  // 32'hfa1efe42;
    ram_cell[    4692] = 32'h0;  // 32'hcf56a773;
    ram_cell[    4693] = 32'h0;  // 32'h288182c2;
    ram_cell[    4694] = 32'h0;  // 32'h32930e9e;
    ram_cell[    4695] = 32'h0;  // 32'he6f74850;
    ram_cell[    4696] = 32'h0;  // 32'h3b76ad4b;
    ram_cell[    4697] = 32'h0;  // 32'h4f62bba2;
    ram_cell[    4698] = 32'h0;  // 32'h0e4486da;
    ram_cell[    4699] = 32'h0;  // 32'h3d04fe2d;
    ram_cell[    4700] = 32'h0;  // 32'hc4d9d209;
    ram_cell[    4701] = 32'h0;  // 32'h065dc2c1;
    ram_cell[    4702] = 32'h0;  // 32'h2d89a408;
    ram_cell[    4703] = 32'h0;  // 32'hb7546081;
    ram_cell[    4704] = 32'h0;  // 32'haea02030;
    ram_cell[    4705] = 32'h0;  // 32'hcdf9ef6f;
    ram_cell[    4706] = 32'h0;  // 32'had261d32;
    ram_cell[    4707] = 32'h0;  // 32'hec0817c0;
    ram_cell[    4708] = 32'h0;  // 32'h638f9526;
    ram_cell[    4709] = 32'h0;  // 32'ha8fbf69b;
    ram_cell[    4710] = 32'h0;  // 32'h389e9a69;
    ram_cell[    4711] = 32'h0;  // 32'hd035d6d1;
    ram_cell[    4712] = 32'h0;  // 32'h14516f3e;
    ram_cell[    4713] = 32'h0;  // 32'h577b85a9;
    ram_cell[    4714] = 32'h0;  // 32'h07af2a28;
    ram_cell[    4715] = 32'h0;  // 32'h05a3dcff;
    ram_cell[    4716] = 32'h0;  // 32'h39723b71;
    ram_cell[    4717] = 32'h0;  // 32'h1020d00e;
    ram_cell[    4718] = 32'h0;  // 32'he4b521d5;
    ram_cell[    4719] = 32'h0;  // 32'h031043e5;
    ram_cell[    4720] = 32'h0;  // 32'h1676b345;
    ram_cell[    4721] = 32'h0;  // 32'hb56b750d;
    ram_cell[    4722] = 32'h0;  // 32'h7bc6347f;
    ram_cell[    4723] = 32'h0;  // 32'heebcb75b;
    ram_cell[    4724] = 32'h0;  // 32'h5b9c4bb0;
    ram_cell[    4725] = 32'h0;  // 32'h58589311;
    ram_cell[    4726] = 32'h0;  // 32'h68933d02;
    ram_cell[    4727] = 32'h0;  // 32'h07b0893e;
    ram_cell[    4728] = 32'h0;  // 32'h11c9f010;
    ram_cell[    4729] = 32'h0;  // 32'h390485c8;
    ram_cell[    4730] = 32'h0;  // 32'h7cd556ee;
    ram_cell[    4731] = 32'h0;  // 32'h0ba0463b;
    ram_cell[    4732] = 32'h0;  // 32'h37d208b8;
    ram_cell[    4733] = 32'h0;  // 32'h6d7d526b;
    ram_cell[    4734] = 32'h0;  // 32'h3327bf8e;
    ram_cell[    4735] = 32'h0;  // 32'hd9571619;
    ram_cell[    4736] = 32'h0;  // 32'hb066026c;
    ram_cell[    4737] = 32'h0;  // 32'he9de9814;
    ram_cell[    4738] = 32'h0;  // 32'hfff1fd09;
    ram_cell[    4739] = 32'h0;  // 32'h4ee12498;
    ram_cell[    4740] = 32'h0;  // 32'h9e2f886b;
    ram_cell[    4741] = 32'h0;  // 32'h1800ab01;
    ram_cell[    4742] = 32'h0;  // 32'hbc6517af;
    ram_cell[    4743] = 32'h0;  // 32'hcc09a913;
    ram_cell[    4744] = 32'h0;  // 32'h30ab48d1;
    ram_cell[    4745] = 32'h0;  // 32'h640508b5;
    ram_cell[    4746] = 32'h0;  // 32'hbb489ff0;
    ram_cell[    4747] = 32'h0;  // 32'he442d594;
    ram_cell[    4748] = 32'h0;  // 32'h6ef50f64;
    ram_cell[    4749] = 32'h0;  // 32'h3aae34c2;
    ram_cell[    4750] = 32'h0;  // 32'hd68f6c2a;
    ram_cell[    4751] = 32'h0;  // 32'hba1aa448;
    ram_cell[    4752] = 32'h0;  // 32'h9205630a;
    ram_cell[    4753] = 32'h0;  // 32'h33d959f2;
    ram_cell[    4754] = 32'h0;  // 32'h56ba74e0;
    ram_cell[    4755] = 32'h0;  // 32'h9eda7cd4;
    ram_cell[    4756] = 32'h0;  // 32'hac955131;
    ram_cell[    4757] = 32'h0;  // 32'h3de9ed29;
    ram_cell[    4758] = 32'h0;  // 32'h4014567e;
    ram_cell[    4759] = 32'h0;  // 32'h58f2eb94;
    ram_cell[    4760] = 32'h0;  // 32'h771505cb;
    ram_cell[    4761] = 32'h0;  // 32'he6f4af8b;
    ram_cell[    4762] = 32'h0;  // 32'h10b34d2f;
    ram_cell[    4763] = 32'h0;  // 32'hef0eb618;
    ram_cell[    4764] = 32'h0;  // 32'hceb6f1cc;
    ram_cell[    4765] = 32'h0;  // 32'h3ebf4f9f;
    ram_cell[    4766] = 32'h0;  // 32'h98eb3fe2;
    ram_cell[    4767] = 32'h0;  // 32'hc4b2e491;
    ram_cell[    4768] = 32'h0;  // 32'h637e8e91;
    ram_cell[    4769] = 32'h0;  // 32'hebc9b8c7;
    ram_cell[    4770] = 32'h0;  // 32'haa40d690;
    ram_cell[    4771] = 32'h0;  // 32'h1fb379dc;
    ram_cell[    4772] = 32'h0;  // 32'h9e82ee70;
    ram_cell[    4773] = 32'h0;  // 32'hff9778dc;
    ram_cell[    4774] = 32'h0;  // 32'hae7deb87;
    ram_cell[    4775] = 32'h0;  // 32'h2a80629b;
    ram_cell[    4776] = 32'h0;  // 32'hc7f2e9f9;
    ram_cell[    4777] = 32'h0;  // 32'hfd16eb4d;
    ram_cell[    4778] = 32'h0;  // 32'ha8ab1d0b;
    ram_cell[    4779] = 32'h0;  // 32'h4b455262;
    ram_cell[    4780] = 32'h0;  // 32'h0f8dce3b;
    ram_cell[    4781] = 32'h0;  // 32'hb52afb33;
    ram_cell[    4782] = 32'h0;  // 32'h93e1a122;
    ram_cell[    4783] = 32'h0;  // 32'h4557d807;
    ram_cell[    4784] = 32'h0;  // 32'hdacfe39b;
    ram_cell[    4785] = 32'h0;  // 32'h3fbfebea;
    ram_cell[    4786] = 32'h0;  // 32'h58cee0a0;
    ram_cell[    4787] = 32'h0;  // 32'h26925943;
    ram_cell[    4788] = 32'h0;  // 32'h84f04fbf;
    ram_cell[    4789] = 32'h0;  // 32'h43ba6ed8;
    ram_cell[    4790] = 32'h0;  // 32'h0a3e498f;
    ram_cell[    4791] = 32'h0;  // 32'hb9db2b2a;
    ram_cell[    4792] = 32'h0;  // 32'ha11234d1;
    ram_cell[    4793] = 32'h0;  // 32'h5388ed08;
    ram_cell[    4794] = 32'h0;  // 32'h79f0b83a;
    ram_cell[    4795] = 32'h0;  // 32'hd82450a7;
    ram_cell[    4796] = 32'h0;  // 32'h2acf6f9a;
    ram_cell[    4797] = 32'h0;  // 32'hc063b615;
    ram_cell[    4798] = 32'h0;  // 32'hde1fc3bb;
    ram_cell[    4799] = 32'h0;  // 32'he182ffb7;
    ram_cell[    4800] = 32'h0;  // 32'hd529bb57;
    ram_cell[    4801] = 32'h0;  // 32'h6817f8be;
    ram_cell[    4802] = 32'h0;  // 32'ha6b48440;
    ram_cell[    4803] = 32'h0;  // 32'h9ae4a46e;
    ram_cell[    4804] = 32'h0;  // 32'h7950edd8;
    ram_cell[    4805] = 32'h0;  // 32'h6f244dfc;
    ram_cell[    4806] = 32'h0;  // 32'h5496b295;
    ram_cell[    4807] = 32'h0;  // 32'hef3c56bb;
    ram_cell[    4808] = 32'h0;  // 32'h290bbea3;
    ram_cell[    4809] = 32'h0;  // 32'h0addf7ad;
    ram_cell[    4810] = 32'h0;  // 32'h36845cf7;
    ram_cell[    4811] = 32'h0;  // 32'h831568d2;
    ram_cell[    4812] = 32'h0;  // 32'hc2a17708;
    ram_cell[    4813] = 32'h0;  // 32'h9d00c26d;
    ram_cell[    4814] = 32'h0;  // 32'h6384e35f;
    ram_cell[    4815] = 32'h0;  // 32'hdda856b4;
    ram_cell[    4816] = 32'h0;  // 32'h57ac184c;
    ram_cell[    4817] = 32'h0;  // 32'h601ed9bf;
    ram_cell[    4818] = 32'h0;  // 32'h4bdab182;
    ram_cell[    4819] = 32'h0;  // 32'hd3becac6;
    ram_cell[    4820] = 32'h0;  // 32'habcac90a;
    ram_cell[    4821] = 32'h0;  // 32'heb26738a;
    ram_cell[    4822] = 32'h0;  // 32'h3a5fd6f1;
    ram_cell[    4823] = 32'h0;  // 32'h841ebb42;
    ram_cell[    4824] = 32'h0;  // 32'he00e4077;
    ram_cell[    4825] = 32'h0;  // 32'hac4883ed;
    ram_cell[    4826] = 32'h0;  // 32'hea9127e8;
    ram_cell[    4827] = 32'h0;  // 32'h85c56fae;
    ram_cell[    4828] = 32'h0;  // 32'h552f195d;
    ram_cell[    4829] = 32'h0;  // 32'h78ae8e4e;
    ram_cell[    4830] = 32'h0;  // 32'h8e3f66cb;
    ram_cell[    4831] = 32'h0;  // 32'h04702f6b;
    ram_cell[    4832] = 32'h0;  // 32'hf7be4169;
    ram_cell[    4833] = 32'h0;  // 32'h17fee7e9;
    ram_cell[    4834] = 32'h0;  // 32'h0215746d;
    ram_cell[    4835] = 32'h0;  // 32'hff9d9b36;
    ram_cell[    4836] = 32'h0;  // 32'h99f30c26;
    ram_cell[    4837] = 32'h0;  // 32'h66514573;
    ram_cell[    4838] = 32'h0;  // 32'h5044ac5e;
    ram_cell[    4839] = 32'h0;  // 32'h0ed11227;
    ram_cell[    4840] = 32'h0;  // 32'hb8dd3bfe;
    ram_cell[    4841] = 32'h0;  // 32'ha73ca7b8;
    ram_cell[    4842] = 32'h0;  // 32'hb4157237;
    ram_cell[    4843] = 32'h0;  // 32'h7eabceb3;
    ram_cell[    4844] = 32'h0;  // 32'h73d326a1;
    ram_cell[    4845] = 32'h0;  // 32'hba484557;
    ram_cell[    4846] = 32'h0;  // 32'h8f24019f;
    ram_cell[    4847] = 32'h0;  // 32'h986e6674;
    ram_cell[    4848] = 32'h0;  // 32'h97f2ade2;
    ram_cell[    4849] = 32'h0;  // 32'h96068d32;
    ram_cell[    4850] = 32'h0;  // 32'h22ed3d0c;
    ram_cell[    4851] = 32'h0;  // 32'h7bd3db60;
    ram_cell[    4852] = 32'h0;  // 32'he925da3d;
    ram_cell[    4853] = 32'h0;  // 32'hf9b61074;
    ram_cell[    4854] = 32'h0;  // 32'ha9c470f7;
    ram_cell[    4855] = 32'h0;  // 32'hd0ec2ed3;
    ram_cell[    4856] = 32'h0;  // 32'hd0825fa1;
    ram_cell[    4857] = 32'h0;  // 32'h40fa5226;
    ram_cell[    4858] = 32'h0;  // 32'h84a2b8ec;
    ram_cell[    4859] = 32'h0;  // 32'h9bb684a0;
    ram_cell[    4860] = 32'h0;  // 32'hfcd7b28d;
    ram_cell[    4861] = 32'h0;  // 32'h79cb3b41;
    ram_cell[    4862] = 32'h0;  // 32'h1e052350;
    ram_cell[    4863] = 32'h0;  // 32'h0099942d;
    ram_cell[    4864] = 32'h0;  // 32'h2293f833;
    ram_cell[    4865] = 32'h0;  // 32'hbf073cd7;
    ram_cell[    4866] = 32'h0;  // 32'ha4ec614b;
    ram_cell[    4867] = 32'h0;  // 32'hd05e6d7a;
    ram_cell[    4868] = 32'h0;  // 32'hacb56975;
    ram_cell[    4869] = 32'h0;  // 32'h9ab8a18c;
    ram_cell[    4870] = 32'h0;  // 32'hed7f5705;
    ram_cell[    4871] = 32'h0;  // 32'h235f7b76;
    ram_cell[    4872] = 32'h0;  // 32'h97b453df;
    ram_cell[    4873] = 32'h0;  // 32'he35c146a;
    ram_cell[    4874] = 32'h0;  // 32'h7ee9e748;
    ram_cell[    4875] = 32'h0;  // 32'h2f2ff9cd;
    ram_cell[    4876] = 32'h0;  // 32'h3f840c30;
    ram_cell[    4877] = 32'h0;  // 32'h365adfc5;
    ram_cell[    4878] = 32'h0;  // 32'hbdc02ad3;
    ram_cell[    4879] = 32'h0;  // 32'h1e0750c6;
    ram_cell[    4880] = 32'h0;  // 32'hc7305077;
    ram_cell[    4881] = 32'h0;  // 32'h2f04e2c9;
    ram_cell[    4882] = 32'h0;  // 32'h5e7b9285;
    ram_cell[    4883] = 32'h0;  // 32'h02522561;
    ram_cell[    4884] = 32'h0;  // 32'hc4eaded5;
    ram_cell[    4885] = 32'h0;  // 32'h890d4680;
    ram_cell[    4886] = 32'h0;  // 32'hc3ac3a8d;
    ram_cell[    4887] = 32'h0;  // 32'h9093876c;
    ram_cell[    4888] = 32'h0;  // 32'h20cb655a;
    ram_cell[    4889] = 32'h0;  // 32'h4c2f8858;
    ram_cell[    4890] = 32'h0;  // 32'h6268cf7a;
    ram_cell[    4891] = 32'h0;  // 32'h43d89f3e;
    ram_cell[    4892] = 32'h0;  // 32'h1fa0b3c4;
    ram_cell[    4893] = 32'h0;  // 32'h582d9817;
    ram_cell[    4894] = 32'h0;  // 32'ha5056f68;
    ram_cell[    4895] = 32'h0;  // 32'hd29425b0;
    ram_cell[    4896] = 32'h0;  // 32'hacb961f1;
    ram_cell[    4897] = 32'h0;  // 32'h97dfdda2;
    ram_cell[    4898] = 32'h0;  // 32'h2dbd474d;
    ram_cell[    4899] = 32'h0;  // 32'h25c70d2c;
    ram_cell[    4900] = 32'h0;  // 32'hb2317caf;
    ram_cell[    4901] = 32'h0;  // 32'h11f1d887;
    ram_cell[    4902] = 32'h0;  // 32'h79336795;
    ram_cell[    4903] = 32'h0;  // 32'h2f4fb776;
    ram_cell[    4904] = 32'h0;  // 32'h8131bf0e;
    ram_cell[    4905] = 32'h0;  // 32'h7e153f8f;
    ram_cell[    4906] = 32'h0;  // 32'h6129dc83;
    ram_cell[    4907] = 32'h0;  // 32'h717f2bd7;
    ram_cell[    4908] = 32'h0;  // 32'h1e2df2cf;
    ram_cell[    4909] = 32'h0;  // 32'h9b0595cd;
    ram_cell[    4910] = 32'h0;  // 32'h8cb25941;
    ram_cell[    4911] = 32'h0;  // 32'he840954b;
    ram_cell[    4912] = 32'h0;  // 32'hcf5f2763;
    ram_cell[    4913] = 32'h0;  // 32'hb6c26638;
    ram_cell[    4914] = 32'h0;  // 32'he3f2615c;
    ram_cell[    4915] = 32'h0;  // 32'h706a11ef;
    ram_cell[    4916] = 32'h0;  // 32'h9d62f823;
    ram_cell[    4917] = 32'h0;  // 32'h6b2eb7fc;
    ram_cell[    4918] = 32'h0;  // 32'h1be4c6d9;
    ram_cell[    4919] = 32'h0;  // 32'hf404a955;
    ram_cell[    4920] = 32'h0;  // 32'he4ffe017;
    ram_cell[    4921] = 32'h0;  // 32'h470db7fd;
    ram_cell[    4922] = 32'h0;  // 32'hd38a0f67;
    ram_cell[    4923] = 32'h0;  // 32'he182eed9;
    ram_cell[    4924] = 32'h0;  // 32'had9359ae;
    ram_cell[    4925] = 32'h0;  // 32'h368ac9a7;
    ram_cell[    4926] = 32'h0;  // 32'h4b1a2f99;
    ram_cell[    4927] = 32'h0;  // 32'h9fea7e0b;
    ram_cell[    4928] = 32'h0;  // 32'ha77c5a64;
    ram_cell[    4929] = 32'h0;  // 32'he478ae11;
    ram_cell[    4930] = 32'h0;  // 32'h1a0eda9c;
    ram_cell[    4931] = 32'h0;  // 32'hf8ee64cc;
    ram_cell[    4932] = 32'h0;  // 32'hf23b983a;
    ram_cell[    4933] = 32'h0;  // 32'hf8601909;
    ram_cell[    4934] = 32'h0;  // 32'h6d769ef9;
    ram_cell[    4935] = 32'h0;  // 32'ha2dc15c1;
    ram_cell[    4936] = 32'h0;  // 32'hcf048fb0;
    ram_cell[    4937] = 32'h0;  // 32'h708f03f8;
    ram_cell[    4938] = 32'h0;  // 32'hfe6358d7;
    ram_cell[    4939] = 32'h0;  // 32'h24db0bd4;
    ram_cell[    4940] = 32'h0;  // 32'h68c17811;
    ram_cell[    4941] = 32'h0;  // 32'hac7e0948;
    ram_cell[    4942] = 32'h0;  // 32'h0e6788c4;
    ram_cell[    4943] = 32'h0;  // 32'h354022b2;
    ram_cell[    4944] = 32'h0;  // 32'hb8a03ba4;
    ram_cell[    4945] = 32'h0;  // 32'h057c7e57;
    ram_cell[    4946] = 32'h0;  // 32'he65f1d6c;
    ram_cell[    4947] = 32'h0;  // 32'h36fbfb12;
    ram_cell[    4948] = 32'h0;  // 32'h6cbd382c;
    ram_cell[    4949] = 32'h0;  // 32'h93b8e1dc;
    ram_cell[    4950] = 32'h0;  // 32'h5eeae606;
    ram_cell[    4951] = 32'h0;  // 32'h7594c305;
    ram_cell[    4952] = 32'h0;  // 32'h64384db2;
    ram_cell[    4953] = 32'h0;  // 32'hbe92db35;
    ram_cell[    4954] = 32'h0;  // 32'hc4e2ee56;
    ram_cell[    4955] = 32'h0;  // 32'hde996a5c;
    ram_cell[    4956] = 32'h0;  // 32'hdff94f58;
    ram_cell[    4957] = 32'h0;  // 32'hef89b1a0;
    ram_cell[    4958] = 32'h0;  // 32'h730d1361;
    ram_cell[    4959] = 32'h0;  // 32'h1520a0fa;
    ram_cell[    4960] = 32'h0;  // 32'h44e80a30;
    ram_cell[    4961] = 32'h0;  // 32'h7b38a0d9;
    ram_cell[    4962] = 32'h0;  // 32'hf254b8d8;
    ram_cell[    4963] = 32'h0;  // 32'h07116dae;
    ram_cell[    4964] = 32'h0;  // 32'h684d5c10;
    ram_cell[    4965] = 32'h0;  // 32'h5864d350;
    ram_cell[    4966] = 32'h0;  // 32'hb8d16279;
    ram_cell[    4967] = 32'h0;  // 32'h76b4d180;
    ram_cell[    4968] = 32'h0;  // 32'h7a41a2d6;
    ram_cell[    4969] = 32'h0;  // 32'h6355d7a6;
    ram_cell[    4970] = 32'h0;  // 32'h128c98c7;
    ram_cell[    4971] = 32'h0;  // 32'hd3473a1a;
    ram_cell[    4972] = 32'h0;  // 32'h9ade7152;
    ram_cell[    4973] = 32'h0;  // 32'h2fce49fe;
    ram_cell[    4974] = 32'h0;  // 32'hb3c7a9cd;
    ram_cell[    4975] = 32'h0;  // 32'hdf11d3ee;
    ram_cell[    4976] = 32'h0;  // 32'h658a6b7c;
    ram_cell[    4977] = 32'h0;  // 32'h0491bc54;
    ram_cell[    4978] = 32'h0;  // 32'h4ce1e27f;
    ram_cell[    4979] = 32'h0;  // 32'h90b50c12;
    ram_cell[    4980] = 32'h0;  // 32'h45888ce5;
    ram_cell[    4981] = 32'h0;  // 32'hee331a0f;
    ram_cell[    4982] = 32'h0;  // 32'hcbc461df;
    ram_cell[    4983] = 32'h0;  // 32'h62bb45f1;
    ram_cell[    4984] = 32'h0;  // 32'hce3c02f4;
    ram_cell[    4985] = 32'h0;  // 32'hc93ecc88;
    ram_cell[    4986] = 32'h0;  // 32'h08bf6e7b;
    ram_cell[    4987] = 32'h0;  // 32'hd6da9aa8;
    ram_cell[    4988] = 32'h0;  // 32'h008bca8a;
    ram_cell[    4989] = 32'h0;  // 32'hd4de82be;
    ram_cell[    4990] = 32'h0;  // 32'hd3f2643f;
    ram_cell[    4991] = 32'h0;  // 32'h74842811;
    ram_cell[    4992] = 32'h0;  // 32'h6b98597e;
    ram_cell[    4993] = 32'h0;  // 32'hca75bb75;
    ram_cell[    4994] = 32'h0;  // 32'hacb69c53;
    ram_cell[    4995] = 32'h0;  // 32'h6bb42736;
    ram_cell[    4996] = 32'h0;  // 32'h7816259b;
    ram_cell[    4997] = 32'h0;  // 32'h94ddbc06;
    ram_cell[    4998] = 32'h0;  // 32'hbec36a30;
    ram_cell[    4999] = 32'h0;  // 32'h4f988525;
    ram_cell[    5000] = 32'h0;  // 32'h736abcde;
    ram_cell[    5001] = 32'h0;  // 32'h62aef779;
    ram_cell[    5002] = 32'h0;  // 32'h30a26fc7;
    ram_cell[    5003] = 32'h0;  // 32'h8e404ba6;
    ram_cell[    5004] = 32'h0;  // 32'h96cc49a8;
    ram_cell[    5005] = 32'h0;  // 32'hd2aca395;
    ram_cell[    5006] = 32'h0;  // 32'h5038826d;
    ram_cell[    5007] = 32'h0;  // 32'hec843eaa;
    ram_cell[    5008] = 32'h0;  // 32'hcc8f3559;
    ram_cell[    5009] = 32'h0;  // 32'hebdd2973;
    ram_cell[    5010] = 32'h0;  // 32'h562d8d34;
    ram_cell[    5011] = 32'h0;  // 32'hdd8efd79;
    ram_cell[    5012] = 32'h0;  // 32'h5b204da9;
    ram_cell[    5013] = 32'h0;  // 32'h16502b30;
    ram_cell[    5014] = 32'h0;  // 32'h0ec50a96;
    ram_cell[    5015] = 32'h0;  // 32'h858ae8ec;
    ram_cell[    5016] = 32'h0;  // 32'h74351c4b;
    ram_cell[    5017] = 32'h0;  // 32'ha8ac2af1;
    ram_cell[    5018] = 32'h0;  // 32'hffdb2ea8;
    ram_cell[    5019] = 32'h0;  // 32'hdfba4d01;
    ram_cell[    5020] = 32'h0;  // 32'h75a9f4b6;
    ram_cell[    5021] = 32'h0;  // 32'hcad7e9cb;
    ram_cell[    5022] = 32'h0;  // 32'h92899070;
    ram_cell[    5023] = 32'h0;  // 32'h930c6919;
    ram_cell[    5024] = 32'h0;  // 32'h43164e96;
    ram_cell[    5025] = 32'h0;  // 32'h976bbbab;
    ram_cell[    5026] = 32'h0;  // 32'h563c02f9;
    ram_cell[    5027] = 32'h0;  // 32'h3f7ab930;
    ram_cell[    5028] = 32'h0;  // 32'hb5254b09;
    ram_cell[    5029] = 32'h0;  // 32'ha16db001;
    ram_cell[    5030] = 32'h0;  // 32'h3022cef0;
    ram_cell[    5031] = 32'h0;  // 32'h0d5b0c0c;
    ram_cell[    5032] = 32'h0;  // 32'h9c998681;
    ram_cell[    5033] = 32'h0;  // 32'hf7217d60;
    ram_cell[    5034] = 32'h0;  // 32'h70f7927f;
    ram_cell[    5035] = 32'h0;  // 32'h6b1e88a6;
    ram_cell[    5036] = 32'h0;  // 32'h1b3ed00a;
    ram_cell[    5037] = 32'h0;  // 32'h0fc1c504;
    ram_cell[    5038] = 32'h0;  // 32'h23978bc1;
    ram_cell[    5039] = 32'h0;  // 32'h80330d95;
    ram_cell[    5040] = 32'h0;  // 32'ha004cc11;
    ram_cell[    5041] = 32'h0;  // 32'h52d9c4d0;
    ram_cell[    5042] = 32'h0;  // 32'hc35923d0;
    ram_cell[    5043] = 32'h0;  // 32'h5f1c0979;
    ram_cell[    5044] = 32'h0;  // 32'h26d5a3a4;
    ram_cell[    5045] = 32'h0;  // 32'hfc03cc0c;
    ram_cell[    5046] = 32'h0;  // 32'h20626fc9;
    ram_cell[    5047] = 32'h0;  // 32'h9e5e52f4;
    ram_cell[    5048] = 32'h0;  // 32'hbbad8fb8;
    ram_cell[    5049] = 32'h0;  // 32'h5b33c77a;
    ram_cell[    5050] = 32'h0;  // 32'h72757789;
    ram_cell[    5051] = 32'h0;  // 32'h2b25b689;
    ram_cell[    5052] = 32'h0;  // 32'h079ccdaf;
    ram_cell[    5053] = 32'h0;  // 32'hde61446f;
    ram_cell[    5054] = 32'h0;  // 32'h1f675832;
    ram_cell[    5055] = 32'h0;  // 32'h1ba348d8;
    ram_cell[    5056] = 32'h0;  // 32'h1f5f8579;
    ram_cell[    5057] = 32'h0;  // 32'h0718f869;
    ram_cell[    5058] = 32'h0;  // 32'h7f74a1c1;
    ram_cell[    5059] = 32'h0;  // 32'hb93c418c;
    ram_cell[    5060] = 32'h0;  // 32'hfcc7ed99;
    ram_cell[    5061] = 32'h0;  // 32'h23df8932;
    ram_cell[    5062] = 32'h0;  // 32'h659c0ca6;
    ram_cell[    5063] = 32'h0;  // 32'hc5fbc64e;
    ram_cell[    5064] = 32'h0;  // 32'hea5e067b;
    ram_cell[    5065] = 32'h0;  // 32'hb7e8bb25;
    ram_cell[    5066] = 32'h0;  // 32'he794d8f2;
    ram_cell[    5067] = 32'h0;  // 32'h5f6d5d55;
    ram_cell[    5068] = 32'h0;  // 32'h54c22dfe;
    ram_cell[    5069] = 32'h0;  // 32'hc8eeb38b;
    ram_cell[    5070] = 32'h0;  // 32'h1206d994;
    ram_cell[    5071] = 32'h0;  // 32'hfeb37357;
    ram_cell[    5072] = 32'h0;  // 32'h27075ee4;
    ram_cell[    5073] = 32'h0;  // 32'hfa061664;
    ram_cell[    5074] = 32'h0;  // 32'h4b865568;
    ram_cell[    5075] = 32'h0;  // 32'h8a3f8e67;
    ram_cell[    5076] = 32'h0;  // 32'h4ac1fe3f;
    ram_cell[    5077] = 32'h0;  // 32'h541018b8;
    ram_cell[    5078] = 32'h0;  // 32'he5a09ec4;
    ram_cell[    5079] = 32'h0;  // 32'h3dcc610e;
    ram_cell[    5080] = 32'h0;  // 32'h02e16aa1;
    ram_cell[    5081] = 32'h0;  // 32'h00a8b2dd;
    ram_cell[    5082] = 32'h0;  // 32'hf94eccc4;
    ram_cell[    5083] = 32'h0;  // 32'h85af8b50;
    ram_cell[    5084] = 32'h0;  // 32'h077bd750;
    ram_cell[    5085] = 32'h0;  // 32'hbeb587a8;
    ram_cell[    5086] = 32'h0;  // 32'h0e921abb;
    ram_cell[    5087] = 32'h0;  // 32'h310a44d7;
    ram_cell[    5088] = 32'h0;  // 32'hacfe0d77;
    ram_cell[    5089] = 32'h0;  // 32'h5caafb2b;
    ram_cell[    5090] = 32'h0;  // 32'h34f68e54;
    ram_cell[    5091] = 32'h0;  // 32'h17d00461;
    ram_cell[    5092] = 32'h0;  // 32'h462941b9;
    ram_cell[    5093] = 32'h0;  // 32'h59ec8506;
    ram_cell[    5094] = 32'h0;  // 32'h46f84425;
    ram_cell[    5095] = 32'h0;  // 32'hd3f588d5;
    ram_cell[    5096] = 32'h0;  // 32'h63a7524f;
    ram_cell[    5097] = 32'h0;  // 32'h2f243067;
    ram_cell[    5098] = 32'h0;  // 32'hb0c57ad3;
    ram_cell[    5099] = 32'h0;  // 32'h478986c8;
    ram_cell[    5100] = 32'h0;  // 32'h2c96ef62;
    ram_cell[    5101] = 32'h0;  // 32'hff68c55b;
    ram_cell[    5102] = 32'h0;  // 32'hda5a350b;
    ram_cell[    5103] = 32'h0;  // 32'he173f225;
    ram_cell[    5104] = 32'h0;  // 32'h4fd3e42e;
    ram_cell[    5105] = 32'h0;  // 32'h3ec4cdc5;
    ram_cell[    5106] = 32'h0;  // 32'haee9c2b1;
    ram_cell[    5107] = 32'h0;  // 32'h4eaaad2d;
    ram_cell[    5108] = 32'h0;  // 32'hacadfb0d;
    ram_cell[    5109] = 32'h0;  // 32'h2ea75304;
    ram_cell[    5110] = 32'h0;  // 32'h980de295;
    ram_cell[    5111] = 32'h0;  // 32'h08451580;
    ram_cell[    5112] = 32'h0;  // 32'h5fa9aa07;
    ram_cell[    5113] = 32'h0;  // 32'h7c17df24;
    ram_cell[    5114] = 32'h0;  // 32'h01dfd715;
    ram_cell[    5115] = 32'h0;  // 32'h831a5291;
    ram_cell[    5116] = 32'h0;  // 32'he2355419;
    ram_cell[    5117] = 32'h0;  // 32'h01672ac1;
    ram_cell[    5118] = 32'h0;  // 32'hba9dbff2;
    ram_cell[    5119] = 32'h0;  // 32'h816c0db9;
    ram_cell[    5120] = 32'h0;  // 32'h92935807;
    ram_cell[    5121] = 32'h0;  // 32'hb51062c7;
    ram_cell[    5122] = 32'h0;  // 32'h5e9bea5a;
    ram_cell[    5123] = 32'h0;  // 32'h495989ce;
    ram_cell[    5124] = 32'h0;  // 32'h27261462;
    ram_cell[    5125] = 32'h0;  // 32'h5b33cd9b;
    ram_cell[    5126] = 32'h0;  // 32'h65cb64cb;
    ram_cell[    5127] = 32'h0;  // 32'ha1dd1b83;
    ram_cell[    5128] = 32'h0;  // 32'h437fd503;
    ram_cell[    5129] = 32'h0;  // 32'h09a09574;
    ram_cell[    5130] = 32'h0;  // 32'h00d421ab;
    ram_cell[    5131] = 32'h0;  // 32'he9afda0c;
    ram_cell[    5132] = 32'h0;  // 32'h19a2cf48;
    ram_cell[    5133] = 32'h0;  // 32'h05068e69;
    ram_cell[    5134] = 32'h0;  // 32'hd93255ff;
    ram_cell[    5135] = 32'h0;  // 32'he4fe6bbe;
    ram_cell[    5136] = 32'h0;  // 32'he782e51f;
    ram_cell[    5137] = 32'h0;  // 32'he17c91c8;
    ram_cell[    5138] = 32'h0;  // 32'he11a8273;
    ram_cell[    5139] = 32'h0;  // 32'hc4501aed;
    ram_cell[    5140] = 32'h0;  // 32'h6ca608c0;
    ram_cell[    5141] = 32'h0;  // 32'h87456682;
    ram_cell[    5142] = 32'h0;  // 32'heab2df72;
    ram_cell[    5143] = 32'h0;  // 32'h93cda64b;
    ram_cell[    5144] = 32'h0;  // 32'h2aee4d12;
    ram_cell[    5145] = 32'h0;  // 32'h4c7da4e8;
    ram_cell[    5146] = 32'h0;  // 32'hae6072d6;
    ram_cell[    5147] = 32'h0;  // 32'ha9258e1e;
    ram_cell[    5148] = 32'h0;  // 32'h3c0b1886;
    ram_cell[    5149] = 32'h0;  // 32'hacb0cadf;
    ram_cell[    5150] = 32'h0;  // 32'h02ea9827;
    ram_cell[    5151] = 32'h0;  // 32'hc914ed1e;
    ram_cell[    5152] = 32'h0;  // 32'h4489a907;
    ram_cell[    5153] = 32'h0;  // 32'h1927d96e;
    ram_cell[    5154] = 32'h0;  // 32'h17e9a6c0;
    ram_cell[    5155] = 32'h0;  // 32'h6caae4dd;
    ram_cell[    5156] = 32'h0;  // 32'h7703fcd8;
    ram_cell[    5157] = 32'h0;  // 32'h74154d07;
    ram_cell[    5158] = 32'h0;  // 32'ha1916cc9;
    ram_cell[    5159] = 32'h0;  // 32'h52e31ec6;
    ram_cell[    5160] = 32'h0;  // 32'h253d5de0;
    ram_cell[    5161] = 32'h0;  // 32'ha964b545;
    ram_cell[    5162] = 32'h0;  // 32'h9cda8640;
    ram_cell[    5163] = 32'h0;  // 32'h60bacfef;
    ram_cell[    5164] = 32'h0;  // 32'h2268a9e7;
    ram_cell[    5165] = 32'h0;  // 32'hdf519300;
    ram_cell[    5166] = 32'h0;  // 32'hc8f5a65e;
    ram_cell[    5167] = 32'h0;  // 32'h2ff66c01;
    ram_cell[    5168] = 32'h0;  // 32'h8d36bebf;
    ram_cell[    5169] = 32'h0;  // 32'hef686f3e;
    ram_cell[    5170] = 32'h0;  // 32'h1d6edcf3;
    ram_cell[    5171] = 32'h0;  // 32'h5f4d5f31;
    ram_cell[    5172] = 32'h0;  // 32'ha9b763c8;
    ram_cell[    5173] = 32'h0;  // 32'h6e54ef82;
    ram_cell[    5174] = 32'h0;  // 32'h6d1768c0;
    ram_cell[    5175] = 32'h0;  // 32'h4d781f13;
    ram_cell[    5176] = 32'h0;  // 32'h359b8383;
    ram_cell[    5177] = 32'h0;  // 32'h7e9d3191;
    ram_cell[    5178] = 32'h0;  // 32'h3720f26e;
    ram_cell[    5179] = 32'h0;  // 32'hef0e52d8;
    ram_cell[    5180] = 32'h0;  // 32'h74c92bc7;
    ram_cell[    5181] = 32'h0;  // 32'hf6e1c35a;
    ram_cell[    5182] = 32'h0;  // 32'h1ff20344;
    ram_cell[    5183] = 32'h0;  // 32'h1eeb6142;
    ram_cell[    5184] = 32'h0;  // 32'h0796751e;
    ram_cell[    5185] = 32'h0;  // 32'hd9cabf40;
    ram_cell[    5186] = 32'h0;  // 32'h3306d9f6;
    ram_cell[    5187] = 32'h0;  // 32'h01a7e82c;
    ram_cell[    5188] = 32'h0;  // 32'h812aff93;
    ram_cell[    5189] = 32'h0;  // 32'h8689b6f7;
    ram_cell[    5190] = 32'h0;  // 32'hd40d14ab;
    ram_cell[    5191] = 32'h0;  // 32'h6d0408c6;
    ram_cell[    5192] = 32'h0;  // 32'hbac356c9;
    ram_cell[    5193] = 32'h0;  // 32'h920fa46b;
    ram_cell[    5194] = 32'h0;  // 32'h67cf9a7d;
    ram_cell[    5195] = 32'h0;  // 32'hd037a7f3;
    ram_cell[    5196] = 32'h0;  // 32'h995fc498;
    ram_cell[    5197] = 32'h0;  // 32'hf9fd6097;
    ram_cell[    5198] = 32'h0;  // 32'hd1f9e05d;
    ram_cell[    5199] = 32'h0;  // 32'h02e3a2d8;
    ram_cell[    5200] = 32'h0;  // 32'hf895a937;
    ram_cell[    5201] = 32'h0;  // 32'h91a87abd;
    ram_cell[    5202] = 32'h0;  // 32'h2ec8fd4c;
    ram_cell[    5203] = 32'h0;  // 32'h62a261b3;
    ram_cell[    5204] = 32'h0;  // 32'h71004510;
    ram_cell[    5205] = 32'h0;  // 32'he0a00e4f;
    ram_cell[    5206] = 32'h0;  // 32'h9d447283;
    ram_cell[    5207] = 32'h0;  // 32'h299e1f8c;
    ram_cell[    5208] = 32'h0;  // 32'h48ce0cd4;
    ram_cell[    5209] = 32'h0;  // 32'h2c8e577d;
    ram_cell[    5210] = 32'h0;  // 32'h340ae875;
    ram_cell[    5211] = 32'h0;  // 32'h6a0276e0;
    ram_cell[    5212] = 32'h0;  // 32'he222df98;
    ram_cell[    5213] = 32'h0;  // 32'h50a04630;
    ram_cell[    5214] = 32'h0;  // 32'h66044b64;
    ram_cell[    5215] = 32'h0;  // 32'h20dcb680;
    ram_cell[    5216] = 32'h0;  // 32'h127ee50f;
    ram_cell[    5217] = 32'h0;  // 32'h00fff11e;
    ram_cell[    5218] = 32'h0;  // 32'h64f20a1c;
    ram_cell[    5219] = 32'h0;  // 32'hc956d4b6;
    ram_cell[    5220] = 32'h0;  // 32'h2b3364e0;
    ram_cell[    5221] = 32'h0;  // 32'h59f447ca;
    ram_cell[    5222] = 32'h0;  // 32'hcfdd77bd;
    ram_cell[    5223] = 32'h0;  // 32'he68c82ea;
    ram_cell[    5224] = 32'h0;  // 32'h8d654f38;
    ram_cell[    5225] = 32'h0;  // 32'hf97c347b;
    ram_cell[    5226] = 32'h0;  // 32'h12efdce5;
    ram_cell[    5227] = 32'h0;  // 32'hcd453cb2;
    ram_cell[    5228] = 32'h0;  // 32'hb41b2d41;
    ram_cell[    5229] = 32'h0;  // 32'h623c25a6;
    ram_cell[    5230] = 32'h0;  // 32'h168387d7;
    ram_cell[    5231] = 32'h0;  // 32'h44567b56;
    ram_cell[    5232] = 32'h0;  // 32'h672fc8fa;
    ram_cell[    5233] = 32'h0;  // 32'hd15573cc;
    ram_cell[    5234] = 32'h0;  // 32'hbda443c3;
    ram_cell[    5235] = 32'h0;  // 32'h46ba8be8;
    ram_cell[    5236] = 32'h0;  // 32'h07a0d5d4;
    ram_cell[    5237] = 32'h0;  // 32'h735513af;
    ram_cell[    5238] = 32'h0;  // 32'hffadc632;
    ram_cell[    5239] = 32'h0;  // 32'ha69ea032;
    ram_cell[    5240] = 32'h0;  // 32'h77cc10b1;
    ram_cell[    5241] = 32'h0;  // 32'h82f98d6b;
    ram_cell[    5242] = 32'h0;  // 32'hb6a88951;
    ram_cell[    5243] = 32'h0;  // 32'h02466269;
    ram_cell[    5244] = 32'h0;  // 32'hb9e589db;
    ram_cell[    5245] = 32'h0;  // 32'hef31de63;
    ram_cell[    5246] = 32'h0;  // 32'he636ff45;
    ram_cell[    5247] = 32'h0;  // 32'h2c856455;
    ram_cell[    5248] = 32'h0;  // 32'hf68170d3;
    ram_cell[    5249] = 32'h0;  // 32'h65001519;
    ram_cell[    5250] = 32'h0;  // 32'h2a3c8411;
    ram_cell[    5251] = 32'h0;  // 32'hd9936aa2;
    ram_cell[    5252] = 32'h0;  // 32'h75f79baa;
    ram_cell[    5253] = 32'h0;  // 32'h60078960;
    ram_cell[    5254] = 32'h0;  // 32'ha7c9f66f;
    ram_cell[    5255] = 32'h0;  // 32'h77973678;
    ram_cell[    5256] = 32'h0;  // 32'hd4c063dc;
    ram_cell[    5257] = 32'h0;  // 32'h374472d0;
    ram_cell[    5258] = 32'h0;  // 32'h4797d15e;
    ram_cell[    5259] = 32'h0;  // 32'h4bbaf9c8;
    ram_cell[    5260] = 32'h0;  // 32'h2c87e2c1;
    ram_cell[    5261] = 32'h0;  // 32'h97d71fd1;
    ram_cell[    5262] = 32'h0;  // 32'h56d2e619;
    ram_cell[    5263] = 32'h0;  // 32'h7c880e8f;
    ram_cell[    5264] = 32'h0;  // 32'h3577acbd;
    ram_cell[    5265] = 32'h0;  // 32'h6e239377;
    ram_cell[    5266] = 32'h0;  // 32'hc5e25736;
    ram_cell[    5267] = 32'h0;  // 32'h163dbf86;
    ram_cell[    5268] = 32'h0;  // 32'hf05968a0;
    ram_cell[    5269] = 32'h0;  // 32'h8a295c92;
    ram_cell[    5270] = 32'h0;  // 32'hed14d493;
    ram_cell[    5271] = 32'h0;  // 32'h53bda9e6;
    ram_cell[    5272] = 32'h0;  // 32'h8c71123f;
    ram_cell[    5273] = 32'h0;  // 32'hbd1e7552;
    ram_cell[    5274] = 32'h0;  // 32'ha3854382;
    ram_cell[    5275] = 32'h0;  // 32'he101a1cc;
    ram_cell[    5276] = 32'h0;  // 32'h8c558400;
    ram_cell[    5277] = 32'h0;  // 32'hb614b9fa;
    ram_cell[    5278] = 32'h0;  // 32'hb3f0db53;
    ram_cell[    5279] = 32'h0;  // 32'h1ab236c5;
    ram_cell[    5280] = 32'h0;  // 32'hb3f89d29;
    ram_cell[    5281] = 32'h0;  // 32'h323e8ef0;
    ram_cell[    5282] = 32'h0;  // 32'hf599d024;
    ram_cell[    5283] = 32'h0;  // 32'h0f03e04e;
    ram_cell[    5284] = 32'h0;  // 32'h57dda51f;
    ram_cell[    5285] = 32'h0;  // 32'h24633850;
    ram_cell[    5286] = 32'h0;  // 32'h90c732ce;
    ram_cell[    5287] = 32'h0;  // 32'h3b3a4a6d;
    ram_cell[    5288] = 32'h0;  // 32'h1f17cb6f;
    ram_cell[    5289] = 32'h0;  // 32'hf72a7aee;
    ram_cell[    5290] = 32'h0;  // 32'h2f800798;
    ram_cell[    5291] = 32'h0;  // 32'ha58c2d21;
    ram_cell[    5292] = 32'h0;  // 32'h7374dcef;
    ram_cell[    5293] = 32'h0;  // 32'h72771089;
    ram_cell[    5294] = 32'h0;  // 32'hab40cf49;
    ram_cell[    5295] = 32'h0;  // 32'h70967e42;
    ram_cell[    5296] = 32'h0;  // 32'h0f0085df;
    ram_cell[    5297] = 32'h0;  // 32'hdd7f71e4;
    ram_cell[    5298] = 32'h0;  // 32'hd8218d8d;
    ram_cell[    5299] = 32'h0;  // 32'h18c63784;
    ram_cell[    5300] = 32'h0;  // 32'h37e1470f;
    ram_cell[    5301] = 32'h0;  // 32'hd1a6f450;
    ram_cell[    5302] = 32'h0;  // 32'h34490079;
    ram_cell[    5303] = 32'h0;  // 32'h3be31c72;
    ram_cell[    5304] = 32'h0;  // 32'he2b6c016;
    ram_cell[    5305] = 32'h0;  // 32'h99f286f2;
    ram_cell[    5306] = 32'h0;  // 32'h2979d587;
    ram_cell[    5307] = 32'h0;  // 32'h250ccba7;
    ram_cell[    5308] = 32'h0;  // 32'he44bf2b1;
    ram_cell[    5309] = 32'h0;  // 32'hc3287813;
    ram_cell[    5310] = 32'h0;  // 32'h1141f6f3;
    ram_cell[    5311] = 32'h0;  // 32'h65d718e0;
    ram_cell[    5312] = 32'h0;  // 32'h533bf5d8;
    ram_cell[    5313] = 32'h0;  // 32'he7dd22c7;
    ram_cell[    5314] = 32'h0;  // 32'hdd95e0af;
    ram_cell[    5315] = 32'h0;  // 32'h2b73d4bc;
    ram_cell[    5316] = 32'h0;  // 32'h0958d639;
    ram_cell[    5317] = 32'h0;  // 32'ha8fbf055;
    ram_cell[    5318] = 32'h0;  // 32'hc6d2ae40;
    ram_cell[    5319] = 32'h0;  // 32'h9a5e074e;
    ram_cell[    5320] = 32'h0;  // 32'h328aeef4;
    ram_cell[    5321] = 32'h0;  // 32'hf1f91d97;
    ram_cell[    5322] = 32'h0;  // 32'hb1d2b845;
    ram_cell[    5323] = 32'h0;  // 32'hf691a88a;
    ram_cell[    5324] = 32'h0;  // 32'h7aef5078;
    ram_cell[    5325] = 32'h0;  // 32'he474a827;
    ram_cell[    5326] = 32'h0;  // 32'hd4844748;
    ram_cell[    5327] = 32'h0;  // 32'h5a698282;
    ram_cell[    5328] = 32'h0;  // 32'hdfd0ea51;
    ram_cell[    5329] = 32'h0;  // 32'hb59d054b;
    ram_cell[    5330] = 32'h0;  // 32'hedc57181;
    ram_cell[    5331] = 32'h0;  // 32'h7eae9756;
    ram_cell[    5332] = 32'h0;  // 32'hddfc6fca;
    ram_cell[    5333] = 32'h0;  // 32'hc903f0a6;
    ram_cell[    5334] = 32'h0;  // 32'hd0ba25e8;
    ram_cell[    5335] = 32'h0;  // 32'h65f9b204;
    ram_cell[    5336] = 32'h0;  // 32'h054695a2;
    ram_cell[    5337] = 32'h0;  // 32'hb01fa164;
    ram_cell[    5338] = 32'h0;  // 32'h8c575299;
    ram_cell[    5339] = 32'h0;  // 32'hb933d5fa;
    ram_cell[    5340] = 32'h0;  // 32'hf19a68f8;
    ram_cell[    5341] = 32'h0;  // 32'hafe582ba;
    ram_cell[    5342] = 32'h0;  // 32'hda529813;
    ram_cell[    5343] = 32'h0;  // 32'h41ff5dea;
    ram_cell[    5344] = 32'h0;  // 32'h3b61deab;
    ram_cell[    5345] = 32'h0;  // 32'h463ed4c1;
    ram_cell[    5346] = 32'h0;  // 32'h7b6e58ff;
    ram_cell[    5347] = 32'h0;  // 32'hc0ffebfd;
    ram_cell[    5348] = 32'h0;  // 32'h130e6597;
    ram_cell[    5349] = 32'h0;  // 32'h1566e9e2;
    ram_cell[    5350] = 32'h0;  // 32'h585c73aa;
    ram_cell[    5351] = 32'h0;  // 32'h4c5c325d;
    ram_cell[    5352] = 32'h0;  // 32'h8b1b3cfd;
    ram_cell[    5353] = 32'h0;  // 32'h07f580fd;
    ram_cell[    5354] = 32'h0;  // 32'h3d207267;
    ram_cell[    5355] = 32'h0;  // 32'h8d9d9525;
    ram_cell[    5356] = 32'h0;  // 32'h3c53166a;
    ram_cell[    5357] = 32'h0;  // 32'hcd03a1fe;
    ram_cell[    5358] = 32'h0;  // 32'hf3e0c08a;
    ram_cell[    5359] = 32'h0;  // 32'ha65119b7;
    ram_cell[    5360] = 32'h0;  // 32'he77b54e5;
    ram_cell[    5361] = 32'h0;  // 32'h9fcac4e6;
    ram_cell[    5362] = 32'h0;  // 32'h217b88dd;
    ram_cell[    5363] = 32'h0;  // 32'h3283a8e1;
    ram_cell[    5364] = 32'h0;  // 32'h3c9cbcba;
    ram_cell[    5365] = 32'h0;  // 32'hf9819993;
    ram_cell[    5366] = 32'h0;  // 32'h660898a3;
    ram_cell[    5367] = 32'h0;  // 32'he70bb219;
    ram_cell[    5368] = 32'h0;  // 32'h3ac0f314;
    ram_cell[    5369] = 32'h0;  // 32'ha2ad4b95;
    ram_cell[    5370] = 32'h0;  // 32'h184c2573;
    ram_cell[    5371] = 32'h0;  // 32'h9f2bad12;
    ram_cell[    5372] = 32'h0;  // 32'h04532a36;
    ram_cell[    5373] = 32'h0;  // 32'h5bcf8b9d;
    ram_cell[    5374] = 32'h0;  // 32'he15e4ddc;
    ram_cell[    5375] = 32'h0;  // 32'h76ab41e2;
    ram_cell[    5376] = 32'h0;  // 32'h45653743;
    ram_cell[    5377] = 32'h0;  // 32'hb8e92fe9;
    ram_cell[    5378] = 32'h0;  // 32'hc7e13e04;
    ram_cell[    5379] = 32'h0;  // 32'he42d1a7a;
    ram_cell[    5380] = 32'h0;  // 32'hb08c11d1;
    ram_cell[    5381] = 32'h0;  // 32'hcdf35dcf;
    ram_cell[    5382] = 32'h0;  // 32'h231c66d1;
    ram_cell[    5383] = 32'h0;  // 32'h77f35de8;
    ram_cell[    5384] = 32'h0;  // 32'hd0363019;
    ram_cell[    5385] = 32'h0;  // 32'h7c086718;
    ram_cell[    5386] = 32'h0;  // 32'hdf448639;
    ram_cell[    5387] = 32'h0;  // 32'he743242b;
    ram_cell[    5388] = 32'h0;  // 32'h95a929f8;
    ram_cell[    5389] = 32'h0;  // 32'h18e51bdb;
    ram_cell[    5390] = 32'h0;  // 32'he42f6b91;
    ram_cell[    5391] = 32'h0;  // 32'h727cdc1a;
    ram_cell[    5392] = 32'h0;  // 32'h9b507fec;
    ram_cell[    5393] = 32'h0;  // 32'h874b83b0;
    ram_cell[    5394] = 32'h0;  // 32'h77ed11b7;
    ram_cell[    5395] = 32'h0;  // 32'hf3386139;
    ram_cell[    5396] = 32'h0;  // 32'hee79b66a;
    ram_cell[    5397] = 32'h0;  // 32'h46766f8e;
    ram_cell[    5398] = 32'h0;  // 32'h05d49ac1;
    ram_cell[    5399] = 32'h0;  // 32'hefe3dfae;
    ram_cell[    5400] = 32'h0;  // 32'h87488e01;
    ram_cell[    5401] = 32'h0;  // 32'h31022a26;
    ram_cell[    5402] = 32'h0;  // 32'ha543d42e;
    ram_cell[    5403] = 32'h0;  // 32'h91f617b9;
    ram_cell[    5404] = 32'h0;  // 32'h09976394;
    ram_cell[    5405] = 32'h0;  // 32'h49c11cd0;
    ram_cell[    5406] = 32'h0;  // 32'hd3184566;
    ram_cell[    5407] = 32'h0;  // 32'h55cde1ea;
    ram_cell[    5408] = 32'h0;  // 32'he4aba583;
    ram_cell[    5409] = 32'h0;  // 32'h1ba10fd2;
    ram_cell[    5410] = 32'h0;  // 32'h9f7ed851;
    ram_cell[    5411] = 32'h0;  // 32'h81f9a1ad;
    ram_cell[    5412] = 32'h0;  // 32'hd3533d58;
    ram_cell[    5413] = 32'h0;  // 32'h5a9a1221;
    ram_cell[    5414] = 32'h0;  // 32'h3c1969fa;
    ram_cell[    5415] = 32'h0;  // 32'h9b51ba5b;
    ram_cell[    5416] = 32'h0;  // 32'h2d0073e5;
    ram_cell[    5417] = 32'h0;  // 32'h5d6a9523;
    ram_cell[    5418] = 32'h0;  // 32'ha8f04baf;
    ram_cell[    5419] = 32'h0;  // 32'h1758ff59;
    ram_cell[    5420] = 32'h0;  // 32'h888e14f6;
    ram_cell[    5421] = 32'h0;  // 32'he0b00973;
    ram_cell[    5422] = 32'h0;  // 32'h50b0365e;
    ram_cell[    5423] = 32'h0;  // 32'h8c34e3c9;
    ram_cell[    5424] = 32'h0;  // 32'hb1f2e994;
    ram_cell[    5425] = 32'h0;  // 32'h5cc4c53a;
    ram_cell[    5426] = 32'h0;  // 32'h2dd6ec40;
    ram_cell[    5427] = 32'h0;  // 32'h0f63938d;
    ram_cell[    5428] = 32'h0;  // 32'hb5407717;
    ram_cell[    5429] = 32'h0;  // 32'h531f9a92;
    ram_cell[    5430] = 32'h0;  // 32'h6196a8c5;
    ram_cell[    5431] = 32'h0;  // 32'h039a800b;
    ram_cell[    5432] = 32'h0;  // 32'h371d20b6;
    ram_cell[    5433] = 32'h0;  // 32'h5e40297a;
    ram_cell[    5434] = 32'h0;  // 32'h85168005;
    ram_cell[    5435] = 32'h0;  // 32'h68c32b21;
    ram_cell[    5436] = 32'h0;  // 32'he5fcdbce;
    ram_cell[    5437] = 32'h0;  // 32'he71c1b4e;
    ram_cell[    5438] = 32'h0;  // 32'h4eaeba63;
    ram_cell[    5439] = 32'h0;  // 32'h45a12708;
    ram_cell[    5440] = 32'h0;  // 32'hd8e0a5bf;
    ram_cell[    5441] = 32'h0;  // 32'h67267d98;
    ram_cell[    5442] = 32'h0;  // 32'hd8d41492;
    ram_cell[    5443] = 32'h0;  // 32'hb8ff4f12;
    ram_cell[    5444] = 32'h0;  // 32'h7f341db4;
    ram_cell[    5445] = 32'h0;  // 32'h7cfc0a58;
    ram_cell[    5446] = 32'h0;  // 32'h5f533a09;
    ram_cell[    5447] = 32'h0;  // 32'h52047dc6;
    ram_cell[    5448] = 32'h0;  // 32'h8160de16;
    ram_cell[    5449] = 32'h0;  // 32'hdd48c645;
    ram_cell[    5450] = 32'h0;  // 32'h116f925f;
    ram_cell[    5451] = 32'h0;  // 32'h7d99944e;
    ram_cell[    5452] = 32'h0;  // 32'h48d1aaab;
    ram_cell[    5453] = 32'h0;  // 32'ha932784c;
    ram_cell[    5454] = 32'h0;  // 32'h41ea8fbc;
    ram_cell[    5455] = 32'h0;  // 32'hd2e18988;
    ram_cell[    5456] = 32'h0;  // 32'h1db70997;
    ram_cell[    5457] = 32'h0;  // 32'hc4dc56a9;
    ram_cell[    5458] = 32'h0;  // 32'hee725a10;
    ram_cell[    5459] = 32'h0;  // 32'hceb374d4;
    ram_cell[    5460] = 32'h0;  // 32'h2171f10e;
    ram_cell[    5461] = 32'h0;  // 32'hd241e3d0;
    ram_cell[    5462] = 32'h0;  // 32'h7bed3e10;
    ram_cell[    5463] = 32'h0;  // 32'h6e23ed0d;
    ram_cell[    5464] = 32'h0;  // 32'h04414ee5;
    ram_cell[    5465] = 32'h0;  // 32'hb9b8082f;
    ram_cell[    5466] = 32'h0;  // 32'h3ed33504;
    ram_cell[    5467] = 32'h0;  // 32'hf7bd3e71;
    ram_cell[    5468] = 32'h0;  // 32'h69e4f193;
    ram_cell[    5469] = 32'h0;  // 32'hc49e76f2;
    ram_cell[    5470] = 32'h0;  // 32'he0ae3cfc;
    ram_cell[    5471] = 32'h0;  // 32'h5435bf0b;
    ram_cell[    5472] = 32'h0;  // 32'had5c5fb7;
    ram_cell[    5473] = 32'h0;  // 32'hcb1a6a0e;
    ram_cell[    5474] = 32'h0;  // 32'h140c9951;
    ram_cell[    5475] = 32'h0;  // 32'h0d6802a5;
    ram_cell[    5476] = 32'h0;  // 32'hda05c611;
    ram_cell[    5477] = 32'h0;  // 32'h4f02b39b;
    ram_cell[    5478] = 32'h0;  // 32'h2c84640b;
    ram_cell[    5479] = 32'h0;  // 32'h18d6c652;
    ram_cell[    5480] = 32'h0;  // 32'hf77d356a;
    ram_cell[    5481] = 32'h0;  // 32'hb9eab86e;
    ram_cell[    5482] = 32'h0;  // 32'h391107e7;
    ram_cell[    5483] = 32'h0;  // 32'ha04c6d96;
    ram_cell[    5484] = 32'h0;  // 32'hb4ca93fb;
    ram_cell[    5485] = 32'h0;  // 32'h2285f08a;
    ram_cell[    5486] = 32'h0;  // 32'h1e4228e2;
    ram_cell[    5487] = 32'h0;  // 32'hab2404e5;
    ram_cell[    5488] = 32'h0;  // 32'h66d9d53b;
    ram_cell[    5489] = 32'h0;  // 32'hfa207451;
    ram_cell[    5490] = 32'h0;  // 32'h51d5a19c;
    ram_cell[    5491] = 32'h0;  // 32'h0d158496;
    ram_cell[    5492] = 32'h0;  // 32'hd8ce63ef;
    ram_cell[    5493] = 32'h0;  // 32'h688642a6;
    ram_cell[    5494] = 32'h0;  // 32'hfb58c14e;
    ram_cell[    5495] = 32'h0;  // 32'h1b4e2bc5;
    ram_cell[    5496] = 32'h0;  // 32'h4cd9ccb4;
    ram_cell[    5497] = 32'h0;  // 32'h29556b2b;
    ram_cell[    5498] = 32'h0;  // 32'h6fecc84b;
    ram_cell[    5499] = 32'h0;  // 32'h4d38e7a8;
    ram_cell[    5500] = 32'h0;  // 32'h857a60d9;
    ram_cell[    5501] = 32'h0;  // 32'h734ee6a9;
    ram_cell[    5502] = 32'h0;  // 32'hec735e02;
    ram_cell[    5503] = 32'h0;  // 32'hf67b3a99;
    ram_cell[    5504] = 32'h0;  // 32'hf1d4aaf9;
    ram_cell[    5505] = 32'h0;  // 32'h36a6b018;
    ram_cell[    5506] = 32'h0;  // 32'h61acd0ab;
    ram_cell[    5507] = 32'h0;  // 32'h5ed5457f;
    ram_cell[    5508] = 32'h0;  // 32'h8ba1c0cc;
    ram_cell[    5509] = 32'h0;  // 32'hae3fb114;
    ram_cell[    5510] = 32'h0;  // 32'h26172a54;
    ram_cell[    5511] = 32'h0;  // 32'h1199e316;
    ram_cell[    5512] = 32'h0;  // 32'hde3b4939;
    ram_cell[    5513] = 32'h0;  // 32'hefc6ba16;
    ram_cell[    5514] = 32'h0;  // 32'h66bbf52f;
    ram_cell[    5515] = 32'h0;  // 32'h8a8d5a99;
    ram_cell[    5516] = 32'h0;  // 32'hce4ab09a;
    ram_cell[    5517] = 32'h0;  // 32'h94a906ef;
    ram_cell[    5518] = 32'h0;  // 32'hd84e1de9;
    ram_cell[    5519] = 32'h0;  // 32'h8ed7794d;
    ram_cell[    5520] = 32'h0;  // 32'h86cde539;
    ram_cell[    5521] = 32'h0;  // 32'h8962ab01;
    ram_cell[    5522] = 32'h0;  // 32'ha30dd297;
    ram_cell[    5523] = 32'h0;  // 32'h80339418;
    ram_cell[    5524] = 32'h0;  // 32'h3aeceb17;
    ram_cell[    5525] = 32'h0;  // 32'h25d6c7ee;
    ram_cell[    5526] = 32'h0;  // 32'hb6beb558;
    ram_cell[    5527] = 32'h0;  // 32'h9ae13790;
    ram_cell[    5528] = 32'h0;  // 32'h65961ecb;
    ram_cell[    5529] = 32'h0;  // 32'h534536ce;
    ram_cell[    5530] = 32'h0;  // 32'h7ec16c24;
    ram_cell[    5531] = 32'h0;  // 32'h02a1abfd;
    ram_cell[    5532] = 32'h0;  // 32'h965d6f03;
    ram_cell[    5533] = 32'h0;  // 32'h761aa0d2;
    ram_cell[    5534] = 32'h0;  // 32'habd881e7;
    ram_cell[    5535] = 32'h0;  // 32'he2d1aba8;
    ram_cell[    5536] = 32'h0;  // 32'h9839af13;
    ram_cell[    5537] = 32'h0;  // 32'hba981b4b;
    ram_cell[    5538] = 32'h0;  // 32'h84e2a19f;
    ram_cell[    5539] = 32'h0;  // 32'h2140cf78;
    ram_cell[    5540] = 32'h0;  // 32'h67f16df6;
    ram_cell[    5541] = 32'h0;  // 32'h3a8d4784;
    ram_cell[    5542] = 32'h0;  // 32'h6b422a92;
    ram_cell[    5543] = 32'h0;  // 32'hf1bb3aa0;
    ram_cell[    5544] = 32'h0;  // 32'h42ff9b34;
    ram_cell[    5545] = 32'h0;  // 32'hb95ab55c;
    ram_cell[    5546] = 32'h0;  // 32'he2830e42;
    ram_cell[    5547] = 32'h0;  // 32'hb89e1967;
    ram_cell[    5548] = 32'h0;  // 32'h4820097c;
    ram_cell[    5549] = 32'h0;  // 32'h816a8ac1;
    ram_cell[    5550] = 32'h0;  // 32'hec758a1b;
    ram_cell[    5551] = 32'h0;  // 32'h60536a3b;
    ram_cell[    5552] = 32'h0;  // 32'h577bfedf;
    ram_cell[    5553] = 32'h0;  // 32'he2b53e8f;
    ram_cell[    5554] = 32'h0;  // 32'h61c7b569;
    ram_cell[    5555] = 32'h0;  // 32'h4e3b622a;
    ram_cell[    5556] = 32'h0;  // 32'hc160293e;
    ram_cell[    5557] = 32'h0;  // 32'hf79844f8;
    ram_cell[    5558] = 32'h0;  // 32'hacf5607c;
    ram_cell[    5559] = 32'h0;  // 32'hf063b893;
    ram_cell[    5560] = 32'h0;  // 32'h1c75df63;
    ram_cell[    5561] = 32'h0;  // 32'hac347001;
    ram_cell[    5562] = 32'h0;  // 32'hd3c4ce3e;
    ram_cell[    5563] = 32'h0;  // 32'hbe378eb1;
    ram_cell[    5564] = 32'h0;  // 32'h677aba41;
    ram_cell[    5565] = 32'h0;  // 32'h2e9c4fb2;
    ram_cell[    5566] = 32'h0;  // 32'hbfa8c368;
    ram_cell[    5567] = 32'h0;  // 32'h111de89a;
    ram_cell[    5568] = 32'h0;  // 32'hfc24d92f;
    ram_cell[    5569] = 32'h0;  // 32'habe27bcf;
    ram_cell[    5570] = 32'h0;  // 32'h3b5d2b00;
    ram_cell[    5571] = 32'h0;  // 32'h8dda684f;
    ram_cell[    5572] = 32'h0;  // 32'h6c10214f;
    ram_cell[    5573] = 32'h0;  // 32'hb16f3452;
    ram_cell[    5574] = 32'h0;  // 32'h434fe6cd;
    ram_cell[    5575] = 32'h0;  // 32'hecc0aa18;
    ram_cell[    5576] = 32'h0;  // 32'h03b65dcf;
    ram_cell[    5577] = 32'h0;  // 32'hd9d24f31;
    ram_cell[    5578] = 32'h0;  // 32'h8b876d00;
    ram_cell[    5579] = 32'h0;  // 32'h59371a58;
    ram_cell[    5580] = 32'h0;  // 32'h25e7ea5d;
    ram_cell[    5581] = 32'h0;  // 32'hf3e0496b;
    ram_cell[    5582] = 32'h0;  // 32'h408070ed;
    ram_cell[    5583] = 32'h0;  // 32'h1d08e501;
    ram_cell[    5584] = 32'h0;  // 32'h503195b9;
    ram_cell[    5585] = 32'h0;  // 32'h2586208b;
    ram_cell[    5586] = 32'h0;  // 32'h0c0e3837;
    ram_cell[    5587] = 32'h0;  // 32'h2dc08c9a;
    ram_cell[    5588] = 32'h0;  // 32'h2955439b;
    ram_cell[    5589] = 32'h0;  // 32'h158692d6;
    ram_cell[    5590] = 32'h0;  // 32'h4f7ae72e;
    ram_cell[    5591] = 32'h0;  // 32'h7d1e2c1b;
    ram_cell[    5592] = 32'h0;  // 32'h1ccbfaae;
    ram_cell[    5593] = 32'h0;  // 32'h4f0ccaf5;
    ram_cell[    5594] = 32'h0;  // 32'h12f89962;
    ram_cell[    5595] = 32'h0;  // 32'h92e28860;
    ram_cell[    5596] = 32'h0;  // 32'h9496ceb5;
    ram_cell[    5597] = 32'h0;  // 32'hcefe8e86;
    ram_cell[    5598] = 32'h0;  // 32'hcdbc9e6d;
    ram_cell[    5599] = 32'h0;  // 32'h9e92e11e;
    ram_cell[    5600] = 32'h0;  // 32'hac664246;
    ram_cell[    5601] = 32'h0;  // 32'h6acc3d17;
    ram_cell[    5602] = 32'h0;  // 32'h3cb90386;
    ram_cell[    5603] = 32'h0;  // 32'h761619c2;
    ram_cell[    5604] = 32'h0;  // 32'h8e51cb5c;
    ram_cell[    5605] = 32'h0;  // 32'he28157a2;
    ram_cell[    5606] = 32'h0;  // 32'h336c8e65;
    ram_cell[    5607] = 32'h0;  // 32'h2d1bca62;
    ram_cell[    5608] = 32'h0;  // 32'h2b02ab4d;
    ram_cell[    5609] = 32'h0;  // 32'h9b6e9a8b;
    ram_cell[    5610] = 32'h0;  // 32'h447e3eaa;
    ram_cell[    5611] = 32'h0;  // 32'hd41a0d4b;
    ram_cell[    5612] = 32'h0;  // 32'h287d9d62;
    ram_cell[    5613] = 32'h0;  // 32'h503a89ee;
    ram_cell[    5614] = 32'h0;  // 32'hbacb9e42;
    ram_cell[    5615] = 32'h0;  // 32'h80b06633;
    ram_cell[    5616] = 32'h0;  // 32'h76db192c;
    ram_cell[    5617] = 32'h0;  // 32'hdaf387a0;
    ram_cell[    5618] = 32'h0;  // 32'hc1a0995a;
    ram_cell[    5619] = 32'h0;  // 32'ha0212718;
    ram_cell[    5620] = 32'h0;  // 32'hb9d1035f;
    ram_cell[    5621] = 32'h0;  // 32'h8121b048;
    ram_cell[    5622] = 32'h0;  // 32'hc0365755;
    ram_cell[    5623] = 32'h0;  // 32'hfc7e0aa9;
    ram_cell[    5624] = 32'h0;  // 32'h0de02e66;
    ram_cell[    5625] = 32'h0;  // 32'h69eaed51;
    ram_cell[    5626] = 32'h0;  // 32'h430b363c;
    ram_cell[    5627] = 32'h0;  // 32'hd5db2d17;
    ram_cell[    5628] = 32'h0;  // 32'h617c51fd;
    ram_cell[    5629] = 32'h0;  // 32'hd7d3e14c;
    ram_cell[    5630] = 32'h0;  // 32'h38d34355;
    ram_cell[    5631] = 32'h0;  // 32'hd44cbf4a;
    ram_cell[    5632] = 32'h0;  // 32'h0e91b5d3;
    ram_cell[    5633] = 32'h0;  // 32'h67192b15;
    ram_cell[    5634] = 32'h0;  // 32'hcd908181;
    ram_cell[    5635] = 32'h0;  // 32'h5b026690;
    ram_cell[    5636] = 32'h0;  // 32'h65d2f8f1;
    ram_cell[    5637] = 32'h0;  // 32'haff644b4;
    ram_cell[    5638] = 32'h0;  // 32'h3661f2a6;
    ram_cell[    5639] = 32'h0;  // 32'h3a4af1f6;
    ram_cell[    5640] = 32'h0;  // 32'h5ae5525b;
    ram_cell[    5641] = 32'h0;  // 32'he6447e25;
    ram_cell[    5642] = 32'h0;  // 32'h2c07b0fb;
    ram_cell[    5643] = 32'h0;  // 32'hce3317a7;
    ram_cell[    5644] = 32'h0;  // 32'h4fae67ca;
    ram_cell[    5645] = 32'h0;  // 32'h5dee5ea2;
    ram_cell[    5646] = 32'h0;  // 32'h74f067a2;
    ram_cell[    5647] = 32'h0;  // 32'hf1e7c447;
    ram_cell[    5648] = 32'h0;  // 32'hf6f5da98;
    ram_cell[    5649] = 32'h0;  // 32'h0f428893;
    ram_cell[    5650] = 32'h0;  // 32'ha5c14487;
    ram_cell[    5651] = 32'h0;  // 32'h5116f832;
    ram_cell[    5652] = 32'h0;  // 32'h3d3244c7;
    ram_cell[    5653] = 32'h0;  // 32'he0c1a25c;
    ram_cell[    5654] = 32'h0;  // 32'h56752ee8;
    ram_cell[    5655] = 32'h0;  // 32'h0a311ece;
    ram_cell[    5656] = 32'h0;  // 32'he81ee29a;
    ram_cell[    5657] = 32'h0;  // 32'h89f1a00d;
    ram_cell[    5658] = 32'h0;  // 32'hdaaab0aa;
    ram_cell[    5659] = 32'h0;  // 32'h262b7e03;
    ram_cell[    5660] = 32'h0;  // 32'had744f5e;
    ram_cell[    5661] = 32'h0;  // 32'h0248db1f;
    ram_cell[    5662] = 32'h0;  // 32'hf4d7001e;
    ram_cell[    5663] = 32'h0;  // 32'h16ef5939;
    ram_cell[    5664] = 32'h0;  // 32'h9bb566f5;
    ram_cell[    5665] = 32'h0;  // 32'h2d175941;
    ram_cell[    5666] = 32'h0;  // 32'he96d695a;
    ram_cell[    5667] = 32'h0;  // 32'hdee064ac;
    ram_cell[    5668] = 32'h0;  // 32'hdc56a417;
    ram_cell[    5669] = 32'h0;  // 32'h3fef3be0;
    ram_cell[    5670] = 32'h0;  // 32'h3b9ae65e;
    ram_cell[    5671] = 32'h0;  // 32'h95d5f1d2;
    ram_cell[    5672] = 32'h0;  // 32'h68c3f1ac;
    ram_cell[    5673] = 32'h0;  // 32'h7f21b8a0;
    ram_cell[    5674] = 32'h0;  // 32'hdee819c1;
    ram_cell[    5675] = 32'h0;  // 32'h199b70c0;
    ram_cell[    5676] = 32'h0;  // 32'h0296e07f;
    ram_cell[    5677] = 32'h0;  // 32'hf808d1f7;
    ram_cell[    5678] = 32'h0;  // 32'ha45f110b;
    ram_cell[    5679] = 32'h0;  // 32'had415ffe;
    ram_cell[    5680] = 32'h0;  // 32'hd9db5afe;
    ram_cell[    5681] = 32'h0;  // 32'h80187cc7;
    ram_cell[    5682] = 32'h0;  // 32'he8c5fc2b;
    ram_cell[    5683] = 32'h0;  // 32'h9e8a98ee;
    ram_cell[    5684] = 32'h0;  // 32'h5feecaca;
    ram_cell[    5685] = 32'h0;  // 32'h202ad4d7;
    ram_cell[    5686] = 32'h0;  // 32'hd2fe45fe;
    ram_cell[    5687] = 32'h0;  // 32'h4d2c1dca;
    ram_cell[    5688] = 32'h0;  // 32'hd84102fd;
    ram_cell[    5689] = 32'h0;  // 32'h766388ab;
    ram_cell[    5690] = 32'h0;  // 32'h0786afda;
    ram_cell[    5691] = 32'h0;  // 32'h8bb5cd19;
    ram_cell[    5692] = 32'h0;  // 32'hcb1c7404;
    ram_cell[    5693] = 32'h0;  // 32'h254716b7;
    ram_cell[    5694] = 32'h0;  // 32'hfec152db;
    ram_cell[    5695] = 32'h0;  // 32'h40142241;
    ram_cell[    5696] = 32'h0;  // 32'h8da2461f;
    ram_cell[    5697] = 32'h0;  // 32'h92503292;
    ram_cell[    5698] = 32'h0;  // 32'h460597fc;
    ram_cell[    5699] = 32'h0;  // 32'he6f1f76b;
    ram_cell[    5700] = 32'h0;  // 32'h94a4f720;
    ram_cell[    5701] = 32'h0;  // 32'h89a57482;
    ram_cell[    5702] = 32'h0;  // 32'hf68ec1c2;
    ram_cell[    5703] = 32'h0;  // 32'h2145147c;
    ram_cell[    5704] = 32'h0;  // 32'h28baa77f;
    ram_cell[    5705] = 32'h0;  // 32'h203dd16c;
    ram_cell[    5706] = 32'h0;  // 32'hc5915eb5;
    ram_cell[    5707] = 32'h0;  // 32'h1dd6d338;
    ram_cell[    5708] = 32'h0;  // 32'h4acea30f;
    ram_cell[    5709] = 32'h0;  // 32'h80bc06a8;
    ram_cell[    5710] = 32'h0;  // 32'h18c15bbe;
    ram_cell[    5711] = 32'h0;  // 32'h51623c01;
    ram_cell[    5712] = 32'h0;  // 32'h87755f54;
    ram_cell[    5713] = 32'h0;  // 32'h1982389f;
    ram_cell[    5714] = 32'h0;  // 32'h740191ec;
    ram_cell[    5715] = 32'h0;  // 32'h83787cc5;
    ram_cell[    5716] = 32'h0;  // 32'hf5c5b29d;
    ram_cell[    5717] = 32'h0;  // 32'h027a1eea;
    ram_cell[    5718] = 32'h0;  // 32'h807a55d2;
    ram_cell[    5719] = 32'h0;  // 32'hb569aa1b;
    ram_cell[    5720] = 32'h0;  // 32'h15ad729f;
    ram_cell[    5721] = 32'h0;  // 32'h9761dc29;
    ram_cell[    5722] = 32'h0;  // 32'hf0a704ee;
    ram_cell[    5723] = 32'h0;  // 32'hb7cb8c8a;
    ram_cell[    5724] = 32'h0;  // 32'h3320598b;
    ram_cell[    5725] = 32'h0;  // 32'h62bcb7a2;
    ram_cell[    5726] = 32'h0;  // 32'h11b5390e;
    ram_cell[    5727] = 32'h0;  // 32'he23fdd35;
    ram_cell[    5728] = 32'h0;  // 32'hb91ae29a;
    ram_cell[    5729] = 32'h0;  // 32'h96e27804;
    ram_cell[    5730] = 32'h0;  // 32'hffb0daf0;
    ram_cell[    5731] = 32'h0;  // 32'hbf4d58e1;
    ram_cell[    5732] = 32'h0;  // 32'h2a92f9b3;
    ram_cell[    5733] = 32'h0;  // 32'h2f9748be;
    ram_cell[    5734] = 32'h0;  // 32'hc46c138a;
    ram_cell[    5735] = 32'h0;  // 32'h6169a4cd;
    ram_cell[    5736] = 32'h0;  // 32'h3ffd46de;
    ram_cell[    5737] = 32'h0;  // 32'h0b621f7b;
    ram_cell[    5738] = 32'h0;  // 32'hb5b2c2d6;
    ram_cell[    5739] = 32'h0;  // 32'hb52cf045;
    ram_cell[    5740] = 32'h0;  // 32'h8430e3c3;
    ram_cell[    5741] = 32'h0;  // 32'h4fc0073c;
    ram_cell[    5742] = 32'h0;  // 32'h398f17c1;
    ram_cell[    5743] = 32'h0;  // 32'ha58b9d15;
    ram_cell[    5744] = 32'h0;  // 32'h8beb8dfe;
    ram_cell[    5745] = 32'h0;  // 32'hcbc83fdc;
    ram_cell[    5746] = 32'h0;  // 32'hb9357584;
    ram_cell[    5747] = 32'h0;  // 32'hac788541;
    ram_cell[    5748] = 32'h0;  // 32'hfb93a7e6;
    ram_cell[    5749] = 32'h0;  // 32'hb6732212;
    ram_cell[    5750] = 32'h0;  // 32'h3cc7256f;
    ram_cell[    5751] = 32'h0;  // 32'h8d81ff6d;
    ram_cell[    5752] = 32'h0;  // 32'h738aa406;
    ram_cell[    5753] = 32'h0;  // 32'h8cf9b5e1;
    ram_cell[    5754] = 32'h0;  // 32'hbd682dfd;
    ram_cell[    5755] = 32'h0;  // 32'hc4143d36;
    ram_cell[    5756] = 32'h0;  // 32'h0abf0728;
    ram_cell[    5757] = 32'h0;  // 32'headf9ee8;
    ram_cell[    5758] = 32'h0;  // 32'hefb619e0;
    ram_cell[    5759] = 32'h0;  // 32'h024589a0;
    ram_cell[    5760] = 32'h0;  // 32'h8fdd7746;
    ram_cell[    5761] = 32'h0;  // 32'hd582e182;
    ram_cell[    5762] = 32'h0;  // 32'haf295bfd;
    ram_cell[    5763] = 32'h0;  // 32'h59c409b9;
    ram_cell[    5764] = 32'h0;  // 32'h44644057;
    ram_cell[    5765] = 32'h0;  // 32'hfcaa5b85;
    ram_cell[    5766] = 32'h0;  // 32'h87237662;
    ram_cell[    5767] = 32'h0;  // 32'h6feaf075;
    ram_cell[    5768] = 32'h0;  // 32'h889d8496;
    ram_cell[    5769] = 32'h0;  // 32'hd3d512e0;
    ram_cell[    5770] = 32'h0;  // 32'h53599ce9;
    ram_cell[    5771] = 32'h0;  // 32'hd016d0c6;
    ram_cell[    5772] = 32'h0;  // 32'ha264dff2;
    ram_cell[    5773] = 32'h0;  // 32'hb9d2947e;
    ram_cell[    5774] = 32'h0;  // 32'h41eae4dc;
    ram_cell[    5775] = 32'h0;  // 32'ha15ac4af;
    ram_cell[    5776] = 32'h0;  // 32'hef9bbc95;
    ram_cell[    5777] = 32'h0;  // 32'hc9040077;
    ram_cell[    5778] = 32'h0;  // 32'haa078d50;
    ram_cell[    5779] = 32'h0;  // 32'h355111f6;
    ram_cell[    5780] = 32'h0;  // 32'h12f117c5;
    ram_cell[    5781] = 32'h0;  // 32'h9e3a4075;
    ram_cell[    5782] = 32'h0;  // 32'hda962cca;
    ram_cell[    5783] = 32'h0;  // 32'h5c88a005;
    ram_cell[    5784] = 32'h0;  // 32'h9783bc5a;
    ram_cell[    5785] = 32'h0;  // 32'h4756a99c;
    ram_cell[    5786] = 32'h0;  // 32'h4c8f0b91;
    ram_cell[    5787] = 32'h0;  // 32'hedfec226;
    ram_cell[    5788] = 32'h0;  // 32'hc60c0b22;
    ram_cell[    5789] = 32'h0;  // 32'h68c7b87b;
    ram_cell[    5790] = 32'h0;  // 32'hf082d7f3;
    ram_cell[    5791] = 32'h0;  // 32'h1b52e1f4;
    ram_cell[    5792] = 32'h0;  // 32'he22027f2;
    ram_cell[    5793] = 32'h0;  // 32'h7ef5610a;
    ram_cell[    5794] = 32'h0;  // 32'ha98f9d77;
    ram_cell[    5795] = 32'h0;  // 32'h2fff1141;
    ram_cell[    5796] = 32'h0;  // 32'h1c8714aa;
    ram_cell[    5797] = 32'h0;  // 32'h8b6d5226;
    ram_cell[    5798] = 32'h0;  // 32'h2f09921e;
    ram_cell[    5799] = 32'h0;  // 32'h1deaa33b;
    ram_cell[    5800] = 32'h0;  // 32'hb0017173;
    ram_cell[    5801] = 32'h0;  // 32'hd9c39630;
    ram_cell[    5802] = 32'h0;  // 32'h3f088c81;
    ram_cell[    5803] = 32'h0;  // 32'h3e92ddd4;
    ram_cell[    5804] = 32'h0;  // 32'h90abc9eb;
    ram_cell[    5805] = 32'h0;  // 32'hd412b6e1;
    ram_cell[    5806] = 32'h0;  // 32'h09c6e0d4;
    ram_cell[    5807] = 32'h0;  // 32'h5b2673e0;
    ram_cell[    5808] = 32'h0;  // 32'hb68808af;
    ram_cell[    5809] = 32'h0;  // 32'h2b5e57ff;
    ram_cell[    5810] = 32'h0;  // 32'hf22c89ad;
    ram_cell[    5811] = 32'h0;  // 32'hf2f5b894;
    ram_cell[    5812] = 32'h0;  // 32'h45a5d398;
    ram_cell[    5813] = 32'h0;  // 32'h3d3e5075;
    ram_cell[    5814] = 32'h0;  // 32'hd329b74e;
    ram_cell[    5815] = 32'h0;  // 32'h432b0a6c;
    ram_cell[    5816] = 32'h0;  // 32'h103445ac;
    ram_cell[    5817] = 32'h0;  // 32'hdb04471b;
    ram_cell[    5818] = 32'h0;  // 32'h81176ae5;
    ram_cell[    5819] = 32'h0;  // 32'h5a16e8eb;
    ram_cell[    5820] = 32'h0;  // 32'hc1f20253;
    ram_cell[    5821] = 32'h0;  // 32'hd2577efe;
    ram_cell[    5822] = 32'h0;  // 32'hf4a9c911;
    ram_cell[    5823] = 32'h0;  // 32'hd3f82b7f;
    ram_cell[    5824] = 32'h0;  // 32'h1329df11;
    ram_cell[    5825] = 32'h0;  // 32'h67ffe12c;
    ram_cell[    5826] = 32'h0;  // 32'h973de0b5;
    ram_cell[    5827] = 32'h0;  // 32'h86cf977f;
    ram_cell[    5828] = 32'h0;  // 32'hbc309112;
    ram_cell[    5829] = 32'h0;  // 32'h292fe715;
    ram_cell[    5830] = 32'h0;  // 32'h364fa329;
    ram_cell[    5831] = 32'h0;  // 32'h52452256;
    ram_cell[    5832] = 32'h0;  // 32'h99c0853c;
    ram_cell[    5833] = 32'h0;  // 32'h52275c68;
    ram_cell[    5834] = 32'h0;  // 32'h962d9e6b;
    ram_cell[    5835] = 32'h0;  // 32'h88d117c3;
    ram_cell[    5836] = 32'h0;  // 32'h77d81a4c;
    ram_cell[    5837] = 32'h0;  // 32'h5d9801ed;
    ram_cell[    5838] = 32'h0;  // 32'h6f30689b;
    ram_cell[    5839] = 32'h0;  // 32'ha8e6679b;
    ram_cell[    5840] = 32'h0;  // 32'h5bb98631;
    ram_cell[    5841] = 32'h0;  // 32'h05923c45;
    ram_cell[    5842] = 32'h0;  // 32'he9fb1236;
    ram_cell[    5843] = 32'h0;  // 32'h6a7224b3;
    ram_cell[    5844] = 32'h0;  // 32'hb461a6d8;
    ram_cell[    5845] = 32'h0;  // 32'hafef69a8;
    ram_cell[    5846] = 32'h0;  // 32'hc3813466;
    ram_cell[    5847] = 32'h0;  // 32'h16bbcfaf;
    ram_cell[    5848] = 32'h0;  // 32'h41431de7;
    ram_cell[    5849] = 32'h0;  // 32'had9f1628;
    ram_cell[    5850] = 32'h0;  // 32'h90b1463b;
    ram_cell[    5851] = 32'h0;  // 32'h2e83d790;
    ram_cell[    5852] = 32'h0;  // 32'ha657eb46;
    ram_cell[    5853] = 32'h0;  // 32'he95620e8;
    ram_cell[    5854] = 32'h0;  // 32'h4e6d1484;
    ram_cell[    5855] = 32'h0;  // 32'h330a349f;
    ram_cell[    5856] = 32'h0;  // 32'h30a1555e;
    ram_cell[    5857] = 32'h0;  // 32'ha7f126e0;
    ram_cell[    5858] = 32'h0;  // 32'hada2d60b;
    ram_cell[    5859] = 32'h0;  // 32'h2bf61e82;
    ram_cell[    5860] = 32'h0;  // 32'he7aa22ea;
    ram_cell[    5861] = 32'h0;  // 32'h3a2dd7b7;
    ram_cell[    5862] = 32'h0;  // 32'h1b1094cb;
    ram_cell[    5863] = 32'h0;  // 32'hb7c43572;
    ram_cell[    5864] = 32'h0;  // 32'hf3326aa8;
    ram_cell[    5865] = 32'h0;  // 32'h36b85655;
    ram_cell[    5866] = 32'h0;  // 32'h982ddace;
    ram_cell[    5867] = 32'h0;  // 32'h97b466fa;
    ram_cell[    5868] = 32'h0;  // 32'h05af294e;
    ram_cell[    5869] = 32'h0;  // 32'hd1ebc99f;
    ram_cell[    5870] = 32'h0;  // 32'hb6855abd;
    ram_cell[    5871] = 32'h0;  // 32'h25445e47;
    ram_cell[    5872] = 32'h0;  // 32'h10647686;
    ram_cell[    5873] = 32'h0;  // 32'hae596162;
    ram_cell[    5874] = 32'h0;  // 32'h647a0f19;
    ram_cell[    5875] = 32'h0;  // 32'hfe055cab;
    ram_cell[    5876] = 32'h0;  // 32'hb1548358;
    ram_cell[    5877] = 32'h0;  // 32'h2cbd018c;
    ram_cell[    5878] = 32'h0;  // 32'hfe59f356;
    ram_cell[    5879] = 32'h0;  // 32'h94f83303;
    ram_cell[    5880] = 32'h0;  // 32'h875a0812;
    ram_cell[    5881] = 32'h0;  // 32'hd7414b53;
    ram_cell[    5882] = 32'h0;  // 32'h0dee92e6;
    ram_cell[    5883] = 32'h0;  // 32'h4ce823a9;
    ram_cell[    5884] = 32'h0;  // 32'h8c611f08;
    ram_cell[    5885] = 32'h0;  // 32'h5d4a241a;
    ram_cell[    5886] = 32'h0;  // 32'h349a9cc8;
    ram_cell[    5887] = 32'h0;  // 32'h3b6dcca5;
    ram_cell[    5888] = 32'h0;  // 32'h78ec9f42;
    ram_cell[    5889] = 32'h0;  // 32'hd65decbe;
    ram_cell[    5890] = 32'h0;  // 32'hf7a7ab9e;
    ram_cell[    5891] = 32'h0;  // 32'hec08cf2b;
    ram_cell[    5892] = 32'h0;  // 32'hc8e09750;
    ram_cell[    5893] = 32'h0;  // 32'hdee4f26f;
    ram_cell[    5894] = 32'h0;  // 32'h7125d080;
    ram_cell[    5895] = 32'h0;  // 32'h1600c89a;
    ram_cell[    5896] = 32'h0;  // 32'hc33f6c48;
    ram_cell[    5897] = 32'h0;  // 32'hc570f5b0;
    ram_cell[    5898] = 32'h0;  // 32'hb7974239;
    ram_cell[    5899] = 32'h0;  // 32'hcf6adee2;
    ram_cell[    5900] = 32'h0;  // 32'h42e02df6;
    ram_cell[    5901] = 32'h0;  // 32'hb64c9778;
    ram_cell[    5902] = 32'h0;  // 32'he6438a07;
    ram_cell[    5903] = 32'h0;  // 32'hbe7895b5;
    ram_cell[    5904] = 32'h0;  // 32'heb5079e8;
    ram_cell[    5905] = 32'h0;  // 32'he0caf791;
    ram_cell[    5906] = 32'h0;  // 32'h533d51ea;
    ram_cell[    5907] = 32'h0;  // 32'hae7051d3;
    ram_cell[    5908] = 32'h0;  // 32'habd37b28;
    ram_cell[    5909] = 32'h0;  // 32'he1b369a4;
    ram_cell[    5910] = 32'h0;  // 32'hbc724086;
    ram_cell[    5911] = 32'h0;  // 32'h4b4b9083;
    ram_cell[    5912] = 32'h0;  // 32'h65046a1d;
    ram_cell[    5913] = 32'h0;  // 32'hbc1d4c5a;
    ram_cell[    5914] = 32'h0;  // 32'h2aae24e2;
    ram_cell[    5915] = 32'h0;  // 32'h75797d6c;
    ram_cell[    5916] = 32'h0;  // 32'h27576f1b;
    ram_cell[    5917] = 32'h0;  // 32'h12a8c489;
    ram_cell[    5918] = 32'h0;  // 32'h92687125;
    ram_cell[    5919] = 32'h0;  // 32'hbe66700e;
    ram_cell[    5920] = 32'h0;  // 32'h7beae183;
    ram_cell[    5921] = 32'h0;  // 32'h90e8de3a;
    ram_cell[    5922] = 32'h0;  // 32'ha3c2a30c;
    ram_cell[    5923] = 32'h0;  // 32'h3e0f2fdd;
    ram_cell[    5924] = 32'h0;  // 32'h5528f13e;
    ram_cell[    5925] = 32'h0;  // 32'h6f831080;
    ram_cell[    5926] = 32'h0;  // 32'h6f4c2733;
    ram_cell[    5927] = 32'h0;  // 32'h2d82706b;
    ram_cell[    5928] = 32'h0;  // 32'h91a513c6;
    ram_cell[    5929] = 32'h0;  // 32'hf257573a;
    ram_cell[    5930] = 32'h0;  // 32'h8413583a;
    ram_cell[    5931] = 32'h0;  // 32'h248691b1;
    ram_cell[    5932] = 32'h0;  // 32'hf98dff1a;
    ram_cell[    5933] = 32'h0;  // 32'hd2990af5;
    ram_cell[    5934] = 32'h0;  // 32'h9e6bd409;
    ram_cell[    5935] = 32'h0;  // 32'h339f79c9;
    ram_cell[    5936] = 32'h0;  // 32'hcdd368dd;
    ram_cell[    5937] = 32'h0;  // 32'h1418035f;
    ram_cell[    5938] = 32'h0;  // 32'he8e67c00;
    ram_cell[    5939] = 32'h0;  // 32'h9ca241bf;
    ram_cell[    5940] = 32'h0;  // 32'h15eedb07;
    ram_cell[    5941] = 32'h0;  // 32'h5a12c123;
    ram_cell[    5942] = 32'h0;  // 32'h16e57e21;
    ram_cell[    5943] = 32'h0;  // 32'h17f536a0;
    ram_cell[    5944] = 32'h0;  // 32'hf61d612d;
    ram_cell[    5945] = 32'h0;  // 32'h041f33c1;
    ram_cell[    5946] = 32'h0;  // 32'hb46720fd;
    ram_cell[    5947] = 32'h0;  // 32'h0964b728;
    ram_cell[    5948] = 32'h0;  // 32'ha05bc1a3;
    ram_cell[    5949] = 32'h0;  // 32'hd2770e85;
    ram_cell[    5950] = 32'h0;  // 32'h9599a76f;
    ram_cell[    5951] = 32'h0;  // 32'hec346c0b;
    ram_cell[    5952] = 32'h0;  // 32'hc7695136;
    ram_cell[    5953] = 32'h0;  // 32'h1b6ec9ec;
    ram_cell[    5954] = 32'h0;  // 32'h8de36b30;
    ram_cell[    5955] = 32'h0;  // 32'h3688b35e;
    ram_cell[    5956] = 32'h0;  // 32'h140d0e76;
    ram_cell[    5957] = 32'h0;  // 32'h82356eb9;
    ram_cell[    5958] = 32'h0;  // 32'h655838f8;
    ram_cell[    5959] = 32'h0;  // 32'hb7fa6718;
    ram_cell[    5960] = 32'h0;  // 32'h8d153a43;
    ram_cell[    5961] = 32'h0;  // 32'h8b27015e;
    ram_cell[    5962] = 32'h0;  // 32'h34169a84;
    ram_cell[    5963] = 32'h0;  // 32'he9d7ee6e;
    ram_cell[    5964] = 32'h0;  // 32'h0c56cbce;
    ram_cell[    5965] = 32'h0;  // 32'h6e272fe0;
    ram_cell[    5966] = 32'h0;  // 32'h88cf653e;
    ram_cell[    5967] = 32'h0;  // 32'h1d732ce8;
    ram_cell[    5968] = 32'h0;  // 32'h225c0887;
    ram_cell[    5969] = 32'h0;  // 32'hc04c5e5b;
    ram_cell[    5970] = 32'h0;  // 32'h8291fae6;
    ram_cell[    5971] = 32'h0;  // 32'ha8c35c6c;
    ram_cell[    5972] = 32'h0;  // 32'hf5523e24;
    ram_cell[    5973] = 32'h0;  // 32'h74cdcd6c;
    ram_cell[    5974] = 32'h0;  // 32'h870607a5;
    ram_cell[    5975] = 32'h0;  // 32'h04e25367;
    ram_cell[    5976] = 32'h0;  // 32'h9e01431d;
    ram_cell[    5977] = 32'h0;  // 32'h165886f0;
    ram_cell[    5978] = 32'h0;  // 32'h981e74d3;
    ram_cell[    5979] = 32'h0;  // 32'hc1c5aa35;
    ram_cell[    5980] = 32'h0;  // 32'ha0532978;
    ram_cell[    5981] = 32'h0;  // 32'ha5122163;
    ram_cell[    5982] = 32'h0;  // 32'h33104f89;
    ram_cell[    5983] = 32'h0;  // 32'h93009b43;
    ram_cell[    5984] = 32'h0;  // 32'h4814a607;
    ram_cell[    5985] = 32'h0;  // 32'hc8b44390;
    ram_cell[    5986] = 32'h0;  // 32'h0fbc37a7;
    ram_cell[    5987] = 32'h0;  // 32'h124bfe33;
    ram_cell[    5988] = 32'h0;  // 32'h4815e1d5;
    ram_cell[    5989] = 32'h0;  // 32'h5cc384a8;
    ram_cell[    5990] = 32'h0;  // 32'h3b1f2b63;
    ram_cell[    5991] = 32'h0;  // 32'hbba62010;
    ram_cell[    5992] = 32'h0;  // 32'hd127cfb5;
    ram_cell[    5993] = 32'h0;  // 32'he3910a5d;
    ram_cell[    5994] = 32'h0;  // 32'he75920f0;
    ram_cell[    5995] = 32'h0;  // 32'heda23f2f;
    ram_cell[    5996] = 32'h0;  // 32'hb4df063d;
    ram_cell[    5997] = 32'h0;  // 32'hc10fbb81;
    ram_cell[    5998] = 32'h0;  // 32'h4372e1de;
    ram_cell[    5999] = 32'h0;  // 32'h4d819767;
    ram_cell[    6000] = 32'h0;  // 32'h47a038cf;
    ram_cell[    6001] = 32'h0;  // 32'h5f8c18d3;
    ram_cell[    6002] = 32'h0;  // 32'h5e498b75;
    ram_cell[    6003] = 32'h0;  // 32'ha5e8b2c5;
    ram_cell[    6004] = 32'h0;  // 32'h78609991;
    ram_cell[    6005] = 32'h0;  // 32'h6d2747c2;
    ram_cell[    6006] = 32'h0;  // 32'he9d3f767;
    ram_cell[    6007] = 32'h0;  // 32'h25450c93;
    ram_cell[    6008] = 32'h0;  // 32'h4e6eb3ed;
    ram_cell[    6009] = 32'h0;  // 32'h0954f808;
    ram_cell[    6010] = 32'h0;  // 32'h275bc88e;
    ram_cell[    6011] = 32'h0;  // 32'h34cded84;
    ram_cell[    6012] = 32'h0;  // 32'hb96b70a2;
    ram_cell[    6013] = 32'h0;  // 32'h57abd35f;
    ram_cell[    6014] = 32'h0;  // 32'h75a81af4;
    ram_cell[    6015] = 32'h0;  // 32'hbf0865a9;
    ram_cell[    6016] = 32'h0;  // 32'h8b2ea363;
    ram_cell[    6017] = 32'h0;  // 32'h7117147c;
    ram_cell[    6018] = 32'h0;  // 32'h0e6ce9c3;
    ram_cell[    6019] = 32'h0;  // 32'hec4d7a23;
    ram_cell[    6020] = 32'h0;  // 32'hde53f8a1;
    ram_cell[    6021] = 32'h0;  // 32'hfe7acf3c;
    ram_cell[    6022] = 32'h0;  // 32'h47413551;
    ram_cell[    6023] = 32'h0;  // 32'h7c16588f;
    ram_cell[    6024] = 32'h0;  // 32'h8f828f9a;
    ram_cell[    6025] = 32'h0;  // 32'h513ec2fa;
    ram_cell[    6026] = 32'h0;  // 32'h16c36534;
    ram_cell[    6027] = 32'h0;  // 32'h2669d7c6;
    ram_cell[    6028] = 32'h0;  // 32'h051d2a76;
    ram_cell[    6029] = 32'h0;  // 32'h80a93771;
    ram_cell[    6030] = 32'h0;  // 32'hb1fa8f03;
    ram_cell[    6031] = 32'h0;  // 32'hfc7530fe;
    ram_cell[    6032] = 32'h0;  // 32'h12cc5d60;
    ram_cell[    6033] = 32'h0;  // 32'h1ef991ff;
    ram_cell[    6034] = 32'h0;  // 32'h517aee7b;
    ram_cell[    6035] = 32'h0;  // 32'h0430f146;
    ram_cell[    6036] = 32'h0;  // 32'hbf845530;
    ram_cell[    6037] = 32'h0;  // 32'he0ba48ce;
    ram_cell[    6038] = 32'h0;  // 32'h84bfdf9c;
    ram_cell[    6039] = 32'h0;  // 32'h15e356b4;
    ram_cell[    6040] = 32'h0;  // 32'h5859c70a;
    ram_cell[    6041] = 32'h0;  // 32'hbbec5696;
    ram_cell[    6042] = 32'h0;  // 32'hef47446c;
    ram_cell[    6043] = 32'h0;  // 32'haeb10921;
    ram_cell[    6044] = 32'h0;  // 32'h8c2b7cbf;
    ram_cell[    6045] = 32'h0;  // 32'hf521d443;
    ram_cell[    6046] = 32'h0;  // 32'h6df38014;
    ram_cell[    6047] = 32'h0;  // 32'heee30f93;
    ram_cell[    6048] = 32'h0;  // 32'h308363f8;
    ram_cell[    6049] = 32'h0;  // 32'ha81a91c6;
    ram_cell[    6050] = 32'h0;  // 32'h72823bb7;
    ram_cell[    6051] = 32'h0;  // 32'h2541bf59;
    ram_cell[    6052] = 32'h0;  // 32'hfcb30e5f;
    ram_cell[    6053] = 32'h0;  // 32'h070d8b58;
    ram_cell[    6054] = 32'h0;  // 32'h1f31a58a;
    ram_cell[    6055] = 32'h0;  // 32'h4665201d;
    ram_cell[    6056] = 32'h0;  // 32'he324f193;
    ram_cell[    6057] = 32'h0;  // 32'hf5b090d6;
    ram_cell[    6058] = 32'h0;  // 32'hc2c72145;
    ram_cell[    6059] = 32'h0;  // 32'hc50ebf69;
    ram_cell[    6060] = 32'h0;  // 32'h6538f73d;
    ram_cell[    6061] = 32'h0;  // 32'hb0b55218;
    ram_cell[    6062] = 32'h0;  // 32'hf4d03ce4;
    ram_cell[    6063] = 32'h0;  // 32'h1e3864cd;
    ram_cell[    6064] = 32'h0;  // 32'h45c596ae;
    ram_cell[    6065] = 32'h0;  // 32'h1df026aa;
    ram_cell[    6066] = 32'h0;  // 32'h37740a30;
    ram_cell[    6067] = 32'h0;  // 32'hc5f5200d;
    ram_cell[    6068] = 32'h0;  // 32'h4020fafd;
    ram_cell[    6069] = 32'h0;  // 32'hbf7e097a;
    ram_cell[    6070] = 32'h0;  // 32'h3e755296;
    ram_cell[    6071] = 32'h0;  // 32'hb3618dfa;
    ram_cell[    6072] = 32'h0;  // 32'hcf516fa2;
    ram_cell[    6073] = 32'h0;  // 32'hec9ba491;
    ram_cell[    6074] = 32'h0;  // 32'ha6911a22;
    ram_cell[    6075] = 32'h0;  // 32'h87df6d0e;
    ram_cell[    6076] = 32'h0;  // 32'h06283b52;
    ram_cell[    6077] = 32'h0;  // 32'h5c47e981;
    ram_cell[    6078] = 32'h0;  // 32'hf1f3d1ef;
    ram_cell[    6079] = 32'h0;  // 32'h6271921a;
    ram_cell[    6080] = 32'h0;  // 32'h375fedea;
    ram_cell[    6081] = 32'h0;  // 32'h1fd52433;
    ram_cell[    6082] = 32'h0;  // 32'h097477b7;
    ram_cell[    6083] = 32'h0;  // 32'hf3d64f97;
    ram_cell[    6084] = 32'h0;  // 32'hb7e18bbb;
    ram_cell[    6085] = 32'h0;  // 32'h1a8d0c84;
    ram_cell[    6086] = 32'h0;  // 32'hca37b55b;
    ram_cell[    6087] = 32'h0;  // 32'h0b9cf2fc;
    ram_cell[    6088] = 32'h0;  // 32'h110d4b92;
    ram_cell[    6089] = 32'h0;  // 32'hd3f052bf;
    ram_cell[    6090] = 32'h0;  // 32'hc536891c;
    ram_cell[    6091] = 32'h0;  // 32'ha319947c;
    ram_cell[    6092] = 32'h0;  // 32'h60a48809;
    ram_cell[    6093] = 32'h0;  // 32'h69bc4f22;
    ram_cell[    6094] = 32'h0;  // 32'h746e1fdd;
    ram_cell[    6095] = 32'h0;  // 32'hca35fc6b;
    ram_cell[    6096] = 32'h0;  // 32'he9feb9fd;
    ram_cell[    6097] = 32'h0;  // 32'h47aaff99;
    ram_cell[    6098] = 32'h0;  // 32'ha663357f;
    ram_cell[    6099] = 32'h0;  // 32'hf2f0ddf9;
    ram_cell[    6100] = 32'h0;  // 32'he0c2f1a5;
    ram_cell[    6101] = 32'h0;  // 32'h1535caaf;
    ram_cell[    6102] = 32'h0;  // 32'h717c13f8;
    ram_cell[    6103] = 32'h0;  // 32'hee6684fc;
    ram_cell[    6104] = 32'h0;  // 32'habb79412;
    ram_cell[    6105] = 32'h0;  // 32'ha40e3ad3;
    ram_cell[    6106] = 32'h0;  // 32'h74332e67;
    ram_cell[    6107] = 32'h0;  // 32'h7a4bbb76;
    ram_cell[    6108] = 32'h0;  // 32'h16bc48e5;
    ram_cell[    6109] = 32'h0;  // 32'h4e93f95e;
    ram_cell[    6110] = 32'h0;  // 32'h34691fc1;
    ram_cell[    6111] = 32'h0;  // 32'hdf0a769a;
    ram_cell[    6112] = 32'h0;  // 32'he5e86499;
    ram_cell[    6113] = 32'h0;  // 32'h735f3568;
    ram_cell[    6114] = 32'h0;  // 32'hdd438e61;
    ram_cell[    6115] = 32'h0;  // 32'hb0593a0f;
    ram_cell[    6116] = 32'h0;  // 32'h0ce5048f;
    ram_cell[    6117] = 32'h0;  // 32'h5f48002c;
    ram_cell[    6118] = 32'h0;  // 32'ha12c394a;
    ram_cell[    6119] = 32'h0;  // 32'h618caa49;
    ram_cell[    6120] = 32'h0;  // 32'hb9721491;
    ram_cell[    6121] = 32'h0;  // 32'h1c1a92ed;
    ram_cell[    6122] = 32'h0;  // 32'h17e7874f;
    ram_cell[    6123] = 32'h0;  // 32'h7bfbfcd1;
    ram_cell[    6124] = 32'h0;  // 32'hd1f5aff4;
    ram_cell[    6125] = 32'h0;  // 32'h79baefca;
    ram_cell[    6126] = 32'h0;  // 32'h493fb7d8;
    ram_cell[    6127] = 32'h0;  // 32'h458d0db4;
    ram_cell[    6128] = 32'h0;  // 32'had6052f4;
    ram_cell[    6129] = 32'h0;  // 32'he7f2b165;
    ram_cell[    6130] = 32'h0;  // 32'heab06829;
    ram_cell[    6131] = 32'h0;  // 32'h86913564;
    ram_cell[    6132] = 32'h0;  // 32'h06244f9f;
    ram_cell[    6133] = 32'h0;  // 32'h06d26859;
    ram_cell[    6134] = 32'h0;  // 32'he6893825;
    ram_cell[    6135] = 32'h0;  // 32'h20de25f8;
    ram_cell[    6136] = 32'h0;  // 32'h8eea07da;
    ram_cell[    6137] = 32'h0;  // 32'h69ef78bb;
    ram_cell[    6138] = 32'h0;  // 32'hd49e2a87;
    ram_cell[    6139] = 32'h0;  // 32'hc610e39b;
    ram_cell[    6140] = 32'h0;  // 32'ha9454160;
    ram_cell[    6141] = 32'h0;  // 32'hcbe6b908;
    ram_cell[    6142] = 32'h0;  // 32'hdd41bdcb;
    ram_cell[    6143] = 32'h0;  // 32'h50d0c305;
    ram_cell[    6144] = 32'h0;  // 32'hb837c7db;
    ram_cell[    6145] = 32'h0;  // 32'h949dd985;
    ram_cell[    6146] = 32'h0;  // 32'h745576ad;
    ram_cell[    6147] = 32'h0;  // 32'h021d806d;
    ram_cell[    6148] = 32'h0;  // 32'h3ff4907b;
    ram_cell[    6149] = 32'h0;  // 32'h74af5a67;
    ram_cell[    6150] = 32'h0;  // 32'hb5712cee;
    ram_cell[    6151] = 32'h0;  // 32'h6afc2a2d;
    ram_cell[    6152] = 32'h0;  // 32'h7d4dcc2b;
    ram_cell[    6153] = 32'h0;  // 32'hf7a1b15f;
    ram_cell[    6154] = 32'h0;  // 32'hf1718d61;
    ram_cell[    6155] = 32'h0;  // 32'h15b6a930;
    ram_cell[    6156] = 32'h0;  // 32'h518da446;
    ram_cell[    6157] = 32'h0;  // 32'h292e3f1a;
    ram_cell[    6158] = 32'h0;  // 32'hae50c172;
    ram_cell[    6159] = 32'h0;  // 32'h759ad7fc;
    ram_cell[    6160] = 32'h0;  // 32'h58ceb046;
    ram_cell[    6161] = 32'h0;  // 32'he92c1ee2;
    ram_cell[    6162] = 32'h0;  // 32'ha1b842d4;
    ram_cell[    6163] = 32'h0;  // 32'h7b1b64c5;
    ram_cell[    6164] = 32'h0;  // 32'h59d26a65;
    ram_cell[    6165] = 32'h0;  // 32'h60fe6974;
    ram_cell[    6166] = 32'h0;  // 32'hbef1689f;
    ram_cell[    6167] = 32'h0;  // 32'ha83748d9;
    ram_cell[    6168] = 32'h0;  // 32'h391b76e1;
    ram_cell[    6169] = 32'h0;  // 32'hc2328ad3;
    ram_cell[    6170] = 32'h0;  // 32'h85611c25;
    ram_cell[    6171] = 32'h0;  // 32'h863ca5ca;
    ram_cell[    6172] = 32'h0;  // 32'haab5ade4;
    ram_cell[    6173] = 32'h0;  // 32'hc0273044;
    ram_cell[    6174] = 32'h0;  // 32'had7e2323;
    ram_cell[    6175] = 32'h0;  // 32'h4b8a62af;
    ram_cell[    6176] = 32'h0;  // 32'hdf0084db;
    ram_cell[    6177] = 32'h0;  // 32'he6f3c704;
    ram_cell[    6178] = 32'h0;  // 32'hab1e4554;
    ram_cell[    6179] = 32'h0;  // 32'h041d94cc;
    ram_cell[    6180] = 32'h0;  // 32'h7ee332fa;
    ram_cell[    6181] = 32'h0;  // 32'h00cad3a9;
    ram_cell[    6182] = 32'h0;  // 32'h450aec71;
    ram_cell[    6183] = 32'h0;  // 32'h9093024c;
    ram_cell[    6184] = 32'h0;  // 32'h6708652b;
    ram_cell[    6185] = 32'h0;  // 32'h8eef841e;
    ram_cell[    6186] = 32'h0;  // 32'h83656199;
    ram_cell[    6187] = 32'h0;  // 32'h95c7b47c;
    ram_cell[    6188] = 32'h0;  // 32'hd5a24f84;
    ram_cell[    6189] = 32'h0;  // 32'he0ea513b;
    ram_cell[    6190] = 32'h0;  // 32'h21e5409b;
    ram_cell[    6191] = 32'h0;  // 32'ha4133b38;
    ram_cell[    6192] = 32'h0;  // 32'h270efecd;
    ram_cell[    6193] = 32'h0;  // 32'h666bf9a4;
    ram_cell[    6194] = 32'h0;  // 32'h83c1e530;
    ram_cell[    6195] = 32'h0;  // 32'h882fb461;
    ram_cell[    6196] = 32'h0;  // 32'h88bda347;
    ram_cell[    6197] = 32'h0;  // 32'he3b423bd;
    ram_cell[    6198] = 32'h0;  // 32'h5c1b27b7;
    ram_cell[    6199] = 32'h0;  // 32'he24ac1d6;
    ram_cell[    6200] = 32'h0;  // 32'h718aee32;
    ram_cell[    6201] = 32'h0;  // 32'hb0be2860;
    ram_cell[    6202] = 32'h0;  // 32'h360cdcad;
    ram_cell[    6203] = 32'h0;  // 32'h69fb43cc;
    ram_cell[    6204] = 32'h0;  // 32'h74ccade9;
    ram_cell[    6205] = 32'h0;  // 32'hbe03d17a;
    ram_cell[    6206] = 32'h0;  // 32'h2a3529f8;
    ram_cell[    6207] = 32'h0;  // 32'h88b86f86;
    ram_cell[    6208] = 32'h0;  // 32'h4be462c2;
    ram_cell[    6209] = 32'h0;  // 32'haa48b7b6;
    ram_cell[    6210] = 32'h0;  // 32'ha50a23e1;
    ram_cell[    6211] = 32'h0;  // 32'hed975dec;
    ram_cell[    6212] = 32'h0;  // 32'hf921ca83;
    ram_cell[    6213] = 32'h0;  // 32'h633da726;
    ram_cell[    6214] = 32'h0;  // 32'hca5f3f4e;
    ram_cell[    6215] = 32'h0;  // 32'h4b1e515e;
    ram_cell[    6216] = 32'h0;  // 32'h359450f3;
    ram_cell[    6217] = 32'h0;  // 32'h82b91699;
    ram_cell[    6218] = 32'h0;  // 32'hc7151844;
    ram_cell[    6219] = 32'h0;  // 32'h1d7a5df8;
    ram_cell[    6220] = 32'h0;  // 32'h2bc50c00;
    ram_cell[    6221] = 32'h0;  // 32'hee3f2052;
    ram_cell[    6222] = 32'h0;  // 32'h2ba6fb40;
    ram_cell[    6223] = 32'h0;  // 32'he7680ec3;
    ram_cell[    6224] = 32'h0;  // 32'h7aca1240;
    ram_cell[    6225] = 32'h0;  // 32'hab0de27a;
    ram_cell[    6226] = 32'h0;  // 32'h37606b82;
    ram_cell[    6227] = 32'h0;  // 32'ha6697856;
    ram_cell[    6228] = 32'h0;  // 32'h7f243b9b;
    ram_cell[    6229] = 32'h0;  // 32'h499fdc71;
    ram_cell[    6230] = 32'h0;  // 32'h19b26ec7;
    ram_cell[    6231] = 32'h0;  // 32'h69636782;
    ram_cell[    6232] = 32'h0;  // 32'hc2e7fa6c;
    ram_cell[    6233] = 32'h0;  // 32'h9936c0e8;
    ram_cell[    6234] = 32'h0;  // 32'h1ae1bf7a;
    ram_cell[    6235] = 32'h0;  // 32'h5e6161c1;
    ram_cell[    6236] = 32'h0;  // 32'habbbe124;
    ram_cell[    6237] = 32'h0;  // 32'he1ab66a4;
    ram_cell[    6238] = 32'h0;  // 32'hb0d16b5d;
    ram_cell[    6239] = 32'h0;  // 32'h219b1072;
    ram_cell[    6240] = 32'h0;  // 32'he86b181e;
    ram_cell[    6241] = 32'h0;  // 32'h0577087c;
    ram_cell[    6242] = 32'h0;  // 32'hb2e6f07d;
    ram_cell[    6243] = 32'h0;  // 32'hd45b0996;
    ram_cell[    6244] = 32'h0;  // 32'h53dd8a27;
    ram_cell[    6245] = 32'h0;  // 32'h933822c0;
    ram_cell[    6246] = 32'h0;  // 32'hfb520eac;
    ram_cell[    6247] = 32'h0;  // 32'h926db7e2;
    ram_cell[    6248] = 32'h0;  // 32'h22226d33;
    ram_cell[    6249] = 32'h0;  // 32'he4415f65;
    ram_cell[    6250] = 32'h0;  // 32'hb07b96e5;
    ram_cell[    6251] = 32'h0;  // 32'hbdc53551;
    ram_cell[    6252] = 32'h0;  // 32'h478b73e7;
    ram_cell[    6253] = 32'h0;  // 32'ha3411b49;
    ram_cell[    6254] = 32'h0;  // 32'hdc281209;
    ram_cell[    6255] = 32'h0;  // 32'h3b8c407d;
    ram_cell[    6256] = 32'h0;  // 32'h3893316c;
    ram_cell[    6257] = 32'h0;  // 32'ha8aebd39;
    ram_cell[    6258] = 32'h0;  // 32'h2bdf219f;
    ram_cell[    6259] = 32'h0;  // 32'h96b48966;
    ram_cell[    6260] = 32'h0;  // 32'hda035ecc;
    ram_cell[    6261] = 32'h0;  // 32'h80bfc84c;
    ram_cell[    6262] = 32'h0;  // 32'h00f3ba4a;
    ram_cell[    6263] = 32'h0;  // 32'h91a0d0c5;
    ram_cell[    6264] = 32'h0;  // 32'h65557d73;
    ram_cell[    6265] = 32'h0;  // 32'hf2501ea9;
    ram_cell[    6266] = 32'h0;  // 32'h07e93e67;
    ram_cell[    6267] = 32'h0;  // 32'h29956907;
    ram_cell[    6268] = 32'h0;  // 32'hd353c6b3;
    ram_cell[    6269] = 32'h0;  // 32'h2953f95b;
    ram_cell[    6270] = 32'h0;  // 32'h140c5171;
    ram_cell[    6271] = 32'h0;  // 32'hd961a436;
    ram_cell[    6272] = 32'h0;  // 32'hb16f785c;
    ram_cell[    6273] = 32'h0;  // 32'h370269ea;
    ram_cell[    6274] = 32'h0;  // 32'hd2c1e8af;
    ram_cell[    6275] = 32'h0;  // 32'ha80d243a;
    ram_cell[    6276] = 32'h0;  // 32'hee46bb1b;
    ram_cell[    6277] = 32'h0;  // 32'h10948e96;
    ram_cell[    6278] = 32'h0;  // 32'h55c2452b;
    ram_cell[    6279] = 32'h0;  // 32'hf930d87d;
    ram_cell[    6280] = 32'h0;  // 32'hd067c59f;
    ram_cell[    6281] = 32'h0;  // 32'he0855a0c;
    ram_cell[    6282] = 32'h0;  // 32'h65919d5a;
    ram_cell[    6283] = 32'h0;  // 32'h2e584b2d;
    ram_cell[    6284] = 32'h0;  // 32'h213515a7;
    ram_cell[    6285] = 32'h0;  // 32'hd69b4f29;
    ram_cell[    6286] = 32'h0;  // 32'hf0a966a4;
    ram_cell[    6287] = 32'h0;  // 32'h7db9f009;
    ram_cell[    6288] = 32'h0;  // 32'heb8366bf;
    ram_cell[    6289] = 32'h0;  // 32'h2d1f42cb;
    ram_cell[    6290] = 32'h0;  // 32'hdef8ad5e;
    ram_cell[    6291] = 32'h0;  // 32'h2a220664;
    ram_cell[    6292] = 32'h0;  // 32'h6dbfa55e;
    ram_cell[    6293] = 32'h0;  // 32'hbf4bc5a4;
    ram_cell[    6294] = 32'h0;  // 32'h91ad6d9d;
    ram_cell[    6295] = 32'h0;  // 32'h8d024dbc;
    ram_cell[    6296] = 32'h0;  // 32'h2e363e68;
    ram_cell[    6297] = 32'h0;  // 32'h45801992;
    ram_cell[    6298] = 32'h0;  // 32'h8578dbe0;
    ram_cell[    6299] = 32'h0;  // 32'hbe70adf2;
    ram_cell[    6300] = 32'h0;  // 32'h5d2655ee;
    ram_cell[    6301] = 32'h0;  // 32'hbe640d95;
    ram_cell[    6302] = 32'h0;  // 32'h1e545012;
    ram_cell[    6303] = 32'h0;  // 32'h908de15c;
    ram_cell[    6304] = 32'h0;  // 32'h3488b9c8;
    ram_cell[    6305] = 32'h0;  // 32'h483d74df;
    ram_cell[    6306] = 32'h0;  // 32'h5c2fc92d;
    ram_cell[    6307] = 32'h0;  // 32'hc4df61a6;
    ram_cell[    6308] = 32'h0;  // 32'h85177408;
    ram_cell[    6309] = 32'h0;  // 32'h72c41e2e;
    ram_cell[    6310] = 32'h0;  // 32'h72883777;
    ram_cell[    6311] = 32'h0;  // 32'h9e83fe73;
    ram_cell[    6312] = 32'h0;  // 32'h93bf68a0;
    ram_cell[    6313] = 32'h0;  // 32'h1e930052;
    ram_cell[    6314] = 32'h0;  // 32'h3b0aa8ef;
    ram_cell[    6315] = 32'h0;  // 32'habfa429d;
    ram_cell[    6316] = 32'h0;  // 32'hbc3868d4;
    ram_cell[    6317] = 32'h0;  // 32'h1766b273;
    ram_cell[    6318] = 32'h0;  // 32'ha51b164e;
    ram_cell[    6319] = 32'h0;  // 32'hdbafe8c8;
    ram_cell[    6320] = 32'h0;  // 32'h7e3a43cd;
    ram_cell[    6321] = 32'h0;  // 32'h69c8121f;
    ram_cell[    6322] = 32'h0;  // 32'had6ece8e;
    ram_cell[    6323] = 32'h0;  // 32'hed6e1058;
    ram_cell[    6324] = 32'h0;  // 32'h229f13d4;
    ram_cell[    6325] = 32'h0;  // 32'h7ab1e5d5;
    ram_cell[    6326] = 32'h0;  // 32'h69e32367;
    ram_cell[    6327] = 32'h0;  // 32'hcfdba0ec;
    ram_cell[    6328] = 32'h0;  // 32'h41441c9d;
    ram_cell[    6329] = 32'h0;  // 32'h5dc7cf70;
    ram_cell[    6330] = 32'h0;  // 32'h525bb169;
    ram_cell[    6331] = 32'h0;  // 32'he4b6829f;
    ram_cell[    6332] = 32'h0;  // 32'h1e0d1ab9;
    ram_cell[    6333] = 32'h0;  // 32'h4c073cb8;
    ram_cell[    6334] = 32'h0;  // 32'h2f4c9f42;
    ram_cell[    6335] = 32'h0;  // 32'h6135e5b0;
    ram_cell[    6336] = 32'h0;  // 32'he13cb582;
    ram_cell[    6337] = 32'h0;  // 32'h70f32f20;
    ram_cell[    6338] = 32'h0;  // 32'hd151beec;
    ram_cell[    6339] = 32'h0;  // 32'h53155b24;
    ram_cell[    6340] = 32'h0;  // 32'h92f60094;
    ram_cell[    6341] = 32'h0;  // 32'h72bd5b3a;
    ram_cell[    6342] = 32'h0;  // 32'hed31a83b;
    ram_cell[    6343] = 32'h0;  // 32'h79ec610b;
    ram_cell[    6344] = 32'h0;  // 32'h6f783d6d;
    ram_cell[    6345] = 32'h0;  // 32'h13dabb3f;
    ram_cell[    6346] = 32'h0;  // 32'h1f151d7d;
    ram_cell[    6347] = 32'h0;  // 32'hbe67c2ad;
    ram_cell[    6348] = 32'h0;  // 32'h2f171e48;
    ram_cell[    6349] = 32'h0;  // 32'h90bb99ed;
    ram_cell[    6350] = 32'h0;  // 32'h06671db4;
    ram_cell[    6351] = 32'h0;  // 32'h2a43b220;
    ram_cell[    6352] = 32'h0;  // 32'h479e7658;
    ram_cell[    6353] = 32'h0;  // 32'h8aaad4d8;
    ram_cell[    6354] = 32'h0;  // 32'h18a017c7;
    ram_cell[    6355] = 32'h0;  // 32'h6cc13963;
    ram_cell[    6356] = 32'h0;  // 32'hc4f2c04b;
    ram_cell[    6357] = 32'h0;  // 32'h39f83532;
    ram_cell[    6358] = 32'h0;  // 32'ha33e2925;
    ram_cell[    6359] = 32'h0;  // 32'h6755f728;
    ram_cell[    6360] = 32'h0;  // 32'hb0435f36;
    ram_cell[    6361] = 32'h0;  // 32'hdc12011e;
    ram_cell[    6362] = 32'h0;  // 32'hb9806ab5;
    ram_cell[    6363] = 32'h0;  // 32'h8081acfc;
    ram_cell[    6364] = 32'h0;  // 32'h4f2569db;
    ram_cell[    6365] = 32'h0;  // 32'hd623c23d;
    ram_cell[    6366] = 32'h0;  // 32'h9a6bb68f;
    ram_cell[    6367] = 32'h0;  // 32'h13ff860b;
    ram_cell[    6368] = 32'h0;  // 32'hb66e87d7;
    ram_cell[    6369] = 32'h0;  // 32'hf12388b0;
    ram_cell[    6370] = 32'h0;  // 32'hcb99d847;
    ram_cell[    6371] = 32'h0;  // 32'hfa868654;
    ram_cell[    6372] = 32'h0;  // 32'h46f4586d;
    ram_cell[    6373] = 32'h0;  // 32'h40c3aab3;
    ram_cell[    6374] = 32'h0;  // 32'h24bd6d16;
    ram_cell[    6375] = 32'h0;  // 32'h6d44906a;
    ram_cell[    6376] = 32'h0;  // 32'h1a7ed837;
    ram_cell[    6377] = 32'h0;  // 32'h4ea07912;
    ram_cell[    6378] = 32'h0;  // 32'he2846959;
    ram_cell[    6379] = 32'h0;  // 32'he5c2f9b7;
    ram_cell[    6380] = 32'h0;  // 32'h8b7cd108;
    ram_cell[    6381] = 32'h0;  // 32'h1fc3a858;
    ram_cell[    6382] = 32'h0;  // 32'hed3c4b95;
    ram_cell[    6383] = 32'h0;  // 32'h1f0b5dfe;
    ram_cell[    6384] = 32'h0;  // 32'h1aef601f;
    ram_cell[    6385] = 32'h0;  // 32'h9677a184;
    ram_cell[    6386] = 32'h0;  // 32'ha166ab52;
    ram_cell[    6387] = 32'h0;  // 32'h30619b5e;
    ram_cell[    6388] = 32'h0;  // 32'hf1e9ef00;
    ram_cell[    6389] = 32'h0;  // 32'hedcc29ce;
    ram_cell[    6390] = 32'h0;  // 32'h5007dfb5;
    ram_cell[    6391] = 32'h0;  // 32'h906044b0;
    ram_cell[    6392] = 32'h0;  // 32'h349517f7;
    ram_cell[    6393] = 32'h0;  // 32'h18aa0333;
    ram_cell[    6394] = 32'h0;  // 32'hdea2e598;
    ram_cell[    6395] = 32'h0;  // 32'h8f88f3ab;
    ram_cell[    6396] = 32'h0;  // 32'hc9fa8834;
    ram_cell[    6397] = 32'h0;  // 32'hfc1af6a0;
    ram_cell[    6398] = 32'h0;  // 32'hd9bbf975;
    ram_cell[    6399] = 32'h0;  // 32'hd6b969a5;
    ram_cell[    6400] = 32'h0;  // 32'h4495a5e8;
    ram_cell[    6401] = 32'h0;  // 32'hd2224d12;
    ram_cell[    6402] = 32'h0;  // 32'h87235da3;
    ram_cell[    6403] = 32'h0;  // 32'h9fad1941;
    ram_cell[    6404] = 32'h0;  // 32'h9606bd3c;
    ram_cell[    6405] = 32'h0;  // 32'h915a7e00;
    ram_cell[    6406] = 32'h0;  // 32'hd9a2fb94;
    ram_cell[    6407] = 32'h0;  // 32'h1483ddbb;
    ram_cell[    6408] = 32'h0;  // 32'h4218adbc;
    ram_cell[    6409] = 32'h0;  // 32'hd54d37d2;
    ram_cell[    6410] = 32'h0;  // 32'h16b6ec02;
    ram_cell[    6411] = 32'h0;  // 32'h1bfc2841;
    ram_cell[    6412] = 32'h0;  // 32'hdf6f4e21;
    ram_cell[    6413] = 32'h0;  // 32'h65e907d2;
    ram_cell[    6414] = 32'h0;  // 32'h84b30597;
    ram_cell[    6415] = 32'h0;  // 32'h06721985;
    ram_cell[    6416] = 32'h0;  // 32'he4d647dc;
    ram_cell[    6417] = 32'h0;  // 32'h337c2d09;
    ram_cell[    6418] = 32'h0;  // 32'h9a01681e;
    ram_cell[    6419] = 32'h0;  // 32'hcf4817cf;
    ram_cell[    6420] = 32'h0;  // 32'h5343ae02;
    ram_cell[    6421] = 32'h0;  // 32'h015239bc;
    ram_cell[    6422] = 32'h0;  // 32'h7d335336;
    ram_cell[    6423] = 32'h0;  // 32'h7db6b67d;
    ram_cell[    6424] = 32'h0;  // 32'h8763e3ab;
    ram_cell[    6425] = 32'h0;  // 32'hc0bad6a1;
    ram_cell[    6426] = 32'h0;  // 32'h0fdd413a;
    ram_cell[    6427] = 32'h0;  // 32'h9a75fa95;
    ram_cell[    6428] = 32'h0;  // 32'h13f343d2;
    ram_cell[    6429] = 32'h0;  // 32'hd025642c;
    ram_cell[    6430] = 32'h0;  // 32'ha23e2ae4;
    ram_cell[    6431] = 32'h0;  // 32'h45158932;
    ram_cell[    6432] = 32'h0;  // 32'h9bab2917;
    ram_cell[    6433] = 32'h0;  // 32'h3d50918a;
    ram_cell[    6434] = 32'h0;  // 32'hb0817036;
    ram_cell[    6435] = 32'h0;  // 32'h30955605;
    ram_cell[    6436] = 32'h0;  // 32'h8fec0785;
    ram_cell[    6437] = 32'h0;  // 32'hf76dfb6e;
    ram_cell[    6438] = 32'h0;  // 32'h6a98ee4c;
    ram_cell[    6439] = 32'h0;  // 32'hedffe969;
    ram_cell[    6440] = 32'h0;  // 32'he43e2f14;
    ram_cell[    6441] = 32'h0;  // 32'h3fa945e3;
    ram_cell[    6442] = 32'h0;  // 32'hc1765fb9;
    ram_cell[    6443] = 32'h0;  // 32'h5e13e6db;
    ram_cell[    6444] = 32'h0;  // 32'h3d9e6358;
    ram_cell[    6445] = 32'h0;  // 32'h76b3edfd;
    ram_cell[    6446] = 32'h0;  // 32'h7651dfd5;
    ram_cell[    6447] = 32'h0;  // 32'h85e266c9;
    ram_cell[    6448] = 32'h0;  // 32'h4ee237b1;
    ram_cell[    6449] = 32'h0;  // 32'h1d6b2f55;
    ram_cell[    6450] = 32'h0;  // 32'h90e46162;
    ram_cell[    6451] = 32'h0;  // 32'h552f34e9;
    ram_cell[    6452] = 32'h0;  // 32'h5eef45d6;
    ram_cell[    6453] = 32'h0;  // 32'h40052b13;
    ram_cell[    6454] = 32'h0;  // 32'hab1d6245;
    ram_cell[    6455] = 32'h0;  // 32'hf4609b50;
    ram_cell[    6456] = 32'h0;  // 32'h663e66c3;
    ram_cell[    6457] = 32'h0;  // 32'h41884ed7;
    ram_cell[    6458] = 32'h0;  // 32'hf22b9e78;
    ram_cell[    6459] = 32'h0;  // 32'h098c2ce2;
    ram_cell[    6460] = 32'h0;  // 32'hece29e9f;
    ram_cell[    6461] = 32'h0;  // 32'h70ab51ec;
    ram_cell[    6462] = 32'h0;  // 32'h529cfeda;
    ram_cell[    6463] = 32'h0;  // 32'h3aa82533;
    ram_cell[    6464] = 32'h0;  // 32'he31289be;
    ram_cell[    6465] = 32'h0;  // 32'h703ccc8b;
    ram_cell[    6466] = 32'h0;  // 32'h6ed6ddd7;
    ram_cell[    6467] = 32'h0;  // 32'h10ea6aab;
    ram_cell[    6468] = 32'h0;  // 32'hca3f9169;
    ram_cell[    6469] = 32'h0;  // 32'ha0ffa2d6;
    ram_cell[    6470] = 32'h0;  // 32'h74a38f0b;
    ram_cell[    6471] = 32'h0;  // 32'h7353b879;
    ram_cell[    6472] = 32'h0;  // 32'h5f05b80c;
    ram_cell[    6473] = 32'h0;  // 32'h27103814;
    ram_cell[    6474] = 32'h0;  // 32'hf1f1d34c;
    ram_cell[    6475] = 32'h0;  // 32'h3169333d;
    ram_cell[    6476] = 32'h0;  // 32'hc627ad78;
    ram_cell[    6477] = 32'h0;  // 32'h7e7580fc;
    ram_cell[    6478] = 32'h0;  // 32'h7e78af35;
    ram_cell[    6479] = 32'h0;  // 32'h1cc88020;
    ram_cell[    6480] = 32'h0;  // 32'h3488bfe4;
    ram_cell[    6481] = 32'h0;  // 32'hf62c8324;
    ram_cell[    6482] = 32'h0;  // 32'h57b1ff7f;
    ram_cell[    6483] = 32'h0;  // 32'hdce1ce43;
    ram_cell[    6484] = 32'h0;  // 32'h1615aea7;
    ram_cell[    6485] = 32'h0;  // 32'h53da4ed4;
    ram_cell[    6486] = 32'h0;  // 32'h530ed045;
    ram_cell[    6487] = 32'h0;  // 32'h1a3a3572;
    ram_cell[    6488] = 32'h0;  // 32'h207d6d17;
    ram_cell[    6489] = 32'h0;  // 32'h3746d4cb;
    ram_cell[    6490] = 32'h0;  // 32'h259f4019;
    ram_cell[    6491] = 32'h0;  // 32'h7521d5e5;
    ram_cell[    6492] = 32'h0;  // 32'h55e19dcf;
    ram_cell[    6493] = 32'h0;  // 32'hcadae361;
    ram_cell[    6494] = 32'h0;  // 32'h7f9541cd;
    ram_cell[    6495] = 32'h0;  // 32'h2fc34188;
    ram_cell[    6496] = 32'h0;  // 32'h01460f62;
    ram_cell[    6497] = 32'h0;  // 32'h42349c6d;
    ram_cell[    6498] = 32'h0;  // 32'hc8e5610b;
    ram_cell[    6499] = 32'h0;  // 32'h9b59f208;
    ram_cell[    6500] = 32'h0;  // 32'hfffcfa88;
    ram_cell[    6501] = 32'h0;  // 32'hcce0513d;
    ram_cell[    6502] = 32'h0;  // 32'hd9cb9169;
    ram_cell[    6503] = 32'h0;  // 32'h92c1da03;
    ram_cell[    6504] = 32'h0;  // 32'hdc2905a6;
    ram_cell[    6505] = 32'h0;  // 32'h93860c9b;
    ram_cell[    6506] = 32'h0;  // 32'h25c8f89a;
    ram_cell[    6507] = 32'h0;  // 32'hbaef7290;
    ram_cell[    6508] = 32'h0;  // 32'hd55022dc;
    ram_cell[    6509] = 32'h0;  // 32'hce15ef59;
    ram_cell[    6510] = 32'h0;  // 32'h0d0a23b2;
    ram_cell[    6511] = 32'h0;  // 32'hdcb4e3d9;
    ram_cell[    6512] = 32'h0;  // 32'h7bb75f42;
    ram_cell[    6513] = 32'h0;  // 32'h8b7ed931;
    ram_cell[    6514] = 32'h0;  // 32'h9132360f;
    ram_cell[    6515] = 32'h0;  // 32'hb201dd6e;
    ram_cell[    6516] = 32'h0;  // 32'hf4d1d8ac;
    ram_cell[    6517] = 32'h0;  // 32'h42c48cb4;
    ram_cell[    6518] = 32'h0;  // 32'h25cc7720;
    ram_cell[    6519] = 32'h0;  // 32'h6adeda1a;
    ram_cell[    6520] = 32'h0;  // 32'h9288d30c;
    ram_cell[    6521] = 32'h0;  // 32'h2f757957;
    ram_cell[    6522] = 32'h0;  // 32'hfc2a94df;
    ram_cell[    6523] = 32'h0;  // 32'h9ab61edd;
    ram_cell[    6524] = 32'h0;  // 32'h08168b0f;
    ram_cell[    6525] = 32'h0;  // 32'h2b43e9f2;
    ram_cell[    6526] = 32'h0;  // 32'h173c7c94;
    ram_cell[    6527] = 32'h0;  // 32'h472273a6;
    ram_cell[    6528] = 32'h0;  // 32'he3fa4bfa;
    ram_cell[    6529] = 32'h0;  // 32'h449c513d;
    ram_cell[    6530] = 32'h0;  // 32'hb480232c;
    ram_cell[    6531] = 32'h0;  // 32'h290a1f49;
    ram_cell[    6532] = 32'h0;  // 32'h2bc87d32;
    ram_cell[    6533] = 32'h0;  // 32'hdac53e6a;
    ram_cell[    6534] = 32'h0;  // 32'h7df57023;
    ram_cell[    6535] = 32'h0;  // 32'h9db32350;
    ram_cell[    6536] = 32'h0;  // 32'hd4b50eee;
    ram_cell[    6537] = 32'h0;  // 32'h9494c46e;
    ram_cell[    6538] = 32'h0;  // 32'h83f77340;
    ram_cell[    6539] = 32'h0;  // 32'h484811f5;
    ram_cell[    6540] = 32'h0;  // 32'h02a8ed8d;
    ram_cell[    6541] = 32'h0;  // 32'hc0b3e79b;
    ram_cell[    6542] = 32'h0;  // 32'haf600d4d;
    ram_cell[    6543] = 32'h0;  // 32'h6a6cff9a;
    ram_cell[    6544] = 32'h0;  // 32'hd247da8e;
    ram_cell[    6545] = 32'h0;  // 32'h990b7c66;
    ram_cell[    6546] = 32'h0;  // 32'hecf1cf0f;
    ram_cell[    6547] = 32'h0;  // 32'h7b49c38b;
    ram_cell[    6548] = 32'h0;  // 32'hcef5dcf6;
    ram_cell[    6549] = 32'h0;  // 32'h3937bb35;
    ram_cell[    6550] = 32'h0;  // 32'ha49c9848;
    ram_cell[    6551] = 32'h0;  // 32'h5bda33ee;
    ram_cell[    6552] = 32'h0;  // 32'h677e2dde;
    ram_cell[    6553] = 32'h0;  // 32'h4e6add10;
    ram_cell[    6554] = 32'h0;  // 32'haf92d8b3;
    ram_cell[    6555] = 32'h0;  // 32'hba3a3c34;
    ram_cell[    6556] = 32'h0;  // 32'h021ae9c5;
    ram_cell[    6557] = 32'h0;  // 32'he0c90a11;
    ram_cell[    6558] = 32'h0;  // 32'h7a45fa86;
    ram_cell[    6559] = 32'h0;  // 32'h20a9035f;
    ram_cell[    6560] = 32'h0;  // 32'h8536a2d3;
    ram_cell[    6561] = 32'h0;  // 32'hf5528d05;
    ram_cell[    6562] = 32'h0;  // 32'h97f811d4;
    ram_cell[    6563] = 32'h0;  // 32'h970424ab;
    ram_cell[    6564] = 32'h0;  // 32'h75ec8d06;
    ram_cell[    6565] = 32'h0;  // 32'he8e66aca;
    ram_cell[    6566] = 32'h0;  // 32'ha3fce89d;
    ram_cell[    6567] = 32'h0;  // 32'h8818f987;
    ram_cell[    6568] = 32'h0;  // 32'h45c864e1;
    ram_cell[    6569] = 32'h0;  // 32'hc2b588f7;
    ram_cell[    6570] = 32'h0;  // 32'h916fabe1;
    ram_cell[    6571] = 32'h0;  // 32'h61d91479;
    ram_cell[    6572] = 32'h0;  // 32'h3fa75612;
    ram_cell[    6573] = 32'h0;  // 32'hebae8d6b;
    ram_cell[    6574] = 32'h0;  // 32'h49b949f1;
    ram_cell[    6575] = 32'h0;  // 32'h9424f54c;
    ram_cell[    6576] = 32'h0;  // 32'h21bd67fc;
    ram_cell[    6577] = 32'h0;  // 32'he9a17117;
    ram_cell[    6578] = 32'h0;  // 32'hccb39eb2;
    ram_cell[    6579] = 32'h0;  // 32'hdb2375e9;
    ram_cell[    6580] = 32'h0;  // 32'h65381303;
    ram_cell[    6581] = 32'h0;  // 32'h399fa5e7;
    ram_cell[    6582] = 32'h0;  // 32'hf89bbdc5;
    ram_cell[    6583] = 32'h0;  // 32'h6af03b8c;
    ram_cell[    6584] = 32'h0;  // 32'h943353fd;
    ram_cell[    6585] = 32'h0;  // 32'ha67fa08e;
    ram_cell[    6586] = 32'h0;  // 32'h896008dd;
    ram_cell[    6587] = 32'h0;  // 32'h8c5fcd8a;
    ram_cell[    6588] = 32'h0;  // 32'h5d601787;
    ram_cell[    6589] = 32'h0;  // 32'hc08c2d33;
    ram_cell[    6590] = 32'h0;  // 32'h801653dc;
    ram_cell[    6591] = 32'h0;  // 32'h5e48217b;
    ram_cell[    6592] = 32'h0;  // 32'hbe50abad;
    ram_cell[    6593] = 32'h0;  // 32'h50666a80;
    ram_cell[    6594] = 32'h0;  // 32'he644d5c5;
    ram_cell[    6595] = 32'h0;  // 32'h9907a7be;
    ram_cell[    6596] = 32'h0;  // 32'h947b2b17;
    ram_cell[    6597] = 32'h0;  // 32'hfc9cb6e4;
    ram_cell[    6598] = 32'h0;  // 32'h6ed9b152;
    ram_cell[    6599] = 32'h0;  // 32'h6827bcf0;
    ram_cell[    6600] = 32'h0;  // 32'hfeb7b737;
    ram_cell[    6601] = 32'h0;  // 32'hd3c53322;
    ram_cell[    6602] = 32'h0;  // 32'hdfcaed65;
    ram_cell[    6603] = 32'h0;  // 32'h9efe208b;
    ram_cell[    6604] = 32'h0;  // 32'hc59929f2;
    ram_cell[    6605] = 32'h0;  // 32'h011de3c6;
    ram_cell[    6606] = 32'h0;  // 32'h1c5a7ffe;
    ram_cell[    6607] = 32'h0;  // 32'h178625fa;
    ram_cell[    6608] = 32'h0;  // 32'h27629a1d;
    ram_cell[    6609] = 32'h0;  // 32'h78ce1e0e;
    ram_cell[    6610] = 32'h0;  // 32'h4b4bacec;
    ram_cell[    6611] = 32'h0;  // 32'h016f78e0;
    ram_cell[    6612] = 32'h0;  // 32'h0591694e;
    ram_cell[    6613] = 32'h0;  // 32'h71994441;
    ram_cell[    6614] = 32'h0;  // 32'ha4da64d5;
    ram_cell[    6615] = 32'h0;  // 32'h07640c9b;
    ram_cell[    6616] = 32'h0;  // 32'h1db056da;
    ram_cell[    6617] = 32'h0;  // 32'h32f7555c;
    ram_cell[    6618] = 32'h0;  // 32'hc8740a9e;
    ram_cell[    6619] = 32'h0;  // 32'h572aa0bb;
    ram_cell[    6620] = 32'h0;  // 32'hf1676caa;
    ram_cell[    6621] = 32'h0;  // 32'hc9d7e6cf;
    ram_cell[    6622] = 32'h0;  // 32'h26a80375;
    ram_cell[    6623] = 32'h0;  // 32'h0b185154;
    ram_cell[    6624] = 32'h0;  // 32'hdf0585d1;
    ram_cell[    6625] = 32'h0;  // 32'hbd56e88a;
    ram_cell[    6626] = 32'h0;  // 32'h0549d7ed;
    ram_cell[    6627] = 32'h0;  // 32'h56d39794;
    ram_cell[    6628] = 32'h0;  // 32'h8f105c19;
    ram_cell[    6629] = 32'h0;  // 32'h529f0e75;
    ram_cell[    6630] = 32'h0;  // 32'h923b8712;
    ram_cell[    6631] = 32'h0;  // 32'hc5456787;
    ram_cell[    6632] = 32'h0;  // 32'he5027e6e;
    ram_cell[    6633] = 32'h0;  // 32'hbcb76724;
    ram_cell[    6634] = 32'h0;  // 32'ha65aa3aa;
    ram_cell[    6635] = 32'h0;  // 32'h0d4854f1;
    ram_cell[    6636] = 32'h0;  // 32'hcbac1328;
    ram_cell[    6637] = 32'h0;  // 32'h384fb87a;
    ram_cell[    6638] = 32'h0;  // 32'h65625f93;
    ram_cell[    6639] = 32'h0;  // 32'hdc98e41d;
    ram_cell[    6640] = 32'h0;  // 32'h7c67358b;
    ram_cell[    6641] = 32'h0;  // 32'he2b3e928;
    ram_cell[    6642] = 32'h0;  // 32'ha8edf667;
    ram_cell[    6643] = 32'h0;  // 32'h3507c201;
    ram_cell[    6644] = 32'h0;  // 32'h7a1b9540;
    ram_cell[    6645] = 32'h0;  // 32'h88ee9e10;
    ram_cell[    6646] = 32'h0;  // 32'h93061db1;
    ram_cell[    6647] = 32'h0;  // 32'hc842cc64;
    ram_cell[    6648] = 32'h0;  // 32'h70f46456;
    ram_cell[    6649] = 32'h0;  // 32'hc3a7e774;
    ram_cell[    6650] = 32'h0;  // 32'h19e7a207;
    ram_cell[    6651] = 32'h0;  // 32'h8813cbce;
    ram_cell[    6652] = 32'h0;  // 32'h7d504a1d;
    ram_cell[    6653] = 32'h0;  // 32'h2d2d16e9;
    ram_cell[    6654] = 32'h0;  // 32'hd365570f;
    ram_cell[    6655] = 32'h0;  // 32'h2a63698f;
    ram_cell[    6656] = 32'h0;  // 32'h4cd58351;
    ram_cell[    6657] = 32'h0;  // 32'hffc8e76e;
    ram_cell[    6658] = 32'h0;  // 32'h8ffe8a53;
    ram_cell[    6659] = 32'h0;  // 32'h21b48743;
    ram_cell[    6660] = 32'h0;  // 32'hf3a23ea8;
    ram_cell[    6661] = 32'h0;  // 32'heea6909e;
    ram_cell[    6662] = 32'h0;  // 32'h1bed7aec;
    ram_cell[    6663] = 32'h0;  // 32'ha105d235;
    ram_cell[    6664] = 32'h0;  // 32'h566b33de;
    ram_cell[    6665] = 32'h0;  // 32'hefa5ed22;
    ram_cell[    6666] = 32'h0;  // 32'h2e35c29d;
    ram_cell[    6667] = 32'h0;  // 32'h735863f9;
    ram_cell[    6668] = 32'h0;  // 32'h0243dda0;
    ram_cell[    6669] = 32'h0;  // 32'hcc2a8d13;
    ram_cell[    6670] = 32'h0;  // 32'h695e6ccd;
    ram_cell[    6671] = 32'h0;  // 32'heb2e84e1;
    ram_cell[    6672] = 32'h0;  // 32'h21709527;
    ram_cell[    6673] = 32'h0;  // 32'h59ff72e8;
    ram_cell[    6674] = 32'h0;  // 32'h0c2ca367;
    ram_cell[    6675] = 32'h0;  // 32'h5513e3e8;
    ram_cell[    6676] = 32'h0;  // 32'h679ad3a9;
    ram_cell[    6677] = 32'h0;  // 32'hd6b65f64;
    ram_cell[    6678] = 32'h0;  // 32'hed2bf268;
    ram_cell[    6679] = 32'h0;  // 32'h6ae53e3e;
    ram_cell[    6680] = 32'h0;  // 32'hb9e27f89;
    ram_cell[    6681] = 32'h0;  // 32'haed48624;
    ram_cell[    6682] = 32'h0;  // 32'h5cdc9b17;
    ram_cell[    6683] = 32'h0;  // 32'h53ed6971;
    ram_cell[    6684] = 32'h0;  // 32'h429b8aa7;
    ram_cell[    6685] = 32'h0;  // 32'h61e86985;
    ram_cell[    6686] = 32'h0;  // 32'hc9e59922;
    ram_cell[    6687] = 32'h0;  // 32'h910201c9;
    ram_cell[    6688] = 32'h0;  // 32'h6f23eae6;
    ram_cell[    6689] = 32'h0;  // 32'h6677dea7;
    ram_cell[    6690] = 32'h0;  // 32'h4ca092ec;
    ram_cell[    6691] = 32'h0;  // 32'h66d3dbf1;
    ram_cell[    6692] = 32'h0;  // 32'hbe67131e;
    ram_cell[    6693] = 32'h0;  // 32'h86d07281;
    ram_cell[    6694] = 32'h0;  // 32'h11b8f609;
    ram_cell[    6695] = 32'h0;  // 32'hc5d00d8b;
    ram_cell[    6696] = 32'h0;  // 32'h530d57e7;
    ram_cell[    6697] = 32'h0;  // 32'h9a20ddc1;
    ram_cell[    6698] = 32'h0;  // 32'hf878967f;
    ram_cell[    6699] = 32'h0;  // 32'hbfa2e447;
    ram_cell[    6700] = 32'h0;  // 32'h9a51e17e;
    ram_cell[    6701] = 32'h0;  // 32'h75c63c4c;
    ram_cell[    6702] = 32'h0;  // 32'h5284c3c4;
    ram_cell[    6703] = 32'h0;  // 32'h52b73b0e;
    ram_cell[    6704] = 32'h0;  // 32'h4ca2c182;
    ram_cell[    6705] = 32'h0;  // 32'hc1b258b5;
    ram_cell[    6706] = 32'h0;  // 32'h7903bdbd;
    ram_cell[    6707] = 32'h0;  // 32'h0cbf0f3f;
    ram_cell[    6708] = 32'h0;  // 32'hf708981a;
    ram_cell[    6709] = 32'h0;  // 32'h893f56b5;
    ram_cell[    6710] = 32'h0;  // 32'h8951863e;
    ram_cell[    6711] = 32'h0;  // 32'hf7cfd486;
    ram_cell[    6712] = 32'h0;  // 32'h2f08bbfe;
    ram_cell[    6713] = 32'h0;  // 32'h76995a46;
    ram_cell[    6714] = 32'h0;  // 32'h68b3c556;
    ram_cell[    6715] = 32'h0;  // 32'h54279dc1;
    ram_cell[    6716] = 32'h0;  // 32'h403d8cf2;
    ram_cell[    6717] = 32'h0;  // 32'hd1fdee7e;
    ram_cell[    6718] = 32'h0;  // 32'h157ab613;
    ram_cell[    6719] = 32'h0;  // 32'h28f234cc;
    ram_cell[    6720] = 32'h0;  // 32'hcb77c6b9;
    ram_cell[    6721] = 32'h0;  // 32'hc7f1fb69;
    ram_cell[    6722] = 32'h0;  // 32'haa2582ee;
    ram_cell[    6723] = 32'h0;  // 32'h91495c08;
    ram_cell[    6724] = 32'h0;  // 32'hab50d741;
    ram_cell[    6725] = 32'h0;  // 32'h7b36fafb;
    ram_cell[    6726] = 32'h0;  // 32'h0b1cb874;
    ram_cell[    6727] = 32'h0;  // 32'hdca7640b;
    ram_cell[    6728] = 32'h0;  // 32'hfd88167e;
    ram_cell[    6729] = 32'h0;  // 32'h7c572718;
    ram_cell[    6730] = 32'h0;  // 32'h2a761637;
    ram_cell[    6731] = 32'h0;  // 32'h88c99c3a;
    ram_cell[    6732] = 32'h0;  // 32'ha032a3a1;
    ram_cell[    6733] = 32'h0;  // 32'hda759bc6;
    ram_cell[    6734] = 32'h0;  // 32'h05647fc0;
    ram_cell[    6735] = 32'h0;  // 32'h94705017;
    ram_cell[    6736] = 32'h0;  // 32'h8c4762ed;
    ram_cell[    6737] = 32'h0;  // 32'h930a2c16;
    ram_cell[    6738] = 32'h0;  // 32'hd47fe53e;
    ram_cell[    6739] = 32'h0;  // 32'h3e1359d3;
    ram_cell[    6740] = 32'h0;  // 32'hac6fb7b6;
    ram_cell[    6741] = 32'h0;  // 32'h441557e1;
    ram_cell[    6742] = 32'h0;  // 32'h5977f2ee;
    ram_cell[    6743] = 32'h0;  // 32'h43f1e6d3;
    ram_cell[    6744] = 32'h0;  // 32'h7ea1c212;
    ram_cell[    6745] = 32'h0;  // 32'h4151adbc;
    ram_cell[    6746] = 32'h0;  // 32'h58877668;
    ram_cell[    6747] = 32'h0;  // 32'hf845c699;
    ram_cell[    6748] = 32'h0;  // 32'h1ab940cf;
    ram_cell[    6749] = 32'h0;  // 32'h3c17c250;
    ram_cell[    6750] = 32'h0;  // 32'he694580b;
    ram_cell[    6751] = 32'h0;  // 32'haecaf84a;
    ram_cell[    6752] = 32'h0;  // 32'hdb826efe;
    ram_cell[    6753] = 32'h0;  // 32'h3fdf9d42;
    ram_cell[    6754] = 32'h0;  // 32'hc60b9a52;
    ram_cell[    6755] = 32'h0;  // 32'hf7547592;
    ram_cell[    6756] = 32'h0;  // 32'h991beedc;
    ram_cell[    6757] = 32'h0;  // 32'h1b214252;
    ram_cell[    6758] = 32'h0;  // 32'he6d18b0b;
    ram_cell[    6759] = 32'h0;  // 32'hea0dd55f;
    ram_cell[    6760] = 32'h0;  // 32'h7c139b31;
    ram_cell[    6761] = 32'h0;  // 32'ha4126d52;
    ram_cell[    6762] = 32'h0;  // 32'h267f9954;
    ram_cell[    6763] = 32'h0;  // 32'hcf2d39f9;
    ram_cell[    6764] = 32'h0;  // 32'h21fa556b;
    ram_cell[    6765] = 32'h0;  // 32'hc823f8a3;
    ram_cell[    6766] = 32'h0;  // 32'h39f61b1f;
    ram_cell[    6767] = 32'h0;  // 32'hcdf3ed7f;
    ram_cell[    6768] = 32'h0;  // 32'h964dfd43;
    ram_cell[    6769] = 32'h0;  // 32'h91b40745;
    ram_cell[    6770] = 32'h0;  // 32'h803cf073;
    ram_cell[    6771] = 32'h0;  // 32'h369fa80f;
    ram_cell[    6772] = 32'h0;  // 32'hc3aaa1bd;
    ram_cell[    6773] = 32'h0;  // 32'h81d7b667;
    ram_cell[    6774] = 32'h0;  // 32'hbff0a91e;
    ram_cell[    6775] = 32'h0;  // 32'h62010f5f;
    ram_cell[    6776] = 32'h0;  // 32'h3c09143b;
    ram_cell[    6777] = 32'h0;  // 32'hed85fb26;
    ram_cell[    6778] = 32'h0;  // 32'h520a0b84;
    ram_cell[    6779] = 32'h0;  // 32'h6333774d;
    ram_cell[    6780] = 32'h0;  // 32'hbb176bf0;
    ram_cell[    6781] = 32'h0;  // 32'h39ba7bac;
    ram_cell[    6782] = 32'h0;  // 32'hfffdd9ca;
    ram_cell[    6783] = 32'h0;  // 32'h6c8acdf3;
    ram_cell[    6784] = 32'h0;  // 32'h9a541fab;
    ram_cell[    6785] = 32'h0;  // 32'h9f69da95;
    ram_cell[    6786] = 32'h0;  // 32'hd3c8cec8;
    ram_cell[    6787] = 32'h0;  // 32'h9c83635a;
    ram_cell[    6788] = 32'h0;  // 32'hebbff47c;
    ram_cell[    6789] = 32'h0;  // 32'h700d7f82;
    ram_cell[    6790] = 32'h0;  // 32'hef45eb66;
    ram_cell[    6791] = 32'h0;  // 32'h2e3a4a62;
    ram_cell[    6792] = 32'h0;  // 32'ha6d6783e;
    ram_cell[    6793] = 32'h0;  // 32'h1f479b09;
    ram_cell[    6794] = 32'h0;  // 32'h2806eee6;
    ram_cell[    6795] = 32'h0;  // 32'hb905c83d;
    ram_cell[    6796] = 32'h0;  // 32'hf5c5a4fe;
    ram_cell[    6797] = 32'h0;  // 32'hdb816fa9;
    ram_cell[    6798] = 32'h0;  // 32'h6a768ed6;
    ram_cell[    6799] = 32'h0;  // 32'h812f36ef;
    ram_cell[    6800] = 32'h0;  // 32'hb51fd505;
    ram_cell[    6801] = 32'h0;  // 32'h3341cd1f;
    ram_cell[    6802] = 32'h0;  // 32'hbdbfed92;
    ram_cell[    6803] = 32'h0;  // 32'hbc5ae1fb;
    ram_cell[    6804] = 32'h0;  // 32'hdd04f7b3;
    ram_cell[    6805] = 32'h0;  // 32'h7d48f8cc;
    ram_cell[    6806] = 32'h0;  // 32'h07b91096;
    ram_cell[    6807] = 32'h0;  // 32'hcd46502d;
    ram_cell[    6808] = 32'h0;  // 32'h855a7b07;
    ram_cell[    6809] = 32'h0;  // 32'h0f1acfdc;
    ram_cell[    6810] = 32'h0;  // 32'h838ab509;
    ram_cell[    6811] = 32'h0;  // 32'h8985e77e;
    ram_cell[    6812] = 32'h0;  // 32'h6e8ae48d;
    ram_cell[    6813] = 32'h0;  // 32'h233bdbf1;
    ram_cell[    6814] = 32'h0;  // 32'hb3de994f;
    ram_cell[    6815] = 32'h0;  // 32'hbab39188;
    ram_cell[    6816] = 32'h0;  // 32'h938c2c05;
    ram_cell[    6817] = 32'h0;  // 32'h1e311f1a;
    ram_cell[    6818] = 32'h0;  // 32'h656c6f40;
    ram_cell[    6819] = 32'h0;  // 32'h614ea102;
    ram_cell[    6820] = 32'h0;  // 32'h4c4ace8c;
    ram_cell[    6821] = 32'h0;  // 32'hc10b5746;
    ram_cell[    6822] = 32'h0;  // 32'h05ea6499;
    ram_cell[    6823] = 32'h0;  // 32'haee971fc;
    ram_cell[    6824] = 32'h0;  // 32'hdb6f1a80;
    ram_cell[    6825] = 32'h0;  // 32'h6855b4f8;
    ram_cell[    6826] = 32'h0;  // 32'hfba27059;
    ram_cell[    6827] = 32'h0;  // 32'h7c633ad1;
    ram_cell[    6828] = 32'h0;  // 32'ha37a706d;
    ram_cell[    6829] = 32'h0;  // 32'h82987005;
    ram_cell[    6830] = 32'h0;  // 32'h6a5dfcda;
    ram_cell[    6831] = 32'h0;  // 32'h980e346a;
    ram_cell[    6832] = 32'h0;  // 32'hec046442;
    ram_cell[    6833] = 32'h0;  // 32'hde8a3f27;
    ram_cell[    6834] = 32'h0;  // 32'ha78cf30c;
    ram_cell[    6835] = 32'h0;  // 32'h9c2d4017;
    ram_cell[    6836] = 32'h0;  // 32'h3f7ca60d;
    ram_cell[    6837] = 32'h0;  // 32'h172c09fe;
    ram_cell[    6838] = 32'h0;  // 32'hdf73196d;
    ram_cell[    6839] = 32'h0;  // 32'hac36c986;
    ram_cell[    6840] = 32'h0;  // 32'h18b78545;
    ram_cell[    6841] = 32'h0;  // 32'hb3cb81d0;
    ram_cell[    6842] = 32'h0;  // 32'h7246f5e5;
    ram_cell[    6843] = 32'h0;  // 32'ha6afc004;
    ram_cell[    6844] = 32'h0;  // 32'h339df688;
    ram_cell[    6845] = 32'h0;  // 32'h39512d16;
    ram_cell[    6846] = 32'h0;  // 32'h978202ea;
    ram_cell[    6847] = 32'h0;  // 32'hf36787e3;
    ram_cell[    6848] = 32'h0;  // 32'hba064ecc;
    ram_cell[    6849] = 32'h0;  // 32'h4a7e100e;
    ram_cell[    6850] = 32'h0;  // 32'h5012d2f2;
    ram_cell[    6851] = 32'h0;  // 32'h8304f7bc;
    ram_cell[    6852] = 32'h0;  // 32'h7b540f67;
    ram_cell[    6853] = 32'h0;  // 32'h03fea4be;
    ram_cell[    6854] = 32'h0;  // 32'he136cc99;
    ram_cell[    6855] = 32'h0;  // 32'h0b3ce4fe;
    ram_cell[    6856] = 32'h0;  // 32'h9d0d7e63;
    ram_cell[    6857] = 32'h0;  // 32'h1165f163;
    ram_cell[    6858] = 32'h0;  // 32'h010c540e;
    ram_cell[    6859] = 32'h0;  // 32'h437a26bb;
    ram_cell[    6860] = 32'h0;  // 32'h6b01dad1;
    ram_cell[    6861] = 32'h0;  // 32'hb333bc64;
    ram_cell[    6862] = 32'h0;  // 32'h38bcfc5a;
    ram_cell[    6863] = 32'h0;  // 32'h656c9f50;
    ram_cell[    6864] = 32'h0;  // 32'h17593781;
    ram_cell[    6865] = 32'h0;  // 32'hf8bd1197;
    ram_cell[    6866] = 32'h0;  // 32'h3e9a6459;
    ram_cell[    6867] = 32'h0;  // 32'h5016880d;
    ram_cell[    6868] = 32'h0;  // 32'h6d19c667;
    ram_cell[    6869] = 32'h0;  // 32'h4c0efd0a;
    ram_cell[    6870] = 32'h0;  // 32'h04dde20f;
    ram_cell[    6871] = 32'h0;  // 32'hbede5634;
    ram_cell[    6872] = 32'h0;  // 32'h67df0c85;
    ram_cell[    6873] = 32'h0;  // 32'h312762f5;
    ram_cell[    6874] = 32'h0;  // 32'h192c5331;
    ram_cell[    6875] = 32'h0;  // 32'hb231178d;
    ram_cell[    6876] = 32'h0;  // 32'h0398f942;
    ram_cell[    6877] = 32'h0;  // 32'ha9c02a45;
    ram_cell[    6878] = 32'h0;  // 32'h8cf2f928;
    ram_cell[    6879] = 32'h0;  // 32'h32678de7;
    ram_cell[    6880] = 32'h0;  // 32'h0ec01e36;
    ram_cell[    6881] = 32'h0;  // 32'ha50476dc;
    ram_cell[    6882] = 32'h0;  // 32'h59006ffe;
    ram_cell[    6883] = 32'h0;  // 32'h4ed9b0da;
    ram_cell[    6884] = 32'h0;  // 32'h31ac85cc;
    ram_cell[    6885] = 32'h0;  // 32'h83bf946a;
    ram_cell[    6886] = 32'h0;  // 32'hc111299d;
    ram_cell[    6887] = 32'h0;  // 32'ha0031008;
    ram_cell[    6888] = 32'h0;  // 32'h77c89111;
    ram_cell[    6889] = 32'h0;  // 32'heb6535ff;
    ram_cell[    6890] = 32'h0;  // 32'hf71d46ca;
    ram_cell[    6891] = 32'h0;  // 32'h2f0fef94;
    ram_cell[    6892] = 32'h0;  // 32'h039522fc;
    ram_cell[    6893] = 32'h0;  // 32'h0ddd098a;
    ram_cell[    6894] = 32'h0;  // 32'h2ea05591;
    ram_cell[    6895] = 32'h0;  // 32'hd67e3210;
    ram_cell[    6896] = 32'h0;  // 32'h13215e3e;
    ram_cell[    6897] = 32'h0;  // 32'hffdcaca3;
    ram_cell[    6898] = 32'h0;  // 32'h3f608562;
    ram_cell[    6899] = 32'h0;  // 32'h65975185;
    ram_cell[    6900] = 32'h0;  // 32'h4b5a5881;
    ram_cell[    6901] = 32'h0;  // 32'hc7aa36b6;
    ram_cell[    6902] = 32'h0;  // 32'hdaeac0d3;
    ram_cell[    6903] = 32'h0;  // 32'h84177442;
    ram_cell[    6904] = 32'h0;  // 32'h5919c86e;
    ram_cell[    6905] = 32'h0;  // 32'h4fb5091b;
    ram_cell[    6906] = 32'h0;  // 32'h1a55afa2;
    ram_cell[    6907] = 32'h0;  // 32'h6a0c65b2;
    ram_cell[    6908] = 32'h0;  // 32'h997ce057;
    ram_cell[    6909] = 32'h0;  // 32'h12b17e16;
    ram_cell[    6910] = 32'h0;  // 32'hffe92f8c;
    ram_cell[    6911] = 32'h0;  // 32'hbb92d2a3;
    ram_cell[    6912] = 32'h0;  // 32'h504db258;
    ram_cell[    6913] = 32'h0;  // 32'he2a2a642;
    ram_cell[    6914] = 32'h0;  // 32'h7cfc7a4e;
    ram_cell[    6915] = 32'h0;  // 32'hd450a798;
    ram_cell[    6916] = 32'h0;  // 32'h46c76946;
    ram_cell[    6917] = 32'h0;  // 32'hb8f4e16b;
    ram_cell[    6918] = 32'h0;  // 32'hbe2ebbd8;
    ram_cell[    6919] = 32'h0;  // 32'h1a2372aa;
    ram_cell[    6920] = 32'h0;  // 32'he455a31e;
    ram_cell[    6921] = 32'h0;  // 32'hb6fca7f5;
    ram_cell[    6922] = 32'h0;  // 32'h344278e8;
    ram_cell[    6923] = 32'h0;  // 32'h35e4ea57;
    ram_cell[    6924] = 32'h0;  // 32'hc96b8cf6;
    ram_cell[    6925] = 32'h0;  // 32'h8ad4a04d;
    ram_cell[    6926] = 32'h0;  // 32'h05029858;
    ram_cell[    6927] = 32'h0;  // 32'h4b2a4425;
    ram_cell[    6928] = 32'h0;  // 32'h1786040b;
    ram_cell[    6929] = 32'h0;  // 32'hf93775e3;
    ram_cell[    6930] = 32'h0;  // 32'h9dc24dae;
    ram_cell[    6931] = 32'h0;  // 32'h1f1e74b7;
    ram_cell[    6932] = 32'h0;  // 32'h732885a5;
    ram_cell[    6933] = 32'h0;  // 32'ha7aee736;
    ram_cell[    6934] = 32'h0;  // 32'hf8128afb;
    ram_cell[    6935] = 32'h0;  // 32'he1bae87d;
    ram_cell[    6936] = 32'h0;  // 32'hcbf22f1d;
    ram_cell[    6937] = 32'h0;  // 32'h125d9a0f;
    ram_cell[    6938] = 32'h0;  // 32'h489d8bd2;
    ram_cell[    6939] = 32'h0;  // 32'h726717c9;
    ram_cell[    6940] = 32'h0;  // 32'h60fc74a3;
    ram_cell[    6941] = 32'h0;  // 32'h76f49d9f;
    ram_cell[    6942] = 32'h0;  // 32'h0e9e25e5;
    ram_cell[    6943] = 32'h0;  // 32'h6fc2da55;
    ram_cell[    6944] = 32'h0;  // 32'h37622a35;
    ram_cell[    6945] = 32'h0;  // 32'hb5558997;
    ram_cell[    6946] = 32'h0;  // 32'h41f18eff;
    ram_cell[    6947] = 32'h0;  // 32'h3d958788;
    ram_cell[    6948] = 32'h0;  // 32'h4cd3dfd9;
    ram_cell[    6949] = 32'h0;  // 32'h6329a060;
    ram_cell[    6950] = 32'h0;  // 32'hd63e2500;
    ram_cell[    6951] = 32'h0;  // 32'h497c8870;
    ram_cell[    6952] = 32'h0;  // 32'he1f1ff73;
    ram_cell[    6953] = 32'h0;  // 32'h60bed967;
    ram_cell[    6954] = 32'h0;  // 32'h62f3adb4;
    ram_cell[    6955] = 32'h0;  // 32'h5e33b7eb;
    ram_cell[    6956] = 32'h0;  // 32'hc9cc4a2c;
    ram_cell[    6957] = 32'h0;  // 32'ha17c8c0f;
    ram_cell[    6958] = 32'h0;  // 32'h04b141f0;
    ram_cell[    6959] = 32'h0;  // 32'hdbb5992d;
    ram_cell[    6960] = 32'h0;  // 32'h0e51e506;
    ram_cell[    6961] = 32'h0;  // 32'h9dd9e862;
    ram_cell[    6962] = 32'h0;  // 32'h7e31df24;
    ram_cell[    6963] = 32'h0;  // 32'h754a2fce;
    ram_cell[    6964] = 32'h0;  // 32'h564d2af1;
    ram_cell[    6965] = 32'h0;  // 32'h53a5327f;
    ram_cell[    6966] = 32'h0;  // 32'hc8628a73;
    ram_cell[    6967] = 32'h0;  // 32'h34e78520;
    ram_cell[    6968] = 32'h0;  // 32'h4f6497d3;
    ram_cell[    6969] = 32'h0;  // 32'hf8e5453a;
    ram_cell[    6970] = 32'h0;  // 32'h5bc2e54f;
    ram_cell[    6971] = 32'h0;  // 32'h0c177e0b;
    ram_cell[    6972] = 32'h0;  // 32'hf8e8b6e5;
    ram_cell[    6973] = 32'h0;  // 32'h3849da5c;
    ram_cell[    6974] = 32'h0;  // 32'h595fdc60;
    ram_cell[    6975] = 32'h0;  // 32'h6a78b38f;
    ram_cell[    6976] = 32'h0;  // 32'hbcfa0b94;
    ram_cell[    6977] = 32'h0;  // 32'hab8db786;
    ram_cell[    6978] = 32'h0;  // 32'h3d4fb903;
    ram_cell[    6979] = 32'h0;  // 32'hf66f348a;
    ram_cell[    6980] = 32'h0;  // 32'h65faa194;
    ram_cell[    6981] = 32'h0;  // 32'ha8fca5ce;
    ram_cell[    6982] = 32'h0;  // 32'h1a3d2591;
    ram_cell[    6983] = 32'h0;  // 32'h98f6e4ab;
    ram_cell[    6984] = 32'h0;  // 32'h207f9f2c;
    ram_cell[    6985] = 32'h0;  // 32'h4706bee8;
    ram_cell[    6986] = 32'h0;  // 32'h98dc9a2a;
    ram_cell[    6987] = 32'h0;  // 32'h9410d293;
    ram_cell[    6988] = 32'h0;  // 32'h83dd5b97;
    ram_cell[    6989] = 32'h0;  // 32'h00a0232c;
    ram_cell[    6990] = 32'h0;  // 32'h90b394d3;
    ram_cell[    6991] = 32'h0;  // 32'h406c9242;
    ram_cell[    6992] = 32'h0;  // 32'he7539f9e;
    ram_cell[    6993] = 32'h0;  // 32'h5eb7f64a;
    ram_cell[    6994] = 32'h0;  // 32'h3b9c8035;
    ram_cell[    6995] = 32'h0;  // 32'h4adb2706;
    ram_cell[    6996] = 32'h0;  // 32'h52998a08;
    ram_cell[    6997] = 32'h0;  // 32'h84ab2177;
    ram_cell[    6998] = 32'h0;  // 32'he898520f;
    ram_cell[    6999] = 32'h0;  // 32'he66360cb;
    ram_cell[    7000] = 32'h0;  // 32'h61956cd3;
    ram_cell[    7001] = 32'h0;  // 32'he449fb81;
    ram_cell[    7002] = 32'h0;  // 32'h1f687202;
    ram_cell[    7003] = 32'h0;  // 32'h4d828add;
    ram_cell[    7004] = 32'h0;  // 32'h142b28c7;
    ram_cell[    7005] = 32'h0;  // 32'hc62f4360;
    ram_cell[    7006] = 32'h0;  // 32'h2ee64e51;
    ram_cell[    7007] = 32'h0;  // 32'h1f2c7c11;
    ram_cell[    7008] = 32'h0;  // 32'hc98f7a9a;
    ram_cell[    7009] = 32'h0;  // 32'hfc4aa396;
    ram_cell[    7010] = 32'h0;  // 32'h8ae3addf;
    ram_cell[    7011] = 32'h0;  // 32'h21cf0621;
    ram_cell[    7012] = 32'h0;  // 32'hb7e733cb;
    ram_cell[    7013] = 32'h0;  // 32'hc596513f;
    ram_cell[    7014] = 32'h0;  // 32'h80d52ec9;
    ram_cell[    7015] = 32'h0;  // 32'h0fefc157;
    ram_cell[    7016] = 32'h0;  // 32'h349dda9e;
    ram_cell[    7017] = 32'h0;  // 32'hb040647a;
    ram_cell[    7018] = 32'h0;  // 32'hdbcf1e24;
    ram_cell[    7019] = 32'h0;  // 32'hdd304446;
    ram_cell[    7020] = 32'h0;  // 32'hf4f23faa;
    ram_cell[    7021] = 32'h0;  // 32'h7d7292ea;
    ram_cell[    7022] = 32'h0;  // 32'h750069c8;
    ram_cell[    7023] = 32'h0;  // 32'h2269e2cd;
    ram_cell[    7024] = 32'h0;  // 32'h03dea3aa;
    ram_cell[    7025] = 32'h0;  // 32'hb9fcdee9;
    ram_cell[    7026] = 32'h0;  // 32'h4b14d930;
    ram_cell[    7027] = 32'h0;  // 32'h6ba9e29e;
    ram_cell[    7028] = 32'h0;  // 32'hc850a475;
    ram_cell[    7029] = 32'h0;  // 32'haf45b8b3;
    ram_cell[    7030] = 32'h0;  // 32'h6dbeb1f0;
    ram_cell[    7031] = 32'h0;  // 32'h433e1601;
    ram_cell[    7032] = 32'h0;  // 32'h77718b9d;
    ram_cell[    7033] = 32'h0;  // 32'hbb6c51c5;
    ram_cell[    7034] = 32'h0;  // 32'h4fa78e5a;
    ram_cell[    7035] = 32'h0;  // 32'h1c3b3a7f;
    ram_cell[    7036] = 32'h0;  // 32'h8ed81526;
    ram_cell[    7037] = 32'h0;  // 32'h7cda5c4f;
    ram_cell[    7038] = 32'h0;  // 32'h676e821f;
    ram_cell[    7039] = 32'h0;  // 32'h7f518de8;
    ram_cell[    7040] = 32'h0;  // 32'h4616d7eb;
    ram_cell[    7041] = 32'h0;  // 32'h4c37c732;
    ram_cell[    7042] = 32'h0;  // 32'hf0af92a2;
    ram_cell[    7043] = 32'h0;  // 32'h3b71c949;
    ram_cell[    7044] = 32'h0;  // 32'h8f0c38e7;
    ram_cell[    7045] = 32'h0;  // 32'h021b776f;
    ram_cell[    7046] = 32'h0;  // 32'h883d27a5;
    ram_cell[    7047] = 32'h0;  // 32'h3e7a85d2;
    ram_cell[    7048] = 32'h0;  // 32'hee95bed8;
    ram_cell[    7049] = 32'h0;  // 32'h8ba1dbcf;
    ram_cell[    7050] = 32'h0;  // 32'h2a8e5e79;
    ram_cell[    7051] = 32'h0;  // 32'h26149f8a;
    ram_cell[    7052] = 32'h0;  // 32'h28c32391;
    ram_cell[    7053] = 32'h0;  // 32'h51e04997;
    ram_cell[    7054] = 32'h0;  // 32'h1ef7bb67;
    ram_cell[    7055] = 32'h0;  // 32'h8e63f117;
    ram_cell[    7056] = 32'h0;  // 32'h5c7883f7;
    ram_cell[    7057] = 32'h0;  // 32'h111f1471;
    ram_cell[    7058] = 32'h0;  // 32'hf3f5bb74;
    ram_cell[    7059] = 32'h0;  // 32'h1c78c239;
    ram_cell[    7060] = 32'h0;  // 32'hc3e45862;
    ram_cell[    7061] = 32'h0;  // 32'h8edb871c;
    ram_cell[    7062] = 32'h0;  // 32'h54ea2902;
    ram_cell[    7063] = 32'h0;  // 32'he6515bf5;
    ram_cell[    7064] = 32'h0;  // 32'hb8e224db;
    ram_cell[    7065] = 32'h0;  // 32'ha7c36cd8;
    ram_cell[    7066] = 32'h0;  // 32'h7cca2fcc;
    ram_cell[    7067] = 32'h0;  // 32'h37434acf;
    ram_cell[    7068] = 32'h0;  // 32'h23fdb09f;
    ram_cell[    7069] = 32'h0;  // 32'he3c79958;
    ram_cell[    7070] = 32'h0;  // 32'h81b0070b;
    ram_cell[    7071] = 32'h0;  // 32'hf30a7374;
    ram_cell[    7072] = 32'h0;  // 32'h8e935cb5;
    ram_cell[    7073] = 32'h0;  // 32'h204d9647;
    ram_cell[    7074] = 32'h0;  // 32'h05be9aa7;
    ram_cell[    7075] = 32'h0;  // 32'h3dd95a66;
    ram_cell[    7076] = 32'h0;  // 32'h2b80298f;
    ram_cell[    7077] = 32'h0;  // 32'hc1b99dcb;
    ram_cell[    7078] = 32'h0;  // 32'h7cd970df;
    ram_cell[    7079] = 32'h0;  // 32'h2704ce9d;
    ram_cell[    7080] = 32'h0;  // 32'hc0cd8830;
    ram_cell[    7081] = 32'h0;  // 32'hf367d36b;
    ram_cell[    7082] = 32'h0;  // 32'h7ea28961;
    ram_cell[    7083] = 32'h0;  // 32'hd57fefd6;
    ram_cell[    7084] = 32'h0;  // 32'hb77bbc3f;
    ram_cell[    7085] = 32'h0;  // 32'h9cfef039;
    ram_cell[    7086] = 32'h0;  // 32'h35e129f9;
    ram_cell[    7087] = 32'h0;  // 32'h9a64403f;
    ram_cell[    7088] = 32'h0;  // 32'hfd1e6c95;
    ram_cell[    7089] = 32'h0;  // 32'h747c3a9f;
    ram_cell[    7090] = 32'h0;  // 32'h67c2e157;
    ram_cell[    7091] = 32'h0;  // 32'h2fc56ae5;
    ram_cell[    7092] = 32'h0;  // 32'h280feb97;
    ram_cell[    7093] = 32'h0;  // 32'h95b471a4;
    ram_cell[    7094] = 32'h0;  // 32'h0b0733dc;
    ram_cell[    7095] = 32'h0;  // 32'h07d4a5c5;
    ram_cell[    7096] = 32'h0;  // 32'hfc60bbea;
    ram_cell[    7097] = 32'h0;  // 32'hdb476350;
    ram_cell[    7098] = 32'h0;  // 32'ha658d12b;
    ram_cell[    7099] = 32'h0;  // 32'h3f98d6df;
    ram_cell[    7100] = 32'h0;  // 32'h603ff75c;
    ram_cell[    7101] = 32'h0;  // 32'h465ad9f3;
    ram_cell[    7102] = 32'h0;  // 32'h5c9b9dab;
    ram_cell[    7103] = 32'h0;  // 32'h8bc4ed31;
    ram_cell[    7104] = 32'h0;  // 32'h5d7ac0db;
    ram_cell[    7105] = 32'h0;  // 32'h3aa413f7;
    ram_cell[    7106] = 32'h0;  // 32'h9cf7e5aa;
    ram_cell[    7107] = 32'h0;  // 32'hb6efcb7d;
    ram_cell[    7108] = 32'h0;  // 32'h0386f0ae;
    ram_cell[    7109] = 32'h0;  // 32'h58daa41e;
    ram_cell[    7110] = 32'h0;  // 32'h35b8f095;
    ram_cell[    7111] = 32'h0;  // 32'h44081e9d;
    ram_cell[    7112] = 32'h0;  // 32'h09221c7c;
    ram_cell[    7113] = 32'h0;  // 32'h317e0ef9;
    ram_cell[    7114] = 32'h0;  // 32'hca4a5a9f;
    ram_cell[    7115] = 32'h0;  // 32'h56f40b49;
    ram_cell[    7116] = 32'h0;  // 32'h3275bfc4;
    ram_cell[    7117] = 32'h0;  // 32'h04653bac;
    ram_cell[    7118] = 32'h0;  // 32'heff6fa95;
    ram_cell[    7119] = 32'h0;  // 32'h82d7dc69;
    ram_cell[    7120] = 32'h0;  // 32'hc4d58d70;
    ram_cell[    7121] = 32'h0;  // 32'h36b8ac79;
    ram_cell[    7122] = 32'h0;  // 32'h74e54f33;
    ram_cell[    7123] = 32'h0;  // 32'hc69697d1;
    ram_cell[    7124] = 32'h0;  // 32'hf0266cc5;
    ram_cell[    7125] = 32'h0;  // 32'hbb4958b3;
    ram_cell[    7126] = 32'h0;  // 32'hccc3ac44;
    ram_cell[    7127] = 32'h0;  // 32'h1946a7a0;
    ram_cell[    7128] = 32'h0;  // 32'hc4419c3e;
    ram_cell[    7129] = 32'h0;  // 32'hf9bbf1c1;
    ram_cell[    7130] = 32'h0;  // 32'hb1043a22;
    ram_cell[    7131] = 32'h0;  // 32'h8705d040;
    ram_cell[    7132] = 32'h0;  // 32'h87961546;
    ram_cell[    7133] = 32'h0;  // 32'h353d77ce;
    ram_cell[    7134] = 32'h0;  // 32'h192e2861;
    ram_cell[    7135] = 32'h0;  // 32'h38f378cb;
    ram_cell[    7136] = 32'h0;  // 32'hd076609b;
    ram_cell[    7137] = 32'h0;  // 32'h49d0fb15;
    ram_cell[    7138] = 32'h0;  // 32'h028ba419;
    ram_cell[    7139] = 32'h0;  // 32'hbc1e17af;
    ram_cell[    7140] = 32'h0;  // 32'hecd4a725;
    ram_cell[    7141] = 32'h0;  // 32'hecba5924;
    ram_cell[    7142] = 32'h0;  // 32'h97a85413;
    ram_cell[    7143] = 32'h0;  // 32'hb271ba8f;
    ram_cell[    7144] = 32'h0;  // 32'h549256d0;
    ram_cell[    7145] = 32'h0;  // 32'h7d777a62;
    ram_cell[    7146] = 32'h0;  // 32'hcd8142e4;
    ram_cell[    7147] = 32'h0;  // 32'hf6e05dea;
    ram_cell[    7148] = 32'h0;  // 32'h76de1a18;
    ram_cell[    7149] = 32'h0;  // 32'he055a662;
    ram_cell[    7150] = 32'h0;  // 32'h0e275bab;
    ram_cell[    7151] = 32'h0;  // 32'hc064eab4;
    ram_cell[    7152] = 32'h0;  // 32'ha6f2787e;
    ram_cell[    7153] = 32'h0;  // 32'h89be72de;
    ram_cell[    7154] = 32'h0;  // 32'h6d353fae;
    ram_cell[    7155] = 32'h0;  // 32'h346d0be2;
    ram_cell[    7156] = 32'h0;  // 32'h9e839c15;
    ram_cell[    7157] = 32'h0;  // 32'hb9670822;
    ram_cell[    7158] = 32'h0;  // 32'h31f7c727;
    ram_cell[    7159] = 32'h0;  // 32'h7a7b48e7;
    ram_cell[    7160] = 32'h0;  // 32'h7fd314c2;
    ram_cell[    7161] = 32'h0;  // 32'hfe2917e9;
    ram_cell[    7162] = 32'h0;  // 32'ha91176af;
    ram_cell[    7163] = 32'h0;  // 32'h8d181fbb;
    ram_cell[    7164] = 32'h0;  // 32'h79919cf8;
    ram_cell[    7165] = 32'h0;  // 32'h5b297580;
    ram_cell[    7166] = 32'h0;  // 32'h9de463c0;
    ram_cell[    7167] = 32'h0;  // 32'h63140c72;
    ram_cell[    7168] = 32'h0;  // 32'h31d7cb0d;
    ram_cell[    7169] = 32'h0;  // 32'hfbe5fd63;
    ram_cell[    7170] = 32'h0;  // 32'h27470159;
    ram_cell[    7171] = 32'h0;  // 32'h3923e659;
    ram_cell[    7172] = 32'h0;  // 32'hcbce29c1;
    ram_cell[    7173] = 32'h0;  // 32'hcd50e37d;
    ram_cell[    7174] = 32'h0;  // 32'h15730045;
    ram_cell[    7175] = 32'h0;  // 32'hdbcb35bf;
    ram_cell[    7176] = 32'h0;  // 32'h1854523e;
    ram_cell[    7177] = 32'h0;  // 32'hda44008f;
    ram_cell[    7178] = 32'h0;  // 32'h163aa22a;
    ram_cell[    7179] = 32'h0;  // 32'h78115368;
    ram_cell[    7180] = 32'h0;  // 32'h6bc073a3;
    ram_cell[    7181] = 32'h0;  // 32'hd96ad21c;
    ram_cell[    7182] = 32'h0;  // 32'h6f8d53cf;
    ram_cell[    7183] = 32'h0;  // 32'h68f065c8;
    ram_cell[    7184] = 32'h0;  // 32'h951a332d;
    ram_cell[    7185] = 32'h0;  // 32'he1a917e4;
    ram_cell[    7186] = 32'h0;  // 32'he608da33;
    ram_cell[    7187] = 32'h0;  // 32'h086c86ee;
    ram_cell[    7188] = 32'h0;  // 32'h8ae50945;
    ram_cell[    7189] = 32'h0;  // 32'h6f6c45d7;
    ram_cell[    7190] = 32'h0;  // 32'h40d16cab;
    ram_cell[    7191] = 32'h0;  // 32'h2fef0668;
    ram_cell[    7192] = 32'h0;  // 32'h914127e1;
    ram_cell[    7193] = 32'h0;  // 32'hc737bb11;
    ram_cell[    7194] = 32'h0;  // 32'h6501c103;
    ram_cell[    7195] = 32'h0;  // 32'h653a3a92;
    ram_cell[    7196] = 32'h0;  // 32'hf4b3a2e1;
    ram_cell[    7197] = 32'h0;  // 32'h57d7a55a;
    ram_cell[    7198] = 32'h0;  // 32'hfb30d8a7;
    ram_cell[    7199] = 32'h0;  // 32'hac245dd1;
    ram_cell[    7200] = 32'h0;  // 32'hfd4215ed;
    ram_cell[    7201] = 32'h0;  // 32'h7a931035;
    ram_cell[    7202] = 32'h0;  // 32'h68774893;
    ram_cell[    7203] = 32'h0;  // 32'h24db5d0e;
    ram_cell[    7204] = 32'h0;  // 32'h374661c1;
    ram_cell[    7205] = 32'h0;  // 32'hcab90907;
    ram_cell[    7206] = 32'h0;  // 32'h8e4374b3;
    ram_cell[    7207] = 32'h0;  // 32'ha250c397;
    ram_cell[    7208] = 32'h0;  // 32'h354b8f04;
    ram_cell[    7209] = 32'h0;  // 32'h3ae09b7b;
    ram_cell[    7210] = 32'h0;  // 32'h02ace6cb;
    ram_cell[    7211] = 32'h0;  // 32'h08bf8d32;
    ram_cell[    7212] = 32'h0;  // 32'h4a0b9b48;
    ram_cell[    7213] = 32'h0;  // 32'h8e1f23f2;
    ram_cell[    7214] = 32'h0;  // 32'he5fc7287;
    ram_cell[    7215] = 32'h0;  // 32'h0e2018ec;
    ram_cell[    7216] = 32'h0;  // 32'h8216a756;
    ram_cell[    7217] = 32'h0;  // 32'hbd5f8e4b;
    ram_cell[    7218] = 32'h0;  // 32'h3cfadeee;
    ram_cell[    7219] = 32'h0;  // 32'h1dbb824e;
    ram_cell[    7220] = 32'h0;  // 32'h67582c55;
    ram_cell[    7221] = 32'h0;  // 32'h3f9ac0df;
    ram_cell[    7222] = 32'h0;  // 32'hf7ce66c9;
    ram_cell[    7223] = 32'h0;  // 32'h1ffd01f7;
    ram_cell[    7224] = 32'h0;  // 32'h9d298943;
    ram_cell[    7225] = 32'h0;  // 32'hb9af00d6;
    ram_cell[    7226] = 32'h0;  // 32'h4166526c;
    ram_cell[    7227] = 32'h0;  // 32'h7f5b91cd;
    ram_cell[    7228] = 32'h0;  // 32'ha8d12539;
    ram_cell[    7229] = 32'h0;  // 32'h0083e8ad;
    ram_cell[    7230] = 32'h0;  // 32'h2252ae81;
    ram_cell[    7231] = 32'h0;  // 32'h857d15a9;
    ram_cell[    7232] = 32'h0;  // 32'h6424fd6e;
    ram_cell[    7233] = 32'h0;  // 32'h51fd3a7c;
    ram_cell[    7234] = 32'h0;  // 32'hc58091ef;
    ram_cell[    7235] = 32'h0;  // 32'h4f2046f4;
    ram_cell[    7236] = 32'h0;  // 32'h8672c428;
    ram_cell[    7237] = 32'h0;  // 32'h7c415ff5;
    ram_cell[    7238] = 32'h0;  // 32'h2aa6cbde;
    ram_cell[    7239] = 32'h0;  // 32'hdb4c6657;
    ram_cell[    7240] = 32'h0;  // 32'he7297fce;
    ram_cell[    7241] = 32'h0;  // 32'hbdba0f5f;
    ram_cell[    7242] = 32'h0;  // 32'h847171c1;
    ram_cell[    7243] = 32'h0;  // 32'h2b59b157;
    ram_cell[    7244] = 32'h0;  // 32'h1b7b4042;
    ram_cell[    7245] = 32'h0;  // 32'h3305c140;
    ram_cell[    7246] = 32'h0;  // 32'h393052e7;
    ram_cell[    7247] = 32'h0;  // 32'h939e0801;
    ram_cell[    7248] = 32'h0;  // 32'haf550796;
    ram_cell[    7249] = 32'h0;  // 32'hf1e6afda;
    ram_cell[    7250] = 32'h0;  // 32'h65b5645a;
    ram_cell[    7251] = 32'h0;  // 32'h66faabbe;
    ram_cell[    7252] = 32'h0;  // 32'h4fe97ffa;
    ram_cell[    7253] = 32'h0;  // 32'h97774d1f;
    ram_cell[    7254] = 32'h0;  // 32'hd45e76fc;
    ram_cell[    7255] = 32'h0;  // 32'h3bb5ec88;
    ram_cell[    7256] = 32'h0;  // 32'h33c1214d;
    ram_cell[    7257] = 32'h0;  // 32'hca14042f;
    ram_cell[    7258] = 32'h0;  // 32'h0bc2b911;
    ram_cell[    7259] = 32'h0;  // 32'h047992c3;
    ram_cell[    7260] = 32'h0;  // 32'hde9f4e47;
    ram_cell[    7261] = 32'h0;  // 32'hb41cd89c;
    ram_cell[    7262] = 32'h0;  // 32'h8e2fb439;
    ram_cell[    7263] = 32'h0;  // 32'h93991bd0;
    ram_cell[    7264] = 32'h0;  // 32'h3fc81cc2;
    ram_cell[    7265] = 32'h0;  // 32'hcf66c988;
    ram_cell[    7266] = 32'h0;  // 32'h0cd8b4ec;
    ram_cell[    7267] = 32'h0;  // 32'h96949dfc;
    ram_cell[    7268] = 32'h0;  // 32'h67469e66;
    ram_cell[    7269] = 32'h0;  // 32'h55fe89f7;
    ram_cell[    7270] = 32'h0;  // 32'he61f6218;
    ram_cell[    7271] = 32'h0;  // 32'he9db86ee;
    ram_cell[    7272] = 32'h0;  // 32'h04cd615c;
    ram_cell[    7273] = 32'h0;  // 32'h5dc5df16;
    ram_cell[    7274] = 32'h0;  // 32'h200a6e5a;
    ram_cell[    7275] = 32'h0;  // 32'h8f73ab96;
    ram_cell[    7276] = 32'h0;  // 32'h7f7b3273;
    ram_cell[    7277] = 32'h0;  // 32'hd84ae627;
    ram_cell[    7278] = 32'h0;  // 32'h9dc72c90;
    ram_cell[    7279] = 32'h0;  // 32'h5780dc18;
    ram_cell[    7280] = 32'h0;  // 32'h0b2c54d3;
    ram_cell[    7281] = 32'h0;  // 32'h192deff0;
    ram_cell[    7282] = 32'h0;  // 32'hb431e0cc;
    ram_cell[    7283] = 32'h0;  // 32'hfe2a5920;
    ram_cell[    7284] = 32'h0;  // 32'hce17a73b;
    ram_cell[    7285] = 32'h0;  // 32'hfa544e46;
    ram_cell[    7286] = 32'h0;  // 32'h76373009;
    ram_cell[    7287] = 32'h0;  // 32'hd27f2bb9;
    ram_cell[    7288] = 32'h0;  // 32'h35e7d54b;
    ram_cell[    7289] = 32'h0;  // 32'h5922adce;
    ram_cell[    7290] = 32'h0;  // 32'h22fbd7c5;
    ram_cell[    7291] = 32'h0;  // 32'h74eae21a;
    ram_cell[    7292] = 32'h0;  // 32'hb90d61c6;
    ram_cell[    7293] = 32'h0;  // 32'h4487d0b0;
    ram_cell[    7294] = 32'h0;  // 32'h96276fa4;
    ram_cell[    7295] = 32'h0;  // 32'ha0f78e64;
    ram_cell[    7296] = 32'h0;  // 32'h5f4e7bac;
    ram_cell[    7297] = 32'h0;  // 32'h73e4bf8d;
    ram_cell[    7298] = 32'h0;  // 32'h7e1f0535;
    ram_cell[    7299] = 32'h0;  // 32'h8ffbb813;
    ram_cell[    7300] = 32'h0;  // 32'hc4d346b9;
    ram_cell[    7301] = 32'h0;  // 32'h3f2b7bc4;
    ram_cell[    7302] = 32'h0;  // 32'hfe82c587;
    ram_cell[    7303] = 32'h0;  // 32'h63567053;
    ram_cell[    7304] = 32'h0;  // 32'hbd65f357;
    ram_cell[    7305] = 32'h0;  // 32'h8b7b55e6;
    ram_cell[    7306] = 32'h0;  // 32'hef181fb3;
    ram_cell[    7307] = 32'h0;  // 32'h4b70c99e;
    ram_cell[    7308] = 32'h0;  // 32'hee132a42;
    ram_cell[    7309] = 32'h0;  // 32'h4679042c;
    ram_cell[    7310] = 32'h0;  // 32'h98ba0479;
    ram_cell[    7311] = 32'h0;  // 32'h7760ed6d;
    ram_cell[    7312] = 32'h0;  // 32'h547647fa;
    ram_cell[    7313] = 32'h0;  // 32'hb0fc7aa5;
    ram_cell[    7314] = 32'h0;  // 32'h56d0b9b9;
    ram_cell[    7315] = 32'h0;  // 32'h8ea025ee;
    ram_cell[    7316] = 32'h0;  // 32'h726f6e16;
    ram_cell[    7317] = 32'h0;  // 32'hd1fbbac0;
    ram_cell[    7318] = 32'h0;  // 32'hecb34bbe;
    ram_cell[    7319] = 32'h0;  // 32'h4e0f9827;
    ram_cell[    7320] = 32'h0;  // 32'hee847f8e;
    ram_cell[    7321] = 32'h0;  // 32'hd07411ad;
    ram_cell[    7322] = 32'h0;  // 32'h47260955;
    ram_cell[    7323] = 32'h0;  // 32'h1639350b;
    ram_cell[    7324] = 32'h0;  // 32'hca71a670;
    ram_cell[    7325] = 32'h0;  // 32'h17ece560;
    ram_cell[    7326] = 32'h0;  // 32'hc25e6824;
    ram_cell[    7327] = 32'h0;  // 32'ha00f6bb8;
    ram_cell[    7328] = 32'h0;  // 32'hb732a962;
    ram_cell[    7329] = 32'h0;  // 32'h458a97db;
    ram_cell[    7330] = 32'h0;  // 32'h0d1ad891;
    ram_cell[    7331] = 32'h0;  // 32'h133d8d70;
    ram_cell[    7332] = 32'h0;  // 32'h717d3548;
    ram_cell[    7333] = 32'h0;  // 32'h51e05b6d;
    ram_cell[    7334] = 32'h0;  // 32'h944fa33c;
    ram_cell[    7335] = 32'h0;  // 32'h52cc0ee3;
    ram_cell[    7336] = 32'h0;  // 32'hf565c630;
    ram_cell[    7337] = 32'h0;  // 32'h9d61ebf6;
    ram_cell[    7338] = 32'h0;  // 32'h0f321e22;
    ram_cell[    7339] = 32'h0;  // 32'hfb6184f6;
    ram_cell[    7340] = 32'h0;  // 32'he19f7ab7;
    ram_cell[    7341] = 32'h0;  // 32'hc4cbb9da;
    ram_cell[    7342] = 32'h0;  // 32'hdaf3a7d1;
    ram_cell[    7343] = 32'h0;  // 32'h5ce4749e;
    ram_cell[    7344] = 32'h0;  // 32'ha29b3e99;
    ram_cell[    7345] = 32'h0;  // 32'he8058cc1;
    ram_cell[    7346] = 32'h0;  // 32'h541605b0;
    ram_cell[    7347] = 32'h0;  // 32'hfbb23460;
    ram_cell[    7348] = 32'h0;  // 32'hb4cb0d0c;
    ram_cell[    7349] = 32'h0;  // 32'h43981d3b;
    ram_cell[    7350] = 32'h0;  // 32'hfaf84cf0;
    ram_cell[    7351] = 32'h0;  // 32'he9cdab55;
    ram_cell[    7352] = 32'h0;  // 32'h7d9d3afe;
    ram_cell[    7353] = 32'h0;  // 32'h2c20bfd3;
    ram_cell[    7354] = 32'h0;  // 32'h3bd69de2;
    ram_cell[    7355] = 32'h0;  // 32'hf7cb56de;
    ram_cell[    7356] = 32'h0;  // 32'hc5266f81;
    ram_cell[    7357] = 32'h0;  // 32'h28938ed0;
    ram_cell[    7358] = 32'h0;  // 32'h634f70d0;
    ram_cell[    7359] = 32'h0;  // 32'h1f518d5b;
    ram_cell[    7360] = 32'h0;  // 32'hd4e7b078;
    ram_cell[    7361] = 32'h0;  // 32'h9950a41a;
    ram_cell[    7362] = 32'h0;  // 32'h592eacc4;
    ram_cell[    7363] = 32'h0;  // 32'h71e27753;
    ram_cell[    7364] = 32'h0;  // 32'h583237a4;
    ram_cell[    7365] = 32'h0;  // 32'h1ccf2ca0;
    ram_cell[    7366] = 32'h0;  // 32'h2e4565b6;
    ram_cell[    7367] = 32'h0;  // 32'h1ad9b22d;
    ram_cell[    7368] = 32'h0;  // 32'hfcc8c0a5;
    ram_cell[    7369] = 32'h0;  // 32'he5c5bce5;
    ram_cell[    7370] = 32'h0;  // 32'h637d97dc;
    ram_cell[    7371] = 32'h0;  // 32'h2964bfa5;
    ram_cell[    7372] = 32'h0;  // 32'h9e97c8ce;
    ram_cell[    7373] = 32'h0;  // 32'hf7899ce2;
    ram_cell[    7374] = 32'h0;  // 32'h733e1cd9;
    ram_cell[    7375] = 32'h0;  // 32'hd2be5dbb;
    ram_cell[    7376] = 32'h0;  // 32'h67a59920;
    ram_cell[    7377] = 32'h0;  // 32'h4c612f93;
    ram_cell[    7378] = 32'h0;  // 32'h61e387a6;
    ram_cell[    7379] = 32'h0;  // 32'h60425a57;
    ram_cell[    7380] = 32'h0;  // 32'h0a75b248;
    ram_cell[    7381] = 32'h0;  // 32'hc2b9b38d;
    ram_cell[    7382] = 32'h0;  // 32'ha94d9b7f;
    ram_cell[    7383] = 32'h0;  // 32'ha376aac4;
    ram_cell[    7384] = 32'h0;  // 32'h1dbbb90a;
    ram_cell[    7385] = 32'h0;  // 32'h2873fde1;
    ram_cell[    7386] = 32'h0;  // 32'h2cc48bc6;
    ram_cell[    7387] = 32'h0;  // 32'hc08229b3;
    ram_cell[    7388] = 32'h0;  // 32'h00145085;
    ram_cell[    7389] = 32'h0;  // 32'h353f7aa3;
    ram_cell[    7390] = 32'h0;  // 32'hae6ebba6;
    ram_cell[    7391] = 32'h0;  // 32'ha6d84324;
    ram_cell[    7392] = 32'h0;  // 32'habd843d9;
    ram_cell[    7393] = 32'h0;  // 32'h9fb044ea;
    ram_cell[    7394] = 32'h0;  // 32'h46a98822;
    ram_cell[    7395] = 32'h0;  // 32'hd0a9ef9b;
    ram_cell[    7396] = 32'h0;  // 32'h675af916;
    ram_cell[    7397] = 32'h0;  // 32'h72c8dd71;
    ram_cell[    7398] = 32'h0;  // 32'h5b41a133;
    ram_cell[    7399] = 32'h0;  // 32'hfcbf7877;
    ram_cell[    7400] = 32'h0;  // 32'h3bc79fa6;
    ram_cell[    7401] = 32'h0;  // 32'h3ca3c1bd;
    ram_cell[    7402] = 32'h0;  // 32'h9cf3e5bb;
    ram_cell[    7403] = 32'h0;  // 32'h3b28afe4;
    ram_cell[    7404] = 32'h0;  // 32'h05e05860;
    ram_cell[    7405] = 32'h0;  // 32'h478e9c2f;
    ram_cell[    7406] = 32'h0;  // 32'h8652ecb4;
    ram_cell[    7407] = 32'h0;  // 32'h58706cd1;
    ram_cell[    7408] = 32'h0;  // 32'h670f9f5f;
    ram_cell[    7409] = 32'h0;  // 32'h242b1ba9;
    ram_cell[    7410] = 32'h0;  // 32'h902cbbc5;
    ram_cell[    7411] = 32'h0;  // 32'h1347eb23;
    ram_cell[    7412] = 32'h0;  // 32'hb14de9da;
    ram_cell[    7413] = 32'h0;  // 32'h3881f722;
    ram_cell[    7414] = 32'h0;  // 32'h34774eff;
    ram_cell[    7415] = 32'h0;  // 32'hd2d64fb1;
    ram_cell[    7416] = 32'h0;  // 32'hf326edcd;
    ram_cell[    7417] = 32'h0;  // 32'h31d76570;
    ram_cell[    7418] = 32'h0;  // 32'ha3dbc919;
    ram_cell[    7419] = 32'h0;  // 32'h818f1028;
    ram_cell[    7420] = 32'h0;  // 32'hc8ca7fe1;
    ram_cell[    7421] = 32'h0;  // 32'h26e27dac;
    ram_cell[    7422] = 32'h0;  // 32'h77d928da;
    ram_cell[    7423] = 32'h0;  // 32'ha7debbb7;
    ram_cell[    7424] = 32'h0;  // 32'h63d2890c;
    ram_cell[    7425] = 32'h0;  // 32'h6bd7ec75;
    ram_cell[    7426] = 32'h0;  // 32'haf842f54;
    ram_cell[    7427] = 32'h0;  // 32'he39d3875;
    ram_cell[    7428] = 32'h0;  // 32'hd2b01000;
    ram_cell[    7429] = 32'h0;  // 32'h2dc62b06;
    ram_cell[    7430] = 32'h0;  // 32'he47fbfd0;
    ram_cell[    7431] = 32'h0;  // 32'hcc005a34;
    ram_cell[    7432] = 32'h0;  // 32'h7c72718b;
    ram_cell[    7433] = 32'h0;  // 32'h53961738;
    ram_cell[    7434] = 32'h0;  // 32'h696f186f;
    ram_cell[    7435] = 32'h0;  // 32'hc1b83579;
    ram_cell[    7436] = 32'h0;  // 32'hed7d7f86;
    ram_cell[    7437] = 32'h0;  // 32'h1905b974;
    ram_cell[    7438] = 32'h0;  // 32'heebd2638;
    ram_cell[    7439] = 32'h0;  // 32'hb9feaaed;
    ram_cell[    7440] = 32'h0;  // 32'h6b515abc;
    ram_cell[    7441] = 32'h0;  // 32'h43629a8a;
    ram_cell[    7442] = 32'h0;  // 32'h3418b5f1;
    ram_cell[    7443] = 32'h0;  // 32'h527d63c8;
    ram_cell[    7444] = 32'h0;  // 32'h90e36499;
    ram_cell[    7445] = 32'h0;  // 32'hbcdc4f18;
    ram_cell[    7446] = 32'h0;  // 32'h4c6e8eca;
    ram_cell[    7447] = 32'h0;  // 32'h18a10593;
    ram_cell[    7448] = 32'h0;  // 32'hcb211e13;
    ram_cell[    7449] = 32'h0;  // 32'h7d811de1;
    ram_cell[    7450] = 32'h0;  // 32'hb3859587;
    ram_cell[    7451] = 32'h0;  // 32'hf3b45ba8;
    ram_cell[    7452] = 32'h0;  // 32'he114f16c;
    ram_cell[    7453] = 32'h0;  // 32'h123dd7c4;
    ram_cell[    7454] = 32'h0;  // 32'hf6746059;
    ram_cell[    7455] = 32'h0;  // 32'hd3604090;
    ram_cell[    7456] = 32'h0;  // 32'hccd14744;
    ram_cell[    7457] = 32'h0;  // 32'h93b5d38f;
    ram_cell[    7458] = 32'h0;  // 32'hca8ccce7;
    ram_cell[    7459] = 32'h0;  // 32'h6b46daaa;
    ram_cell[    7460] = 32'h0;  // 32'h6b3d6d6a;
    ram_cell[    7461] = 32'h0;  // 32'h3a0ac7e2;
    ram_cell[    7462] = 32'h0;  // 32'h26e9a89b;
    ram_cell[    7463] = 32'h0;  // 32'h8c530b30;
    ram_cell[    7464] = 32'h0;  // 32'hf0d64736;
    ram_cell[    7465] = 32'h0;  // 32'h89f6cec3;
    ram_cell[    7466] = 32'h0;  // 32'h38a1ce78;
    ram_cell[    7467] = 32'h0;  // 32'hcc7ce6eb;
    ram_cell[    7468] = 32'h0;  // 32'hf5db3262;
    ram_cell[    7469] = 32'h0;  // 32'hd39087e5;
    ram_cell[    7470] = 32'h0;  // 32'h475120e5;
    ram_cell[    7471] = 32'h0;  // 32'he7db732b;
    ram_cell[    7472] = 32'h0;  // 32'hb44a7792;
    ram_cell[    7473] = 32'h0;  // 32'hb5fb55e8;
    ram_cell[    7474] = 32'h0;  // 32'h9aa772f7;
    ram_cell[    7475] = 32'h0;  // 32'haebf1626;
    ram_cell[    7476] = 32'h0;  // 32'hd3529aa4;
    ram_cell[    7477] = 32'h0;  // 32'he8dea6dd;
    ram_cell[    7478] = 32'h0;  // 32'hf476ddd3;
    ram_cell[    7479] = 32'h0;  // 32'hd7869c9c;
    ram_cell[    7480] = 32'h0;  // 32'h3f9e6c5f;
    ram_cell[    7481] = 32'h0;  // 32'h55a3eb18;
    ram_cell[    7482] = 32'h0;  // 32'he9b89bbb;
    ram_cell[    7483] = 32'h0;  // 32'h43b94d5b;
    ram_cell[    7484] = 32'h0;  // 32'h95bd3bcd;
    ram_cell[    7485] = 32'h0;  // 32'h03b70026;
    ram_cell[    7486] = 32'h0;  // 32'h3d38c77e;
    ram_cell[    7487] = 32'h0;  // 32'h1f68ab22;
    ram_cell[    7488] = 32'h0;  // 32'h48872358;
    ram_cell[    7489] = 32'h0;  // 32'ha1c9597f;
    ram_cell[    7490] = 32'h0;  // 32'hcb9f3dd4;
    ram_cell[    7491] = 32'h0;  // 32'h1a614779;
    ram_cell[    7492] = 32'h0;  // 32'he40d7cca;
    ram_cell[    7493] = 32'h0;  // 32'ha7359244;
    ram_cell[    7494] = 32'h0;  // 32'hcbf97b9b;
    ram_cell[    7495] = 32'h0;  // 32'h72e7c703;
    ram_cell[    7496] = 32'h0;  // 32'h7d5c08ca;
    ram_cell[    7497] = 32'h0;  // 32'h49b2ba8d;
    ram_cell[    7498] = 32'h0;  // 32'h6b30d07e;
    ram_cell[    7499] = 32'h0;  // 32'h33f6d717;
    ram_cell[    7500] = 32'h0;  // 32'h840f21f6;
    ram_cell[    7501] = 32'h0;  // 32'hf1f2b069;
    ram_cell[    7502] = 32'h0;  // 32'h89237377;
    ram_cell[    7503] = 32'h0;  // 32'hdb8867f3;
    ram_cell[    7504] = 32'h0;  // 32'hb09f8682;
    ram_cell[    7505] = 32'h0;  // 32'h83f8849b;
    ram_cell[    7506] = 32'h0;  // 32'h4516fa6f;
    ram_cell[    7507] = 32'h0;  // 32'h6608a77e;
    ram_cell[    7508] = 32'h0;  // 32'h9c1e1028;
    ram_cell[    7509] = 32'h0;  // 32'h4049cf4e;
    ram_cell[    7510] = 32'h0;  // 32'h80a074cc;
    ram_cell[    7511] = 32'h0;  // 32'h45ef97d7;
    ram_cell[    7512] = 32'h0;  // 32'h93455d8d;
    ram_cell[    7513] = 32'h0;  // 32'h6e30df01;
    ram_cell[    7514] = 32'h0;  // 32'hf7c4cfb6;
    ram_cell[    7515] = 32'h0;  // 32'he01eb0d7;
    ram_cell[    7516] = 32'h0;  // 32'h91871e4d;
    ram_cell[    7517] = 32'h0;  // 32'h2dab5b99;
    ram_cell[    7518] = 32'h0;  // 32'h361531d8;
    ram_cell[    7519] = 32'h0;  // 32'h0f97830d;
    ram_cell[    7520] = 32'h0;  // 32'hd74098a8;
    ram_cell[    7521] = 32'h0;  // 32'h5c8f6925;
    ram_cell[    7522] = 32'h0;  // 32'hb371b213;
    ram_cell[    7523] = 32'h0;  // 32'h02faf212;
    ram_cell[    7524] = 32'h0;  // 32'hbe1d7a48;
    ram_cell[    7525] = 32'h0;  // 32'h7f393437;
    ram_cell[    7526] = 32'h0;  // 32'hebbf557e;
    ram_cell[    7527] = 32'h0;  // 32'hefe7c70e;
    ram_cell[    7528] = 32'h0;  // 32'h051d7c55;
    ram_cell[    7529] = 32'h0;  // 32'he874822f;
    ram_cell[    7530] = 32'h0;  // 32'h2b233b29;
    ram_cell[    7531] = 32'h0;  // 32'ha81ec699;
    ram_cell[    7532] = 32'h0;  // 32'hf0066ff6;
    ram_cell[    7533] = 32'h0;  // 32'h21daaa18;
    ram_cell[    7534] = 32'h0;  // 32'h48c1c8bc;
    ram_cell[    7535] = 32'h0;  // 32'hbcf90b8a;
    ram_cell[    7536] = 32'h0;  // 32'hd683276e;
    ram_cell[    7537] = 32'h0;  // 32'h85d0cc61;
    ram_cell[    7538] = 32'h0;  // 32'h0ae0683d;
    ram_cell[    7539] = 32'h0;  // 32'h1b110d2f;
    ram_cell[    7540] = 32'h0;  // 32'h95a4fe07;
    ram_cell[    7541] = 32'h0;  // 32'h650a4664;
    ram_cell[    7542] = 32'h0;  // 32'h445ee404;
    ram_cell[    7543] = 32'h0;  // 32'h2dbafbb9;
    ram_cell[    7544] = 32'h0;  // 32'h1a3badd8;
    ram_cell[    7545] = 32'h0;  // 32'h85c67827;
    ram_cell[    7546] = 32'h0;  // 32'h12af29d3;
    ram_cell[    7547] = 32'h0;  // 32'h7265bae4;
    ram_cell[    7548] = 32'h0;  // 32'hb5883248;
    ram_cell[    7549] = 32'h0;  // 32'he16b218c;
    ram_cell[    7550] = 32'h0;  // 32'h0393a401;
    ram_cell[    7551] = 32'h0;  // 32'h6b5bb5bb;
    ram_cell[    7552] = 32'h0;  // 32'hffc0e867;
    ram_cell[    7553] = 32'h0;  // 32'h25a27afc;
    ram_cell[    7554] = 32'h0;  // 32'h7d54e590;
    ram_cell[    7555] = 32'h0;  // 32'h7f70b79a;
    ram_cell[    7556] = 32'h0;  // 32'h3d59ad73;
    ram_cell[    7557] = 32'h0;  // 32'h95cb32e4;
    ram_cell[    7558] = 32'h0;  // 32'h6959e0de;
    ram_cell[    7559] = 32'h0;  // 32'ha731301b;
    ram_cell[    7560] = 32'h0;  // 32'h956022a6;
    ram_cell[    7561] = 32'h0;  // 32'hde56a2fa;
    ram_cell[    7562] = 32'h0;  // 32'h4e18edfa;
    ram_cell[    7563] = 32'h0;  // 32'h169d3bde;
    ram_cell[    7564] = 32'h0;  // 32'h6be34475;
    ram_cell[    7565] = 32'h0;  // 32'h87e12a71;
    ram_cell[    7566] = 32'h0;  // 32'h5f7c7c98;
    ram_cell[    7567] = 32'h0;  // 32'h48bbfa9b;
    ram_cell[    7568] = 32'h0;  // 32'h0a67933b;
    ram_cell[    7569] = 32'h0;  // 32'hc573f917;
    ram_cell[    7570] = 32'h0;  // 32'h744df87b;
    ram_cell[    7571] = 32'h0;  // 32'h1b2c8b37;
    ram_cell[    7572] = 32'h0;  // 32'h1d394db1;
    ram_cell[    7573] = 32'h0;  // 32'hc45b4966;
    ram_cell[    7574] = 32'h0;  // 32'hf8e67ccd;
    ram_cell[    7575] = 32'h0;  // 32'h7ab2b320;
    ram_cell[    7576] = 32'h0;  // 32'he4832cc6;
    ram_cell[    7577] = 32'h0;  // 32'h336a5eef;
    ram_cell[    7578] = 32'h0;  // 32'hf3d9fe1a;
    ram_cell[    7579] = 32'h0;  // 32'hdfbb2911;
    ram_cell[    7580] = 32'h0;  // 32'hc146bc48;
    ram_cell[    7581] = 32'h0;  // 32'hf2494b15;
    ram_cell[    7582] = 32'h0;  // 32'h14a73451;
    ram_cell[    7583] = 32'h0;  // 32'hd22b537d;
    ram_cell[    7584] = 32'h0;  // 32'h0bac798c;
    ram_cell[    7585] = 32'h0;  // 32'h84fb9fee;
    ram_cell[    7586] = 32'h0;  // 32'h978ac326;
    ram_cell[    7587] = 32'h0;  // 32'h761a39bf;
    ram_cell[    7588] = 32'h0;  // 32'h3c8971f9;
    ram_cell[    7589] = 32'h0;  // 32'hf19d6a3c;
    ram_cell[    7590] = 32'h0;  // 32'h7824c7ad;
    ram_cell[    7591] = 32'h0;  // 32'h16884041;
    ram_cell[    7592] = 32'h0;  // 32'h242add17;
    ram_cell[    7593] = 32'h0;  // 32'hdde313b2;
    ram_cell[    7594] = 32'h0;  // 32'hf6dc1863;
    ram_cell[    7595] = 32'h0;  // 32'h46c2604f;
    ram_cell[    7596] = 32'h0;  // 32'h575473cc;
    ram_cell[    7597] = 32'h0;  // 32'h8499a817;
    ram_cell[    7598] = 32'h0;  // 32'h2fdaa518;
    ram_cell[    7599] = 32'h0;  // 32'h595a1942;
    ram_cell[    7600] = 32'h0;  // 32'hd312a917;
    ram_cell[    7601] = 32'h0;  // 32'h0495d282;
    ram_cell[    7602] = 32'h0;  // 32'h8be75f64;
    ram_cell[    7603] = 32'h0;  // 32'h109b8064;
    ram_cell[    7604] = 32'h0;  // 32'h7a3e65d0;
    ram_cell[    7605] = 32'h0;  // 32'h12798469;
    ram_cell[    7606] = 32'h0;  // 32'h9aac9f44;
    ram_cell[    7607] = 32'h0;  // 32'h40db7955;
    ram_cell[    7608] = 32'h0;  // 32'h9d23a567;
    ram_cell[    7609] = 32'h0;  // 32'h05213061;
    ram_cell[    7610] = 32'h0;  // 32'h26193006;
    ram_cell[    7611] = 32'h0;  // 32'h722007b6;
    ram_cell[    7612] = 32'h0;  // 32'h1001556e;
    ram_cell[    7613] = 32'h0;  // 32'h8ee1218b;
    ram_cell[    7614] = 32'h0;  // 32'h060f4776;
    ram_cell[    7615] = 32'h0;  // 32'h81690ec5;
    ram_cell[    7616] = 32'h0;  // 32'h466f00bd;
    ram_cell[    7617] = 32'h0;  // 32'hac898af2;
    ram_cell[    7618] = 32'h0;  // 32'h00b079b7;
    ram_cell[    7619] = 32'h0;  // 32'h36735409;
    ram_cell[    7620] = 32'h0;  // 32'h4ee8c719;
    ram_cell[    7621] = 32'h0;  // 32'h6b8e6656;
    ram_cell[    7622] = 32'h0;  // 32'h350c1630;
    ram_cell[    7623] = 32'h0;  // 32'h329058cb;
    ram_cell[    7624] = 32'h0;  // 32'h2c722078;
    ram_cell[    7625] = 32'h0;  // 32'h44d0584d;
    ram_cell[    7626] = 32'h0;  // 32'h77216540;
    ram_cell[    7627] = 32'h0;  // 32'hcb67329f;
    ram_cell[    7628] = 32'h0;  // 32'h3efc2815;
    ram_cell[    7629] = 32'h0;  // 32'h0600f305;
    ram_cell[    7630] = 32'h0;  // 32'h9f713d6d;
    ram_cell[    7631] = 32'h0;  // 32'h5dfc2551;
    ram_cell[    7632] = 32'h0;  // 32'h8b35a21d;
    ram_cell[    7633] = 32'h0;  // 32'h0b0c3d91;
    ram_cell[    7634] = 32'h0;  // 32'hc476bc02;
    ram_cell[    7635] = 32'h0;  // 32'hbe6af43e;
    ram_cell[    7636] = 32'h0;  // 32'h3cb2e966;
    ram_cell[    7637] = 32'h0;  // 32'hf372a322;
    ram_cell[    7638] = 32'h0;  // 32'h0d56b493;
    ram_cell[    7639] = 32'h0;  // 32'h1dfa0c05;
    ram_cell[    7640] = 32'h0;  // 32'hcecd994b;
    ram_cell[    7641] = 32'h0;  // 32'h1f421529;
    ram_cell[    7642] = 32'h0;  // 32'hbb346984;
    ram_cell[    7643] = 32'h0;  // 32'h8a0fcada;
    ram_cell[    7644] = 32'h0;  // 32'h46704fc7;
    ram_cell[    7645] = 32'h0;  // 32'h09aea9d0;
    ram_cell[    7646] = 32'h0;  // 32'h76f383ce;
    ram_cell[    7647] = 32'h0;  // 32'h222d97fa;
    ram_cell[    7648] = 32'h0;  // 32'h1246afb3;
    ram_cell[    7649] = 32'h0;  // 32'hc4ec1bb7;
    ram_cell[    7650] = 32'h0;  // 32'h4d17bf34;
    ram_cell[    7651] = 32'h0;  // 32'h8601be96;
    ram_cell[    7652] = 32'h0;  // 32'h8d1da1b1;
    ram_cell[    7653] = 32'h0;  // 32'h482a29d0;
    ram_cell[    7654] = 32'h0;  // 32'h2c55a9fa;
    ram_cell[    7655] = 32'h0;  // 32'h4275efaa;
    ram_cell[    7656] = 32'h0;  // 32'h4b609ebf;
    ram_cell[    7657] = 32'h0;  // 32'h616a8425;
    ram_cell[    7658] = 32'h0;  // 32'hfe3c4acc;
    ram_cell[    7659] = 32'h0;  // 32'hd7d7bf59;
    ram_cell[    7660] = 32'h0;  // 32'h23a139a1;
    ram_cell[    7661] = 32'h0;  // 32'h051adc18;
    ram_cell[    7662] = 32'h0;  // 32'h468fb8da;
    ram_cell[    7663] = 32'h0;  // 32'h304bc9e4;
    ram_cell[    7664] = 32'h0;  // 32'h7f085597;
    ram_cell[    7665] = 32'h0;  // 32'ha245ab89;
    ram_cell[    7666] = 32'h0;  // 32'h2950bbb2;
    ram_cell[    7667] = 32'h0;  // 32'h6342a4ee;
    ram_cell[    7668] = 32'h0;  // 32'h0c40252f;
    ram_cell[    7669] = 32'h0;  // 32'h795e8f55;
    ram_cell[    7670] = 32'h0;  // 32'haa7d1d37;
    ram_cell[    7671] = 32'h0;  // 32'h8d2ef4cc;
    ram_cell[    7672] = 32'h0;  // 32'h6580ca02;
    ram_cell[    7673] = 32'h0;  // 32'h1c0170dd;
    ram_cell[    7674] = 32'h0;  // 32'h3f1a74af;
    ram_cell[    7675] = 32'h0;  // 32'hcc784262;
    ram_cell[    7676] = 32'h0;  // 32'h00cb665c;
    ram_cell[    7677] = 32'h0;  // 32'he988844b;
    ram_cell[    7678] = 32'h0;  // 32'hf081553c;
    ram_cell[    7679] = 32'h0;  // 32'h5f7ebc48;
    ram_cell[    7680] = 32'h0;  // 32'h19e03799;
    ram_cell[    7681] = 32'h0;  // 32'h679a4fd2;
    ram_cell[    7682] = 32'h0;  // 32'h8f53c3e1;
    ram_cell[    7683] = 32'h0;  // 32'h8522e458;
    ram_cell[    7684] = 32'h0;  // 32'hdd4d79e5;
    ram_cell[    7685] = 32'h0;  // 32'hc7dfc697;
    ram_cell[    7686] = 32'h0;  // 32'h6b603331;
    ram_cell[    7687] = 32'h0;  // 32'hc28e14fb;
    ram_cell[    7688] = 32'h0;  // 32'h9dfa6b0b;
    ram_cell[    7689] = 32'h0;  // 32'h02c1d656;
    ram_cell[    7690] = 32'h0;  // 32'h690b271f;
    ram_cell[    7691] = 32'h0;  // 32'hd06e212a;
    ram_cell[    7692] = 32'h0;  // 32'h8f6adf00;
    ram_cell[    7693] = 32'h0;  // 32'h753c01e9;
    ram_cell[    7694] = 32'h0;  // 32'h626220e0;
    ram_cell[    7695] = 32'h0;  // 32'h74aec908;
    ram_cell[    7696] = 32'h0;  // 32'h7e44dce1;
    ram_cell[    7697] = 32'h0;  // 32'h666f9e42;
    ram_cell[    7698] = 32'h0;  // 32'h73cd2ab1;
    ram_cell[    7699] = 32'h0;  // 32'h74a2cc8d;
    ram_cell[    7700] = 32'h0;  // 32'hfcfb1a10;
    ram_cell[    7701] = 32'h0;  // 32'hf7d412fb;
    ram_cell[    7702] = 32'h0;  // 32'h3cd50970;
    ram_cell[    7703] = 32'h0;  // 32'h09607523;
    ram_cell[    7704] = 32'h0;  // 32'h5931664b;
    ram_cell[    7705] = 32'h0;  // 32'he6be4131;
    ram_cell[    7706] = 32'h0;  // 32'h1cbb0b16;
    ram_cell[    7707] = 32'h0;  // 32'h3b6b9090;
    ram_cell[    7708] = 32'h0;  // 32'h442ae64e;
    ram_cell[    7709] = 32'h0;  // 32'h84ba6dd9;
    ram_cell[    7710] = 32'h0;  // 32'hb3f60de2;
    ram_cell[    7711] = 32'h0;  // 32'h52bb8ed8;
    ram_cell[    7712] = 32'h0;  // 32'h3f72cce1;
    ram_cell[    7713] = 32'h0;  // 32'h2bd661ad;
    ram_cell[    7714] = 32'h0;  // 32'h8ec60a35;
    ram_cell[    7715] = 32'h0;  // 32'h1b8d72dc;
    ram_cell[    7716] = 32'h0;  // 32'hc154a90a;
    ram_cell[    7717] = 32'h0;  // 32'h14dfd4be;
    ram_cell[    7718] = 32'h0;  // 32'h47a9cb77;
    ram_cell[    7719] = 32'h0;  // 32'hdec62ec9;
    ram_cell[    7720] = 32'h0;  // 32'hfb66595e;
    ram_cell[    7721] = 32'h0;  // 32'h635cd8fc;
    ram_cell[    7722] = 32'h0;  // 32'hc509ae62;
    ram_cell[    7723] = 32'h0;  // 32'h96d15794;
    ram_cell[    7724] = 32'h0;  // 32'h98c3deec;
    ram_cell[    7725] = 32'h0;  // 32'hc48b4ba7;
    ram_cell[    7726] = 32'h0;  // 32'h05cec9a2;
    ram_cell[    7727] = 32'h0;  // 32'h330a720e;
    ram_cell[    7728] = 32'h0;  // 32'h21b8efb9;
    ram_cell[    7729] = 32'h0;  // 32'h40bda401;
    ram_cell[    7730] = 32'h0;  // 32'h180a1635;
    ram_cell[    7731] = 32'h0;  // 32'h8bd9321f;
    ram_cell[    7732] = 32'h0;  // 32'hf2ce0090;
    ram_cell[    7733] = 32'h0;  // 32'h833c6dbf;
    ram_cell[    7734] = 32'h0;  // 32'he751ff19;
    ram_cell[    7735] = 32'h0;  // 32'hff68f57c;
    ram_cell[    7736] = 32'h0;  // 32'h2a6d621f;
    ram_cell[    7737] = 32'h0;  // 32'ha5c61adf;
    ram_cell[    7738] = 32'h0;  // 32'h8f205bec;
    ram_cell[    7739] = 32'h0;  // 32'h83fc46ab;
    ram_cell[    7740] = 32'h0;  // 32'hc96bf894;
    ram_cell[    7741] = 32'h0;  // 32'h0af82541;
    ram_cell[    7742] = 32'h0;  // 32'h230dbe4d;
    ram_cell[    7743] = 32'h0;  // 32'hbc9c60dc;
    ram_cell[    7744] = 32'h0;  // 32'h34f49267;
    ram_cell[    7745] = 32'h0;  // 32'h795357d1;
    ram_cell[    7746] = 32'h0;  // 32'h04c0303f;
    ram_cell[    7747] = 32'h0;  // 32'h2284269b;
    ram_cell[    7748] = 32'h0;  // 32'hfef246c7;
    ram_cell[    7749] = 32'h0;  // 32'h42f7ce1a;
    ram_cell[    7750] = 32'h0;  // 32'h28704d14;
    ram_cell[    7751] = 32'h0;  // 32'h1ef57c6e;
    ram_cell[    7752] = 32'h0;  // 32'h8e43cf1e;
    ram_cell[    7753] = 32'h0;  // 32'h5244d54a;
    ram_cell[    7754] = 32'h0;  // 32'h1db5ba85;
    ram_cell[    7755] = 32'h0;  // 32'h4a44aa02;
    ram_cell[    7756] = 32'h0;  // 32'h8f91e8df;
    ram_cell[    7757] = 32'h0;  // 32'h3d03a3fe;
    ram_cell[    7758] = 32'h0;  // 32'h32bc7964;
    ram_cell[    7759] = 32'h0;  // 32'hb44461b4;
    ram_cell[    7760] = 32'h0;  // 32'hb461c784;
    ram_cell[    7761] = 32'h0;  // 32'h4437e4c2;
    ram_cell[    7762] = 32'h0;  // 32'haeb1b247;
    ram_cell[    7763] = 32'h0;  // 32'h180d3675;
    ram_cell[    7764] = 32'h0;  // 32'h13d4feab;
    ram_cell[    7765] = 32'h0;  // 32'h664a5785;
    ram_cell[    7766] = 32'h0;  // 32'h1badf248;
    ram_cell[    7767] = 32'h0;  // 32'h37b45c48;
    ram_cell[    7768] = 32'h0;  // 32'haf9a2536;
    ram_cell[    7769] = 32'h0;  // 32'he1137aec;
    ram_cell[    7770] = 32'h0;  // 32'had7f5a79;
    ram_cell[    7771] = 32'h0;  // 32'hbfe6e675;
    ram_cell[    7772] = 32'h0;  // 32'hc756daba;
    ram_cell[    7773] = 32'h0;  // 32'hd859a31a;
    ram_cell[    7774] = 32'h0;  // 32'h9db1dfdf;
    ram_cell[    7775] = 32'h0;  // 32'hd4406f0a;
    ram_cell[    7776] = 32'h0;  // 32'ha6e1980d;
    ram_cell[    7777] = 32'h0;  // 32'h77786ba7;
    ram_cell[    7778] = 32'h0;  // 32'h529df127;
    ram_cell[    7779] = 32'h0;  // 32'h94886ba2;
    ram_cell[    7780] = 32'h0;  // 32'h84c7a644;
    ram_cell[    7781] = 32'h0;  // 32'h46d96c07;
    ram_cell[    7782] = 32'h0;  // 32'h9cd9becc;
    ram_cell[    7783] = 32'h0;  // 32'hc1d470d0;
    ram_cell[    7784] = 32'h0;  // 32'h29788f86;
    ram_cell[    7785] = 32'h0;  // 32'h636205f5;
    ram_cell[    7786] = 32'h0;  // 32'hdafd66de;
    ram_cell[    7787] = 32'h0;  // 32'h83537d6b;
    ram_cell[    7788] = 32'h0;  // 32'hbb4ca67c;
    ram_cell[    7789] = 32'h0;  // 32'hf07b5269;
    ram_cell[    7790] = 32'h0;  // 32'h9ac51ddc;
    ram_cell[    7791] = 32'h0;  // 32'he2a3b52e;
    ram_cell[    7792] = 32'h0;  // 32'h1e4a9daf;
    ram_cell[    7793] = 32'h0;  // 32'h942dc8de;
    ram_cell[    7794] = 32'h0;  // 32'h9ae33334;
    ram_cell[    7795] = 32'h0;  // 32'he50f851f;
    ram_cell[    7796] = 32'h0;  // 32'h06e995ac;
    ram_cell[    7797] = 32'h0;  // 32'h87896f92;
    ram_cell[    7798] = 32'h0;  // 32'hcb747126;
    ram_cell[    7799] = 32'h0;  // 32'he146013a;
    ram_cell[    7800] = 32'h0;  // 32'h29e40b2f;
    ram_cell[    7801] = 32'h0;  // 32'h513e1ceb;
    ram_cell[    7802] = 32'h0;  // 32'hbf5edd91;
    ram_cell[    7803] = 32'h0;  // 32'h8a7cbcd2;
    ram_cell[    7804] = 32'h0;  // 32'h4b24f434;
    ram_cell[    7805] = 32'h0;  // 32'h1b8929b4;
    ram_cell[    7806] = 32'h0;  // 32'h8b760978;
    ram_cell[    7807] = 32'h0;  // 32'h399b34dd;
    ram_cell[    7808] = 32'h0;  // 32'h427fc7a0;
    ram_cell[    7809] = 32'h0;  // 32'h8a67b01f;
    ram_cell[    7810] = 32'h0;  // 32'h9fbca46d;
    ram_cell[    7811] = 32'h0;  // 32'h969e66ca;
    ram_cell[    7812] = 32'h0;  // 32'h8b17e8b2;
    ram_cell[    7813] = 32'h0;  // 32'h3fd99218;
    ram_cell[    7814] = 32'h0;  // 32'h8f79cf39;
    ram_cell[    7815] = 32'h0;  // 32'hb5f17503;
    ram_cell[    7816] = 32'h0;  // 32'hb591cbe6;
    ram_cell[    7817] = 32'h0;  // 32'hd2b94637;
    ram_cell[    7818] = 32'h0;  // 32'h0dfb48a8;
    ram_cell[    7819] = 32'h0;  // 32'h687f8051;
    ram_cell[    7820] = 32'h0;  // 32'h48230c7a;
    ram_cell[    7821] = 32'h0;  // 32'h97ecbfe8;
    ram_cell[    7822] = 32'h0;  // 32'h850f4a3d;
    ram_cell[    7823] = 32'h0;  // 32'hce62c9a3;
    ram_cell[    7824] = 32'h0;  // 32'h85d61ce0;
    ram_cell[    7825] = 32'h0;  // 32'h2502f04c;
    ram_cell[    7826] = 32'h0;  // 32'h21786dc0;
    ram_cell[    7827] = 32'h0;  // 32'h4e4e60a8;
    ram_cell[    7828] = 32'h0;  // 32'hbf19fc4d;
    ram_cell[    7829] = 32'h0;  // 32'ha0218582;
    ram_cell[    7830] = 32'h0;  // 32'h0de60d18;
    ram_cell[    7831] = 32'h0;  // 32'hacf21f26;
    ram_cell[    7832] = 32'h0;  // 32'h2db9c15b;
    ram_cell[    7833] = 32'h0;  // 32'heb79ffe7;
    ram_cell[    7834] = 32'h0;  // 32'h014eb964;
    ram_cell[    7835] = 32'h0;  // 32'h30367cf8;
    ram_cell[    7836] = 32'h0;  // 32'h72b7d227;
    ram_cell[    7837] = 32'h0;  // 32'ha07f41d9;
    ram_cell[    7838] = 32'h0;  // 32'hf591f7ca;
    ram_cell[    7839] = 32'h0;  // 32'h404ad63e;
    ram_cell[    7840] = 32'h0;  // 32'h8fe14de9;
    ram_cell[    7841] = 32'h0;  // 32'hc390adaa;
    ram_cell[    7842] = 32'h0;  // 32'h51c386a9;
    ram_cell[    7843] = 32'h0;  // 32'h6cfdcb55;
    ram_cell[    7844] = 32'h0;  // 32'h55921aee;
    ram_cell[    7845] = 32'h0;  // 32'hec3cf807;
    ram_cell[    7846] = 32'h0;  // 32'hf02169de;
    ram_cell[    7847] = 32'h0;  // 32'hdd83a84d;
    ram_cell[    7848] = 32'h0;  // 32'h2da605a2;
    ram_cell[    7849] = 32'h0;  // 32'h351a3c65;
    ram_cell[    7850] = 32'h0;  // 32'h934eb728;
    ram_cell[    7851] = 32'h0;  // 32'h0f6c67ad;
    ram_cell[    7852] = 32'h0;  // 32'h5ec70add;
    ram_cell[    7853] = 32'h0;  // 32'h0461d4a7;
    ram_cell[    7854] = 32'h0;  // 32'ha404abc5;
    ram_cell[    7855] = 32'h0;  // 32'h40a81fd4;
    ram_cell[    7856] = 32'h0;  // 32'hb4e2f435;
    ram_cell[    7857] = 32'h0;  // 32'hca9c8ed2;
    ram_cell[    7858] = 32'h0;  // 32'hcf1bc0e7;
    ram_cell[    7859] = 32'h0;  // 32'h40e336d1;
    ram_cell[    7860] = 32'h0;  // 32'h56feb14a;
    ram_cell[    7861] = 32'h0;  // 32'he407c688;
    ram_cell[    7862] = 32'h0;  // 32'h614fcbc0;
    ram_cell[    7863] = 32'h0;  // 32'he9d9bb24;
    ram_cell[    7864] = 32'h0;  // 32'h2491c501;
    ram_cell[    7865] = 32'h0;  // 32'h63a6bd29;
    ram_cell[    7866] = 32'h0;  // 32'ha8eea535;
    ram_cell[    7867] = 32'h0;  // 32'h50ee6237;
    ram_cell[    7868] = 32'h0;  // 32'h73444ff5;
    ram_cell[    7869] = 32'h0;  // 32'h917fcf75;
    ram_cell[    7870] = 32'h0;  // 32'h00bd360c;
    ram_cell[    7871] = 32'h0;  // 32'hf180f361;
    ram_cell[    7872] = 32'h0;  // 32'h2f317bac;
    ram_cell[    7873] = 32'h0;  // 32'ha9fc259e;
    ram_cell[    7874] = 32'h0;  // 32'h8502095e;
    ram_cell[    7875] = 32'h0;  // 32'h58e5f799;
    ram_cell[    7876] = 32'h0;  // 32'hb4c2f1df;
    ram_cell[    7877] = 32'h0;  // 32'h7ebc8ce0;
    ram_cell[    7878] = 32'h0;  // 32'h4f370020;
    ram_cell[    7879] = 32'h0;  // 32'h4bc4e437;
    ram_cell[    7880] = 32'h0;  // 32'h4e89a315;
    ram_cell[    7881] = 32'h0;  // 32'haa2731b1;
    ram_cell[    7882] = 32'h0;  // 32'h444e5fb9;
    ram_cell[    7883] = 32'h0;  // 32'hf17cb295;
    ram_cell[    7884] = 32'h0;  // 32'hb8db885a;
    ram_cell[    7885] = 32'h0;  // 32'h018c1835;
    ram_cell[    7886] = 32'h0;  // 32'h059fa1f5;
    ram_cell[    7887] = 32'h0;  // 32'h5bba6a52;
    ram_cell[    7888] = 32'h0;  // 32'h10f928c1;
    ram_cell[    7889] = 32'h0;  // 32'h1a808ed4;
    ram_cell[    7890] = 32'h0;  // 32'h2eac8811;
    ram_cell[    7891] = 32'h0;  // 32'ha6d557c3;
    ram_cell[    7892] = 32'h0;  // 32'he791a04d;
    ram_cell[    7893] = 32'h0;  // 32'h139d7a49;
    ram_cell[    7894] = 32'h0;  // 32'h8a61b89a;
    ram_cell[    7895] = 32'h0;  // 32'h9153f493;
    ram_cell[    7896] = 32'h0;  // 32'hcf39ca65;
    ram_cell[    7897] = 32'h0;  // 32'h054096ef;
    ram_cell[    7898] = 32'h0;  // 32'h33f46652;
    ram_cell[    7899] = 32'h0;  // 32'hc019468c;
    ram_cell[    7900] = 32'h0;  // 32'hc49bcd49;
    ram_cell[    7901] = 32'h0;  // 32'h410584ac;
    ram_cell[    7902] = 32'h0;  // 32'h72ec7f92;
    ram_cell[    7903] = 32'h0;  // 32'h4ea96bbb;
    ram_cell[    7904] = 32'h0;  // 32'h27b6c97e;
    ram_cell[    7905] = 32'h0;  // 32'hf0bd6843;
    ram_cell[    7906] = 32'h0;  // 32'h8019af81;
    ram_cell[    7907] = 32'h0;  // 32'hd6bf3dc5;
    ram_cell[    7908] = 32'h0;  // 32'h6053671d;
    ram_cell[    7909] = 32'h0;  // 32'h96d01fb9;
    ram_cell[    7910] = 32'h0;  // 32'he5aae660;
    ram_cell[    7911] = 32'h0;  // 32'he4f4ab4b;
    ram_cell[    7912] = 32'h0;  // 32'h43c7f616;
    ram_cell[    7913] = 32'h0;  // 32'he14e256c;
    ram_cell[    7914] = 32'h0;  // 32'hdf97437b;
    ram_cell[    7915] = 32'h0;  // 32'hbb576672;
    ram_cell[    7916] = 32'h0;  // 32'hb9b2e818;
    ram_cell[    7917] = 32'h0;  // 32'hf3049194;
    ram_cell[    7918] = 32'h0;  // 32'h0f5ec834;
    ram_cell[    7919] = 32'h0;  // 32'he0a0e38b;
    ram_cell[    7920] = 32'h0;  // 32'h8c74bd03;
    ram_cell[    7921] = 32'h0;  // 32'h8a6c96bd;
    ram_cell[    7922] = 32'h0;  // 32'hc68b8663;
    ram_cell[    7923] = 32'h0;  // 32'hd840fede;
    ram_cell[    7924] = 32'h0;  // 32'h55db9057;
    ram_cell[    7925] = 32'h0;  // 32'hcb822f33;
    ram_cell[    7926] = 32'h0;  // 32'h5e754001;
    ram_cell[    7927] = 32'h0;  // 32'h480e6bd7;
    ram_cell[    7928] = 32'h0;  // 32'h3e894cb1;
    ram_cell[    7929] = 32'h0;  // 32'h2ebbabf8;
    ram_cell[    7930] = 32'h0;  // 32'h2f2d9049;
    ram_cell[    7931] = 32'h0;  // 32'h2061b71b;
    ram_cell[    7932] = 32'h0;  // 32'h484ea067;
    ram_cell[    7933] = 32'h0;  // 32'h6a41673f;
    ram_cell[    7934] = 32'h0;  // 32'hfe4e8a61;
    ram_cell[    7935] = 32'h0;  // 32'h5b1db809;
    ram_cell[    7936] = 32'h0;  // 32'h12a58afa;
    ram_cell[    7937] = 32'h0;  // 32'hd297aa81;
    ram_cell[    7938] = 32'h0;  // 32'h9b7b2868;
    ram_cell[    7939] = 32'h0;  // 32'h5b40195e;
    ram_cell[    7940] = 32'h0;  // 32'h8e9d9910;
    ram_cell[    7941] = 32'h0;  // 32'hf6721c48;
    ram_cell[    7942] = 32'h0;  // 32'hfdd3c169;
    ram_cell[    7943] = 32'h0;  // 32'h62ccb655;
    ram_cell[    7944] = 32'h0;  // 32'he1b6ce21;
    ram_cell[    7945] = 32'h0;  // 32'h55fee53d;
    ram_cell[    7946] = 32'h0;  // 32'h48b74172;
    ram_cell[    7947] = 32'h0;  // 32'hf0f99430;
    ram_cell[    7948] = 32'h0;  // 32'hc952348f;
    ram_cell[    7949] = 32'h0;  // 32'h9e5a3006;
    ram_cell[    7950] = 32'h0;  // 32'he6fb02f7;
    ram_cell[    7951] = 32'h0;  // 32'hadcb3444;
    ram_cell[    7952] = 32'h0;  // 32'ha659fcab;
    ram_cell[    7953] = 32'h0;  // 32'h29ffd310;
    ram_cell[    7954] = 32'h0;  // 32'h4aee9e81;
    ram_cell[    7955] = 32'h0;  // 32'hdfab9a4f;
    ram_cell[    7956] = 32'h0;  // 32'h22a0a02f;
    ram_cell[    7957] = 32'h0;  // 32'h6a2e083d;
    ram_cell[    7958] = 32'h0;  // 32'hb7b936f3;
    ram_cell[    7959] = 32'h0;  // 32'hc914887c;
    ram_cell[    7960] = 32'h0;  // 32'hc7ab9019;
    ram_cell[    7961] = 32'h0;  // 32'hb3e6cd8b;
    ram_cell[    7962] = 32'h0;  // 32'h97b2dd77;
    ram_cell[    7963] = 32'h0;  // 32'hed1099dd;
    ram_cell[    7964] = 32'h0;  // 32'h9625db5c;
    ram_cell[    7965] = 32'h0;  // 32'hc1996720;
    ram_cell[    7966] = 32'h0;  // 32'h745b0973;
    ram_cell[    7967] = 32'h0;  // 32'h4c1a8826;
    ram_cell[    7968] = 32'h0;  // 32'h416f91c0;
    ram_cell[    7969] = 32'h0;  // 32'hdbee969e;
    ram_cell[    7970] = 32'h0;  // 32'h0782b573;
    ram_cell[    7971] = 32'h0;  // 32'hb96f18f9;
    ram_cell[    7972] = 32'h0;  // 32'hfb08e6c5;
    ram_cell[    7973] = 32'h0;  // 32'h0f3a3d80;
    ram_cell[    7974] = 32'h0;  // 32'h35621e17;
    ram_cell[    7975] = 32'h0;  // 32'hc44f1a3c;
    ram_cell[    7976] = 32'h0;  // 32'hfc49f6c4;
    ram_cell[    7977] = 32'h0;  // 32'h7f0e1b57;
    ram_cell[    7978] = 32'h0;  // 32'h93554b7b;
    ram_cell[    7979] = 32'h0;  // 32'he2913aca;
    ram_cell[    7980] = 32'h0;  // 32'hf848e7ea;
    ram_cell[    7981] = 32'h0;  // 32'h5447a445;
    ram_cell[    7982] = 32'h0;  // 32'h364c39cc;
    ram_cell[    7983] = 32'h0;  // 32'he8a56de4;
    ram_cell[    7984] = 32'h0;  // 32'h5c04b32b;
    ram_cell[    7985] = 32'h0;  // 32'h11991083;
    ram_cell[    7986] = 32'h0;  // 32'hf76af161;
    ram_cell[    7987] = 32'h0;  // 32'haba8c497;
    ram_cell[    7988] = 32'h0;  // 32'hf4c641a3;
    ram_cell[    7989] = 32'h0;  // 32'hdb2e342b;
    ram_cell[    7990] = 32'h0;  // 32'h6d61783a;
    ram_cell[    7991] = 32'h0;  // 32'h8e4514b2;
    ram_cell[    7992] = 32'h0;  // 32'h8241ca9b;
    ram_cell[    7993] = 32'h0;  // 32'h1420bf6a;
    ram_cell[    7994] = 32'h0;  // 32'hd4c4ab1c;
    ram_cell[    7995] = 32'h0;  // 32'h4363fd28;
    ram_cell[    7996] = 32'h0;  // 32'h377abb5b;
    ram_cell[    7997] = 32'h0;  // 32'h1ceb1072;
    ram_cell[    7998] = 32'h0;  // 32'he9d909e4;
    ram_cell[    7999] = 32'h0;  // 32'h0005e3db;
    ram_cell[    8000] = 32'h0;  // 32'hf09f85f3;
    ram_cell[    8001] = 32'h0;  // 32'h7be0ccd0;
    ram_cell[    8002] = 32'h0;  // 32'hf2b54d42;
    ram_cell[    8003] = 32'h0;  // 32'h094fdd77;
    ram_cell[    8004] = 32'h0;  // 32'hb8a6da55;
    ram_cell[    8005] = 32'h0;  // 32'h4322599e;
    ram_cell[    8006] = 32'h0;  // 32'hd1752035;
    ram_cell[    8007] = 32'h0;  // 32'h68947fcc;
    ram_cell[    8008] = 32'h0;  // 32'h4fec6490;
    ram_cell[    8009] = 32'h0;  // 32'h2d577405;
    ram_cell[    8010] = 32'h0;  // 32'h5a3c0e8a;
    ram_cell[    8011] = 32'h0;  // 32'h97d8fae5;
    ram_cell[    8012] = 32'h0;  // 32'h1d8e8dbf;
    ram_cell[    8013] = 32'h0;  // 32'he6b0ce7a;
    ram_cell[    8014] = 32'h0;  // 32'h1341dc7a;
    ram_cell[    8015] = 32'h0;  // 32'h0889a18d;
    ram_cell[    8016] = 32'h0;  // 32'h592e4d96;
    ram_cell[    8017] = 32'h0;  // 32'hfafaa5d3;
    ram_cell[    8018] = 32'h0;  // 32'hb08d5ddb;
    ram_cell[    8019] = 32'h0;  // 32'h1dee5549;
    ram_cell[    8020] = 32'h0;  // 32'h44c54bd6;
    ram_cell[    8021] = 32'h0;  // 32'h5826a3b4;
    ram_cell[    8022] = 32'h0;  // 32'h7bceb205;
    ram_cell[    8023] = 32'h0;  // 32'h1a768431;
    ram_cell[    8024] = 32'h0;  // 32'h85963527;
    ram_cell[    8025] = 32'h0;  // 32'h12583bf5;
    ram_cell[    8026] = 32'h0;  // 32'hc629a83f;
    ram_cell[    8027] = 32'h0;  // 32'h2b1a0a8a;
    ram_cell[    8028] = 32'h0;  // 32'hf48984c2;
    ram_cell[    8029] = 32'h0;  // 32'h568a99ee;
    ram_cell[    8030] = 32'h0;  // 32'h6c91edf1;
    ram_cell[    8031] = 32'h0;  // 32'h042781e4;
    ram_cell[    8032] = 32'h0;  // 32'hf58e0b65;
    ram_cell[    8033] = 32'h0;  // 32'h912afcd1;
    ram_cell[    8034] = 32'h0;  // 32'hafc0d002;
    ram_cell[    8035] = 32'h0;  // 32'hdc73863c;
    ram_cell[    8036] = 32'h0;  // 32'h915354f0;
    ram_cell[    8037] = 32'h0;  // 32'h42a5c672;
    ram_cell[    8038] = 32'h0;  // 32'h9195d7e1;
    ram_cell[    8039] = 32'h0;  // 32'hc626b087;
    ram_cell[    8040] = 32'h0;  // 32'he17342e2;
    ram_cell[    8041] = 32'h0;  // 32'h7c6ea57a;
    ram_cell[    8042] = 32'h0;  // 32'hed5bed93;
    ram_cell[    8043] = 32'h0;  // 32'h7ef62668;
    ram_cell[    8044] = 32'h0;  // 32'hbcd61fdd;
    ram_cell[    8045] = 32'h0;  // 32'h2ad4d92a;
    ram_cell[    8046] = 32'h0;  // 32'h2b391438;
    ram_cell[    8047] = 32'h0;  // 32'ha46ccd7a;
    ram_cell[    8048] = 32'h0;  // 32'h7d012afb;
    ram_cell[    8049] = 32'h0;  // 32'hcdc41d78;
    ram_cell[    8050] = 32'h0;  // 32'h6985a1a4;
    ram_cell[    8051] = 32'h0;  // 32'h6ea33bf1;
    ram_cell[    8052] = 32'h0;  // 32'h4fbd8caa;
    ram_cell[    8053] = 32'h0;  // 32'h23b843cc;
    ram_cell[    8054] = 32'h0;  // 32'h001eaece;
    ram_cell[    8055] = 32'h0;  // 32'hcf654a2e;
    ram_cell[    8056] = 32'h0;  // 32'hed29faca;
    ram_cell[    8057] = 32'h0;  // 32'h04997cfd;
    ram_cell[    8058] = 32'h0;  // 32'ha5e4951d;
    ram_cell[    8059] = 32'h0;  // 32'hc78b9907;
    ram_cell[    8060] = 32'h0;  // 32'hcb5655e3;
    ram_cell[    8061] = 32'h0;  // 32'h17bf0827;
    ram_cell[    8062] = 32'h0;  // 32'h86f157fc;
    ram_cell[    8063] = 32'h0;  // 32'hb60ceb66;
    ram_cell[    8064] = 32'h0;  // 32'hb2284796;
    ram_cell[    8065] = 32'h0;  // 32'h20c64241;
    ram_cell[    8066] = 32'h0;  // 32'hbbc119b5;
    ram_cell[    8067] = 32'h0;  // 32'habb58a30;
    ram_cell[    8068] = 32'h0;  // 32'h76454595;
    ram_cell[    8069] = 32'h0;  // 32'h8e5b9911;
    ram_cell[    8070] = 32'h0;  // 32'h7b3dd05d;
    ram_cell[    8071] = 32'h0;  // 32'hc1e40ae1;
    ram_cell[    8072] = 32'h0;  // 32'h05d8c131;
    ram_cell[    8073] = 32'h0;  // 32'he1c6cc54;
    ram_cell[    8074] = 32'h0;  // 32'h03ce0cc2;
    ram_cell[    8075] = 32'h0;  // 32'h1ae2de6d;
    ram_cell[    8076] = 32'h0;  // 32'h30b6b0ad;
    ram_cell[    8077] = 32'h0;  // 32'he41c45a3;
    ram_cell[    8078] = 32'h0;  // 32'h9051ea6d;
    ram_cell[    8079] = 32'h0;  // 32'hb7ce90d5;
    ram_cell[    8080] = 32'h0;  // 32'h29d20714;
    ram_cell[    8081] = 32'h0;  // 32'h042c6c23;
    ram_cell[    8082] = 32'h0;  // 32'h182ac056;
    ram_cell[    8083] = 32'h0;  // 32'ha2f987b0;
    ram_cell[    8084] = 32'h0;  // 32'h3d30edda;
    ram_cell[    8085] = 32'h0;  // 32'hdd6d07f4;
    ram_cell[    8086] = 32'h0;  // 32'hcaef9ec5;
    ram_cell[    8087] = 32'h0;  // 32'hf4474859;
    ram_cell[    8088] = 32'h0;  // 32'ha722ad6d;
    ram_cell[    8089] = 32'h0;  // 32'h79b403f0;
    ram_cell[    8090] = 32'h0;  // 32'h148303bb;
    ram_cell[    8091] = 32'h0;  // 32'he36beac9;
    ram_cell[    8092] = 32'h0;  // 32'habcbb64c;
    ram_cell[    8093] = 32'h0;  // 32'h82b5f95f;
    ram_cell[    8094] = 32'h0;  // 32'h16184310;
    ram_cell[    8095] = 32'h0;  // 32'hc1086041;
    ram_cell[    8096] = 32'h0;  // 32'h710c0f27;
    ram_cell[    8097] = 32'h0;  // 32'h68882162;
    ram_cell[    8098] = 32'h0;  // 32'h618b439e;
    ram_cell[    8099] = 32'h0;  // 32'h017b3800;
    ram_cell[    8100] = 32'h0;  // 32'h9e4a957d;
    ram_cell[    8101] = 32'h0;  // 32'hb301e8a5;
    ram_cell[    8102] = 32'h0;  // 32'h4eabef00;
    ram_cell[    8103] = 32'h0;  // 32'hd4b0074f;
    ram_cell[    8104] = 32'h0;  // 32'h4fc17701;
    ram_cell[    8105] = 32'h0;  // 32'h55c3737e;
    ram_cell[    8106] = 32'h0;  // 32'h3efa1bd6;
    ram_cell[    8107] = 32'h0;  // 32'h49728174;
    ram_cell[    8108] = 32'h0;  // 32'h5c72bde4;
    ram_cell[    8109] = 32'h0;  // 32'h6b44046d;
    ram_cell[    8110] = 32'h0;  // 32'h1f6c51a2;
    ram_cell[    8111] = 32'h0;  // 32'hd4755ebe;
    ram_cell[    8112] = 32'h0;  // 32'h37fb3300;
    ram_cell[    8113] = 32'h0;  // 32'hedc0ac2e;
    ram_cell[    8114] = 32'h0;  // 32'ha69a2dea;
    ram_cell[    8115] = 32'h0;  // 32'h14375116;
    ram_cell[    8116] = 32'h0;  // 32'ha71829a0;
    ram_cell[    8117] = 32'h0;  // 32'h812d5a37;
    ram_cell[    8118] = 32'h0;  // 32'h9015a4e9;
    ram_cell[    8119] = 32'h0;  // 32'h9c010e35;
    ram_cell[    8120] = 32'h0;  // 32'hc0ef6a7f;
    ram_cell[    8121] = 32'h0;  // 32'h5c0bb79e;
    ram_cell[    8122] = 32'h0;  // 32'h8164fde4;
    ram_cell[    8123] = 32'h0;  // 32'hd7f6885b;
    ram_cell[    8124] = 32'h0;  // 32'he49ded14;
    ram_cell[    8125] = 32'h0;  // 32'h7621e75a;
    ram_cell[    8126] = 32'h0;  // 32'h19d0aa32;
    ram_cell[    8127] = 32'h0;  // 32'hcd9ae76c;
    ram_cell[    8128] = 32'h0;  // 32'h382715a7;
    ram_cell[    8129] = 32'h0;  // 32'h10ba96a9;
    ram_cell[    8130] = 32'h0;  // 32'he8412c88;
    ram_cell[    8131] = 32'h0;  // 32'h40c0a61f;
    ram_cell[    8132] = 32'h0;  // 32'h1943e03f;
    ram_cell[    8133] = 32'h0;  // 32'h1be0cd02;
    ram_cell[    8134] = 32'h0;  // 32'h4140f6a1;
    ram_cell[    8135] = 32'h0;  // 32'hfbb1a323;
    ram_cell[    8136] = 32'h0;  // 32'h47966abc;
    ram_cell[    8137] = 32'h0;  // 32'ha0f68c52;
    ram_cell[    8138] = 32'h0;  // 32'hb817bba2;
    ram_cell[    8139] = 32'h0;  // 32'h13b59f75;
    ram_cell[    8140] = 32'h0;  // 32'h49292ca1;
    ram_cell[    8141] = 32'h0;  // 32'hae66f5b3;
    ram_cell[    8142] = 32'h0;  // 32'h637cba41;
    ram_cell[    8143] = 32'h0;  // 32'h491fefbe;
    ram_cell[    8144] = 32'h0;  // 32'h3124f602;
    ram_cell[    8145] = 32'h0;  // 32'h9ee9ac8c;
    ram_cell[    8146] = 32'h0;  // 32'hee3e8fdd;
    ram_cell[    8147] = 32'h0;  // 32'h90ab854c;
    ram_cell[    8148] = 32'h0;  // 32'hd79bd306;
    ram_cell[    8149] = 32'h0;  // 32'h51cbdcef;
    ram_cell[    8150] = 32'h0;  // 32'hb6c087da;
    ram_cell[    8151] = 32'h0;  // 32'h73bb9411;
    ram_cell[    8152] = 32'h0;  // 32'he2e69cf2;
    ram_cell[    8153] = 32'h0;  // 32'hcdb89ae8;
    ram_cell[    8154] = 32'h0;  // 32'h1766d61c;
    ram_cell[    8155] = 32'h0;  // 32'h846c42a6;
    ram_cell[    8156] = 32'h0;  // 32'h1f53bbb1;
    ram_cell[    8157] = 32'h0;  // 32'hb628a4b7;
    ram_cell[    8158] = 32'h0;  // 32'h33935195;
    ram_cell[    8159] = 32'h0;  // 32'h70b5bcb1;
    ram_cell[    8160] = 32'h0;  // 32'h055b7007;
    ram_cell[    8161] = 32'h0;  // 32'hf24d42ce;
    ram_cell[    8162] = 32'h0;  // 32'h02f53ff4;
    ram_cell[    8163] = 32'h0;  // 32'h79f32b5e;
    ram_cell[    8164] = 32'h0;  // 32'h4110f9d7;
    ram_cell[    8165] = 32'h0;  // 32'h35a813ee;
    ram_cell[    8166] = 32'h0;  // 32'h3011d8ad;
    ram_cell[    8167] = 32'h0;  // 32'hf6128aeb;
    ram_cell[    8168] = 32'h0;  // 32'hd68dbcd4;
    ram_cell[    8169] = 32'h0;  // 32'hac31bb70;
    ram_cell[    8170] = 32'h0;  // 32'h09016bfb;
    ram_cell[    8171] = 32'h0;  // 32'h968cb46e;
    ram_cell[    8172] = 32'h0;  // 32'h7c77b74e;
    ram_cell[    8173] = 32'h0;  // 32'hcf75cc4e;
    ram_cell[    8174] = 32'h0;  // 32'hdfd9dfe7;
    ram_cell[    8175] = 32'h0;  // 32'hac24e806;
    ram_cell[    8176] = 32'h0;  // 32'hae086e69;
    ram_cell[    8177] = 32'h0;  // 32'h5d69509c;
    ram_cell[    8178] = 32'h0;  // 32'h4518b32a;
    ram_cell[    8179] = 32'h0;  // 32'h97663742;
    ram_cell[    8180] = 32'h0;  // 32'h56b19ac9;
    ram_cell[    8181] = 32'h0;  // 32'h0b36a2f0;
    ram_cell[    8182] = 32'h0;  // 32'hdd92decb;
    ram_cell[    8183] = 32'h0;  // 32'h08e8a660;
    ram_cell[    8184] = 32'h0;  // 32'h814763ba;
    ram_cell[    8185] = 32'h0;  // 32'he91036ad;
    ram_cell[    8186] = 32'h0;  // 32'h186e53af;
    ram_cell[    8187] = 32'h0;  // 32'h181cbdf8;
    ram_cell[    8188] = 32'h0;  // 32'haccd5dbf;
    ram_cell[    8189] = 32'h0;  // 32'hbcdddc27;
    ram_cell[    8190] = 32'h0;  // 32'h5599a6db;
    ram_cell[    8191] = 32'h0;  // 32'h60f39552;
    ram_cell[    8192] = 32'h0;  // 32'hf28942f0;
    ram_cell[    8193] = 32'h0;  // 32'h1aea4508;
    ram_cell[    8194] = 32'h0;  // 32'h0dd1f909;
    ram_cell[    8195] = 32'h0;  // 32'hbdf33f3d;
    ram_cell[    8196] = 32'h0;  // 32'he7a22b42;
    ram_cell[    8197] = 32'h0;  // 32'h10bc121e;
    ram_cell[    8198] = 32'h0;  // 32'ha08a3ab5;
    ram_cell[    8199] = 32'h0;  // 32'h2c014c54;
    ram_cell[    8200] = 32'h0;  // 32'h1be60f2d;
    ram_cell[    8201] = 32'h0;  // 32'h5c83c46f;
    ram_cell[    8202] = 32'h0;  // 32'h8344a965;
    ram_cell[    8203] = 32'h0;  // 32'h0c04a1d3;
    ram_cell[    8204] = 32'h0;  // 32'h0b8dc4eb;
    ram_cell[    8205] = 32'h0;  // 32'h7d16104c;
    ram_cell[    8206] = 32'h0;  // 32'hd6b3efba;
    ram_cell[    8207] = 32'h0;  // 32'h6a4fb9e9;
    ram_cell[    8208] = 32'h0;  // 32'hb8a55646;
    ram_cell[    8209] = 32'h0;  // 32'h7a13b8c7;
    ram_cell[    8210] = 32'h0;  // 32'h3d1a78c7;
    ram_cell[    8211] = 32'h0;  // 32'h22e10de8;
    ram_cell[    8212] = 32'h0;  // 32'h8e4e1b07;
    ram_cell[    8213] = 32'h0;  // 32'h3ab2c39a;
    ram_cell[    8214] = 32'h0;  // 32'hb449bffd;
    ram_cell[    8215] = 32'h0;  // 32'h9bacd7d8;
    ram_cell[    8216] = 32'h0;  // 32'hd286577e;
    ram_cell[    8217] = 32'h0;  // 32'hf34d99f4;
    ram_cell[    8218] = 32'h0;  // 32'h54ee2871;
    ram_cell[    8219] = 32'h0;  // 32'hbe7f5aec;
    ram_cell[    8220] = 32'h0;  // 32'h53969b61;
    ram_cell[    8221] = 32'h0;  // 32'ha7bb54d6;
    ram_cell[    8222] = 32'h0;  // 32'h5e1d1deb;
    ram_cell[    8223] = 32'h0;  // 32'h1159aac1;
    ram_cell[    8224] = 32'h0;  // 32'hb2009d14;
    ram_cell[    8225] = 32'h0;  // 32'hebf5c0d8;
    ram_cell[    8226] = 32'h0;  // 32'h406aa657;
    ram_cell[    8227] = 32'h0;  // 32'h60695a34;
    ram_cell[    8228] = 32'h0;  // 32'h387dcd92;
    ram_cell[    8229] = 32'h0;  // 32'h1ee059dd;
    ram_cell[    8230] = 32'h0;  // 32'h6e01ddd5;
    ram_cell[    8231] = 32'h0;  // 32'h04ded1d8;
    ram_cell[    8232] = 32'h0;  // 32'h83842ba4;
    ram_cell[    8233] = 32'h0;  // 32'h82a8c448;
    ram_cell[    8234] = 32'h0;  // 32'h97aa7ed8;
    ram_cell[    8235] = 32'h0;  // 32'hd2863a16;
    ram_cell[    8236] = 32'h0;  // 32'h157648ce;
    ram_cell[    8237] = 32'h0;  // 32'hec98ee3d;
    ram_cell[    8238] = 32'h0;  // 32'h40ec7175;
    ram_cell[    8239] = 32'h0;  // 32'h66f0b2ea;
    ram_cell[    8240] = 32'h0;  // 32'h6aa5401e;
    ram_cell[    8241] = 32'h0;  // 32'h6b86d2e1;
    ram_cell[    8242] = 32'h0;  // 32'h624e35bb;
    ram_cell[    8243] = 32'h0;  // 32'h7676224b;
    ram_cell[    8244] = 32'h0;  // 32'hb233496d;
    ram_cell[    8245] = 32'h0;  // 32'h7a681603;
    ram_cell[    8246] = 32'h0;  // 32'hea527755;
    ram_cell[    8247] = 32'h0;  // 32'h88813e3b;
    ram_cell[    8248] = 32'h0;  // 32'ha5f6a773;
    ram_cell[    8249] = 32'h0;  // 32'hee869c72;
    ram_cell[    8250] = 32'h0;  // 32'h1b8f7e40;
    ram_cell[    8251] = 32'h0;  // 32'hfb5cd104;
    ram_cell[    8252] = 32'h0;  // 32'h2aed8c67;
    ram_cell[    8253] = 32'h0;  // 32'h918958c4;
    ram_cell[    8254] = 32'h0;  // 32'h334eab95;
    ram_cell[    8255] = 32'h0;  // 32'hc014d15a;
    ram_cell[    8256] = 32'h0;  // 32'hadb06b6f;
    ram_cell[    8257] = 32'h0;  // 32'hab826fac;
    ram_cell[    8258] = 32'h0;  // 32'haf365bd1;
    ram_cell[    8259] = 32'h0;  // 32'he88e2ad4;
    ram_cell[    8260] = 32'h0;  // 32'hcd94ad73;
    ram_cell[    8261] = 32'h0;  // 32'hf1f38f4c;
    ram_cell[    8262] = 32'h0;  // 32'hc91ac1ee;
    ram_cell[    8263] = 32'h0;  // 32'h011e193b;
    ram_cell[    8264] = 32'h0;  // 32'h18e460be;
    ram_cell[    8265] = 32'h0;  // 32'hf3a37ab2;
    ram_cell[    8266] = 32'h0;  // 32'hb41c0bf3;
    ram_cell[    8267] = 32'h0;  // 32'ha09ad4d9;
    ram_cell[    8268] = 32'h0;  // 32'ha943170a;
    ram_cell[    8269] = 32'h0;  // 32'ha44d9242;
    ram_cell[    8270] = 32'h0;  // 32'h492d8cde;
    ram_cell[    8271] = 32'h0;  // 32'h91c04784;
    ram_cell[    8272] = 32'h0;  // 32'h04502d31;
    ram_cell[    8273] = 32'h0;  // 32'hbb0c8b91;
    ram_cell[    8274] = 32'h0;  // 32'h426a74c5;
    ram_cell[    8275] = 32'h0;  // 32'h0430722b;
    ram_cell[    8276] = 32'h0;  // 32'h44f636f1;
    ram_cell[    8277] = 32'h0;  // 32'h48014825;
    ram_cell[    8278] = 32'h0;  // 32'hbadf794c;
    ram_cell[    8279] = 32'h0;  // 32'hf9f7c186;
    ram_cell[    8280] = 32'h0;  // 32'h844eb56a;
    ram_cell[    8281] = 32'h0;  // 32'hfec26498;
    ram_cell[    8282] = 32'h0;  // 32'h7d61ad3f;
    ram_cell[    8283] = 32'h0;  // 32'h9cb0bbd5;
    ram_cell[    8284] = 32'h0;  // 32'h59455aec;
    ram_cell[    8285] = 32'h0;  // 32'h0b82d6e8;
    ram_cell[    8286] = 32'h0;  // 32'hbe9c76a4;
    ram_cell[    8287] = 32'h0;  // 32'he85b9b91;
    ram_cell[    8288] = 32'h0;  // 32'hf074e521;
    ram_cell[    8289] = 32'h0;  // 32'hf1d87e7f;
    ram_cell[    8290] = 32'h0;  // 32'hc64c5580;
    ram_cell[    8291] = 32'h0;  // 32'h5c34ade2;
    ram_cell[    8292] = 32'h0;  // 32'h4736c804;
    ram_cell[    8293] = 32'h0;  // 32'h3f15e458;
    ram_cell[    8294] = 32'h0;  // 32'h72c9123f;
    ram_cell[    8295] = 32'h0;  // 32'heb5e47e1;
    ram_cell[    8296] = 32'h0;  // 32'hf275ef0c;
    ram_cell[    8297] = 32'h0;  // 32'h65c135e0;
    ram_cell[    8298] = 32'h0;  // 32'h187a2dea;
    ram_cell[    8299] = 32'h0;  // 32'h6257e01d;
    ram_cell[    8300] = 32'h0;  // 32'h8c243c8c;
    ram_cell[    8301] = 32'h0;  // 32'h2fdec5e8;
    ram_cell[    8302] = 32'h0;  // 32'h11d75a21;
    ram_cell[    8303] = 32'h0;  // 32'h7bb1586e;
    ram_cell[    8304] = 32'h0;  // 32'h1a1a71c7;
    ram_cell[    8305] = 32'h0;  // 32'h361bea84;
    ram_cell[    8306] = 32'h0;  // 32'h321f0ea7;
    ram_cell[    8307] = 32'h0;  // 32'hdfa7e7f1;
    ram_cell[    8308] = 32'h0;  // 32'hd9d61fc9;
    ram_cell[    8309] = 32'h0;  // 32'he616282a;
    ram_cell[    8310] = 32'h0;  // 32'h9a54c796;
    ram_cell[    8311] = 32'h0;  // 32'h3bf19f8a;
    ram_cell[    8312] = 32'h0;  // 32'hd3f621a3;
    ram_cell[    8313] = 32'h0;  // 32'h63351855;
    ram_cell[    8314] = 32'h0;  // 32'hba0ee28d;
    ram_cell[    8315] = 32'h0;  // 32'h82d1dfa3;
    ram_cell[    8316] = 32'h0;  // 32'hb54e5911;
    ram_cell[    8317] = 32'h0;  // 32'hc2ca2a94;
    ram_cell[    8318] = 32'h0;  // 32'h1c1a64bf;
    ram_cell[    8319] = 32'h0;  // 32'h9d385d88;
    ram_cell[    8320] = 32'h0;  // 32'h5d8d9c3a;
    ram_cell[    8321] = 32'h0;  // 32'h5c896243;
    ram_cell[    8322] = 32'h0;  // 32'h0283a8c6;
    ram_cell[    8323] = 32'h0;  // 32'h0f125d83;
    ram_cell[    8324] = 32'h0;  // 32'h948d455b;
    ram_cell[    8325] = 32'h0;  // 32'h53ed5b58;
    ram_cell[    8326] = 32'h0;  // 32'hbca321cc;
    ram_cell[    8327] = 32'h0;  // 32'h004cfac6;
    ram_cell[    8328] = 32'h0;  // 32'hdf25e018;
    ram_cell[    8329] = 32'h0;  // 32'hf731643d;
    ram_cell[    8330] = 32'h0;  // 32'h2caf3000;
    ram_cell[    8331] = 32'h0;  // 32'h96fb9da2;
    ram_cell[    8332] = 32'h0;  // 32'h5126146b;
    ram_cell[    8333] = 32'h0;  // 32'h5eb77dd2;
    ram_cell[    8334] = 32'h0;  // 32'h9a7b4ebc;
    ram_cell[    8335] = 32'h0;  // 32'h96ead57e;
    ram_cell[    8336] = 32'h0;  // 32'hcd945c9a;
    ram_cell[    8337] = 32'h0;  // 32'h80cf4452;
    ram_cell[    8338] = 32'h0;  // 32'heb0fa9c8;
    ram_cell[    8339] = 32'h0;  // 32'h5c0ec044;
    ram_cell[    8340] = 32'h0;  // 32'ha74f831b;
    ram_cell[    8341] = 32'h0;  // 32'hfe536160;
    ram_cell[    8342] = 32'h0;  // 32'haac136c2;
    ram_cell[    8343] = 32'h0;  // 32'h4acdc959;
    ram_cell[    8344] = 32'h0;  // 32'h4eb47aa6;
    ram_cell[    8345] = 32'h0;  // 32'h40c4cb26;
    ram_cell[    8346] = 32'h0;  // 32'h14ce5232;
    ram_cell[    8347] = 32'h0;  // 32'h4a834dd6;
    ram_cell[    8348] = 32'h0;  // 32'h0dabf3af;
    ram_cell[    8349] = 32'h0;  // 32'h2dd10911;
    ram_cell[    8350] = 32'h0;  // 32'h956d6e06;
    ram_cell[    8351] = 32'h0;  // 32'he0f8f397;
    ram_cell[    8352] = 32'h0;  // 32'h10bbbd83;
    ram_cell[    8353] = 32'h0;  // 32'ha3ede77c;
    ram_cell[    8354] = 32'h0;  // 32'he53d65c2;
    ram_cell[    8355] = 32'h0;  // 32'hfff5b5c1;
    ram_cell[    8356] = 32'h0;  // 32'he56ccc6c;
    ram_cell[    8357] = 32'h0;  // 32'h09e66df0;
    ram_cell[    8358] = 32'h0;  // 32'h5ccd2df2;
    ram_cell[    8359] = 32'h0;  // 32'h70b133b9;
    ram_cell[    8360] = 32'h0;  // 32'ha732b08a;
    ram_cell[    8361] = 32'h0;  // 32'hfcadb19b;
    ram_cell[    8362] = 32'h0;  // 32'hde0cf45c;
    ram_cell[    8363] = 32'h0;  // 32'h6e4e9e9a;
    ram_cell[    8364] = 32'h0;  // 32'hd3ac76f5;
    ram_cell[    8365] = 32'h0;  // 32'hd5d0288c;
    ram_cell[    8366] = 32'h0;  // 32'hba30f4a4;
    ram_cell[    8367] = 32'h0;  // 32'h7a63a25e;
    ram_cell[    8368] = 32'h0;  // 32'hcac32e1a;
    ram_cell[    8369] = 32'h0;  // 32'hbb64ee7e;
    ram_cell[    8370] = 32'h0;  // 32'h5d0443a1;
    ram_cell[    8371] = 32'h0;  // 32'h53a9b5be;
    ram_cell[    8372] = 32'h0;  // 32'h07f4a7f7;
    ram_cell[    8373] = 32'h0;  // 32'h7430f4ee;
    ram_cell[    8374] = 32'h0;  // 32'h156c1388;
    ram_cell[    8375] = 32'h0;  // 32'hab12515e;
    ram_cell[    8376] = 32'h0;  // 32'h2e075bdc;
    ram_cell[    8377] = 32'h0;  // 32'hc528ab4e;
    ram_cell[    8378] = 32'h0;  // 32'h23baabc7;
    ram_cell[    8379] = 32'h0;  // 32'h99fc0d95;
    ram_cell[    8380] = 32'h0;  // 32'hb3446598;
    ram_cell[    8381] = 32'h0;  // 32'hff0450aa;
    ram_cell[    8382] = 32'h0;  // 32'h709f1d73;
    ram_cell[    8383] = 32'h0;  // 32'he998aa5d;
    ram_cell[    8384] = 32'h0;  // 32'h4a1013d4;
    ram_cell[    8385] = 32'h0;  // 32'hd07399e6;
    ram_cell[    8386] = 32'h0;  // 32'h3f13ce0b;
    ram_cell[    8387] = 32'h0;  // 32'h5369c68d;
    ram_cell[    8388] = 32'h0;  // 32'h561182d6;
    ram_cell[    8389] = 32'h0;  // 32'hc161bb88;
    ram_cell[    8390] = 32'h0;  // 32'hbad4aa33;
    ram_cell[    8391] = 32'h0;  // 32'h48a4aa2e;
    ram_cell[    8392] = 32'h0;  // 32'h327a2b7d;
    ram_cell[    8393] = 32'h0;  // 32'h84c80d98;
    ram_cell[    8394] = 32'h0;  // 32'h3084cb1f;
    ram_cell[    8395] = 32'h0;  // 32'h23f24626;
    ram_cell[    8396] = 32'h0;  // 32'h71df9f4e;
    ram_cell[    8397] = 32'h0;  // 32'h372e2663;
    ram_cell[    8398] = 32'h0;  // 32'hf1cd1bb5;
    ram_cell[    8399] = 32'h0;  // 32'h7e663bfb;
    ram_cell[    8400] = 32'h0;  // 32'h0255ed65;
    ram_cell[    8401] = 32'h0;  // 32'h425828a3;
    ram_cell[    8402] = 32'h0;  // 32'hf97dd115;
    ram_cell[    8403] = 32'h0;  // 32'hbb67e5e5;
    ram_cell[    8404] = 32'h0;  // 32'hadfc2389;
    ram_cell[    8405] = 32'h0;  // 32'h42403660;
    ram_cell[    8406] = 32'h0;  // 32'h7d2f9cd7;
    ram_cell[    8407] = 32'h0;  // 32'h3f32e85c;
    ram_cell[    8408] = 32'h0;  // 32'h601c10e8;
    ram_cell[    8409] = 32'h0;  // 32'hc94b34aa;
    ram_cell[    8410] = 32'h0;  // 32'h69680f3d;
    ram_cell[    8411] = 32'h0;  // 32'h3fa5a1df;
    ram_cell[    8412] = 32'h0;  // 32'h11a68454;
    ram_cell[    8413] = 32'h0;  // 32'h28115df9;
    ram_cell[    8414] = 32'h0;  // 32'h093b2cc9;
    ram_cell[    8415] = 32'h0;  // 32'h55682867;
    ram_cell[    8416] = 32'h0;  // 32'hf2c21b0d;
    ram_cell[    8417] = 32'h0;  // 32'hbcebaaf8;
    ram_cell[    8418] = 32'h0;  // 32'hb13646ca;
    ram_cell[    8419] = 32'h0;  // 32'h3529c2fa;
    ram_cell[    8420] = 32'h0;  // 32'he5f5286a;
    ram_cell[    8421] = 32'h0;  // 32'hea382e2f;
    ram_cell[    8422] = 32'h0;  // 32'hd99e4995;
    ram_cell[    8423] = 32'h0;  // 32'hb0d04fbf;
    ram_cell[    8424] = 32'h0;  // 32'h804adaec;
    ram_cell[    8425] = 32'h0;  // 32'hdfe2977c;
    ram_cell[    8426] = 32'h0;  // 32'h8cf4a118;
    ram_cell[    8427] = 32'h0;  // 32'h7ea2b518;
    ram_cell[    8428] = 32'h0;  // 32'h242ac68a;
    ram_cell[    8429] = 32'h0;  // 32'h2a196bda;
    ram_cell[    8430] = 32'h0;  // 32'ha8b657ad;
    ram_cell[    8431] = 32'h0;  // 32'h9c05650f;
    ram_cell[    8432] = 32'h0;  // 32'h87817ef1;
    ram_cell[    8433] = 32'h0;  // 32'hf4d27e9b;
    ram_cell[    8434] = 32'h0;  // 32'hb772f755;
    ram_cell[    8435] = 32'h0;  // 32'h942d7908;
    ram_cell[    8436] = 32'h0;  // 32'hdc578598;
    ram_cell[    8437] = 32'h0;  // 32'hda496f32;
    ram_cell[    8438] = 32'h0;  // 32'h90f70c38;
    ram_cell[    8439] = 32'h0;  // 32'h156de00f;
    ram_cell[    8440] = 32'h0;  // 32'h7dc98438;
    ram_cell[    8441] = 32'h0;  // 32'h25674c1c;
    ram_cell[    8442] = 32'h0;  // 32'hc6e5b4ad;
    ram_cell[    8443] = 32'h0;  // 32'hef98e052;
    ram_cell[    8444] = 32'h0;  // 32'hbfdadb51;
    ram_cell[    8445] = 32'h0;  // 32'h83d26c20;
    ram_cell[    8446] = 32'h0;  // 32'h5cb04180;
    ram_cell[    8447] = 32'h0;  // 32'hb146d345;
    ram_cell[    8448] = 32'h0;  // 32'h3f35b486;
    ram_cell[    8449] = 32'h0;  // 32'hfcf2944e;
    ram_cell[    8450] = 32'h0;  // 32'ha8bcf339;
    ram_cell[    8451] = 32'h0;  // 32'h89f26fd9;
    ram_cell[    8452] = 32'h0;  // 32'h68c97183;
    ram_cell[    8453] = 32'h0;  // 32'h9c055021;
    ram_cell[    8454] = 32'h0;  // 32'ha804c1fe;
    ram_cell[    8455] = 32'h0;  // 32'h2d7bd2d1;
    ram_cell[    8456] = 32'h0;  // 32'hcaa2ab17;
    ram_cell[    8457] = 32'h0;  // 32'he34cee0a;
    ram_cell[    8458] = 32'h0;  // 32'h54eb74bf;
    ram_cell[    8459] = 32'h0;  // 32'h91850d5b;
    ram_cell[    8460] = 32'h0;  // 32'hf936d57e;
    ram_cell[    8461] = 32'h0;  // 32'hcd495f36;
    ram_cell[    8462] = 32'h0;  // 32'hdee607fa;
    ram_cell[    8463] = 32'h0;  // 32'hc476b92a;
    ram_cell[    8464] = 32'h0;  // 32'h35a804c5;
    ram_cell[    8465] = 32'h0;  // 32'h23d6a15c;
    ram_cell[    8466] = 32'h0;  // 32'h8f735daf;
    ram_cell[    8467] = 32'h0;  // 32'hf1fddb0f;
    ram_cell[    8468] = 32'h0;  // 32'h6e6a8ddc;
    ram_cell[    8469] = 32'h0;  // 32'h213d848f;
    ram_cell[    8470] = 32'h0;  // 32'h2de41bc3;
    ram_cell[    8471] = 32'h0;  // 32'h391bf491;
    ram_cell[    8472] = 32'h0;  // 32'hcd912208;
    ram_cell[    8473] = 32'h0;  // 32'hb32151f0;
    ram_cell[    8474] = 32'h0;  // 32'hf4b9db31;
    ram_cell[    8475] = 32'h0;  // 32'hc89bc3f1;
    ram_cell[    8476] = 32'h0;  // 32'h58683597;
    ram_cell[    8477] = 32'h0;  // 32'ha5972f2a;
    ram_cell[    8478] = 32'h0;  // 32'h932d0d52;
    ram_cell[    8479] = 32'h0;  // 32'hcd2af721;
    ram_cell[    8480] = 32'h0;  // 32'h7e403f0d;
    ram_cell[    8481] = 32'h0;  // 32'h316b9244;
    ram_cell[    8482] = 32'h0;  // 32'h7a60dc33;
    ram_cell[    8483] = 32'h0;  // 32'h6efd4d68;
    ram_cell[    8484] = 32'h0;  // 32'h5407a7ee;
    ram_cell[    8485] = 32'h0;  // 32'h4e63823d;
    ram_cell[    8486] = 32'h0;  // 32'h15b4b9fb;
    ram_cell[    8487] = 32'h0;  // 32'h361fa8e7;
    ram_cell[    8488] = 32'h0;  // 32'hf041f256;
    ram_cell[    8489] = 32'h0;  // 32'ha56196e5;
    ram_cell[    8490] = 32'h0;  // 32'h029f9900;
    ram_cell[    8491] = 32'h0;  // 32'hf24f578f;
    ram_cell[    8492] = 32'h0;  // 32'hcf013207;
    ram_cell[    8493] = 32'h0;  // 32'h0de9f49f;
    ram_cell[    8494] = 32'h0;  // 32'hbd40f92c;
    ram_cell[    8495] = 32'h0;  // 32'ha39cb16b;
    ram_cell[    8496] = 32'h0;  // 32'he3b65033;
    ram_cell[    8497] = 32'h0;  // 32'hc58cbef8;
    ram_cell[    8498] = 32'h0;  // 32'h820975b7;
    ram_cell[    8499] = 32'h0;  // 32'hc86cd423;
    ram_cell[    8500] = 32'h0;  // 32'hd6f844f5;
    ram_cell[    8501] = 32'h0;  // 32'h49ac035e;
    ram_cell[    8502] = 32'h0;  // 32'h185e2237;
    ram_cell[    8503] = 32'h0;  // 32'hdacd8774;
    ram_cell[    8504] = 32'h0;  // 32'hf576459b;
    ram_cell[    8505] = 32'h0;  // 32'h4ff2a489;
    ram_cell[    8506] = 32'h0;  // 32'h92dbd60b;
    ram_cell[    8507] = 32'h0;  // 32'hc169c270;
    ram_cell[    8508] = 32'h0;  // 32'h3fa6188d;
    ram_cell[    8509] = 32'h0;  // 32'he71ef71c;
    ram_cell[    8510] = 32'h0;  // 32'h9f3e41d7;
    ram_cell[    8511] = 32'h0;  // 32'heb7144d0;
    ram_cell[    8512] = 32'h0;  // 32'h40208f2b;
    ram_cell[    8513] = 32'h0;  // 32'h9325e1f9;
    ram_cell[    8514] = 32'h0;  // 32'hce1a0145;
    ram_cell[    8515] = 32'h0;  // 32'h9af0f244;
    ram_cell[    8516] = 32'h0;  // 32'h7d35f2b9;
    ram_cell[    8517] = 32'h0;  // 32'hcbe14163;
    ram_cell[    8518] = 32'h0;  // 32'h47fe50d4;
    ram_cell[    8519] = 32'h0;  // 32'hf3698bd7;
    ram_cell[    8520] = 32'h0;  // 32'h09a924dc;
    ram_cell[    8521] = 32'h0;  // 32'h0c0d0c7d;
    ram_cell[    8522] = 32'h0;  // 32'h7a22e24b;
    ram_cell[    8523] = 32'h0;  // 32'he1f5f98a;
    ram_cell[    8524] = 32'h0;  // 32'hb6607ba0;
    ram_cell[    8525] = 32'h0;  // 32'h29cd0cd8;
    ram_cell[    8526] = 32'h0;  // 32'h9fd42188;
    ram_cell[    8527] = 32'h0;  // 32'h74a94d2c;
    ram_cell[    8528] = 32'h0;  // 32'h81bd502d;
    ram_cell[    8529] = 32'h0;  // 32'h7a0698e5;
    ram_cell[    8530] = 32'h0;  // 32'h171715b6;
    ram_cell[    8531] = 32'h0;  // 32'he8ad2afe;
    ram_cell[    8532] = 32'h0;  // 32'hc322c4a0;
    ram_cell[    8533] = 32'h0;  // 32'h6891a415;
    ram_cell[    8534] = 32'h0;  // 32'h78ee0391;
    ram_cell[    8535] = 32'h0;  // 32'hd6f63e18;
    ram_cell[    8536] = 32'h0;  // 32'h74eadaa1;
    ram_cell[    8537] = 32'h0;  // 32'h9eee64d3;
    ram_cell[    8538] = 32'h0;  // 32'h741af39f;
    ram_cell[    8539] = 32'h0;  // 32'hc5741faa;
    ram_cell[    8540] = 32'h0;  // 32'h1c2420e5;
    ram_cell[    8541] = 32'h0;  // 32'h74266373;
    ram_cell[    8542] = 32'h0;  // 32'hf01384c7;
    ram_cell[    8543] = 32'h0;  // 32'h201bc585;
    ram_cell[    8544] = 32'h0;  // 32'h7777bef7;
    ram_cell[    8545] = 32'h0;  // 32'h5cf7bf5f;
    ram_cell[    8546] = 32'h0;  // 32'hde4219b0;
    ram_cell[    8547] = 32'h0;  // 32'h1d382ce6;
    ram_cell[    8548] = 32'h0;  // 32'haf7ecf24;
    ram_cell[    8549] = 32'h0;  // 32'h63d3b2eb;
    ram_cell[    8550] = 32'h0;  // 32'h533e9d50;
    ram_cell[    8551] = 32'h0;  // 32'h0ea43d9a;
    ram_cell[    8552] = 32'h0;  // 32'h6930388f;
    ram_cell[    8553] = 32'h0;  // 32'h6e9545ee;
    ram_cell[    8554] = 32'h0;  // 32'hc295dbd0;
    ram_cell[    8555] = 32'h0;  // 32'h505cbc8f;
    ram_cell[    8556] = 32'h0;  // 32'h15680579;
    ram_cell[    8557] = 32'h0;  // 32'h357c59d4;
    ram_cell[    8558] = 32'h0;  // 32'hdb5d135b;
    ram_cell[    8559] = 32'h0;  // 32'h4f5332db;
    ram_cell[    8560] = 32'h0;  // 32'h8e656bad;
    ram_cell[    8561] = 32'h0;  // 32'h0ba9c304;
    ram_cell[    8562] = 32'h0;  // 32'hd1d6e40f;
    ram_cell[    8563] = 32'h0;  // 32'h31fccfe5;
    ram_cell[    8564] = 32'h0;  // 32'h53ce2eaa;
    ram_cell[    8565] = 32'h0;  // 32'h742fe9b5;
    ram_cell[    8566] = 32'h0;  // 32'h3d163046;
    ram_cell[    8567] = 32'h0;  // 32'h4df03815;
    ram_cell[    8568] = 32'h0;  // 32'h337b5dfe;
    ram_cell[    8569] = 32'h0;  // 32'h23006c0c;
    ram_cell[    8570] = 32'h0;  // 32'h32f9a30e;
    ram_cell[    8571] = 32'h0;  // 32'h33c7d7bd;
    ram_cell[    8572] = 32'h0;  // 32'h4fed4911;
    ram_cell[    8573] = 32'h0;  // 32'h6bf6daa1;
    ram_cell[    8574] = 32'h0;  // 32'h4bd97459;
    ram_cell[    8575] = 32'h0;  // 32'h7596df8a;
    ram_cell[    8576] = 32'h0;  // 32'h99f7e8ac;
    ram_cell[    8577] = 32'h0;  // 32'h34ea8d68;
    ram_cell[    8578] = 32'h0;  // 32'h9e233511;
    ram_cell[    8579] = 32'h0;  // 32'heef5506d;
    ram_cell[    8580] = 32'h0;  // 32'hd506896c;
    ram_cell[    8581] = 32'h0;  // 32'hf2f03f07;
    ram_cell[    8582] = 32'h0;  // 32'h52ca1e2f;
    ram_cell[    8583] = 32'h0;  // 32'h9927c2ea;
    ram_cell[    8584] = 32'h0;  // 32'h5a6ee8eb;
    ram_cell[    8585] = 32'h0;  // 32'hfd651df7;
    ram_cell[    8586] = 32'h0;  // 32'h67bcf923;
    ram_cell[    8587] = 32'h0;  // 32'h6118df55;
    ram_cell[    8588] = 32'h0;  // 32'hba89bcb8;
    ram_cell[    8589] = 32'h0;  // 32'h62c3bf59;
    ram_cell[    8590] = 32'h0;  // 32'h4377af29;
    ram_cell[    8591] = 32'h0;  // 32'hb988f7f7;
    ram_cell[    8592] = 32'h0;  // 32'h0b6cdb09;
    ram_cell[    8593] = 32'h0;  // 32'he4104ce6;
    ram_cell[    8594] = 32'h0;  // 32'he522f005;
    ram_cell[    8595] = 32'h0;  // 32'h86235ad8;
    ram_cell[    8596] = 32'h0;  // 32'h872a7e60;
    ram_cell[    8597] = 32'h0;  // 32'ha1042a75;
    ram_cell[    8598] = 32'h0;  // 32'hb83457af;
    ram_cell[    8599] = 32'h0;  // 32'hd58bb730;
    ram_cell[    8600] = 32'h0;  // 32'h0d3a15eb;
    ram_cell[    8601] = 32'h0;  // 32'h9872ea08;
    ram_cell[    8602] = 32'h0;  // 32'ha24f46cb;
    ram_cell[    8603] = 32'h0;  // 32'hc5df901c;
    ram_cell[    8604] = 32'h0;  // 32'h15dfd06c;
    ram_cell[    8605] = 32'h0;  // 32'hfe53016c;
    ram_cell[    8606] = 32'h0;  // 32'hecf48c93;
    ram_cell[    8607] = 32'h0;  // 32'he6ab60f6;
    ram_cell[    8608] = 32'h0;  // 32'h88709204;
    ram_cell[    8609] = 32'h0;  // 32'hd0896020;
    ram_cell[    8610] = 32'h0;  // 32'hf620a1dd;
    ram_cell[    8611] = 32'h0;  // 32'ha0def9f6;
    ram_cell[    8612] = 32'h0;  // 32'h8320203f;
    ram_cell[    8613] = 32'h0;  // 32'hfa5fa0d6;
    ram_cell[    8614] = 32'h0;  // 32'h4cb05ed5;
    ram_cell[    8615] = 32'h0;  // 32'hfacd3a17;
    ram_cell[    8616] = 32'h0;  // 32'hdabad46b;
    ram_cell[    8617] = 32'h0;  // 32'h76c3f555;
    ram_cell[    8618] = 32'h0;  // 32'he3a9ba40;
    ram_cell[    8619] = 32'h0;  // 32'h5f83875e;
    ram_cell[    8620] = 32'h0;  // 32'h09001f30;
    ram_cell[    8621] = 32'h0;  // 32'h207431a7;
    ram_cell[    8622] = 32'h0;  // 32'h3a182a48;
    ram_cell[    8623] = 32'h0;  // 32'hf9337986;
    ram_cell[    8624] = 32'h0;  // 32'hd6f6e3ac;
    ram_cell[    8625] = 32'h0;  // 32'h8d45e4b2;
    ram_cell[    8626] = 32'h0;  // 32'h55dfd9e5;
    ram_cell[    8627] = 32'h0;  // 32'hd9362313;
    ram_cell[    8628] = 32'h0;  // 32'h32972ee0;
    ram_cell[    8629] = 32'h0;  // 32'h9542cbdc;
    ram_cell[    8630] = 32'h0;  // 32'h36ffcc15;
    ram_cell[    8631] = 32'h0;  // 32'h2ea70975;
    ram_cell[    8632] = 32'h0;  // 32'h04178be8;
    ram_cell[    8633] = 32'h0;  // 32'h28ec6262;
    ram_cell[    8634] = 32'h0;  // 32'hf303f501;
    ram_cell[    8635] = 32'h0;  // 32'hc9d2ac99;
    ram_cell[    8636] = 32'h0;  // 32'h43365e51;
    ram_cell[    8637] = 32'h0;  // 32'h361a1df4;
    ram_cell[    8638] = 32'h0;  // 32'hd0e5a5b9;
    ram_cell[    8639] = 32'h0;  // 32'h576b0938;
    ram_cell[    8640] = 32'h0;  // 32'hb118298b;
    ram_cell[    8641] = 32'h0;  // 32'h60de52ab;
    ram_cell[    8642] = 32'h0;  // 32'h0ea6382f;
    ram_cell[    8643] = 32'h0;  // 32'hac7d4297;
    ram_cell[    8644] = 32'h0;  // 32'h61101e74;
    ram_cell[    8645] = 32'h0;  // 32'he869ad24;
    ram_cell[    8646] = 32'h0;  // 32'hd0194434;
    ram_cell[    8647] = 32'h0;  // 32'h9e7bcfc3;
    ram_cell[    8648] = 32'h0;  // 32'h5ca341fc;
    ram_cell[    8649] = 32'h0;  // 32'h28e6f354;
    ram_cell[    8650] = 32'h0;  // 32'he9f6fae5;
    ram_cell[    8651] = 32'h0;  // 32'h88664d48;
    ram_cell[    8652] = 32'h0;  // 32'h026e6dad;
    ram_cell[    8653] = 32'h0;  // 32'h00126048;
    ram_cell[    8654] = 32'h0;  // 32'h04ed1b11;
    ram_cell[    8655] = 32'h0;  // 32'hc78d90f1;
    ram_cell[    8656] = 32'h0;  // 32'hf30ed269;
    ram_cell[    8657] = 32'h0;  // 32'he71bd180;
    ram_cell[    8658] = 32'h0;  // 32'h768de29f;
    ram_cell[    8659] = 32'h0;  // 32'h2eaa547d;
    ram_cell[    8660] = 32'h0;  // 32'had8a0fc8;
    ram_cell[    8661] = 32'h0;  // 32'h1a39d134;
    ram_cell[    8662] = 32'h0;  // 32'ha777743d;
    ram_cell[    8663] = 32'h0;  // 32'h5bf2d870;
    ram_cell[    8664] = 32'h0;  // 32'h92f5beb9;
    ram_cell[    8665] = 32'h0;  // 32'h99791c7c;
    ram_cell[    8666] = 32'h0;  // 32'h7419862c;
    ram_cell[    8667] = 32'h0;  // 32'h48ab971d;
    ram_cell[    8668] = 32'h0;  // 32'h32596c6b;
    ram_cell[    8669] = 32'h0;  // 32'h8ee18d9f;
    ram_cell[    8670] = 32'h0;  // 32'h076207a5;
    ram_cell[    8671] = 32'h0;  // 32'hf14a3c85;
    ram_cell[    8672] = 32'h0;  // 32'hd4604066;
    ram_cell[    8673] = 32'h0;  // 32'h875f5a18;
    ram_cell[    8674] = 32'h0;  // 32'h620e4bea;
    ram_cell[    8675] = 32'h0;  // 32'hb78208c1;
    ram_cell[    8676] = 32'h0;  // 32'hdff8eaa8;
    ram_cell[    8677] = 32'h0;  // 32'hf5193157;
    ram_cell[    8678] = 32'h0;  // 32'h6d56a78b;
    ram_cell[    8679] = 32'h0;  // 32'h68d5a359;
    ram_cell[    8680] = 32'h0;  // 32'h93a5c083;
    ram_cell[    8681] = 32'h0;  // 32'h5c5e08dd;
    ram_cell[    8682] = 32'h0;  // 32'h70c8185c;
    ram_cell[    8683] = 32'h0;  // 32'h9facdded;
    ram_cell[    8684] = 32'h0;  // 32'hecf5a1e4;
    ram_cell[    8685] = 32'h0;  // 32'h152dd276;
    ram_cell[    8686] = 32'h0;  // 32'h868c264b;
    ram_cell[    8687] = 32'h0;  // 32'h68d733d1;
    ram_cell[    8688] = 32'h0;  // 32'h2e408e93;
    ram_cell[    8689] = 32'h0;  // 32'hdd4180a8;
    ram_cell[    8690] = 32'h0;  // 32'hcfe3ecad;
    ram_cell[    8691] = 32'h0;  // 32'hff7445a7;
    ram_cell[    8692] = 32'h0;  // 32'ha682bcf4;
    ram_cell[    8693] = 32'h0;  // 32'hf55b5a36;
    ram_cell[    8694] = 32'h0;  // 32'h35bea9e8;
    ram_cell[    8695] = 32'h0;  // 32'h6fcd77cd;
    ram_cell[    8696] = 32'h0;  // 32'h5d8e9d94;
    ram_cell[    8697] = 32'h0;  // 32'hf95dbd4a;
    ram_cell[    8698] = 32'h0;  // 32'h0943e895;
    ram_cell[    8699] = 32'h0;  // 32'hfda3798d;
    ram_cell[    8700] = 32'h0;  // 32'h1bfb973c;
    ram_cell[    8701] = 32'h0;  // 32'he03be9ab;
    ram_cell[    8702] = 32'h0;  // 32'hfd5275c0;
    ram_cell[    8703] = 32'h0;  // 32'h5542d46e;
    ram_cell[    8704] = 32'h0;  // 32'hdeb6dd66;
    ram_cell[    8705] = 32'h0;  // 32'h373712db;
    ram_cell[    8706] = 32'h0;  // 32'hecc8bfb0;
    ram_cell[    8707] = 32'h0;  // 32'he96dd6dc;
    ram_cell[    8708] = 32'h0;  // 32'h9e16d6d3;
    ram_cell[    8709] = 32'h0;  // 32'h70bb49a0;
    ram_cell[    8710] = 32'h0;  // 32'h3e02dd65;
    ram_cell[    8711] = 32'h0;  // 32'h58f53a6d;
    ram_cell[    8712] = 32'h0;  // 32'h2a02960c;
    ram_cell[    8713] = 32'h0;  // 32'h2dd57efe;
    ram_cell[    8714] = 32'h0;  // 32'h919fb798;
    ram_cell[    8715] = 32'h0;  // 32'hbca48277;
    ram_cell[    8716] = 32'h0;  // 32'h663135e2;
    ram_cell[    8717] = 32'h0;  // 32'h59f3795d;
    ram_cell[    8718] = 32'h0;  // 32'h96279719;
    ram_cell[    8719] = 32'h0;  // 32'h5e320e82;
    ram_cell[    8720] = 32'h0;  // 32'hba615874;
    ram_cell[    8721] = 32'h0;  // 32'h211df739;
    ram_cell[    8722] = 32'h0;  // 32'hf1dc8da5;
    ram_cell[    8723] = 32'h0;  // 32'he68e86e8;
    ram_cell[    8724] = 32'h0;  // 32'hc524b466;
    ram_cell[    8725] = 32'h0;  // 32'h8ce07c7a;
    ram_cell[    8726] = 32'h0;  // 32'h646a7a5a;
    ram_cell[    8727] = 32'h0;  // 32'hea53c3b7;
    ram_cell[    8728] = 32'h0;  // 32'ha3492605;
    ram_cell[    8729] = 32'h0;  // 32'h476117d4;
    ram_cell[    8730] = 32'h0;  // 32'hba47cb59;
    ram_cell[    8731] = 32'h0;  // 32'hd4b33dc8;
    ram_cell[    8732] = 32'h0;  // 32'h812d3e22;
    ram_cell[    8733] = 32'h0;  // 32'h4e2ba986;
    ram_cell[    8734] = 32'h0;  // 32'hecc5c3c5;
    ram_cell[    8735] = 32'h0;  // 32'he674eb74;
    ram_cell[    8736] = 32'h0;  // 32'h267045ca;
    ram_cell[    8737] = 32'h0;  // 32'ha4b478e7;
    ram_cell[    8738] = 32'h0;  // 32'hf312e224;
    ram_cell[    8739] = 32'h0;  // 32'h0b67d5a2;
    ram_cell[    8740] = 32'h0;  // 32'h01960a09;
    ram_cell[    8741] = 32'h0;  // 32'hdc4e6680;
    ram_cell[    8742] = 32'h0;  // 32'hd3c7acea;
    ram_cell[    8743] = 32'h0;  // 32'haf27a902;
    ram_cell[    8744] = 32'h0;  // 32'h580da126;
    ram_cell[    8745] = 32'h0;  // 32'h555324b6;
    ram_cell[    8746] = 32'h0;  // 32'h71a1155c;
    ram_cell[    8747] = 32'h0;  // 32'hc5257739;
    ram_cell[    8748] = 32'h0;  // 32'hcdc27a8e;
    ram_cell[    8749] = 32'h0;  // 32'h530af351;
    ram_cell[    8750] = 32'h0;  // 32'h17be80ff;
    ram_cell[    8751] = 32'h0;  // 32'hfd13a8c8;
    ram_cell[    8752] = 32'h0;  // 32'ha11bcbe8;
    ram_cell[    8753] = 32'h0;  // 32'h9a9e944b;
    ram_cell[    8754] = 32'h0;  // 32'hdddf259f;
    ram_cell[    8755] = 32'h0;  // 32'h180f2a3f;
    ram_cell[    8756] = 32'h0;  // 32'h25f9dc62;
    ram_cell[    8757] = 32'h0;  // 32'h875bcfa2;
    ram_cell[    8758] = 32'h0;  // 32'h69eb3dfd;
    ram_cell[    8759] = 32'h0;  // 32'hb06ed7f5;
    ram_cell[    8760] = 32'h0;  // 32'hf2641aae;
    ram_cell[    8761] = 32'h0;  // 32'hf198013e;
    ram_cell[    8762] = 32'h0;  // 32'h026e9594;
    ram_cell[    8763] = 32'h0;  // 32'h5f3a7f41;
    ram_cell[    8764] = 32'h0;  // 32'h6471aaa8;
    ram_cell[    8765] = 32'h0;  // 32'heb97f530;
    ram_cell[    8766] = 32'h0;  // 32'h29507f09;
    ram_cell[    8767] = 32'h0;  // 32'he6c30e92;
    ram_cell[    8768] = 32'h0;  // 32'h362c154d;
    ram_cell[    8769] = 32'h0;  // 32'hc89d831c;
    ram_cell[    8770] = 32'h0;  // 32'hef1008b3;
    ram_cell[    8771] = 32'h0;  // 32'hc0934768;
    ram_cell[    8772] = 32'h0;  // 32'h1c533425;
    ram_cell[    8773] = 32'h0;  // 32'h7351a808;
    ram_cell[    8774] = 32'h0;  // 32'h9d5e38c8;
    ram_cell[    8775] = 32'h0;  // 32'h3ad5c5c1;
    ram_cell[    8776] = 32'h0;  // 32'h98bdf79f;
    ram_cell[    8777] = 32'h0;  // 32'h61defead;
    ram_cell[    8778] = 32'h0;  // 32'h07e29dbe;
    ram_cell[    8779] = 32'h0;  // 32'h9a4dcb85;
    ram_cell[    8780] = 32'h0;  // 32'hc4a7b030;
    ram_cell[    8781] = 32'h0;  // 32'h32791572;
    ram_cell[    8782] = 32'h0;  // 32'h228216ef;
    ram_cell[    8783] = 32'h0;  // 32'he07734dd;
    ram_cell[    8784] = 32'h0;  // 32'hb3690745;
    ram_cell[    8785] = 32'h0;  // 32'hcb14e6bd;
    ram_cell[    8786] = 32'h0;  // 32'h856714b3;
    ram_cell[    8787] = 32'h0;  // 32'h0278e84f;
    ram_cell[    8788] = 32'h0;  // 32'hd0b9f482;
    ram_cell[    8789] = 32'h0;  // 32'h4989a875;
    ram_cell[    8790] = 32'h0;  // 32'haf5af0ed;
    ram_cell[    8791] = 32'h0;  // 32'h7608f2ab;
    ram_cell[    8792] = 32'h0;  // 32'h22b97a26;
    ram_cell[    8793] = 32'h0;  // 32'h8229d36b;
    ram_cell[    8794] = 32'h0;  // 32'hc559b34d;
    ram_cell[    8795] = 32'h0;  // 32'h943ff78a;
    ram_cell[    8796] = 32'h0;  // 32'ha13ab8b9;
    ram_cell[    8797] = 32'h0;  // 32'h59ee1938;
    ram_cell[    8798] = 32'h0;  // 32'h40bb94c8;
    ram_cell[    8799] = 32'h0;  // 32'h398047ef;
    ram_cell[    8800] = 32'h0;  // 32'h5eae6174;
    ram_cell[    8801] = 32'h0;  // 32'h8b8794bb;
    ram_cell[    8802] = 32'h0;  // 32'h5607efee;
    ram_cell[    8803] = 32'h0;  // 32'hec1ad8b4;
    ram_cell[    8804] = 32'h0;  // 32'h3f87bc78;
    ram_cell[    8805] = 32'h0;  // 32'h9da178f2;
    ram_cell[    8806] = 32'h0;  // 32'hcef1230f;
    ram_cell[    8807] = 32'h0;  // 32'h68f959f0;
    ram_cell[    8808] = 32'h0;  // 32'h9a8fd5f6;
    ram_cell[    8809] = 32'h0;  // 32'hdf739326;
    ram_cell[    8810] = 32'h0;  // 32'he7aa732c;
    ram_cell[    8811] = 32'h0;  // 32'h4a0ad712;
    ram_cell[    8812] = 32'h0;  // 32'h0e62f429;
    ram_cell[    8813] = 32'h0;  // 32'he22c6bb1;
    ram_cell[    8814] = 32'h0;  // 32'h66c734d2;
    ram_cell[    8815] = 32'h0;  // 32'h2937f92b;
    ram_cell[    8816] = 32'h0;  // 32'h70c35bc6;
    ram_cell[    8817] = 32'h0;  // 32'h2c6b271e;
    ram_cell[    8818] = 32'h0;  // 32'h70bae390;
    ram_cell[    8819] = 32'h0;  // 32'heb874ed0;
    ram_cell[    8820] = 32'h0;  // 32'h64d07b53;
    ram_cell[    8821] = 32'h0;  // 32'h23b1be6c;
    ram_cell[    8822] = 32'h0;  // 32'hb065a8c0;
    ram_cell[    8823] = 32'h0;  // 32'h5b54bbb6;
    ram_cell[    8824] = 32'h0;  // 32'h34fe9294;
    ram_cell[    8825] = 32'h0;  // 32'h9fe7a60e;
    ram_cell[    8826] = 32'h0;  // 32'h72b78997;
    ram_cell[    8827] = 32'h0;  // 32'h297ec9b4;
    ram_cell[    8828] = 32'h0;  // 32'h9c9140d4;
    ram_cell[    8829] = 32'h0;  // 32'h3058cd6f;
    ram_cell[    8830] = 32'h0;  // 32'h31a55816;
    ram_cell[    8831] = 32'h0;  // 32'hd3fe437f;
    ram_cell[    8832] = 32'h0;  // 32'h548b0fbb;
    ram_cell[    8833] = 32'h0;  // 32'h35389c93;
    ram_cell[    8834] = 32'h0;  // 32'hb84171d1;
    ram_cell[    8835] = 32'h0;  // 32'h6df6b69c;
    ram_cell[    8836] = 32'h0;  // 32'h0a6b5d04;
    ram_cell[    8837] = 32'h0;  // 32'hd3af925b;
    ram_cell[    8838] = 32'h0;  // 32'h7246f413;
    ram_cell[    8839] = 32'h0;  // 32'h293c7659;
    ram_cell[    8840] = 32'h0;  // 32'h2c4d8b18;
    ram_cell[    8841] = 32'h0;  // 32'ha354b322;
    ram_cell[    8842] = 32'h0;  // 32'hc8760c7a;
    ram_cell[    8843] = 32'h0;  // 32'he0fef332;
    ram_cell[    8844] = 32'h0;  // 32'h9cbec6e2;
    ram_cell[    8845] = 32'h0;  // 32'h4fea5e18;
    ram_cell[    8846] = 32'h0;  // 32'hbbe63955;
    ram_cell[    8847] = 32'h0;  // 32'h2835b857;
    ram_cell[    8848] = 32'h0;  // 32'h319e595a;
    ram_cell[    8849] = 32'h0;  // 32'h65376464;
    ram_cell[    8850] = 32'h0;  // 32'h265d535c;
    ram_cell[    8851] = 32'h0;  // 32'hc266e517;
    ram_cell[    8852] = 32'h0;  // 32'h9765eb00;
    ram_cell[    8853] = 32'h0;  // 32'h406c5d30;
    ram_cell[    8854] = 32'h0;  // 32'h72b9a2fe;
    ram_cell[    8855] = 32'h0;  // 32'h2571b95c;
    ram_cell[    8856] = 32'h0;  // 32'h5efd00cf;
    ram_cell[    8857] = 32'h0;  // 32'h8f50ad59;
    ram_cell[    8858] = 32'h0;  // 32'h7acaec84;
    ram_cell[    8859] = 32'h0;  // 32'h780d80e1;
    ram_cell[    8860] = 32'h0;  // 32'h1f6556df;
    ram_cell[    8861] = 32'h0;  // 32'hf6b66414;
    ram_cell[    8862] = 32'h0;  // 32'hf6221ac7;
    ram_cell[    8863] = 32'h0;  // 32'h46f67cd5;
    ram_cell[    8864] = 32'h0;  // 32'h870e7589;
    ram_cell[    8865] = 32'h0;  // 32'hf33eab0e;
    ram_cell[    8866] = 32'h0;  // 32'he63edd4d;
    ram_cell[    8867] = 32'h0;  // 32'h1e8316fe;
    ram_cell[    8868] = 32'h0;  // 32'h5672e4b6;
    ram_cell[    8869] = 32'h0;  // 32'h4b08cb18;
    ram_cell[    8870] = 32'h0;  // 32'h8511608b;
    ram_cell[    8871] = 32'h0;  // 32'h124a5851;
    ram_cell[    8872] = 32'h0;  // 32'hcd9479f8;
    ram_cell[    8873] = 32'h0;  // 32'h76030130;
    ram_cell[    8874] = 32'h0;  // 32'hbedfb4d4;
    ram_cell[    8875] = 32'h0;  // 32'hd136e420;
    ram_cell[    8876] = 32'h0;  // 32'h67daaeea;
    ram_cell[    8877] = 32'h0;  // 32'hecb55354;
    ram_cell[    8878] = 32'h0;  // 32'h75e204e0;
    ram_cell[    8879] = 32'h0;  // 32'h02414949;
    ram_cell[    8880] = 32'h0;  // 32'h72fe168c;
    ram_cell[    8881] = 32'h0;  // 32'h1ff6a68d;
    ram_cell[    8882] = 32'h0;  // 32'hce688d8a;
    ram_cell[    8883] = 32'h0;  // 32'h935ecb28;
    ram_cell[    8884] = 32'h0;  // 32'h831496d4;
    ram_cell[    8885] = 32'h0;  // 32'h5cc1f025;
    ram_cell[    8886] = 32'h0;  // 32'hc134a805;
    ram_cell[    8887] = 32'h0;  // 32'h4deb8e8e;
    ram_cell[    8888] = 32'h0;  // 32'h170e2d9a;
    ram_cell[    8889] = 32'h0;  // 32'h14bc720a;
    ram_cell[    8890] = 32'h0;  // 32'hc80fd4c4;
    ram_cell[    8891] = 32'h0;  // 32'hef363972;
    ram_cell[    8892] = 32'h0;  // 32'h6c9c9ccc;
    ram_cell[    8893] = 32'h0;  // 32'hd4f11aab;
    ram_cell[    8894] = 32'h0;  // 32'he9e52839;
    ram_cell[    8895] = 32'h0;  // 32'h406c194f;
    ram_cell[    8896] = 32'h0;  // 32'h433bd071;
    ram_cell[    8897] = 32'h0;  // 32'h80439488;
    ram_cell[    8898] = 32'h0;  // 32'h8a2f7593;
    ram_cell[    8899] = 32'h0;  // 32'h84dcb4ad;
    ram_cell[    8900] = 32'h0;  // 32'h5f041eed;
    ram_cell[    8901] = 32'h0;  // 32'h2a7518ce;
    ram_cell[    8902] = 32'h0;  // 32'hee023d9f;
    ram_cell[    8903] = 32'h0;  // 32'h8777bb84;
    ram_cell[    8904] = 32'h0;  // 32'h177d9562;
    ram_cell[    8905] = 32'h0;  // 32'h0ac34a26;
    ram_cell[    8906] = 32'h0;  // 32'h131a0ceb;
    ram_cell[    8907] = 32'h0;  // 32'h9ba368e5;
    ram_cell[    8908] = 32'h0;  // 32'h49798966;
    ram_cell[    8909] = 32'h0;  // 32'h3500542c;
    ram_cell[    8910] = 32'h0;  // 32'hbc6f33c8;
    ram_cell[    8911] = 32'h0;  // 32'h00eb37ea;
    ram_cell[    8912] = 32'h0;  // 32'h7319e2c5;
    ram_cell[    8913] = 32'h0;  // 32'h1b18114a;
    ram_cell[    8914] = 32'h0;  // 32'ha0e5fd21;
    ram_cell[    8915] = 32'h0;  // 32'hb5222628;
    ram_cell[    8916] = 32'h0;  // 32'h07f3b656;
    ram_cell[    8917] = 32'h0;  // 32'hc689b56d;
    ram_cell[    8918] = 32'h0;  // 32'h2e18af41;
    ram_cell[    8919] = 32'h0;  // 32'h44784128;
    ram_cell[    8920] = 32'h0;  // 32'h960f21a2;
    ram_cell[    8921] = 32'h0;  // 32'hf9d17749;
    ram_cell[    8922] = 32'h0;  // 32'h8a6a6fb0;
    ram_cell[    8923] = 32'h0;  // 32'hf6228fc6;
    ram_cell[    8924] = 32'h0;  // 32'h3fa7140e;
    ram_cell[    8925] = 32'h0;  // 32'hbc3b236d;
    ram_cell[    8926] = 32'h0;  // 32'h5d81c249;
    ram_cell[    8927] = 32'h0;  // 32'hfb38cd77;
    ram_cell[    8928] = 32'h0;  // 32'hb04b3d24;
    ram_cell[    8929] = 32'h0;  // 32'h4a635498;
    ram_cell[    8930] = 32'h0;  // 32'hc1884e01;
    ram_cell[    8931] = 32'h0;  // 32'h61e3886f;
    ram_cell[    8932] = 32'h0;  // 32'hab4b51cd;
    ram_cell[    8933] = 32'h0;  // 32'ha997e551;
    ram_cell[    8934] = 32'h0;  // 32'h910d554a;
    ram_cell[    8935] = 32'h0;  // 32'h1f077f46;
    ram_cell[    8936] = 32'h0;  // 32'h091109e0;
    ram_cell[    8937] = 32'h0;  // 32'h1d629ee3;
    ram_cell[    8938] = 32'h0;  // 32'h98ae0e64;
    ram_cell[    8939] = 32'h0;  // 32'hf0a817df;
    ram_cell[    8940] = 32'h0;  // 32'h87378bc5;
    ram_cell[    8941] = 32'h0;  // 32'h9f88c33c;
    ram_cell[    8942] = 32'h0;  // 32'h806e3590;
    ram_cell[    8943] = 32'h0;  // 32'h8e04fa0d;
    ram_cell[    8944] = 32'h0;  // 32'h6cb485c8;
    ram_cell[    8945] = 32'h0;  // 32'hbb525c02;
    ram_cell[    8946] = 32'h0;  // 32'hbb0cbe6e;
    ram_cell[    8947] = 32'h0;  // 32'hbde29154;
    ram_cell[    8948] = 32'h0;  // 32'h997139fe;
    ram_cell[    8949] = 32'h0;  // 32'h6f3df22d;
    ram_cell[    8950] = 32'h0;  // 32'hda01bade;
    ram_cell[    8951] = 32'h0;  // 32'hfd2fb307;
    ram_cell[    8952] = 32'h0;  // 32'hb74533f9;
    ram_cell[    8953] = 32'h0;  // 32'hc747703f;
    ram_cell[    8954] = 32'h0;  // 32'he927876f;
    ram_cell[    8955] = 32'h0;  // 32'h140df303;
    ram_cell[    8956] = 32'h0;  // 32'h7ec07ff7;
    ram_cell[    8957] = 32'h0;  // 32'hac09732b;
    ram_cell[    8958] = 32'h0;  // 32'h65622c5a;
    ram_cell[    8959] = 32'h0;  // 32'h53291774;
    ram_cell[    8960] = 32'h0;  // 32'h0c1fdf9d;
    ram_cell[    8961] = 32'h0;  // 32'hd6e5be92;
    ram_cell[    8962] = 32'h0;  // 32'hf04287c4;
    ram_cell[    8963] = 32'h0;  // 32'hdcb9d500;
    ram_cell[    8964] = 32'h0;  // 32'h60d432c6;
    ram_cell[    8965] = 32'h0;  // 32'h06242256;
    ram_cell[    8966] = 32'h0;  // 32'h3ee19bc4;
    ram_cell[    8967] = 32'h0;  // 32'hc0e6a4ce;
    ram_cell[    8968] = 32'h0;  // 32'h45415559;
    ram_cell[    8969] = 32'h0;  // 32'h7b9674a7;
    ram_cell[    8970] = 32'h0;  // 32'h7f3de185;
    ram_cell[    8971] = 32'h0;  // 32'h568db241;
    ram_cell[    8972] = 32'h0;  // 32'h8d7338d5;
    ram_cell[    8973] = 32'h0;  // 32'h20251a3a;
    ram_cell[    8974] = 32'h0;  // 32'h1b78edd2;
    ram_cell[    8975] = 32'h0;  // 32'hb408fa5f;
    ram_cell[    8976] = 32'h0;  // 32'hbc0af66d;
    ram_cell[    8977] = 32'h0;  // 32'he5e378cb;
    ram_cell[    8978] = 32'h0;  // 32'h46487a7a;
    ram_cell[    8979] = 32'h0;  // 32'hfb4bb7a3;
    ram_cell[    8980] = 32'h0;  // 32'hc9d760d4;
    ram_cell[    8981] = 32'h0;  // 32'h8d51ca33;
    ram_cell[    8982] = 32'h0;  // 32'hc800e39c;
    ram_cell[    8983] = 32'h0;  // 32'h9e603800;
    ram_cell[    8984] = 32'h0;  // 32'h59e20548;
    ram_cell[    8985] = 32'h0;  // 32'ha0e19d4d;
    ram_cell[    8986] = 32'h0;  // 32'h3256e293;
    ram_cell[    8987] = 32'h0;  // 32'hb685a1b6;
    ram_cell[    8988] = 32'h0;  // 32'hddbe6a19;
    ram_cell[    8989] = 32'h0;  // 32'h55c1a846;
    ram_cell[    8990] = 32'h0;  // 32'hf33b5d2a;
    ram_cell[    8991] = 32'h0;  // 32'h0ba12070;
    ram_cell[    8992] = 32'h0;  // 32'h94802285;
    ram_cell[    8993] = 32'h0;  // 32'h034a729b;
    ram_cell[    8994] = 32'h0;  // 32'h77815321;
    ram_cell[    8995] = 32'h0;  // 32'h3d11963e;
    ram_cell[    8996] = 32'h0;  // 32'h778fac9c;
    ram_cell[    8997] = 32'h0;  // 32'h2721a5e2;
    ram_cell[    8998] = 32'h0;  // 32'h76c6dc9e;
    ram_cell[    8999] = 32'h0;  // 32'h3f553180;
    ram_cell[    9000] = 32'h0;  // 32'h7143bd85;
    ram_cell[    9001] = 32'h0;  // 32'h1b5c8229;
    ram_cell[    9002] = 32'h0;  // 32'hbf73a128;
    ram_cell[    9003] = 32'h0;  // 32'hc369837d;
    ram_cell[    9004] = 32'h0;  // 32'h61e360ce;
    ram_cell[    9005] = 32'h0;  // 32'hd1affe9e;
    ram_cell[    9006] = 32'h0;  // 32'hb34c2e50;
    ram_cell[    9007] = 32'h0;  // 32'hf820ad5a;
    ram_cell[    9008] = 32'h0;  // 32'h1b385283;
    ram_cell[    9009] = 32'h0;  // 32'h2664cf7c;
    ram_cell[    9010] = 32'h0;  // 32'hdd4b0ff4;
    ram_cell[    9011] = 32'h0;  // 32'h568ce673;
    ram_cell[    9012] = 32'h0;  // 32'h8db1bf00;
    ram_cell[    9013] = 32'h0;  // 32'h4b8f877b;
    ram_cell[    9014] = 32'h0;  // 32'hcebfaecc;
    ram_cell[    9015] = 32'h0;  // 32'h415f196c;
    ram_cell[    9016] = 32'h0;  // 32'h7142731f;
    ram_cell[    9017] = 32'h0;  // 32'h97b6aec1;
    ram_cell[    9018] = 32'h0;  // 32'hac9f5f0e;
    ram_cell[    9019] = 32'h0;  // 32'h073785d1;
    ram_cell[    9020] = 32'h0;  // 32'hf6cc1401;
    ram_cell[    9021] = 32'h0;  // 32'h6ffcc5e4;
    ram_cell[    9022] = 32'h0;  // 32'h57df03c7;
    ram_cell[    9023] = 32'h0;  // 32'h0be561a1;
    ram_cell[    9024] = 32'h0;  // 32'h678557d7;
    ram_cell[    9025] = 32'h0;  // 32'h2cdf9f54;
    ram_cell[    9026] = 32'h0;  // 32'h732a8e4e;
    ram_cell[    9027] = 32'h0;  // 32'h3bc47595;
    ram_cell[    9028] = 32'h0;  // 32'h4a863e0e;
    ram_cell[    9029] = 32'h0;  // 32'h88057d42;
    ram_cell[    9030] = 32'h0;  // 32'hcd85e76b;
    ram_cell[    9031] = 32'h0;  // 32'h68c0e0d2;
    ram_cell[    9032] = 32'h0;  // 32'hc371c1d6;
    ram_cell[    9033] = 32'h0;  // 32'h6ee9cc13;
    ram_cell[    9034] = 32'h0;  // 32'h78d379f7;
    ram_cell[    9035] = 32'h0;  // 32'h1e14f3c4;
    ram_cell[    9036] = 32'h0;  // 32'h87cf4f2e;
    ram_cell[    9037] = 32'h0;  // 32'h0af543e8;
    ram_cell[    9038] = 32'h0;  // 32'hc60d9c5a;
    ram_cell[    9039] = 32'h0;  // 32'hf325ad55;
    ram_cell[    9040] = 32'h0;  // 32'hf446e8f6;
    ram_cell[    9041] = 32'h0;  // 32'h4fcd4903;
    ram_cell[    9042] = 32'h0;  // 32'hd5da331f;
    ram_cell[    9043] = 32'h0;  // 32'h8d9c57c1;
    ram_cell[    9044] = 32'h0;  // 32'h4440576b;
    ram_cell[    9045] = 32'h0;  // 32'h4b7b8128;
    ram_cell[    9046] = 32'h0;  // 32'h590e189d;
    ram_cell[    9047] = 32'h0;  // 32'h20c79f20;
    ram_cell[    9048] = 32'h0;  // 32'hab7d60af;
    ram_cell[    9049] = 32'h0;  // 32'he65e3a2b;
    ram_cell[    9050] = 32'h0;  // 32'h60a55695;
    ram_cell[    9051] = 32'h0;  // 32'hf47acff9;
    ram_cell[    9052] = 32'h0;  // 32'h6d913f84;
    ram_cell[    9053] = 32'h0;  // 32'h272aaf0d;
    ram_cell[    9054] = 32'h0;  // 32'hbdebda85;
    ram_cell[    9055] = 32'h0;  // 32'hda78318a;
    ram_cell[    9056] = 32'h0;  // 32'h4cbe4f47;
    ram_cell[    9057] = 32'h0;  // 32'h4293f7a9;
    ram_cell[    9058] = 32'h0;  // 32'h896b6d81;
    ram_cell[    9059] = 32'h0;  // 32'h8be41254;
    ram_cell[    9060] = 32'h0;  // 32'hf1de9f66;
    ram_cell[    9061] = 32'h0;  // 32'h66b05f48;
    ram_cell[    9062] = 32'h0;  // 32'hcc3bdb16;
    ram_cell[    9063] = 32'h0;  // 32'h6eec7401;
    ram_cell[    9064] = 32'h0;  // 32'h344e7150;
    ram_cell[    9065] = 32'h0;  // 32'h5a3e6c3c;
    ram_cell[    9066] = 32'h0;  // 32'hf8b2f982;
    ram_cell[    9067] = 32'h0;  // 32'h681bc137;
    ram_cell[    9068] = 32'h0;  // 32'h8cbdae14;
    ram_cell[    9069] = 32'h0;  // 32'hae29ba74;
    ram_cell[    9070] = 32'h0;  // 32'ha8ffb3c6;
    ram_cell[    9071] = 32'h0;  // 32'h4aa0e2c7;
    ram_cell[    9072] = 32'h0;  // 32'h1e11413b;
    ram_cell[    9073] = 32'h0;  // 32'h9f79d5e4;
    ram_cell[    9074] = 32'h0;  // 32'ha6737186;
    ram_cell[    9075] = 32'h0;  // 32'h85f07311;
    ram_cell[    9076] = 32'h0;  // 32'h71cf8540;
    ram_cell[    9077] = 32'h0;  // 32'h75564fe0;
    ram_cell[    9078] = 32'h0;  // 32'h52dd665e;
    ram_cell[    9079] = 32'h0;  // 32'hfcf783f2;
    ram_cell[    9080] = 32'h0;  // 32'h632676f8;
    ram_cell[    9081] = 32'h0;  // 32'h26c1522c;
    ram_cell[    9082] = 32'h0;  // 32'h40131157;
    ram_cell[    9083] = 32'h0;  // 32'h0c7ed959;
    ram_cell[    9084] = 32'h0;  // 32'hc9f2e53d;
    ram_cell[    9085] = 32'h0;  // 32'head99e98;
    ram_cell[    9086] = 32'h0;  // 32'h24f13756;
    ram_cell[    9087] = 32'h0;  // 32'h97f29f03;
    ram_cell[    9088] = 32'h0;  // 32'h99c26927;
    ram_cell[    9089] = 32'h0;  // 32'h27d76056;
    ram_cell[    9090] = 32'h0;  // 32'he9b243c0;
    ram_cell[    9091] = 32'h0;  // 32'h199b66a6;
    ram_cell[    9092] = 32'h0;  // 32'h7d1b3f36;
    ram_cell[    9093] = 32'h0;  // 32'he245906a;
    ram_cell[    9094] = 32'h0;  // 32'ha31fc004;
    ram_cell[    9095] = 32'h0;  // 32'hb4273e55;
    ram_cell[    9096] = 32'h0;  // 32'hc69051ee;
    ram_cell[    9097] = 32'h0;  // 32'h2ecbbbc2;
    ram_cell[    9098] = 32'h0;  // 32'h5f2ff972;
    ram_cell[    9099] = 32'h0;  // 32'h10a474ad;
    ram_cell[    9100] = 32'h0;  // 32'h6bcc1c20;
    ram_cell[    9101] = 32'h0;  // 32'hf2d9f171;
    ram_cell[    9102] = 32'h0;  // 32'he108986c;
    ram_cell[    9103] = 32'h0;  // 32'he34b2f31;
    ram_cell[    9104] = 32'h0;  // 32'h21dd9f3a;
    ram_cell[    9105] = 32'h0;  // 32'h1fd3afe5;
    ram_cell[    9106] = 32'h0;  // 32'h0d5ef557;
    ram_cell[    9107] = 32'h0;  // 32'h5f75f181;
    ram_cell[    9108] = 32'h0;  // 32'he13201a5;
    ram_cell[    9109] = 32'h0;  // 32'hf18c3c15;
    ram_cell[    9110] = 32'h0;  // 32'hed233856;
    ram_cell[    9111] = 32'h0;  // 32'had006e81;
    ram_cell[    9112] = 32'h0;  // 32'hba29ec0a;
    ram_cell[    9113] = 32'h0;  // 32'h7d5336c9;
    ram_cell[    9114] = 32'h0;  // 32'hc1de9086;
    ram_cell[    9115] = 32'h0;  // 32'hcbc60f73;
    ram_cell[    9116] = 32'h0;  // 32'h3f1e42cc;
    ram_cell[    9117] = 32'h0;  // 32'h8ba645dc;
    ram_cell[    9118] = 32'h0;  // 32'had694b51;
    ram_cell[    9119] = 32'h0;  // 32'ha87c1b6b;
    ram_cell[    9120] = 32'h0;  // 32'ha049e752;
    ram_cell[    9121] = 32'h0;  // 32'h7fd24e0f;
    ram_cell[    9122] = 32'h0;  // 32'h281742a4;
    ram_cell[    9123] = 32'h0;  // 32'hf2c6ecf0;
    ram_cell[    9124] = 32'h0;  // 32'h3867160a;
    ram_cell[    9125] = 32'h0;  // 32'hc0b408db;
    ram_cell[    9126] = 32'h0;  // 32'hb06161ee;
    ram_cell[    9127] = 32'h0;  // 32'h1b6fc348;
    ram_cell[    9128] = 32'h0;  // 32'h49878f96;
    ram_cell[    9129] = 32'h0;  // 32'hcb6a8264;
    ram_cell[    9130] = 32'h0;  // 32'h7c2ca5ec;
    ram_cell[    9131] = 32'h0;  // 32'h0c769698;
    ram_cell[    9132] = 32'h0;  // 32'hdec2855c;
    ram_cell[    9133] = 32'h0;  // 32'h3c4613b1;
    ram_cell[    9134] = 32'h0;  // 32'h6127a75d;
    ram_cell[    9135] = 32'h0;  // 32'h2a318e62;
    ram_cell[    9136] = 32'h0;  // 32'h2bbd3bcb;
    ram_cell[    9137] = 32'h0;  // 32'h40390c99;
    ram_cell[    9138] = 32'h0;  // 32'h2ad029cf;
    ram_cell[    9139] = 32'h0;  // 32'ha27adc58;
    ram_cell[    9140] = 32'h0;  // 32'h7db43d10;
    ram_cell[    9141] = 32'h0;  // 32'h12d410e2;
    ram_cell[    9142] = 32'h0;  // 32'h9ba7582e;
    ram_cell[    9143] = 32'h0;  // 32'h6bb6c252;
    ram_cell[    9144] = 32'h0;  // 32'hadea2ec4;
    ram_cell[    9145] = 32'h0;  // 32'h13d43468;
    ram_cell[    9146] = 32'h0;  // 32'hf0035f46;
    ram_cell[    9147] = 32'h0;  // 32'hb7694817;
    ram_cell[    9148] = 32'h0;  // 32'h600ba9b4;
    ram_cell[    9149] = 32'h0;  // 32'haef75f74;
    ram_cell[    9150] = 32'h0;  // 32'hd9c6c902;
    ram_cell[    9151] = 32'h0;  // 32'heff60ba7;
    ram_cell[    9152] = 32'h0;  // 32'hdc6030ee;
    ram_cell[    9153] = 32'h0;  // 32'hf0eed3a3;
    ram_cell[    9154] = 32'h0;  // 32'hf8ac8029;
    ram_cell[    9155] = 32'h0;  // 32'h5fa81e5c;
    ram_cell[    9156] = 32'h0;  // 32'h5c9e7575;
    ram_cell[    9157] = 32'h0;  // 32'hc55d3377;
    ram_cell[    9158] = 32'h0;  // 32'h2d3a9bd8;
    ram_cell[    9159] = 32'h0;  // 32'h1e68e019;
    ram_cell[    9160] = 32'h0;  // 32'h7b712e3e;
    ram_cell[    9161] = 32'h0;  // 32'h57de6df4;
    ram_cell[    9162] = 32'h0;  // 32'hcc37f029;
    ram_cell[    9163] = 32'h0;  // 32'h1df12279;
    ram_cell[    9164] = 32'h0;  // 32'hfba28700;
    ram_cell[    9165] = 32'h0;  // 32'hb73fc653;
    ram_cell[    9166] = 32'h0;  // 32'h595f0e51;
    ram_cell[    9167] = 32'h0;  // 32'he6f84a09;
    ram_cell[    9168] = 32'h0;  // 32'h850c4702;
    ram_cell[    9169] = 32'h0;  // 32'ha80dabeb;
    ram_cell[    9170] = 32'h0;  // 32'hd8cd2f72;
    ram_cell[    9171] = 32'h0;  // 32'h583698fa;
    ram_cell[    9172] = 32'h0;  // 32'hc32d0dbf;
    ram_cell[    9173] = 32'h0;  // 32'hf04b14dc;
    ram_cell[    9174] = 32'h0;  // 32'h47d4ec34;
    ram_cell[    9175] = 32'h0;  // 32'h855395b4;
    ram_cell[    9176] = 32'h0;  // 32'h5c86ccc2;
    ram_cell[    9177] = 32'h0;  // 32'h82657fa8;
    ram_cell[    9178] = 32'h0;  // 32'h8e2ffb8b;
    ram_cell[    9179] = 32'h0;  // 32'h4e03ebd8;
    ram_cell[    9180] = 32'h0;  // 32'h754dcb1d;
    ram_cell[    9181] = 32'h0;  // 32'h55cec9c8;
    ram_cell[    9182] = 32'h0;  // 32'h3a8820cd;
    ram_cell[    9183] = 32'h0;  // 32'hc34b755f;
    ram_cell[    9184] = 32'h0;  // 32'h9991e4cf;
    ram_cell[    9185] = 32'h0;  // 32'h1ca58f52;
    ram_cell[    9186] = 32'h0;  // 32'h450484ea;
    ram_cell[    9187] = 32'h0;  // 32'hc8886831;
    ram_cell[    9188] = 32'h0;  // 32'h84157858;
    ram_cell[    9189] = 32'h0;  // 32'h190a8f97;
    ram_cell[    9190] = 32'h0;  // 32'h26b9efab;
    ram_cell[    9191] = 32'h0;  // 32'hd0533a3b;
    ram_cell[    9192] = 32'h0;  // 32'hbeecd530;
    ram_cell[    9193] = 32'h0;  // 32'h62a7f31a;
    ram_cell[    9194] = 32'h0;  // 32'h98a1b7f2;
    ram_cell[    9195] = 32'h0;  // 32'h8867168a;
    ram_cell[    9196] = 32'h0;  // 32'h50975eee;
    ram_cell[    9197] = 32'h0;  // 32'h1e91cf86;
    ram_cell[    9198] = 32'h0;  // 32'h1dbeaa6e;
    ram_cell[    9199] = 32'h0;  // 32'hfc4422cb;
    ram_cell[    9200] = 32'h0;  // 32'hd515ce66;
    ram_cell[    9201] = 32'h0;  // 32'hd01e1363;
    ram_cell[    9202] = 32'h0;  // 32'h8187bd3b;
    ram_cell[    9203] = 32'h0;  // 32'h60d74f08;
    ram_cell[    9204] = 32'h0;  // 32'h3e3bcd96;
    ram_cell[    9205] = 32'h0;  // 32'hd32ddc27;
    ram_cell[    9206] = 32'h0;  // 32'h1e32ced6;
    ram_cell[    9207] = 32'h0;  // 32'h4ebdf9bf;
    ram_cell[    9208] = 32'h0;  // 32'ha5c9234d;
    ram_cell[    9209] = 32'h0;  // 32'hfa3e9bc7;
    ram_cell[    9210] = 32'h0;  // 32'h4f8d013a;
    ram_cell[    9211] = 32'h0;  // 32'h16984432;
    ram_cell[    9212] = 32'h0;  // 32'h07bb28ea;
    ram_cell[    9213] = 32'h0;  // 32'hc13d6f08;
    ram_cell[    9214] = 32'h0;  // 32'h87061849;
    ram_cell[    9215] = 32'h0;  // 32'h9530f4a1;
    ram_cell[    9216] = 32'h0;  // 32'h72bafafa;
    ram_cell[    9217] = 32'h0;  // 32'hd4978ee7;
    ram_cell[    9218] = 32'h0;  // 32'he27c7f71;
    ram_cell[    9219] = 32'h0;  // 32'hc5dd7115;
    ram_cell[    9220] = 32'h0;  // 32'h8d6c070a;
    ram_cell[    9221] = 32'h0;  // 32'h838f208e;
    ram_cell[    9222] = 32'h0;  // 32'h7d1a3fd6;
    ram_cell[    9223] = 32'h0;  // 32'h30254a31;
    ram_cell[    9224] = 32'h0;  // 32'h3336c527;
    ram_cell[    9225] = 32'h0;  // 32'hf093aed5;
    ram_cell[    9226] = 32'h0;  // 32'hc57d955e;
    ram_cell[    9227] = 32'h0;  // 32'hbefec59d;
    ram_cell[    9228] = 32'h0;  // 32'h2c066e34;
    ram_cell[    9229] = 32'h0;  // 32'h9166b853;
    ram_cell[    9230] = 32'h0;  // 32'h3992fad2;
    ram_cell[    9231] = 32'h0;  // 32'h577e7ece;
    ram_cell[    9232] = 32'h0;  // 32'h6361bb56;
    ram_cell[    9233] = 32'h0;  // 32'ha1bcdf14;
    ram_cell[    9234] = 32'h0;  // 32'h70c68b63;
    ram_cell[    9235] = 32'h0;  // 32'ha3318933;
    ram_cell[    9236] = 32'h0;  // 32'hdf7211d9;
    ram_cell[    9237] = 32'h0;  // 32'ha8efe040;
    ram_cell[    9238] = 32'h0;  // 32'h9a5195bb;
    ram_cell[    9239] = 32'h0;  // 32'h1d96b0fd;
    ram_cell[    9240] = 32'h0;  // 32'h870b5fae;
    ram_cell[    9241] = 32'h0;  // 32'h9eaed8e6;
    ram_cell[    9242] = 32'h0;  // 32'he0c4d388;
    ram_cell[    9243] = 32'h0;  // 32'h0594addd;
    ram_cell[    9244] = 32'h0;  // 32'hfc636ef9;
    ram_cell[    9245] = 32'h0;  // 32'hfa4c483a;
    ram_cell[    9246] = 32'h0;  // 32'h2a1f5f5a;
    ram_cell[    9247] = 32'h0;  // 32'hd938e38a;
    ram_cell[    9248] = 32'h0;  // 32'hea91d375;
    ram_cell[    9249] = 32'h0;  // 32'h4642d1ce;
    ram_cell[    9250] = 32'h0;  // 32'hc33f27f7;
    ram_cell[    9251] = 32'h0;  // 32'hbe58e23e;
    ram_cell[    9252] = 32'h0;  // 32'hb893bab2;
    ram_cell[    9253] = 32'h0;  // 32'h9a3082f1;
    ram_cell[    9254] = 32'h0;  // 32'h9dd61803;
    ram_cell[    9255] = 32'h0;  // 32'h4f93d091;
    ram_cell[    9256] = 32'h0;  // 32'h160a8663;
    ram_cell[    9257] = 32'h0;  // 32'h007e98c6;
    ram_cell[    9258] = 32'h0;  // 32'h6dd35f1a;
    ram_cell[    9259] = 32'h0;  // 32'h736b044b;
    ram_cell[    9260] = 32'h0;  // 32'h5ef9a670;
    ram_cell[    9261] = 32'h0;  // 32'h529781c5;
    ram_cell[    9262] = 32'h0;  // 32'hbde89de9;
    ram_cell[    9263] = 32'h0;  // 32'h72112ab4;
    ram_cell[    9264] = 32'h0;  // 32'hc28cbcab;
    ram_cell[    9265] = 32'h0;  // 32'h959557ae;
    ram_cell[    9266] = 32'h0;  // 32'h21c3d3c4;
    ram_cell[    9267] = 32'h0;  // 32'hfc0d98da;
    ram_cell[    9268] = 32'h0;  // 32'hf11a5aae;
    ram_cell[    9269] = 32'h0;  // 32'hac86a8cc;
    ram_cell[    9270] = 32'h0;  // 32'hf096bd38;
    ram_cell[    9271] = 32'h0;  // 32'hb46f5250;
    ram_cell[    9272] = 32'h0;  // 32'he8f9a0d8;
    ram_cell[    9273] = 32'h0;  // 32'h994f01f8;
    ram_cell[    9274] = 32'h0;  // 32'h22d49967;
    ram_cell[    9275] = 32'h0;  // 32'h5b2ed85c;
    ram_cell[    9276] = 32'h0;  // 32'h198829d1;
    ram_cell[    9277] = 32'h0;  // 32'h73ac8940;
    ram_cell[    9278] = 32'h0;  // 32'h4db8a120;
    ram_cell[    9279] = 32'h0;  // 32'h96055c77;
    ram_cell[    9280] = 32'h0;  // 32'h4e9d7777;
    ram_cell[    9281] = 32'h0;  // 32'h6e987656;
    ram_cell[    9282] = 32'h0;  // 32'h9064d652;
    ram_cell[    9283] = 32'h0;  // 32'h754972cc;
    ram_cell[    9284] = 32'h0;  // 32'h947dce9a;
    ram_cell[    9285] = 32'h0;  // 32'hefcc0c94;
    ram_cell[    9286] = 32'h0;  // 32'h395a4e04;
    ram_cell[    9287] = 32'h0;  // 32'h76484f1d;
    ram_cell[    9288] = 32'h0;  // 32'h59057e39;
    ram_cell[    9289] = 32'h0;  // 32'hb316f5af;
    ram_cell[    9290] = 32'h0;  // 32'h6eb054a4;
    ram_cell[    9291] = 32'h0;  // 32'h739e7057;
    ram_cell[    9292] = 32'h0;  // 32'hcfba3157;
    ram_cell[    9293] = 32'h0;  // 32'h1b8030ee;
    ram_cell[    9294] = 32'h0;  // 32'h9687e85d;
    ram_cell[    9295] = 32'h0;  // 32'h3a518ee1;
    ram_cell[    9296] = 32'h0;  // 32'heda28f56;
    ram_cell[    9297] = 32'h0;  // 32'h0c83fbf3;
    ram_cell[    9298] = 32'h0;  // 32'hc7f94575;
    ram_cell[    9299] = 32'h0;  // 32'ha48deddc;
    ram_cell[    9300] = 32'h0;  // 32'h71da1955;
    ram_cell[    9301] = 32'h0;  // 32'hc3a68ac2;
    ram_cell[    9302] = 32'h0;  // 32'h8c6a9194;
    ram_cell[    9303] = 32'h0;  // 32'h6018620f;
    ram_cell[    9304] = 32'h0;  // 32'hbf486c31;
    ram_cell[    9305] = 32'h0;  // 32'hc25a6a24;
    ram_cell[    9306] = 32'h0;  // 32'h239b858b;
    ram_cell[    9307] = 32'h0;  // 32'hf42bf73e;
    ram_cell[    9308] = 32'h0;  // 32'h1b60dd0b;
    ram_cell[    9309] = 32'h0;  // 32'h5bbcd8d8;
    ram_cell[    9310] = 32'h0;  // 32'h01e972d3;
    ram_cell[    9311] = 32'h0;  // 32'h6a838b07;
    ram_cell[    9312] = 32'h0;  // 32'h878df9ad;
    ram_cell[    9313] = 32'h0;  // 32'h23457d01;
    ram_cell[    9314] = 32'h0;  // 32'hb087be2a;
    ram_cell[    9315] = 32'h0;  // 32'hc4cdd7b9;
    ram_cell[    9316] = 32'h0;  // 32'hea02f05d;
    ram_cell[    9317] = 32'h0;  // 32'heb7f11bf;
    ram_cell[    9318] = 32'h0;  // 32'h8c032a1b;
    ram_cell[    9319] = 32'h0;  // 32'hdcc9c068;
    ram_cell[    9320] = 32'h0;  // 32'h536e2df3;
    ram_cell[    9321] = 32'h0;  // 32'hcaf499a9;
    ram_cell[    9322] = 32'h0;  // 32'h3dc12e12;
    ram_cell[    9323] = 32'h0;  // 32'h48859d19;
    ram_cell[    9324] = 32'h0;  // 32'h497d1cdc;
    ram_cell[    9325] = 32'h0;  // 32'h71fa4bcd;
    ram_cell[    9326] = 32'h0;  // 32'h1806253e;
    ram_cell[    9327] = 32'h0;  // 32'h916e57dc;
    ram_cell[    9328] = 32'h0;  // 32'h483dfb8c;
    ram_cell[    9329] = 32'h0;  // 32'h58d6a1d7;
    ram_cell[    9330] = 32'h0;  // 32'h9f190c1b;
    ram_cell[    9331] = 32'h0;  // 32'hecfaa575;
    ram_cell[    9332] = 32'h0;  // 32'h5a9d5b65;
    ram_cell[    9333] = 32'h0;  // 32'h836a4374;
    ram_cell[    9334] = 32'h0;  // 32'h277b1187;
    ram_cell[    9335] = 32'h0;  // 32'h7d5f2eaf;
    ram_cell[    9336] = 32'h0;  // 32'ha24cb4d0;
    ram_cell[    9337] = 32'h0;  // 32'hb3e6772e;
    ram_cell[    9338] = 32'h0;  // 32'hd8f39c8b;
    ram_cell[    9339] = 32'h0;  // 32'h482a73a0;
    ram_cell[    9340] = 32'h0;  // 32'h1c6ce8e9;
    ram_cell[    9341] = 32'h0;  // 32'hce2d3ede;
    ram_cell[    9342] = 32'h0;  // 32'h0561398b;
    ram_cell[    9343] = 32'h0;  // 32'h7aec5ad9;
    ram_cell[    9344] = 32'h0;  // 32'he24f5d90;
    ram_cell[    9345] = 32'h0;  // 32'h8bc6728a;
    ram_cell[    9346] = 32'h0;  // 32'h75b02f88;
    ram_cell[    9347] = 32'h0;  // 32'h0850ebf7;
    ram_cell[    9348] = 32'h0;  // 32'h497495e5;
    ram_cell[    9349] = 32'h0;  // 32'h84ec06c5;
    ram_cell[    9350] = 32'h0;  // 32'h346582cb;
    ram_cell[    9351] = 32'h0;  // 32'hd05a9fe0;
    ram_cell[    9352] = 32'h0;  // 32'h984f5c21;
    ram_cell[    9353] = 32'h0;  // 32'hd5b0057e;
    ram_cell[    9354] = 32'h0;  // 32'h6db37310;
    ram_cell[    9355] = 32'h0;  // 32'h9995afed;
    ram_cell[    9356] = 32'h0;  // 32'ha5d6bb9c;
    ram_cell[    9357] = 32'h0;  // 32'h258313a2;
    ram_cell[    9358] = 32'h0;  // 32'h02c60cb8;
    ram_cell[    9359] = 32'h0;  // 32'hdf2ec571;
    ram_cell[    9360] = 32'h0;  // 32'hc515a0aa;
    ram_cell[    9361] = 32'h0;  // 32'h63f75b6e;
    ram_cell[    9362] = 32'h0;  // 32'h8eadf277;
    ram_cell[    9363] = 32'h0;  // 32'h9a708448;
    ram_cell[    9364] = 32'h0;  // 32'heab3c0db;
    ram_cell[    9365] = 32'h0;  // 32'he64668e9;
    ram_cell[    9366] = 32'h0;  // 32'h2205ca39;
    ram_cell[    9367] = 32'h0;  // 32'h12f7aec8;
    ram_cell[    9368] = 32'h0;  // 32'h4281d9d0;
    ram_cell[    9369] = 32'h0;  // 32'h9aff101a;
    ram_cell[    9370] = 32'h0;  // 32'h94336e62;
    ram_cell[    9371] = 32'h0;  // 32'h3d02d8af;
    ram_cell[    9372] = 32'h0;  // 32'hb6d8af75;
    ram_cell[    9373] = 32'h0;  // 32'hcea7a2d3;
    ram_cell[    9374] = 32'h0;  // 32'haedfec8f;
    ram_cell[    9375] = 32'h0;  // 32'h96a357d4;
    ram_cell[    9376] = 32'h0;  // 32'h188b7b43;
    ram_cell[    9377] = 32'h0;  // 32'h36981e32;
    ram_cell[    9378] = 32'h0;  // 32'h4497914b;
    ram_cell[    9379] = 32'h0;  // 32'h5011483b;
    ram_cell[    9380] = 32'h0;  // 32'hd8ece520;
    ram_cell[    9381] = 32'h0;  // 32'had40d599;
    ram_cell[    9382] = 32'h0;  // 32'hc4e70b5e;
    ram_cell[    9383] = 32'h0;  // 32'h0a00f362;
    ram_cell[    9384] = 32'h0;  // 32'h0ebf9c4c;
    ram_cell[    9385] = 32'h0;  // 32'h30a4390d;
    ram_cell[    9386] = 32'h0;  // 32'hcc6226dc;
    ram_cell[    9387] = 32'h0;  // 32'h06f988bf;
    ram_cell[    9388] = 32'h0;  // 32'h1e6483dc;
    ram_cell[    9389] = 32'h0;  // 32'hfeda4261;
    ram_cell[    9390] = 32'h0;  // 32'h7b3cb6a3;
    ram_cell[    9391] = 32'h0;  // 32'h2e191bcc;
    ram_cell[    9392] = 32'h0;  // 32'h06f6f258;
    ram_cell[    9393] = 32'h0;  // 32'h8e464bfb;
    ram_cell[    9394] = 32'h0;  // 32'h3838c2f5;
    ram_cell[    9395] = 32'h0;  // 32'h65c0db03;
    ram_cell[    9396] = 32'h0;  // 32'h2600e4b0;
    ram_cell[    9397] = 32'h0;  // 32'h4aea098d;
    ram_cell[    9398] = 32'h0;  // 32'h33f207b3;
    ram_cell[    9399] = 32'h0;  // 32'h44122729;
    ram_cell[    9400] = 32'h0;  // 32'hb94801a1;
    ram_cell[    9401] = 32'h0;  // 32'hf40af526;
    ram_cell[    9402] = 32'h0;  // 32'h647d93a0;
    ram_cell[    9403] = 32'h0;  // 32'ha153b524;
    ram_cell[    9404] = 32'h0;  // 32'h70d1376f;
    ram_cell[    9405] = 32'h0;  // 32'hffef62f5;
    ram_cell[    9406] = 32'h0;  // 32'h4d2ebc89;
    ram_cell[    9407] = 32'h0;  // 32'h4b4eef75;
    ram_cell[    9408] = 32'h0;  // 32'h93a2f896;
    ram_cell[    9409] = 32'h0;  // 32'hb15fecb6;
    ram_cell[    9410] = 32'h0;  // 32'h43480875;
    ram_cell[    9411] = 32'h0;  // 32'h59e2d819;
    ram_cell[    9412] = 32'h0;  // 32'h6299b27a;
    ram_cell[    9413] = 32'h0;  // 32'h23eaf006;
    ram_cell[    9414] = 32'h0;  // 32'h316df5fd;
    ram_cell[    9415] = 32'h0;  // 32'he3a80400;
    ram_cell[    9416] = 32'h0;  // 32'h48a0c37d;
    ram_cell[    9417] = 32'h0;  // 32'hd934448d;
    ram_cell[    9418] = 32'h0;  // 32'h1da5e8ca;
    ram_cell[    9419] = 32'h0;  // 32'hfa92e243;
    ram_cell[    9420] = 32'h0;  // 32'h7c6e2ba5;
    ram_cell[    9421] = 32'h0;  // 32'hfefa19d1;
    ram_cell[    9422] = 32'h0;  // 32'h25b933e7;
    ram_cell[    9423] = 32'h0;  // 32'h41d0fff9;
    ram_cell[    9424] = 32'h0;  // 32'hf4756f35;
    ram_cell[    9425] = 32'h0;  // 32'h7ee4c18f;
    ram_cell[    9426] = 32'h0;  // 32'h143afec1;
    ram_cell[    9427] = 32'h0;  // 32'hcbda8142;
    ram_cell[    9428] = 32'h0;  // 32'hef7f4f63;
    ram_cell[    9429] = 32'h0;  // 32'haf50e346;
    ram_cell[    9430] = 32'h0;  // 32'hd41c0819;
    ram_cell[    9431] = 32'h0;  // 32'h1ebcb62f;
    ram_cell[    9432] = 32'h0;  // 32'he9f9a681;
    ram_cell[    9433] = 32'h0;  // 32'he2fb1027;
    ram_cell[    9434] = 32'h0;  // 32'h72d5203d;
    ram_cell[    9435] = 32'h0;  // 32'hbd8b678c;
    ram_cell[    9436] = 32'h0;  // 32'hb9a6a53a;
    ram_cell[    9437] = 32'h0;  // 32'h26b91783;
    ram_cell[    9438] = 32'h0;  // 32'h0cff2a2f;
    ram_cell[    9439] = 32'h0;  // 32'ha251be8d;
    ram_cell[    9440] = 32'h0;  // 32'hd59c8ead;
    ram_cell[    9441] = 32'h0;  // 32'ha4d2612b;
    ram_cell[    9442] = 32'h0;  // 32'h7c9a549d;
    ram_cell[    9443] = 32'h0;  // 32'h409c6289;
    ram_cell[    9444] = 32'h0;  // 32'h9d5db3dd;
    ram_cell[    9445] = 32'h0;  // 32'h92752e8b;
    ram_cell[    9446] = 32'h0;  // 32'h0a4a3ba8;
    ram_cell[    9447] = 32'h0;  // 32'h71356857;
    ram_cell[    9448] = 32'h0;  // 32'h44e35f68;
    ram_cell[    9449] = 32'h0;  // 32'h961c519f;
    ram_cell[    9450] = 32'h0;  // 32'hb7cf39f4;
    ram_cell[    9451] = 32'h0;  // 32'hb2df51ee;
    ram_cell[    9452] = 32'h0;  // 32'hceaf6255;
    ram_cell[    9453] = 32'h0;  // 32'he86922dd;
    ram_cell[    9454] = 32'h0;  // 32'h6e465f5e;
    ram_cell[    9455] = 32'h0;  // 32'hfb05a880;
    ram_cell[    9456] = 32'h0;  // 32'hf7ae62b7;
    ram_cell[    9457] = 32'h0;  // 32'hee3bb54c;
    ram_cell[    9458] = 32'h0;  // 32'he1474312;
    ram_cell[    9459] = 32'h0;  // 32'hf6efebf8;
    ram_cell[    9460] = 32'h0;  // 32'h8bd51171;
    ram_cell[    9461] = 32'h0;  // 32'h7bc935c0;
    ram_cell[    9462] = 32'h0;  // 32'h05a50112;
    ram_cell[    9463] = 32'h0;  // 32'h37847a46;
    ram_cell[    9464] = 32'h0;  // 32'h1eb7c7d5;
    ram_cell[    9465] = 32'h0;  // 32'h1147f241;
    ram_cell[    9466] = 32'h0;  // 32'h9be02910;
    ram_cell[    9467] = 32'h0;  // 32'ha14fa796;
    ram_cell[    9468] = 32'h0;  // 32'h9f36c9ab;
    ram_cell[    9469] = 32'h0;  // 32'h2f870024;
    ram_cell[    9470] = 32'h0;  // 32'hdc824f54;
    ram_cell[    9471] = 32'h0;  // 32'h8539415f;
    ram_cell[    9472] = 32'h0;  // 32'ha041133a;
    ram_cell[    9473] = 32'h0;  // 32'h900da921;
    ram_cell[    9474] = 32'h0;  // 32'h25e20417;
    ram_cell[    9475] = 32'h0;  // 32'h3317438e;
    ram_cell[    9476] = 32'h0;  // 32'hfcaa6372;
    ram_cell[    9477] = 32'h0;  // 32'hd6e13cb7;
    ram_cell[    9478] = 32'h0;  // 32'haa66e503;
    ram_cell[    9479] = 32'h0;  // 32'hcdcdf731;
    ram_cell[    9480] = 32'h0;  // 32'h1ab92a66;
    ram_cell[    9481] = 32'h0;  // 32'ha83d3d14;
    ram_cell[    9482] = 32'h0;  // 32'heb327a45;
    ram_cell[    9483] = 32'h0;  // 32'h0f0bc094;
    ram_cell[    9484] = 32'h0;  // 32'hacad1059;
    ram_cell[    9485] = 32'h0;  // 32'h2e6d51bb;
    ram_cell[    9486] = 32'h0;  // 32'h568c7e31;
    ram_cell[    9487] = 32'h0;  // 32'h5da80eac;
    ram_cell[    9488] = 32'h0;  // 32'h4e9e0b96;
    ram_cell[    9489] = 32'h0;  // 32'h3e522d4d;
    ram_cell[    9490] = 32'h0;  // 32'h04773846;
    ram_cell[    9491] = 32'h0;  // 32'h1706e021;
    ram_cell[    9492] = 32'h0;  // 32'h7d287bbb;
    ram_cell[    9493] = 32'h0;  // 32'hd18d6fd2;
    ram_cell[    9494] = 32'h0;  // 32'hf4ac5bf4;
    ram_cell[    9495] = 32'h0;  // 32'hb7804e20;
    ram_cell[    9496] = 32'h0;  // 32'h28186b3b;
    ram_cell[    9497] = 32'h0;  // 32'haa5a851f;
    ram_cell[    9498] = 32'h0;  // 32'ha312b521;
    ram_cell[    9499] = 32'h0;  // 32'h54d89d8e;
    ram_cell[    9500] = 32'h0;  // 32'h355b33d9;
    ram_cell[    9501] = 32'h0;  // 32'hcaf2016f;
    ram_cell[    9502] = 32'h0;  // 32'h37b68234;
    ram_cell[    9503] = 32'h0;  // 32'h33821ad5;
    ram_cell[    9504] = 32'h0;  // 32'h7fe66726;
    ram_cell[    9505] = 32'h0;  // 32'h0696fc69;
    ram_cell[    9506] = 32'h0;  // 32'h708c8171;
    ram_cell[    9507] = 32'h0;  // 32'h7f41d6ee;
    ram_cell[    9508] = 32'h0;  // 32'hf8d4d8b9;
    ram_cell[    9509] = 32'h0;  // 32'hf2664bd8;
    ram_cell[    9510] = 32'h0;  // 32'h36bafac4;
    ram_cell[    9511] = 32'h0;  // 32'h4ccd207f;
    ram_cell[    9512] = 32'h0;  // 32'h57f46c7d;
    ram_cell[    9513] = 32'h0;  // 32'hfcca82de;
    ram_cell[    9514] = 32'h0;  // 32'hc0890559;
    ram_cell[    9515] = 32'h0;  // 32'h1c67ebb6;
    ram_cell[    9516] = 32'h0;  // 32'h64303ed2;
    ram_cell[    9517] = 32'h0;  // 32'h920129ba;
    ram_cell[    9518] = 32'h0;  // 32'h957fa5ba;
    ram_cell[    9519] = 32'h0;  // 32'h64df507e;
    ram_cell[    9520] = 32'h0;  // 32'hd8961109;
    ram_cell[    9521] = 32'h0;  // 32'h160b4be5;
    ram_cell[    9522] = 32'h0;  // 32'hed9bae67;
    ram_cell[    9523] = 32'h0;  // 32'h961a4966;
    ram_cell[    9524] = 32'h0;  // 32'h2490241d;
    ram_cell[    9525] = 32'h0;  // 32'h0213a8e1;
    ram_cell[    9526] = 32'h0;  // 32'h1256cec8;
    ram_cell[    9527] = 32'h0;  // 32'h9589ef27;
    ram_cell[    9528] = 32'h0;  // 32'hb32c73ae;
    ram_cell[    9529] = 32'h0;  // 32'hcf449bcd;
    ram_cell[    9530] = 32'h0;  // 32'h34431d24;
    ram_cell[    9531] = 32'h0;  // 32'h6f9b8eb5;
    ram_cell[    9532] = 32'h0;  // 32'hc467eb71;
    ram_cell[    9533] = 32'h0;  // 32'h9ff954f5;
    ram_cell[    9534] = 32'h0;  // 32'h291e0178;
    ram_cell[    9535] = 32'h0;  // 32'ha67e535b;
    ram_cell[    9536] = 32'h0;  // 32'hdaf8672d;
    ram_cell[    9537] = 32'h0;  // 32'h31af4f78;
    ram_cell[    9538] = 32'h0;  // 32'he782e4b4;
    ram_cell[    9539] = 32'h0;  // 32'hd754bd4a;
    ram_cell[    9540] = 32'h0;  // 32'h5a44bae3;
    ram_cell[    9541] = 32'h0;  // 32'h58841408;
    ram_cell[    9542] = 32'h0;  // 32'ha262cd3d;
    ram_cell[    9543] = 32'h0;  // 32'h02d788ab;
    ram_cell[    9544] = 32'h0;  // 32'h765ea831;
    ram_cell[    9545] = 32'h0;  // 32'h0965ad68;
    ram_cell[    9546] = 32'h0;  // 32'h9b7a1263;
    ram_cell[    9547] = 32'h0;  // 32'ha05d103e;
    ram_cell[    9548] = 32'h0;  // 32'h2a6d9a53;
    ram_cell[    9549] = 32'h0;  // 32'he84227e5;
    ram_cell[    9550] = 32'h0;  // 32'h3fee1174;
    ram_cell[    9551] = 32'h0;  // 32'h8655a08b;
    ram_cell[    9552] = 32'h0;  // 32'h0c76ea0f;
    ram_cell[    9553] = 32'h0;  // 32'h64ec685f;
    ram_cell[    9554] = 32'h0;  // 32'h8315acf1;
    ram_cell[    9555] = 32'h0;  // 32'hc20a9858;
    ram_cell[    9556] = 32'h0;  // 32'hed476d01;
    ram_cell[    9557] = 32'h0;  // 32'h27ee0a1d;
    ram_cell[    9558] = 32'h0;  // 32'h23b16a52;
    ram_cell[    9559] = 32'h0;  // 32'h066aece7;
    ram_cell[    9560] = 32'h0;  // 32'hd1d3675b;
    ram_cell[    9561] = 32'h0;  // 32'h6e171238;
    ram_cell[    9562] = 32'h0;  // 32'hf3d42223;
    ram_cell[    9563] = 32'h0;  // 32'h8f77bc41;
    ram_cell[    9564] = 32'h0;  // 32'h998e90a7;
    ram_cell[    9565] = 32'h0;  // 32'he3a65664;
    ram_cell[    9566] = 32'h0;  // 32'h62c75a6e;
    ram_cell[    9567] = 32'h0;  // 32'h75013b8b;
    ram_cell[    9568] = 32'h0;  // 32'h2610fa1c;
    ram_cell[    9569] = 32'h0;  // 32'hefd804a9;
    ram_cell[    9570] = 32'h0;  // 32'h3c6ee827;
    ram_cell[    9571] = 32'h0;  // 32'h7e24a6f6;
    ram_cell[    9572] = 32'h0;  // 32'he89b1450;
    ram_cell[    9573] = 32'h0;  // 32'h9d863cc2;
    ram_cell[    9574] = 32'h0;  // 32'hc6afbaf2;
    ram_cell[    9575] = 32'h0;  // 32'h55c5d4d1;
    ram_cell[    9576] = 32'h0;  // 32'hb04e5c87;
    ram_cell[    9577] = 32'h0;  // 32'hb1e4b2b3;
    ram_cell[    9578] = 32'h0;  // 32'h431aece9;
    ram_cell[    9579] = 32'h0;  // 32'ha2fae6ba;
    ram_cell[    9580] = 32'h0;  // 32'hbe5a68b9;
    ram_cell[    9581] = 32'h0;  // 32'hb8199ce0;
    ram_cell[    9582] = 32'h0;  // 32'ha874fa86;
    ram_cell[    9583] = 32'h0;  // 32'hb943e9a6;
    ram_cell[    9584] = 32'h0;  // 32'hf2421b3f;
    ram_cell[    9585] = 32'h0;  // 32'hba0508b6;
    ram_cell[    9586] = 32'h0;  // 32'hfdfbbe17;
    ram_cell[    9587] = 32'h0;  // 32'hb674e34d;
    ram_cell[    9588] = 32'h0;  // 32'h777a91e2;
    ram_cell[    9589] = 32'h0;  // 32'hdcfc94ad;
    ram_cell[    9590] = 32'h0;  // 32'hefd0435a;
    ram_cell[    9591] = 32'h0;  // 32'hdd9eed8d;
    ram_cell[    9592] = 32'h0;  // 32'hfbda903c;
    ram_cell[    9593] = 32'h0;  // 32'h2982b0ef;
    ram_cell[    9594] = 32'h0;  // 32'ha619de38;
    ram_cell[    9595] = 32'h0;  // 32'h4989ad14;
    ram_cell[    9596] = 32'h0;  // 32'h811b2810;
    ram_cell[    9597] = 32'h0;  // 32'h5ce64259;
    ram_cell[    9598] = 32'h0;  // 32'h17a6680a;
    ram_cell[    9599] = 32'h0;  // 32'heb9112ad;
    ram_cell[    9600] = 32'h0;  // 32'h025fa839;
    ram_cell[    9601] = 32'h0;  // 32'h0c73a43f;
    ram_cell[    9602] = 32'h0;  // 32'h964f1c4a;
    ram_cell[    9603] = 32'h0;  // 32'h277bd4d7;
    ram_cell[    9604] = 32'h0;  // 32'h9ec9739f;
    ram_cell[    9605] = 32'h0;  // 32'h6d86e928;
    ram_cell[    9606] = 32'h0;  // 32'h919373c1;
    ram_cell[    9607] = 32'h0;  // 32'he7ed4b0d;
    ram_cell[    9608] = 32'h0;  // 32'h35a85d8d;
    ram_cell[    9609] = 32'h0;  // 32'h930533a5;
    ram_cell[    9610] = 32'h0;  // 32'hbd0ae513;
    ram_cell[    9611] = 32'h0;  // 32'h4e402ae3;
    ram_cell[    9612] = 32'h0;  // 32'h5e7e44d6;
    ram_cell[    9613] = 32'h0;  // 32'h333868bf;
    ram_cell[    9614] = 32'h0;  // 32'hac95f6b2;
    ram_cell[    9615] = 32'h0;  // 32'hebcb1a07;
    ram_cell[    9616] = 32'h0;  // 32'h903c1e93;
    ram_cell[    9617] = 32'h0;  // 32'h12457fd0;
    ram_cell[    9618] = 32'h0;  // 32'hf9624b72;
    ram_cell[    9619] = 32'h0;  // 32'h856d8906;
    ram_cell[    9620] = 32'h0;  // 32'h1f497d55;
    ram_cell[    9621] = 32'h0;  // 32'hbfd4b8cc;
    ram_cell[    9622] = 32'h0;  // 32'h4c1b88f8;
    ram_cell[    9623] = 32'h0;  // 32'h6b8b4034;
    ram_cell[    9624] = 32'h0;  // 32'hecf198f5;
    ram_cell[    9625] = 32'h0;  // 32'ha89721db;
    ram_cell[    9626] = 32'h0;  // 32'hfc37c4fd;
    ram_cell[    9627] = 32'h0;  // 32'h9e1a25c9;
    ram_cell[    9628] = 32'h0;  // 32'h03f7c453;
    ram_cell[    9629] = 32'h0;  // 32'hbf543469;
    ram_cell[    9630] = 32'h0;  // 32'h02477f17;
    ram_cell[    9631] = 32'h0;  // 32'h8a1de822;
    ram_cell[    9632] = 32'h0;  // 32'h1cf39313;
    ram_cell[    9633] = 32'h0;  // 32'hc1e1c797;
    ram_cell[    9634] = 32'h0;  // 32'h8165821f;
    ram_cell[    9635] = 32'h0;  // 32'hbc21e12d;
    ram_cell[    9636] = 32'h0;  // 32'h64931e89;
    ram_cell[    9637] = 32'h0;  // 32'hd2d6cae7;
    ram_cell[    9638] = 32'h0;  // 32'hb6815f65;
    ram_cell[    9639] = 32'h0;  // 32'hd86a9ab7;
    ram_cell[    9640] = 32'h0;  // 32'h9871238d;
    ram_cell[    9641] = 32'h0;  // 32'h8bdbc6b5;
    ram_cell[    9642] = 32'h0;  // 32'hf2fca65e;
    ram_cell[    9643] = 32'h0;  // 32'h707c0aa4;
    ram_cell[    9644] = 32'h0;  // 32'h9eacae2a;
    ram_cell[    9645] = 32'h0;  // 32'hc7cca24c;
    ram_cell[    9646] = 32'h0;  // 32'haa0bda42;
    ram_cell[    9647] = 32'h0;  // 32'h3e7354ea;
    ram_cell[    9648] = 32'h0;  // 32'h19c09e0c;
    ram_cell[    9649] = 32'h0;  // 32'h9a3f3c81;
    ram_cell[    9650] = 32'h0;  // 32'h8b21654e;
    ram_cell[    9651] = 32'h0;  // 32'h748f6cfc;
    ram_cell[    9652] = 32'h0;  // 32'hf63d97ef;
    ram_cell[    9653] = 32'h0;  // 32'h2e16c19f;
    ram_cell[    9654] = 32'h0;  // 32'h067b90fa;
    ram_cell[    9655] = 32'h0;  // 32'h33bc5594;
    ram_cell[    9656] = 32'h0;  // 32'ha1ebd747;
    ram_cell[    9657] = 32'h0;  // 32'hd9f5e645;
    ram_cell[    9658] = 32'h0;  // 32'h81d64bc9;
    ram_cell[    9659] = 32'h0;  // 32'he8c70639;
    ram_cell[    9660] = 32'h0;  // 32'h45721a83;
    ram_cell[    9661] = 32'h0;  // 32'h57e6b1ea;
    ram_cell[    9662] = 32'h0;  // 32'hb39c777d;
    ram_cell[    9663] = 32'h0;  // 32'ha694aebf;
    ram_cell[    9664] = 32'h0;  // 32'h2cf1c391;
    ram_cell[    9665] = 32'h0;  // 32'h1054e630;
    ram_cell[    9666] = 32'h0;  // 32'h5a7827c0;
    ram_cell[    9667] = 32'h0;  // 32'h753f3d61;
    ram_cell[    9668] = 32'h0;  // 32'hc3a33790;
    ram_cell[    9669] = 32'h0;  // 32'hd463857e;
    ram_cell[    9670] = 32'h0;  // 32'h1ba41a80;
    ram_cell[    9671] = 32'h0;  // 32'h05c88bd7;
    ram_cell[    9672] = 32'h0;  // 32'hc4b1d667;
    ram_cell[    9673] = 32'h0;  // 32'h7de4ede9;
    ram_cell[    9674] = 32'h0;  // 32'h458e126a;
    ram_cell[    9675] = 32'h0;  // 32'h17e938a8;
    ram_cell[    9676] = 32'h0;  // 32'h07a96663;
    ram_cell[    9677] = 32'h0;  // 32'hf5c663e9;
    ram_cell[    9678] = 32'h0;  // 32'h44f979f6;
    ram_cell[    9679] = 32'h0;  // 32'hc746a0b8;
    ram_cell[    9680] = 32'h0;  // 32'ha04b709f;
    ram_cell[    9681] = 32'h0;  // 32'h6c9ba2db;
    ram_cell[    9682] = 32'h0;  // 32'hdea7d452;
    ram_cell[    9683] = 32'h0;  // 32'h767ca5ed;
    ram_cell[    9684] = 32'h0;  // 32'h4a568656;
    ram_cell[    9685] = 32'h0;  // 32'h115a6a3f;
    ram_cell[    9686] = 32'h0;  // 32'hbeffa7e9;
    ram_cell[    9687] = 32'h0;  // 32'hf83e8663;
    ram_cell[    9688] = 32'h0;  // 32'h1610e2fd;
    ram_cell[    9689] = 32'h0;  // 32'h121ad59e;
    ram_cell[    9690] = 32'h0;  // 32'h9fa42b5a;
    ram_cell[    9691] = 32'h0;  // 32'h4d37e2ec;
    ram_cell[    9692] = 32'h0;  // 32'hc5738e35;
    ram_cell[    9693] = 32'h0;  // 32'h8f7f5fd5;
    ram_cell[    9694] = 32'h0;  // 32'hbdba6174;
    ram_cell[    9695] = 32'h0;  // 32'h62f7151d;
    ram_cell[    9696] = 32'h0;  // 32'h88037688;
    ram_cell[    9697] = 32'h0;  // 32'h5feef86b;
    ram_cell[    9698] = 32'h0;  // 32'hec4f9560;
    ram_cell[    9699] = 32'h0;  // 32'h8db6aef1;
    ram_cell[    9700] = 32'h0;  // 32'hcbad346a;
    ram_cell[    9701] = 32'h0;  // 32'h7229e23d;
    ram_cell[    9702] = 32'h0;  // 32'h3c0a6535;
    ram_cell[    9703] = 32'h0;  // 32'hf8c29a94;
    ram_cell[    9704] = 32'h0;  // 32'hfe1dc197;
    ram_cell[    9705] = 32'h0;  // 32'h5df4a8cc;
    ram_cell[    9706] = 32'h0;  // 32'h250c65c5;
    ram_cell[    9707] = 32'h0;  // 32'h8384b640;
    ram_cell[    9708] = 32'h0;  // 32'h4b42fd8e;
    ram_cell[    9709] = 32'h0;  // 32'h89e8bbfe;
    ram_cell[    9710] = 32'h0;  // 32'h8aaab8c9;
    ram_cell[    9711] = 32'h0;  // 32'hdef32cd8;
    ram_cell[    9712] = 32'h0;  // 32'h7b64100f;
    ram_cell[    9713] = 32'h0;  // 32'h70f0dc12;
    ram_cell[    9714] = 32'h0;  // 32'h43f99cb5;
    ram_cell[    9715] = 32'h0;  // 32'hf5144647;
    ram_cell[    9716] = 32'h0;  // 32'h44b962bc;
    ram_cell[    9717] = 32'h0;  // 32'h935d6289;
    ram_cell[    9718] = 32'h0;  // 32'hb8bff116;
    ram_cell[    9719] = 32'h0;  // 32'h38591118;
    ram_cell[    9720] = 32'h0;  // 32'h772c54e9;
    ram_cell[    9721] = 32'h0;  // 32'h1044b3f6;
    ram_cell[    9722] = 32'h0;  // 32'h26f5c165;
    ram_cell[    9723] = 32'h0;  // 32'h34c5fecf;
    ram_cell[    9724] = 32'h0;  // 32'h4afac252;
    ram_cell[    9725] = 32'h0;  // 32'he6e91bc6;
    ram_cell[    9726] = 32'h0;  // 32'hb21e7113;
    ram_cell[    9727] = 32'h0;  // 32'h032bd5b8;
    ram_cell[    9728] = 32'h0;  // 32'hdb5648a5;
    ram_cell[    9729] = 32'h0;  // 32'hf39e50a2;
    ram_cell[    9730] = 32'h0;  // 32'hc75bdfba;
    ram_cell[    9731] = 32'h0;  // 32'h9b9cd725;
    ram_cell[    9732] = 32'h0;  // 32'h1b0ebc0d;
    ram_cell[    9733] = 32'h0;  // 32'hd188f1d5;
    ram_cell[    9734] = 32'h0;  // 32'hbc9a6ee2;
    ram_cell[    9735] = 32'h0;  // 32'hf2332265;
    ram_cell[    9736] = 32'h0;  // 32'h0b1af63c;
    ram_cell[    9737] = 32'h0;  // 32'h9247e28f;
    ram_cell[    9738] = 32'h0;  // 32'h20f32913;
    ram_cell[    9739] = 32'h0;  // 32'ha14ebd50;
    ram_cell[    9740] = 32'h0;  // 32'h1e5a1b70;
    ram_cell[    9741] = 32'h0;  // 32'h79b97f40;
    ram_cell[    9742] = 32'h0;  // 32'h53ce38ab;
    ram_cell[    9743] = 32'h0;  // 32'h71f4005f;
    ram_cell[    9744] = 32'h0;  // 32'h48c56388;
    ram_cell[    9745] = 32'h0;  // 32'hcfce41b0;
    ram_cell[    9746] = 32'h0;  // 32'h38a9e990;
    ram_cell[    9747] = 32'h0;  // 32'h3e2da3a1;
    ram_cell[    9748] = 32'h0;  // 32'h4f852dd4;
    ram_cell[    9749] = 32'h0;  // 32'h265af7d4;
    ram_cell[    9750] = 32'h0;  // 32'h6eb9ddb4;
    ram_cell[    9751] = 32'h0;  // 32'h0f671f3c;
    ram_cell[    9752] = 32'h0;  // 32'hd6e3cb2e;
    ram_cell[    9753] = 32'h0;  // 32'he4a0dfc8;
    ram_cell[    9754] = 32'h0;  // 32'h2f468525;
    ram_cell[    9755] = 32'h0;  // 32'hbcb15de0;
    ram_cell[    9756] = 32'h0;  // 32'haf22d24e;
    ram_cell[    9757] = 32'h0;  // 32'he70fa350;
    ram_cell[    9758] = 32'h0;  // 32'h554d2dfc;
    ram_cell[    9759] = 32'h0;  // 32'h6074ee41;
    ram_cell[    9760] = 32'h0;  // 32'hf92e2458;
    ram_cell[    9761] = 32'h0;  // 32'h399069b5;
    ram_cell[    9762] = 32'h0;  // 32'heb8e1e86;
    ram_cell[    9763] = 32'h0;  // 32'hab0ae98a;
    ram_cell[    9764] = 32'h0;  // 32'hc4548059;
    ram_cell[    9765] = 32'h0;  // 32'h8631cb21;
    ram_cell[    9766] = 32'h0;  // 32'h963addb3;
    ram_cell[    9767] = 32'h0;  // 32'hdf8782bd;
    ram_cell[    9768] = 32'h0;  // 32'h2b25ac14;
    ram_cell[    9769] = 32'h0;  // 32'hb8de509b;
    ram_cell[    9770] = 32'h0;  // 32'h2c21b4ee;
    ram_cell[    9771] = 32'h0;  // 32'hd0c31a39;
    ram_cell[    9772] = 32'h0;  // 32'hb5912e02;
    ram_cell[    9773] = 32'h0;  // 32'h5d27191b;
    ram_cell[    9774] = 32'h0;  // 32'he8c86edb;
    ram_cell[    9775] = 32'h0;  // 32'h545928bf;
    ram_cell[    9776] = 32'h0;  // 32'h079f03a9;
    ram_cell[    9777] = 32'h0;  // 32'h1847b935;
    ram_cell[    9778] = 32'h0;  // 32'h778ef2e9;
    ram_cell[    9779] = 32'h0;  // 32'h2adf96cf;
    ram_cell[    9780] = 32'h0;  // 32'h98ce5f18;
    ram_cell[    9781] = 32'h0;  // 32'h82d8782e;
    ram_cell[    9782] = 32'h0;  // 32'hc53890fd;
    ram_cell[    9783] = 32'h0;  // 32'h3c5ed6cd;
    ram_cell[    9784] = 32'h0;  // 32'h962951a4;
    ram_cell[    9785] = 32'h0;  // 32'h5e7e22ad;
    ram_cell[    9786] = 32'h0;  // 32'h0b1df87b;
    ram_cell[    9787] = 32'h0;  // 32'hd4d7e68a;
    ram_cell[    9788] = 32'h0;  // 32'h358fc41c;
    ram_cell[    9789] = 32'h0;  // 32'h8ba08181;
    ram_cell[    9790] = 32'h0;  // 32'hef00df49;
    ram_cell[    9791] = 32'h0;  // 32'h4c1070ff;
    ram_cell[    9792] = 32'h0;  // 32'h92f3af46;
    ram_cell[    9793] = 32'h0;  // 32'h60b79ca1;
    ram_cell[    9794] = 32'h0;  // 32'h253d0a78;
    ram_cell[    9795] = 32'h0;  // 32'hc4af75e8;
    ram_cell[    9796] = 32'h0;  // 32'h0fb2265a;
    ram_cell[    9797] = 32'h0;  // 32'hbf5a0ffd;
    ram_cell[    9798] = 32'h0;  // 32'h064ad4f3;
    ram_cell[    9799] = 32'h0;  // 32'h0e760f8d;
    ram_cell[    9800] = 32'h0;  // 32'hcfbd7277;
    ram_cell[    9801] = 32'h0;  // 32'h0e1e7957;
    ram_cell[    9802] = 32'h0;  // 32'h43955741;
    ram_cell[    9803] = 32'h0;  // 32'he8d9fbad;
    ram_cell[    9804] = 32'h0;  // 32'he6664c9c;
    ram_cell[    9805] = 32'h0;  // 32'h7f282824;
    ram_cell[    9806] = 32'h0;  // 32'h6dee4286;
    ram_cell[    9807] = 32'h0;  // 32'ha9bf8143;
    ram_cell[    9808] = 32'h0;  // 32'hc17f9a6e;
    ram_cell[    9809] = 32'h0;  // 32'ha7905a17;
    ram_cell[    9810] = 32'h0;  // 32'hfa814462;
    ram_cell[    9811] = 32'h0;  // 32'h03519d87;
    ram_cell[    9812] = 32'h0;  // 32'h12bc820a;
    ram_cell[    9813] = 32'h0;  // 32'he31c4793;
    ram_cell[    9814] = 32'h0;  // 32'h3b3c67e9;
    ram_cell[    9815] = 32'h0;  // 32'hb49edd44;
    ram_cell[    9816] = 32'h0;  // 32'h5dab3c5e;
    ram_cell[    9817] = 32'h0;  // 32'h145339d3;
    ram_cell[    9818] = 32'h0;  // 32'hb8fe0a01;
    ram_cell[    9819] = 32'h0;  // 32'h80fa1e4f;
    ram_cell[    9820] = 32'h0;  // 32'hfd7e4766;
    ram_cell[    9821] = 32'h0;  // 32'h1b6a9acb;
    ram_cell[    9822] = 32'h0;  // 32'h6483a774;
    ram_cell[    9823] = 32'h0;  // 32'h74513c48;
    ram_cell[    9824] = 32'h0;  // 32'h61b33106;
    ram_cell[    9825] = 32'h0;  // 32'hbfdf37d9;
    ram_cell[    9826] = 32'h0;  // 32'h8becff04;
    ram_cell[    9827] = 32'h0;  // 32'hd7bc28a7;
    ram_cell[    9828] = 32'h0;  // 32'h94b7e5f9;
    ram_cell[    9829] = 32'h0;  // 32'h3ca40169;
    ram_cell[    9830] = 32'h0;  // 32'h3cb38ca3;
    ram_cell[    9831] = 32'h0;  // 32'h0c21573a;
    ram_cell[    9832] = 32'h0;  // 32'hf67bdddc;
    ram_cell[    9833] = 32'h0;  // 32'hbe7cbb66;
    ram_cell[    9834] = 32'h0;  // 32'hfdde10ed;
    ram_cell[    9835] = 32'h0;  // 32'ha91002d2;
    ram_cell[    9836] = 32'h0;  // 32'hdb66b376;
    ram_cell[    9837] = 32'h0;  // 32'h2d7ca104;
    ram_cell[    9838] = 32'h0;  // 32'h1ba0508c;
    ram_cell[    9839] = 32'h0;  // 32'h97831e02;
    ram_cell[    9840] = 32'h0;  // 32'h22a4d578;
    ram_cell[    9841] = 32'h0;  // 32'h63e3ab33;
    ram_cell[    9842] = 32'h0;  // 32'h5311c059;
    ram_cell[    9843] = 32'h0;  // 32'h1c8f4ba5;
    ram_cell[    9844] = 32'h0;  // 32'haa7a4612;
    ram_cell[    9845] = 32'h0;  // 32'hbf557079;
    ram_cell[    9846] = 32'h0;  // 32'h27d469ee;
    ram_cell[    9847] = 32'h0;  // 32'h4d54b26a;
    ram_cell[    9848] = 32'h0;  // 32'haa307f98;
    ram_cell[    9849] = 32'h0;  // 32'h2dea66dd;
    ram_cell[    9850] = 32'h0;  // 32'hf2847c22;
    ram_cell[    9851] = 32'h0;  // 32'h7716a662;
    ram_cell[    9852] = 32'h0;  // 32'h030fc5b4;
    ram_cell[    9853] = 32'h0;  // 32'h1b7b7ac8;
    ram_cell[    9854] = 32'h0;  // 32'h6de81a1d;
    ram_cell[    9855] = 32'h0;  // 32'h74cfcf99;
    ram_cell[    9856] = 32'h0;  // 32'h58d075f2;
    ram_cell[    9857] = 32'h0;  // 32'h748f1fd9;
    ram_cell[    9858] = 32'h0;  // 32'h0785952e;
    ram_cell[    9859] = 32'h0;  // 32'h5cfd04e4;
    ram_cell[    9860] = 32'h0;  // 32'hcfa13619;
    ram_cell[    9861] = 32'h0;  // 32'h59b86509;
    ram_cell[    9862] = 32'h0;  // 32'h679e3f3f;
    ram_cell[    9863] = 32'h0;  // 32'h96e9bb39;
    ram_cell[    9864] = 32'h0;  // 32'h92ce5a12;
    ram_cell[    9865] = 32'h0;  // 32'hc210eae6;
    ram_cell[    9866] = 32'h0;  // 32'h1d3f2592;
    ram_cell[    9867] = 32'h0;  // 32'hd1f864be;
    ram_cell[    9868] = 32'h0;  // 32'hfed2f1c2;
    ram_cell[    9869] = 32'h0;  // 32'hfa585fab;
    ram_cell[    9870] = 32'h0;  // 32'h33436980;
    ram_cell[    9871] = 32'h0;  // 32'h3877a813;
    ram_cell[    9872] = 32'h0;  // 32'h3ceb7932;
    ram_cell[    9873] = 32'h0;  // 32'hb1617911;
    ram_cell[    9874] = 32'h0;  // 32'h563df42f;
    ram_cell[    9875] = 32'h0;  // 32'h6b0a6652;
    ram_cell[    9876] = 32'h0;  // 32'h2bec09c8;
    ram_cell[    9877] = 32'h0;  // 32'h04f9eb88;
    ram_cell[    9878] = 32'h0;  // 32'h98a990df;
    ram_cell[    9879] = 32'h0;  // 32'ha1bdf320;
    ram_cell[    9880] = 32'h0;  // 32'h2704e134;
    ram_cell[    9881] = 32'h0;  // 32'hf7bd1b24;
    ram_cell[    9882] = 32'h0;  // 32'h70093b5a;
    ram_cell[    9883] = 32'h0;  // 32'h6a45eef9;
    ram_cell[    9884] = 32'h0;  // 32'h9515b2d7;
    ram_cell[    9885] = 32'h0;  // 32'ha87e7a46;
    ram_cell[    9886] = 32'h0;  // 32'hcb8a4ec0;
    ram_cell[    9887] = 32'h0;  // 32'hf5ca68f9;
    ram_cell[    9888] = 32'h0;  // 32'h8c049067;
    ram_cell[    9889] = 32'h0;  // 32'h3a656685;
    ram_cell[    9890] = 32'h0;  // 32'ha51279d5;
    ram_cell[    9891] = 32'h0;  // 32'h08c6449b;
    ram_cell[    9892] = 32'h0;  // 32'h7afc807f;
    ram_cell[    9893] = 32'h0;  // 32'hbadd5786;
    ram_cell[    9894] = 32'h0;  // 32'h745ae2da;
    ram_cell[    9895] = 32'h0;  // 32'h9a5cc5a1;
    ram_cell[    9896] = 32'h0;  // 32'hd3a9bee2;
    ram_cell[    9897] = 32'h0;  // 32'h1ff6d08e;
    ram_cell[    9898] = 32'h0;  // 32'hc14255d6;
    ram_cell[    9899] = 32'h0;  // 32'hfa24091d;
    ram_cell[    9900] = 32'h0;  // 32'h0ae8da8a;
    ram_cell[    9901] = 32'h0;  // 32'h1d4f7529;
    ram_cell[    9902] = 32'h0;  // 32'h0a42f9a8;
    ram_cell[    9903] = 32'h0;  // 32'h8a29522e;
    ram_cell[    9904] = 32'h0;  // 32'h18851c7f;
    ram_cell[    9905] = 32'h0;  // 32'h250807ae;
    ram_cell[    9906] = 32'h0;  // 32'hd948b6a4;
    ram_cell[    9907] = 32'h0;  // 32'h615e0492;
    ram_cell[    9908] = 32'h0;  // 32'he7a25c14;
    ram_cell[    9909] = 32'h0;  // 32'h275a9ea9;
    ram_cell[    9910] = 32'h0;  // 32'hfff3105f;
    ram_cell[    9911] = 32'h0;  // 32'h491c7b1e;
    ram_cell[    9912] = 32'h0;  // 32'hfff28770;
    ram_cell[    9913] = 32'h0;  // 32'hada601a0;
    ram_cell[    9914] = 32'h0;  // 32'h4fc88f3a;
    ram_cell[    9915] = 32'h0;  // 32'h2c11187a;
    ram_cell[    9916] = 32'h0;  // 32'hb9dcfb53;
    ram_cell[    9917] = 32'h0;  // 32'h00db3295;
    ram_cell[    9918] = 32'h0;  // 32'hb054048e;
    ram_cell[    9919] = 32'h0;  // 32'hdec082a6;
    ram_cell[    9920] = 32'h0;  // 32'h158c8cb9;
    ram_cell[    9921] = 32'h0;  // 32'h73c3df6c;
    ram_cell[    9922] = 32'h0;  // 32'hfa86f7db;
    ram_cell[    9923] = 32'h0;  // 32'h255a4b99;
    ram_cell[    9924] = 32'h0;  // 32'h992e9250;
    ram_cell[    9925] = 32'h0;  // 32'hba8811be;
    ram_cell[    9926] = 32'h0;  // 32'h1982acfd;
    ram_cell[    9927] = 32'h0;  // 32'h0decd1ff;
    ram_cell[    9928] = 32'h0;  // 32'h5670b692;
    ram_cell[    9929] = 32'h0;  // 32'ha7b87a02;
    ram_cell[    9930] = 32'h0;  // 32'h6556940b;
    ram_cell[    9931] = 32'h0;  // 32'ha3bd8f67;
    ram_cell[    9932] = 32'h0;  // 32'haa065b44;
    ram_cell[    9933] = 32'h0;  // 32'hfc496791;
    ram_cell[    9934] = 32'h0;  // 32'hdf92009b;
    ram_cell[    9935] = 32'h0;  // 32'h3f0d8a8f;
    ram_cell[    9936] = 32'h0;  // 32'h75e31d5c;
    ram_cell[    9937] = 32'h0;  // 32'h18a90748;
    ram_cell[    9938] = 32'h0;  // 32'h2a901876;
    ram_cell[    9939] = 32'h0;  // 32'h9dcac66e;
    ram_cell[    9940] = 32'h0;  // 32'hace86936;
    ram_cell[    9941] = 32'h0;  // 32'hdefb2e19;
    ram_cell[    9942] = 32'h0;  // 32'ha773db68;
    ram_cell[    9943] = 32'h0;  // 32'h16a88afd;
    ram_cell[    9944] = 32'h0;  // 32'ha5468398;
    ram_cell[    9945] = 32'h0;  // 32'hf1042ffd;
    ram_cell[    9946] = 32'h0;  // 32'h2ed4cad2;
    ram_cell[    9947] = 32'h0;  // 32'hecb93924;
    ram_cell[    9948] = 32'h0;  // 32'hbd673528;
    ram_cell[    9949] = 32'h0;  // 32'h3fccb072;
    ram_cell[    9950] = 32'h0;  // 32'h6296768a;
    ram_cell[    9951] = 32'h0;  // 32'hde2a9ba2;
    ram_cell[    9952] = 32'h0;  // 32'h0fab4e91;
    ram_cell[    9953] = 32'h0;  // 32'ha2961ca0;
    ram_cell[    9954] = 32'h0;  // 32'h75ae2bb4;
    ram_cell[    9955] = 32'h0;  // 32'h8f2ab94d;
    ram_cell[    9956] = 32'h0;  // 32'hc2e81a7f;
    ram_cell[    9957] = 32'h0;  // 32'h17830ce4;
    ram_cell[    9958] = 32'h0;  // 32'hb34079fb;
    ram_cell[    9959] = 32'h0;  // 32'hf5f3850f;
    ram_cell[    9960] = 32'h0;  // 32'he2f07646;
    ram_cell[    9961] = 32'h0;  // 32'he4d83d43;
    ram_cell[    9962] = 32'h0;  // 32'h8d812c2f;
    ram_cell[    9963] = 32'h0;  // 32'h0af3a23b;
    ram_cell[    9964] = 32'h0;  // 32'h18663c4a;
    ram_cell[    9965] = 32'h0;  // 32'h60836a92;
    ram_cell[    9966] = 32'h0;  // 32'h320d53ca;
    ram_cell[    9967] = 32'h0;  // 32'h4d06c7f4;
    ram_cell[    9968] = 32'h0;  // 32'h639175b6;
    ram_cell[    9969] = 32'h0;  // 32'hdc1429a7;
    ram_cell[    9970] = 32'h0;  // 32'h61c2087b;
    ram_cell[    9971] = 32'h0;  // 32'h93a59757;
    ram_cell[    9972] = 32'h0;  // 32'ha83ac178;
    ram_cell[    9973] = 32'h0;  // 32'ha935f8bd;
    ram_cell[    9974] = 32'h0;  // 32'h290800c6;
    ram_cell[    9975] = 32'h0;  // 32'h604a3611;
    ram_cell[    9976] = 32'h0;  // 32'hb7a69937;
    ram_cell[    9977] = 32'h0;  // 32'h9b446d61;
    ram_cell[    9978] = 32'h0;  // 32'h3a48d84a;
    ram_cell[    9979] = 32'h0;  // 32'hfd81108f;
    ram_cell[    9980] = 32'h0;  // 32'h16cc2737;
    ram_cell[    9981] = 32'h0;  // 32'h0469272f;
    ram_cell[    9982] = 32'h0;  // 32'h6ce5ffc6;
    ram_cell[    9983] = 32'h0;  // 32'h5b2f9c66;
    ram_cell[    9984] = 32'h0;  // 32'h236a1f31;
    ram_cell[    9985] = 32'h0;  // 32'h1c91e446;
    ram_cell[    9986] = 32'h0;  // 32'h5035b251;
    ram_cell[    9987] = 32'h0;  // 32'hc2c83766;
    ram_cell[    9988] = 32'h0;  // 32'h1a4abfb1;
    ram_cell[    9989] = 32'h0;  // 32'h38c5a18e;
    ram_cell[    9990] = 32'h0;  // 32'h08f7621e;
    ram_cell[    9991] = 32'h0;  // 32'h53dc3642;
    ram_cell[    9992] = 32'h0;  // 32'hf699de4f;
    ram_cell[    9993] = 32'h0;  // 32'h56d4dfca;
    ram_cell[    9994] = 32'h0;  // 32'h6cc2436c;
    ram_cell[    9995] = 32'h0;  // 32'he7b1531e;
    ram_cell[    9996] = 32'h0;  // 32'hde408d2d;
    ram_cell[    9997] = 32'h0;  // 32'hb3195f82;
    ram_cell[    9998] = 32'h0;  // 32'he51019d3;
    ram_cell[    9999] = 32'h0;  // 32'hc014ae52;
    ram_cell[   10000] = 32'h0;  // 32'h8bc852f0;
    ram_cell[   10001] = 32'h0;  // 32'h09f55dbb;
    ram_cell[   10002] = 32'h0;  // 32'hf4e05c6c;
    ram_cell[   10003] = 32'h0;  // 32'h78c8663f;
    ram_cell[   10004] = 32'h0;  // 32'h252454f6;
    ram_cell[   10005] = 32'h0;  // 32'he871b113;
    ram_cell[   10006] = 32'h0;  // 32'h92e51df6;
    ram_cell[   10007] = 32'h0;  // 32'hfb0dbaa2;
    ram_cell[   10008] = 32'h0;  // 32'h2678599c;
    ram_cell[   10009] = 32'h0;  // 32'h35b8528d;
    ram_cell[   10010] = 32'h0;  // 32'h42c9c10b;
    ram_cell[   10011] = 32'h0;  // 32'h2c59892f;
    ram_cell[   10012] = 32'h0;  // 32'h52d036a7;
    ram_cell[   10013] = 32'h0;  // 32'h68db1552;
    ram_cell[   10014] = 32'h0;  // 32'h3dd6d8c9;
    ram_cell[   10015] = 32'h0;  // 32'hdb2ebb8f;
    ram_cell[   10016] = 32'h0;  // 32'hbbe5fc9e;
    ram_cell[   10017] = 32'h0;  // 32'hf080831e;
    ram_cell[   10018] = 32'h0;  // 32'h2f5053ed;
    ram_cell[   10019] = 32'h0;  // 32'hf380f623;
    ram_cell[   10020] = 32'h0;  // 32'hfd406009;
    ram_cell[   10021] = 32'h0;  // 32'h108d7118;
    ram_cell[   10022] = 32'h0;  // 32'he4150494;
    ram_cell[   10023] = 32'h0;  // 32'h49331e60;
    ram_cell[   10024] = 32'h0;  // 32'h094ea6b3;
    ram_cell[   10025] = 32'h0;  // 32'h0e7eb698;
    ram_cell[   10026] = 32'h0;  // 32'h1a4b47fc;
    ram_cell[   10027] = 32'h0;  // 32'h2721f55e;
    ram_cell[   10028] = 32'h0;  // 32'hd6bf5d69;
    ram_cell[   10029] = 32'h0;  // 32'hd8552b67;
    ram_cell[   10030] = 32'h0;  // 32'h506bcccb;
    ram_cell[   10031] = 32'h0;  // 32'h134dd92e;
    ram_cell[   10032] = 32'h0;  // 32'h58a6e367;
    ram_cell[   10033] = 32'h0;  // 32'h255d1ee2;
    ram_cell[   10034] = 32'h0;  // 32'h3f27e25e;
    ram_cell[   10035] = 32'h0;  // 32'h968503cc;
    ram_cell[   10036] = 32'h0;  // 32'h3fac90c9;
    ram_cell[   10037] = 32'h0;  // 32'h3d73bbf8;
    ram_cell[   10038] = 32'h0;  // 32'h54923a43;
    ram_cell[   10039] = 32'h0;  // 32'h3ec92611;
    ram_cell[   10040] = 32'h0;  // 32'h84486089;
    ram_cell[   10041] = 32'h0;  // 32'h852fe935;
    ram_cell[   10042] = 32'h0;  // 32'hf2643a14;
    ram_cell[   10043] = 32'h0;  // 32'h9b30d7d4;
    ram_cell[   10044] = 32'h0;  // 32'h517796aa;
    ram_cell[   10045] = 32'h0;  // 32'h6e847866;
    ram_cell[   10046] = 32'h0;  // 32'h41623cb8;
    ram_cell[   10047] = 32'h0;  // 32'h134c9297;
    ram_cell[   10048] = 32'h0;  // 32'h885a6b72;
    ram_cell[   10049] = 32'h0;  // 32'h078591d6;
    ram_cell[   10050] = 32'h0;  // 32'hf7d56b22;
    ram_cell[   10051] = 32'h0;  // 32'hf80d4524;
    ram_cell[   10052] = 32'h0;  // 32'h319ad304;
    ram_cell[   10053] = 32'h0;  // 32'hbf4c2d9c;
    ram_cell[   10054] = 32'h0;  // 32'h519e2c79;
    ram_cell[   10055] = 32'h0;  // 32'ha0fd8388;
    ram_cell[   10056] = 32'h0;  // 32'h2d9a4770;
    ram_cell[   10057] = 32'h0;  // 32'h7114102f;
    ram_cell[   10058] = 32'h0;  // 32'hc764e9d5;
    ram_cell[   10059] = 32'h0;  // 32'he97a5f7c;
    ram_cell[   10060] = 32'h0;  // 32'hc7c8a3c7;
    ram_cell[   10061] = 32'h0;  // 32'h66082711;
    ram_cell[   10062] = 32'h0;  // 32'h83e2c02f;
    ram_cell[   10063] = 32'h0;  // 32'h14007a9e;
    ram_cell[   10064] = 32'h0;  // 32'h0f44689a;
    ram_cell[   10065] = 32'h0;  // 32'h6aae75b7;
    ram_cell[   10066] = 32'h0;  // 32'h52d04423;
    ram_cell[   10067] = 32'h0;  // 32'hdb3728be;
    ram_cell[   10068] = 32'h0;  // 32'h83bac4a6;
    ram_cell[   10069] = 32'h0;  // 32'h4875a8a3;
    ram_cell[   10070] = 32'h0;  // 32'h70411e76;
    ram_cell[   10071] = 32'h0;  // 32'h837a0760;
    ram_cell[   10072] = 32'h0;  // 32'h68f00f05;
    ram_cell[   10073] = 32'h0;  // 32'h99ae33cd;
    ram_cell[   10074] = 32'h0;  // 32'h8ba9e98e;
    ram_cell[   10075] = 32'h0;  // 32'haf1f2510;
    ram_cell[   10076] = 32'h0;  // 32'hc818f0b0;
    ram_cell[   10077] = 32'h0;  // 32'h093d21d3;
    ram_cell[   10078] = 32'h0;  // 32'h73a38207;
    ram_cell[   10079] = 32'h0;  // 32'h07c85796;
    ram_cell[   10080] = 32'h0;  // 32'h193c1490;
    ram_cell[   10081] = 32'h0;  // 32'h4ff15a25;
    ram_cell[   10082] = 32'h0;  // 32'he0c876d1;
    ram_cell[   10083] = 32'h0;  // 32'hf5b51f46;
    ram_cell[   10084] = 32'h0;  // 32'h79fa6b37;
    ram_cell[   10085] = 32'h0;  // 32'he52b6cbe;
    ram_cell[   10086] = 32'h0;  // 32'h05a579a4;
    ram_cell[   10087] = 32'h0;  // 32'hc2e91e48;
    ram_cell[   10088] = 32'h0;  // 32'hc91fae7b;
    ram_cell[   10089] = 32'h0;  // 32'h9cb5a9c1;
    ram_cell[   10090] = 32'h0;  // 32'h14292e96;
    ram_cell[   10091] = 32'h0;  // 32'h4f7bf999;
    ram_cell[   10092] = 32'h0;  // 32'ha209334d;
    ram_cell[   10093] = 32'h0;  // 32'hbf50cd38;
    ram_cell[   10094] = 32'h0;  // 32'h8c8267e6;
    ram_cell[   10095] = 32'h0;  // 32'hbe9ed9a0;
    ram_cell[   10096] = 32'h0;  // 32'h451d97f5;
    ram_cell[   10097] = 32'h0;  // 32'h068e2160;
    ram_cell[   10098] = 32'h0;  // 32'hfccd8df7;
    ram_cell[   10099] = 32'h0;  // 32'h59c79c1d;
    ram_cell[   10100] = 32'h0;  // 32'h817e53b4;
    ram_cell[   10101] = 32'h0;  // 32'h0f4331a5;
    ram_cell[   10102] = 32'h0;  // 32'h010a2b62;
    ram_cell[   10103] = 32'h0;  // 32'hc18ffe83;
    ram_cell[   10104] = 32'h0;  // 32'h45ba8da5;
    ram_cell[   10105] = 32'h0;  // 32'h48be6acb;
    ram_cell[   10106] = 32'h0;  // 32'h1a316465;
    ram_cell[   10107] = 32'h0;  // 32'h28b3bc79;
    ram_cell[   10108] = 32'h0;  // 32'ha0e2de1d;
    ram_cell[   10109] = 32'h0;  // 32'h88ae80b1;
    ram_cell[   10110] = 32'h0;  // 32'h928e97c1;
    ram_cell[   10111] = 32'h0;  // 32'h1b8c1ae8;
    ram_cell[   10112] = 32'h0;  // 32'h261591a0;
    ram_cell[   10113] = 32'h0;  // 32'h87d4b79d;
    ram_cell[   10114] = 32'h0;  // 32'h27f7b980;
    ram_cell[   10115] = 32'h0;  // 32'h7f956a1b;
    ram_cell[   10116] = 32'h0;  // 32'hd0ac2490;
    ram_cell[   10117] = 32'h0;  // 32'h2ac001a0;
    ram_cell[   10118] = 32'h0;  // 32'h64252c08;
    ram_cell[   10119] = 32'h0;  // 32'h19c4961a;
    ram_cell[   10120] = 32'h0;  // 32'h913caf00;
    ram_cell[   10121] = 32'h0;  // 32'h817e3fbd;
    ram_cell[   10122] = 32'h0;  // 32'h98b1bcba;
    ram_cell[   10123] = 32'h0;  // 32'h7241583b;
    ram_cell[   10124] = 32'h0;  // 32'h834ef4b5;
    ram_cell[   10125] = 32'h0;  // 32'h12b716fe;
    ram_cell[   10126] = 32'h0;  // 32'h1adad97b;
    ram_cell[   10127] = 32'h0;  // 32'hffc673b9;
    ram_cell[   10128] = 32'h0;  // 32'hf9c396ef;
    ram_cell[   10129] = 32'h0;  // 32'h15ddda24;
    ram_cell[   10130] = 32'h0;  // 32'hf97b2cfc;
    ram_cell[   10131] = 32'h0;  // 32'h866af7f7;
    ram_cell[   10132] = 32'h0;  // 32'h976686ae;
    ram_cell[   10133] = 32'h0;  // 32'hc6b486c4;
    ram_cell[   10134] = 32'h0;  // 32'h6b3cfe83;
    ram_cell[   10135] = 32'h0;  // 32'hb8faeef5;
    ram_cell[   10136] = 32'h0;  // 32'h53635407;
    ram_cell[   10137] = 32'h0;  // 32'h2af94848;
    ram_cell[   10138] = 32'h0;  // 32'h8c041fda;
    ram_cell[   10139] = 32'h0;  // 32'haa34a9d0;
    ram_cell[   10140] = 32'h0;  // 32'h9c97be2d;
    ram_cell[   10141] = 32'h0;  // 32'h9973ac63;
    ram_cell[   10142] = 32'h0;  // 32'h98e36f13;
    ram_cell[   10143] = 32'h0;  // 32'h6941c39b;
    ram_cell[   10144] = 32'h0;  // 32'hfcb42cde;
    ram_cell[   10145] = 32'h0;  // 32'h2c5d8121;
    ram_cell[   10146] = 32'h0;  // 32'h02877433;
    ram_cell[   10147] = 32'h0;  // 32'h0b4856cd;
    ram_cell[   10148] = 32'h0;  // 32'h4cd8a2a3;
    ram_cell[   10149] = 32'h0;  // 32'h4e952324;
    ram_cell[   10150] = 32'h0;  // 32'hf32ced20;
    ram_cell[   10151] = 32'h0;  // 32'hdfcac8ef;
    ram_cell[   10152] = 32'h0;  // 32'hfdb8b8da;
    ram_cell[   10153] = 32'h0;  // 32'h49df6677;
    ram_cell[   10154] = 32'h0;  // 32'hd4c79da1;
    ram_cell[   10155] = 32'h0;  // 32'hd23bcf09;
    ram_cell[   10156] = 32'h0;  // 32'h4e347d61;
    ram_cell[   10157] = 32'h0;  // 32'h2d4ca56b;
    ram_cell[   10158] = 32'h0;  // 32'hfeb93ed2;
    ram_cell[   10159] = 32'h0;  // 32'h1934df76;
    ram_cell[   10160] = 32'h0;  // 32'h5d90d031;
    ram_cell[   10161] = 32'h0;  // 32'hf0b98125;
    ram_cell[   10162] = 32'h0;  // 32'h9df907ef;
    ram_cell[   10163] = 32'h0;  // 32'h1f9ab581;
    ram_cell[   10164] = 32'h0;  // 32'h360dbc46;
    ram_cell[   10165] = 32'h0;  // 32'he82a8eb0;
    ram_cell[   10166] = 32'h0;  // 32'h4d5b3355;
    ram_cell[   10167] = 32'h0;  // 32'h65cb1ccc;
    ram_cell[   10168] = 32'h0;  // 32'h476e19fa;
    ram_cell[   10169] = 32'h0;  // 32'h0b223448;
    ram_cell[   10170] = 32'h0;  // 32'h302a876b;
    ram_cell[   10171] = 32'h0;  // 32'hf50c2b23;
    ram_cell[   10172] = 32'h0;  // 32'hb1ae601b;
    ram_cell[   10173] = 32'h0;  // 32'he6dc4e71;
    ram_cell[   10174] = 32'h0;  // 32'h20f952c1;
    ram_cell[   10175] = 32'h0;  // 32'hac855bd3;
    ram_cell[   10176] = 32'h0;  // 32'hf483e819;
    ram_cell[   10177] = 32'h0;  // 32'h3e3eb09a;
    ram_cell[   10178] = 32'h0;  // 32'hc1c1d48f;
    ram_cell[   10179] = 32'h0;  // 32'hb87fc28c;
    ram_cell[   10180] = 32'h0;  // 32'h66eeaae1;
    ram_cell[   10181] = 32'h0;  // 32'h6343429d;
    ram_cell[   10182] = 32'h0;  // 32'hdb0d6359;
    ram_cell[   10183] = 32'h0;  // 32'h8d360ecd;
    ram_cell[   10184] = 32'h0;  // 32'h3d1caf68;
    ram_cell[   10185] = 32'h0;  // 32'h7c14a2ea;
    ram_cell[   10186] = 32'h0;  // 32'h42fde899;
    ram_cell[   10187] = 32'h0;  // 32'h5ad7a999;
    ram_cell[   10188] = 32'h0;  // 32'h909b6ff4;
    ram_cell[   10189] = 32'h0;  // 32'hd98f5af9;
    ram_cell[   10190] = 32'h0;  // 32'ha8403037;
    ram_cell[   10191] = 32'h0;  // 32'hf951fdef;
    ram_cell[   10192] = 32'h0;  // 32'h1823583c;
    ram_cell[   10193] = 32'h0;  // 32'h10361cd5;
    ram_cell[   10194] = 32'h0;  // 32'h61763041;
    ram_cell[   10195] = 32'h0;  // 32'h575c8727;
    ram_cell[   10196] = 32'h0;  // 32'h527e5f73;
    ram_cell[   10197] = 32'h0;  // 32'he937f69e;
    ram_cell[   10198] = 32'h0;  // 32'h05cbb22a;
    ram_cell[   10199] = 32'h0;  // 32'hee0aa95b;
    ram_cell[   10200] = 32'h0;  // 32'h32cb500a;
    ram_cell[   10201] = 32'h0;  // 32'h0596ef4e;
    ram_cell[   10202] = 32'h0;  // 32'hd93a83c7;
    ram_cell[   10203] = 32'h0;  // 32'hc5a6546c;
    ram_cell[   10204] = 32'h0;  // 32'hf4a87128;
    ram_cell[   10205] = 32'h0;  // 32'h15cf9d37;
    ram_cell[   10206] = 32'h0;  // 32'h016dfc4c;
    ram_cell[   10207] = 32'h0;  // 32'h89c22af4;
    ram_cell[   10208] = 32'h0;  // 32'hc3cbb9f5;
    ram_cell[   10209] = 32'h0;  // 32'hb67b56f7;
    ram_cell[   10210] = 32'h0;  // 32'hd94f6fdf;
    ram_cell[   10211] = 32'h0;  // 32'h1a8c8e36;
    ram_cell[   10212] = 32'h0;  // 32'h2fa874c7;
    ram_cell[   10213] = 32'h0;  // 32'h5423a342;
    ram_cell[   10214] = 32'h0;  // 32'hf90fe7c0;
    ram_cell[   10215] = 32'h0;  // 32'h5fbff3b8;
    ram_cell[   10216] = 32'h0;  // 32'h46f6d821;
    ram_cell[   10217] = 32'h0;  // 32'h469f1ce6;
    ram_cell[   10218] = 32'h0;  // 32'h39e65ff2;
    ram_cell[   10219] = 32'h0;  // 32'h9ccf4803;
    ram_cell[   10220] = 32'h0;  // 32'hec52954b;
    ram_cell[   10221] = 32'h0;  // 32'h0a566907;
    ram_cell[   10222] = 32'h0;  // 32'h04e53174;
    ram_cell[   10223] = 32'h0;  // 32'hb13080b5;
    ram_cell[   10224] = 32'h0;  // 32'h54aa4a5d;
    ram_cell[   10225] = 32'h0;  // 32'he3d49b33;
    ram_cell[   10226] = 32'h0;  // 32'h205f690b;
    ram_cell[   10227] = 32'h0;  // 32'hef1ad4bf;
    ram_cell[   10228] = 32'h0;  // 32'h6d9d1e69;
    ram_cell[   10229] = 32'h0;  // 32'h44af9cdd;
    ram_cell[   10230] = 32'h0;  // 32'he0a2e3c9;
    ram_cell[   10231] = 32'h0;  // 32'h4c6a8acf;
    ram_cell[   10232] = 32'h0;  // 32'h75dfbc30;
    ram_cell[   10233] = 32'h0;  // 32'heb10de8c;
    ram_cell[   10234] = 32'h0;  // 32'h36049da1;
    ram_cell[   10235] = 32'h0;  // 32'hfa73a6ea;
    ram_cell[   10236] = 32'h0;  // 32'h3903acba;
    ram_cell[   10237] = 32'h0;  // 32'hef6249aa;
    ram_cell[   10238] = 32'h0;  // 32'h6fde42e4;
    ram_cell[   10239] = 32'h0;  // 32'h76b42a76;
    ram_cell[   10240] = 32'h0;  // 32'hdad6c210;
    ram_cell[   10241] = 32'h0;  // 32'h7432edc2;
    ram_cell[   10242] = 32'h0;  // 32'h50d442da;
    ram_cell[   10243] = 32'h0;  // 32'h12441834;
    ram_cell[   10244] = 32'h0;  // 32'h3614c101;
    ram_cell[   10245] = 32'h0;  // 32'h3295d3b9;
    ram_cell[   10246] = 32'h0;  // 32'h73d75110;
    ram_cell[   10247] = 32'h0;  // 32'hbfb96c6d;
    ram_cell[   10248] = 32'h0;  // 32'hf4191c04;
    ram_cell[   10249] = 32'h0;  // 32'h3f6f3264;
    ram_cell[   10250] = 32'h0;  // 32'hf08dcef1;
    ram_cell[   10251] = 32'h0;  // 32'h7e1d02a5;
    ram_cell[   10252] = 32'h0;  // 32'hc02ea8b7;
    ram_cell[   10253] = 32'h0;  // 32'had312a1b;
    ram_cell[   10254] = 32'h0;  // 32'hbee7c2da;
    ram_cell[   10255] = 32'h0;  // 32'hc2331e46;
    ram_cell[   10256] = 32'h0;  // 32'h18fc7e1d;
    ram_cell[   10257] = 32'h0;  // 32'h635260cb;
    ram_cell[   10258] = 32'h0;  // 32'hce6cd7b6;
    ram_cell[   10259] = 32'h0;  // 32'h2214b865;
    ram_cell[   10260] = 32'h0;  // 32'hc2f03c8d;
    ram_cell[   10261] = 32'h0;  // 32'h619fb08a;
    ram_cell[   10262] = 32'h0;  // 32'h92733d79;
    ram_cell[   10263] = 32'h0;  // 32'h36784d0c;
    ram_cell[   10264] = 32'h0;  // 32'h5553f344;
    ram_cell[   10265] = 32'h0;  // 32'hbc66c734;
    ram_cell[   10266] = 32'h0;  // 32'h3c6c9d1f;
    ram_cell[   10267] = 32'h0;  // 32'h7a853560;
    ram_cell[   10268] = 32'h0;  // 32'hf003f474;
    ram_cell[   10269] = 32'h0;  // 32'h3fe95a2c;
    ram_cell[   10270] = 32'h0;  // 32'hf61ac24e;
    ram_cell[   10271] = 32'h0;  // 32'h87fe3e3d;
    ram_cell[   10272] = 32'h0;  // 32'h6c51a9d6;
    ram_cell[   10273] = 32'h0;  // 32'h3877d432;
    ram_cell[   10274] = 32'h0;  // 32'hd21453a3;
    ram_cell[   10275] = 32'h0;  // 32'h7f6d8932;
    ram_cell[   10276] = 32'h0;  // 32'h2ed97bc6;
    ram_cell[   10277] = 32'h0;  // 32'h47fea90a;
    ram_cell[   10278] = 32'h0;  // 32'h4c4023b9;
    ram_cell[   10279] = 32'h0;  // 32'h53e3daae;
    ram_cell[   10280] = 32'h0;  // 32'h6a1d9e68;
    ram_cell[   10281] = 32'h0;  // 32'hc2d6d2df;
    ram_cell[   10282] = 32'h0;  // 32'h0923939a;
    ram_cell[   10283] = 32'h0;  // 32'h283b34f9;
    ram_cell[   10284] = 32'h0;  // 32'h9bd117fc;
    ram_cell[   10285] = 32'h0;  // 32'h01df291c;
    ram_cell[   10286] = 32'h0;  // 32'h5814f01b;
    ram_cell[   10287] = 32'h0;  // 32'haea99129;
    ram_cell[   10288] = 32'h0;  // 32'h980356d3;
    ram_cell[   10289] = 32'h0;  // 32'h0d15d328;
    ram_cell[   10290] = 32'h0;  // 32'hc147d437;
    ram_cell[   10291] = 32'h0;  // 32'h2c8cd6ab;
    ram_cell[   10292] = 32'h0;  // 32'h8fd8261c;
    ram_cell[   10293] = 32'h0;  // 32'h586e33ce;
    ram_cell[   10294] = 32'h0;  // 32'h0e99e8af;
    ram_cell[   10295] = 32'h0;  // 32'h3c7bc842;
    ram_cell[   10296] = 32'h0;  // 32'h54e8463a;
    ram_cell[   10297] = 32'h0;  // 32'hed01be82;
    ram_cell[   10298] = 32'h0;  // 32'hf2f3cde0;
    ram_cell[   10299] = 32'h0;  // 32'h0a135801;
    ram_cell[   10300] = 32'h0;  // 32'h6adab801;
    ram_cell[   10301] = 32'h0;  // 32'h6d3b29f9;
    ram_cell[   10302] = 32'h0;  // 32'h7aca5e19;
    ram_cell[   10303] = 32'h0;  // 32'ha0ec7d8e;
    ram_cell[   10304] = 32'h0;  // 32'h16554302;
    ram_cell[   10305] = 32'h0;  // 32'h5743088e;
    ram_cell[   10306] = 32'h0;  // 32'h588f6b80;
    ram_cell[   10307] = 32'h0;  // 32'h1618139e;
    ram_cell[   10308] = 32'h0;  // 32'h42dd56ec;
    ram_cell[   10309] = 32'h0;  // 32'h74aff401;
    ram_cell[   10310] = 32'h0;  // 32'h70aa622a;
    ram_cell[   10311] = 32'h0;  // 32'h423a64b0;
    ram_cell[   10312] = 32'h0;  // 32'h0d74ec91;
    ram_cell[   10313] = 32'h0;  // 32'h41d553d5;
    ram_cell[   10314] = 32'h0;  // 32'h25a7c89f;
    ram_cell[   10315] = 32'h0;  // 32'hd596fc38;
    ram_cell[   10316] = 32'h0;  // 32'hd91ff68d;
    ram_cell[   10317] = 32'h0;  // 32'h2ea65137;
    ram_cell[   10318] = 32'h0;  // 32'hf122a923;
    ram_cell[   10319] = 32'h0;  // 32'h696c1f0e;
    ram_cell[   10320] = 32'h0;  // 32'h9ef37e3c;
    ram_cell[   10321] = 32'h0;  // 32'h3db15868;
    ram_cell[   10322] = 32'h0;  // 32'h91ee7b9e;
    ram_cell[   10323] = 32'h0;  // 32'ha1c0da82;
    ram_cell[   10324] = 32'h0;  // 32'he1657e47;
    ram_cell[   10325] = 32'h0;  // 32'hf9b0bf3f;
    ram_cell[   10326] = 32'h0;  // 32'h94afeebe;
    ram_cell[   10327] = 32'h0;  // 32'h8f8a825d;
    ram_cell[   10328] = 32'h0;  // 32'hdc7feb3b;
    ram_cell[   10329] = 32'h0;  // 32'h765e62bf;
    ram_cell[   10330] = 32'h0;  // 32'h58ae7025;
    ram_cell[   10331] = 32'h0;  // 32'hfaaf3730;
    ram_cell[   10332] = 32'h0;  // 32'hbf6cc97e;
    ram_cell[   10333] = 32'h0;  // 32'h31913b89;
    ram_cell[   10334] = 32'h0;  // 32'h09832a00;
    ram_cell[   10335] = 32'h0;  // 32'hcfd0a632;
    ram_cell[   10336] = 32'h0;  // 32'h5ca85fb1;
    ram_cell[   10337] = 32'h0;  // 32'haa300aa6;
    ram_cell[   10338] = 32'h0;  // 32'hc5580849;
    ram_cell[   10339] = 32'h0;  // 32'hfaf7dd65;
    ram_cell[   10340] = 32'h0;  // 32'h8bec8b61;
    ram_cell[   10341] = 32'h0;  // 32'hcffd9e00;
    ram_cell[   10342] = 32'h0;  // 32'h58ba4bfa;
    ram_cell[   10343] = 32'h0;  // 32'h9ff96a98;
    ram_cell[   10344] = 32'h0;  // 32'h717f9936;
    ram_cell[   10345] = 32'h0;  // 32'hc9b9d73f;
    ram_cell[   10346] = 32'h0;  // 32'hecc41a0e;
    ram_cell[   10347] = 32'h0;  // 32'h95fa1d69;
    ram_cell[   10348] = 32'h0;  // 32'h88ef78d0;
    ram_cell[   10349] = 32'h0;  // 32'h56226629;
    ram_cell[   10350] = 32'h0;  // 32'hb63e016c;
    ram_cell[   10351] = 32'h0;  // 32'h3b1f4382;
    ram_cell[   10352] = 32'h0;  // 32'h239afe6f;
    ram_cell[   10353] = 32'h0;  // 32'h5e256536;
    ram_cell[   10354] = 32'h0;  // 32'hb378e741;
    ram_cell[   10355] = 32'h0;  // 32'h34b2d8b7;
    ram_cell[   10356] = 32'h0;  // 32'hfb8f9b5f;
    ram_cell[   10357] = 32'h0;  // 32'h3464ddfc;
    ram_cell[   10358] = 32'h0;  // 32'h82292797;
    ram_cell[   10359] = 32'h0;  // 32'h7908f13f;
    ram_cell[   10360] = 32'h0;  // 32'hfeac470b;
    ram_cell[   10361] = 32'h0;  // 32'hd8495c06;
    ram_cell[   10362] = 32'h0;  // 32'hf3b5f79e;
    ram_cell[   10363] = 32'h0;  // 32'h057c1d54;
    ram_cell[   10364] = 32'h0;  // 32'hf2fdd7d7;
    ram_cell[   10365] = 32'h0;  // 32'h016f2140;
    ram_cell[   10366] = 32'h0;  // 32'h1ffe1fa2;
    ram_cell[   10367] = 32'h0;  // 32'h94ba3413;
    ram_cell[   10368] = 32'h0;  // 32'hba6b2ba4;
    ram_cell[   10369] = 32'h0;  // 32'h401dcf2b;
    ram_cell[   10370] = 32'h0;  // 32'h2bcdf31b;
    ram_cell[   10371] = 32'h0;  // 32'h14caca86;
    ram_cell[   10372] = 32'h0;  // 32'h01abc040;
    ram_cell[   10373] = 32'h0;  // 32'heca4417c;
    ram_cell[   10374] = 32'h0;  // 32'h1ece94b0;
    ram_cell[   10375] = 32'h0;  // 32'h0bf237db;
    ram_cell[   10376] = 32'h0;  // 32'hb88c1ef5;
    ram_cell[   10377] = 32'h0;  // 32'h37567469;
    ram_cell[   10378] = 32'h0;  // 32'hf340ffbc;
    ram_cell[   10379] = 32'h0;  // 32'hbb93f557;
    ram_cell[   10380] = 32'h0;  // 32'h7cddde79;
    ram_cell[   10381] = 32'h0;  // 32'haca11c58;
    ram_cell[   10382] = 32'h0;  // 32'he24e813c;
    ram_cell[   10383] = 32'h0;  // 32'h248468e6;
    ram_cell[   10384] = 32'h0;  // 32'hdf35428b;
    ram_cell[   10385] = 32'h0;  // 32'h4cc7dc76;
    ram_cell[   10386] = 32'h0;  // 32'haa05f189;
    ram_cell[   10387] = 32'h0;  // 32'h12ecd7e3;
    ram_cell[   10388] = 32'h0;  // 32'hed3de4e2;
    ram_cell[   10389] = 32'h0;  // 32'hf499d313;
    ram_cell[   10390] = 32'h0;  // 32'hd70e31ab;
    ram_cell[   10391] = 32'h0;  // 32'h7fd3723b;
    ram_cell[   10392] = 32'h0;  // 32'h8f8ea75f;
    ram_cell[   10393] = 32'h0;  // 32'hed8f80a4;
    ram_cell[   10394] = 32'h0;  // 32'hfc262458;
    ram_cell[   10395] = 32'h0;  // 32'h43ba9364;
    ram_cell[   10396] = 32'h0;  // 32'h3af1164c;
    ram_cell[   10397] = 32'h0;  // 32'h34783ffb;
    ram_cell[   10398] = 32'h0;  // 32'hcfbe5dbc;
    ram_cell[   10399] = 32'h0;  // 32'h8283516f;
    ram_cell[   10400] = 32'h0;  // 32'h217cddfa;
    ram_cell[   10401] = 32'h0;  // 32'h2840a838;
    ram_cell[   10402] = 32'h0;  // 32'hdec6d0cf;
    ram_cell[   10403] = 32'h0;  // 32'hc73dabe9;
    ram_cell[   10404] = 32'h0;  // 32'h50a0fdb7;
    ram_cell[   10405] = 32'h0;  // 32'h8a30cb78;
    ram_cell[   10406] = 32'h0;  // 32'h42a655b9;
    ram_cell[   10407] = 32'h0;  // 32'h3289c410;
    ram_cell[   10408] = 32'h0;  // 32'h99948bc2;
    ram_cell[   10409] = 32'h0;  // 32'hd3db7837;
    ram_cell[   10410] = 32'h0;  // 32'hcc4d2205;
    ram_cell[   10411] = 32'h0;  // 32'h717982b4;
    ram_cell[   10412] = 32'h0;  // 32'heaf48103;
    ram_cell[   10413] = 32'h0;  // 32'hdcfbfcfe;
    ram_cell[   10414] = 32'h0;  // 32'h4dadf0a0;
    ram_cell[   10415] = 32'h0;  // 32'h87260e2b;
    ram_cell[   10416] = 32'h0;  // 32'h66dd436f;
    ram_cell[   10417] = 32'h0;  // 32'h81f09f45;
    ram_cell[   10418] = 32'h0;  // 32'h9e9d0487;
    ram_cell[   10419] = 32'h0;  // 32'h6ffcad21;
    ram_cell[   10420] = 32'h0;  // 32'h16aa42e5;
    ram_cell[   10421] = 32'h0;  // 32'hdae3ea33;
    ram_cell[   10422] = 32'h0;  // 32'h8400be2c;
    ram_cell[   10423] = 32'h0;  // 32'he6de39e5;
    ram_cell[   10424] = 32'h0;  // 32'h79734360;
    ram_cell[   10425] = 32'h0;  // 32'hc8454893;
    ram_cell[   10426] = 32'h0;  // 32'hed786653;
    ram_cell[   10427] = 32'h0;  // 32'hbdbaf1e7;
    ram_cell[   10428] = 32'h0;  // 32'hb5091445;
    ram_cell[   10429] = 32'h0;  // 32'hbe17e743;
    ram_cell[   10430] = 32'h0;  // 32'h5fbd0279;
    ram_cell[   10431] = 32'h0;  // 32'h9ad934f9;
    ram_cell[   10432] = 32'h0;  // 32'h435085f3;
    ram_cell[   10433] = 32'h0;  // 32'h965a64bf;
    ram_cell[   10434] = 32'h0;  // 32'hc369a920;
    ram_cell[   10435] = 32'h0;  // 32'h77418b0b;
    ram_cell[   10436] = 32'h0;  // 32'h069a308a;
    ram_cell[   10437] = 32'h0;  // 32'h4c54ac40;
    ram_cell[   10438] = 32'h0;  // 32'hb4c406ee;
    ram_cell[   10439] = 32'h0;  // 32'h58b38287;
    ram_cell[   10440] = 32'h0;  // 32'h61384924;
    ram_cell[   10441] = 32'h0;  // 32'h5c570b06;
    ram_cell[   10442] = 32'h0;  // 32'he11951e5;
    ram_cell[   10443] = 32'h0;  // 32'he6dc0cd8;
    ram_cell[   10444] = 32'h0;  // 32'h1d12bc12;
    ram_cell[   10445] = 32'h0;  // 32'h7c2c74a1;
    ram_cell[   10446] = 32'h0;  // 32'h0e40044b;
    ram_cell[   10447] = 32'h0;  // 32'hb8891107;
    ram_cell[   10448] = 32'h0;  // 32'h88779403;
    ram_cell[   10449] = 32'h0;  // 32'h206599f7;
    ram_cell[   10450] = 32'h0;  // 32'hda6fd715;
    ram_cell[   10451] = 32'h0;  // 32'hf2548d39;
    ram_cell[   10452] = 32'h0;  // 32'h3b9a836c;
    ram_cell[   10453] = 32'h0;  // 32'heb9ce2cc;
    ram_cell[   10454] = 32'h0;  // 32'h105ed7ae;
    ram_cell[   10455] = 32'h0;  // 32'h34e16bb9;
    ram_cell[   10456] = 32'h0;  // 32'h82e810e1;
    ram_cell[   10457] = 32'h0;  // 32'h3f863280;
    ram_cell[   10458] = 32'h0;  // 32'h3f4a0bfa;
    ram_cell[   10459] = 32'h0;  // 32'h6d618524;
    ram_cell[   10460] = 32'h0;  // 32'h29f20f0c;
    ram_cell[   10461] = 32'h0;  // 32'h8fdba767;
    ram_cell[   10462] = 32'h0;  // 32'h4ffc2bd8;
    ram_cell[   10463] = 32'h0;  // 32'h403b0bf8;
    ram_cell[   10464] = 32'h0;  // 32'h7712a052;
    ram_cell[   10465] = 32'h0;  // 32'h504ad1d5;
    ram_cell[   10466] = 32'h0;  // 32'h80b2bf46;
    ram_cell[   10467] = 32'h0;  // 32'hf46fd528;
    ram_cell[   10468] = 32'h0;  // 32'hb0d25ec9;
    ram_cell[   10469] = 32'h0;  // 32'hc87d5315;
    ram_cell[   10470] = 32'h0;  // 32'h61aff8f0;
    ram_cell[   10471] = 32'h0;  // 32'h6167e352;
    ram_cell[   10472] = 32'h0;  // 32'ha88955c6;
    ram_cell[   10473] = 32'h0;  // 32'hd8417b54;
    ram_cell[   10474] = 32'h0;  // 32'h69325cff;
    ram_cell[   10475] = 32'h0;  // 32'hf7994bbf;
    ram_cell[   10476] = 32'h0;  // 32'hc068090d;
    ram_cell[   10477] = 32'h0;  // 32'h4f525300;
    ram_cell[   10478] = 32'h0;  // 32'h0d23a207;
    ram_cell[   10479] = 32'h0;  // 32'h068fe435;
    ram_cell[   10480] = 32'h0;  // 32'h03a8679b;
    ram_cell[   10481] = 32'h0;  // 32'h8a32a5ed;
    ram_cell[   10482] = 32'h0;  // 32'h0b3f5890;
    ram_cell[   10483] = 32'h0;  // 32'hd80357f7;
    ram_cell[   10484] = 32'h0;  // 32'h690156d2;
    ram_cell[   10485] = 32'h0;  // 32'h9a7e5782;
    ram_cell[   10486] = 32'h0;  // 32'h1e41a2d9;
    ram_cell[   10487] = 32'h0;  // 32'h0014c9f8;
    ram_cell[   10488] = 32'h0;  // 32'hcc9a6361;
    ram_cell[   10489] = 32'h0;  // 32'h067b668e;
    ram_cell[   10490] = 32'h0;  // 32'h1453724d;
    ram_cell[   10491] = 32'h0;  // 32'h790d9f4f;
    ram_cell[   10492] = 32'h0;  // 32'h851c5b0e;
    ram_cell[   10493] = 32'h0;  // 32'h2c791fbc;
    ram_cell[   10494] = 32'h0;  // 32'ha2abd560;
    ram_cell[   10495] = 32'h0;  // 32'ha45dc3c8;
    ram_cell[   10496] = 32'h0;  // 32'ha2c61bfb;
    ram_cell[   10497] = 32'h0;  // 32'h1c93dbaa;
    ram_cell[   10498] = 32'h0;  // 32'h4fd362e2;
    ram_cell[   10499] = 32'h0;  // 32'h3303b93d;
    ram_cell[   10500] = 32'h0;  // 32'h3b428d74;
    ram_cell[   10501] = 32'h0;  // 32'h08415c39;
    ram_cell[   10502] = 32'h0;  // 32'h6ac22027;
    ram_cell[   10503] = 32'h0;  // 32'h382a0af3;
    ram_cell[   10504] = 32'h0;  // 32'h77fd09b3;
    ram_cell[   10505] = 32'h0;  // 32'had8a615c;
    ram_cell[   10506] = 32'h0;  // 32'h4e5b4fe0;
    ram_cell[   10507] = 32'h0;  // 32'h4ca09115;
    ram_cell[   10508] = 32'h0;  // 32'h622e1584;
    ram_cell[   10509] = 32'h0;  // 32'h7b4ad927;
    ram_cell[   10510] = 32'h0;  // 32'hf4d36e29;
    ram_cell[   10511] = 32'h0;  // 32'hced35eae;
    ram_cell[   10512] = 32'h0;  // 32'h3ff300f9;
    ram_cell[   10513] = 32'h0;  // 32'he64a7a49;
    ram_cell[   10514] = 32'h0;  // 32'hd3f79a8e;
    ram_cell[   10515] = 32'h0;  // 32'h20d3f6da;
    ram_cell[   10516] = 32'h0;  // 32'h2fba1a07;
    ram_cell[   10517] = 32'h0;  // 32'h9f25e467;
    ram_cell[   10518] = 32'h0;  // 32'h71328ebc;
    ram_cell[   10519] = 32'h0;  // 32'h191a641c;
    ram_cell[   10520] = 32'h0;  // 32'h5c53a22d;
    ram_cell[   10521] = 32'h0;  // 32'he6c1e5fd;
    ram_cell[   10522] = 32'h0;  // 32'h14480985;
    ram_cell[   10523] = 32'h0;  // 32'hfa43fd02;
    ram_cell[   10524] = 32'h0;  // 32'h26f8d343;
    ram_cell[   10525] = 32'h0;  // 32'h0b4cbe4c;
    ram_cell[   10526] = 32'h0;  // 32'h812b4f17;
    ram_cell[   10527] = 32'h0;  // 32'hc7dea0ac;
    ram_cell[   10528] = 32'h0;  // 32'hd8a0c6c3;
    ram_cell[   10529] = 32'h0;  // 32'hcdc054ab;
    ram_cell[   10530] = 32'h0;  // 32'h981ee929;
    ram_cell[   10531] = 32'h0;  // 32'h7270085f;
    ram_cell[   10532] = 32'h0;  // 32'h56519d81;
    ram_cell[   10533] = 32'h0;  // 32'hbad9cf49;
    ram_cell[   10534] = 32'h0;  // 32'h59e73387;
    ram_cell[   10535] = 32'h0;  // 32'h69d556ee;
    ram_cell[   10536] = 32'h0;  // 32'h109a2359;
    ram_cell[   10537] = 32'h0;  // 32'h6133cb02;
    ram_cell[   10538] = 32'h0;  // 32'h74917fe2;
    ram_cell[   10539] = 32'h0;  // 32'hf62b98de;
    ram_cell[   10540] = 32'h0;  // 32'h0b628e14;
    ram_cell[   10541] = 32'h0;  // 32'h17d6b0e7;
    ram_cell[   10542] = 32'h0;  // 32'hf0b92318;
    ram_cell[   10543] = 32'h0;  // 32'h338f35f1;
    ram_cell[   10544] = 32'h0;  // 32'h7adbd70c;
    ram_cell[   10545] = 32'h0;  // 32'hda2cb7ce;
    ram_cell[   10546] = 32'h0;  // 32'haa2d665a;
    ram_cell[   10547] = 32'h0;  // 32'h4ccb872f;
    ram_cell[   10548] = 32'h0;  // 32'h471f2329;
    ram_cell[   10549] = 32'h0;  // 32'h9a92a529;
    ram_cell[   10550] = 32'h0;  // 32'h43718311;
    ram_cell[   10551] = 32'h0;  // 32'h617eecbe;
    ram_cell[   10552] = 32'h0;  // 32'h630f7028;
    ram_cell[   10553] = 32'h0;  // 32'hd141c9c1;
    ram_cell[   10554] = 32'h0;  // 32'h6a94d9f9;
    ram_cell[   10555] = 32'h0;  // 32'h1f546af3;
    ram_cell[   10556] = 32'h0;  // 32'h3f8d014c;
    ram_cell[   10557] = 32'h0;  // 32'hbabda20b;
    ram_cell[   10558] = 32'h0;  // 32'h9f92aed9;
    ram_cell[   10559] = 32'h0;  // 32'h004325d3;
    ram_cell[   10560] = 32'h0;  // 32'h0509fc5a;
    ram_cell[   10561] = 32'h0;  // 32'h1ecd323e;
    ram_cell[   10562] = 32'h0;  // 32'ha525abaf;
    ram_cell[   10563] = 32'h0;  // 32'h57ccb565;
    ram_cell[   10564] = 32'h0;  // 32'h011855f8;
    ram_cell[   10565] = 32'h0;  // 32'hb842ccd5;
    ram_cell[   10566] = 32'h0;  // 32'h055a52dc;
    ram_cell[   10567] = 32'h0;  // 32'h0bafd045;
    ram_cell[   10568] = 32'h0;  // 32'h76e4d1f9;
    ram_cell[   10569] = 32'h0;  // 32'h1e107f98;
    ram_cell[   10570] = 32'h0;  // 32'hdfa1b496;
    ram_cell[   10571] = 32'h0;  // 32'hf326a1f8;
    ram_cell[   10572] = 32'h0;  // 32'h08045eaf;
    ram_cell[   10573] = 32'h0;  // 32'hb29fc28e;
    ram_cell[   10574] = 32'h0;  // 32'h40594b4c;
    ram_cell[   10575] = 32'h0;  // 32'hccede4ee;
    ram_cell[   10576] = 32'h0;  // 32'hf8870ea6;
    ram_cell[   10577] = 32'h0;  // 32'h545e46c5;
    ram_cell[   10578] = 32'h0;  // 32'h3e35ba9d;
    ram_cell[   10579] = 32'h0;  // 32'hf942fff5;
    ram_cell[   10580] = 32'h0;  // 32'h17c3171b;
    ram_cell[   10581] = 32'h0;  // 32'h628b283f;
    ram_cell[   10582] = 32'h0;  // 32'h1ebc2d3f;
    ram_cell[   10583] = 32'h0;  // 32'h090096ea;
    ram_cell[   10584] = 32'h0;  // 32'hb9b2f9e9;
    ram_cell[   10585] = 32'h0;  // 32'h465c80ce;
    ram_cell[   10586] = 32'h0;  // 32'h39d528fd;
    ram_cell[   10587] = 32'h0;  // 32'h703bb77d;
    ram_cell[   10588] = 32'h0;  // 32'h62f3f48f;
    ram_cell[   10589] = 32'h0;  // 32'h8a4bec35;
    ram_cell[   10590] = 32'h0;  // 32'h4fe39426;
    ram_cell[   10591] = 32'h0;  // 32'hf7601ad5;
    ram_cell[   10592] = 32'h0;  // 32'hea21799d;
    ram_cell[   10593] = 32'h0;  // 32'hc48a1be2;
    ram_cell[   10594] = 32'h0;  // 32'h83f004f4;
    ram_cell[   10595] = 32'h0;  // 32'h72dffb98;
    ram_cell[   10596] = 32'h0;  // 32'h788e83e8;
    ram_cell[   10597] = 32'h0;  // 32'h235160f4;
    ram_cell[   10598] = 32'h0;  // 32'hf96159ce;
    ram_cell[   10599] = 32'h0;  // 32'h8e76f207;
    ram_cell[   10600] = 32'h0;  // 32'he5da26b6;
    ram_cell[   10601] = 32'h0;  // 32'h2a8fa9ed;
    ram_cell[   10602] = 32'h0;  // 32'hdd6d8b34;
    ram_cell[   10603] = 32'h0;  // 32'hf7ce16b6;
    ram_cell[   10604] = 32'h0;  // 32'h993aea04;
    ram_cell[   10605] = 32'h0;  // 32'hef27412a;
    ram_cell[   10606] = 32'h0;  // 32'h6ed55faf;
    ram_cell[   10607] = 32'h0;  // 32'h6ca6d530;
    ram_cell[   10608] = 32'h0;  // 32'h7cc97af9;
    ram_cell[   10609] = 32'h0;  // 32'h0227b670;
    ram_cell[   10610] = 32'h0;  // 32'ha98f09db;
    ram_cell[   10611] = 32'h0;  // 32'h075ff6d9;
    ram_cell[   10612] = 32'h0;  // 32'hd067adcc;
    ram_cell[   10613] = 32'h0;  // 32'h944675bd;
    ram_cell[   10614] = 32'h0;  // 32'h87dd39ba;
    ram_cell[   10615] = 32'h0;  // 32'h63a51a17;
    ram_cell[   10616] = 32'h0;  // 32'h99b4cdfd;
    ram_cell[   10617] = 32'h0;  // 32'ha5bc8d45;
    ram_cell[   10618] = 32'h0;  // 32'hbd16db69;
    ram_cell[   10619] = 32'h0;  // 32'hb8e13fed;
    ram_cell[   10620] = 32'h0;  // 32'h3ad7bab4;
    ram_cell[   10621] = 32'h0;  // 32'hd0e204a2;
    ram_cell[   10622] = 32'h0;  // 32'h1c65ea2c;
    ram_cell[   10623] = 32'h0;  // 32'h661e6629;
    ram_cell[   10624] = 32'h0;  // 32'h7f0908a9;
    ram_cell[   10625] = 32'h0;  // 32'h53324459;
    ram_cell[   10626] = 32'h0;  // 32'hf959a00c;
    ram_cell[   10627] = 32'h0;  // 32'h0b57fdc5;
    ram_cell[   10628] = 32'h0;  // 32'hbe8764ba;
    ram_cell[   10629] = 32'h0;  // 32'hc7d7ad96;
    ram_cell[   10630] = 32'h0;  // 32'h4713da5d;
    ram_cell[   10631] = 32'h0;  // 32'hbb4f9f85;
    ram_cell[   10632] = 32'h0;  // 32'h0aee5f44;
    ram_cell[   10633] = 32'h0;  // 32'h24c41255;
    ram_cell[   10634] = 32'h0;  // 32'h5a82a432;
    ram_cell[   10635] = 32'h0;  // 32'h33247e26;
    ram_cell[   10636] = 32'h0;  // 32'h7366770d;
    ram_cell[   10637] = 32'h0;  // 32'hfd74c5d5;
    ram_cell[   10638] = 32'h0;  // 32'h890b9a16;
    ram_cell[   10639] = 32'h0;  // 32'hdfdb37d0;
    ram_cell[   10640] = 32'h0;  // 32'he5f96317;
    ram_cell[   10641] = 32'h0;  // 32'h1d1b2a42;
    ram_cell[   10642] = 32'h0;  // 32'h17b10302;
    ram_cell[   10643] = 32'h0;  // 32'h06aacf1c;
    ram_cell[   10644] = 32'h0;  // 32'h8908e8da;
    ram_cell[   10645] = 32'h0;  // 32'hdfccc74f;
    ram_cell[   10646] = 32'h0;  // 32'h21d15897;
    ram_cell[   10647] = 32'h0;  // 32'h191cc583;
    ram_cell[   10648] = 32'h0;  // 32'h65619f60;
    ram_cell[   10649] = 32'h0;  // 32'h985230df;
    ram_cell[   10650] = 32'h0;  // 32'h3d7c8da2;
    ram_cell[   10651] = 32'h0;  // 32'h456dfc04;
    ram_cell[   10652] = 32'h0;  // 32'hd8d73a94;
    ram_cell[   10653] = 32'h0;  // 32'hbf81f026;
    ram_cell[   10654] = 32'h0;  // 32'hc29abf4c;
    ram_cell[   10655] = 32'h0;  // 32'hbdf2ba44;
    ram_cell[   10656] = 32'h0;  // 32'hb97fab9c;
    ram_cell[   10657] = 32'h0;  // 32'hdb203304;
    ram_cell[   10658] = 32'h0;  // 32'ha82a3fe4;
    ram_cell[   10659] = 32'h0;  // 32'ha02b2a3f;
    ram_cell[   10660] = 32'h0;  // 32'hcda048d8;
    ram_cell[   10661] = 32'h0;  // 32'hda88c54b;
    ram_cell[   10662] = 32'h0;  // 32'h74a77777;
    ram_cell[   10663] = 32'h0;  // 32'h3d1772cf;
    ram_cell[   10664] = 32'h0;  // 32'he450a028;
    ram_cell[   10665] = 32'h0;  // 32'h2ea55789;
    ram_cell[   10666] = 32'h0;  // 32'h47be15fb;
    ram_cell[   10667] = 32'h0;  // 32'ha8bf72b8;
    ram_cell[   10668] = 32'h0;  // 32'h12538cec;
    ram_cell[   10669] = 32'h0;  // 32'h3b2f9c0f;
    ram_cell[   10670] = 32'h0;  // 32'hd1ac0164;
    ram_cell[   10671] = 32'h0;  // 32'h8a1464bd;
    ram_cell[   10672] = 32'h0;  // 32'he6b13c6c;
    ram_cell[   10673] = 32'h0;  // 32'hb698257b;
    ram_cell[   10674] = 32'h0;  // 32'hb83006ab;
    ram_cell[   10675] = 32'h0;  // 32'h16ae8b09;
    ram_cell[   10676] = 32'h0;  // 32'h93b39271;
    ram_cell[   10677] = 32'h0;  // 32'h9640bf9d;
    ram_cell[   10678] = 32'h0;  // 32'hf029f1ea;
    ram_cell[   10679] = 32'h0;  // 32'h2daed79f;
    ram_cell[   10680] = 32'h0;  // 32'hc52b27dc;
    ram_cell[   10681] = 32'h0;  // 32'ha35c92bd;
    ram_cell[   10682] = 32'h0;  // 32'h4f879cb3;
    ram_cell[   10683] = 32'h0;  // 32'h9f4b9eac;
    ram_cell[   10684] = 32'h0;  // 32'h1c2b6121;
    ram_cell[   10685] = 32'h0;  // 32'h7683444b;
    ram_cell[   10686] = 32'h0;  // 32'h7103ee58;
    ram_cell[   10687] = 32'h0;  // 32'h1cd08669;
    ram_cell[   10688] = 32'h0;  // 32'h73dd7e22;
    ram_cell[   10689] = 32'h0;  // 32'hba9a46e1;
    ram_cell[   10690] = 32'h0;  // 32'hc00d906e;
    ram_cell[   10691] = 32'h0;  // 32'h66304fdd;
    ram_cell[   10692] = 32'h0;  // 32'h27931ddd;
    ram_cell[   10693] = 32'h0;  // 32'hdfe94901;
    ram_cell[   10694] = 32'h0;  // 32'h54a229d4;
    ram_cell[   10695] = 32'h0;  // 32'hf7931661;
    ram_cell[   10696] = 32'h0;  // 32'h86f29807;
    ram_cell[   10697] = 32'h0;  // 32'h083652a3;
    ram_cell[   10698] = 32'h0;  // 32'heb8b939c;
    ram_cell[   10699] = 32'h0;  // 32'h9046a2bf;
    ram_cell[   10700] = 32'h0;  // 32'h23fa5459;
    ram_cell[   10701] = 32'h0;  // 32'h8c7b0e61;
    ram_cell[   10702] = 32'h0;  // 32'h01fd3168;
    ram_cell[   10703] = 32'h0;  // 32'h95d986b1;
    ram_cell[   10704] = 32'h0;  // 32'hfbefdd56;
    ram_cell[   10705] = 32'h0;  // 32'h3d493fbc;
    ram_cell[   10706] = 32'h0;  // 32'hd79195bf;
    ram_cell[   10707] = 32'h0;  // 32'hab5bef9c;
    ram_cell[   10708] = 32'h0;  // 32'h5e8dd475;
    ram_cell[   10709] = 32'h0;  // 32'he7bdae41;
    ram_cell[   10710] = 32'h0;  // 32'h92a35796;
    ram_cell[   10711] = 32'h0;  // 32'hc418f9aa;
    ram_cell[   10712] = 32'h0;  // 32'he3e5f40a;
    ram_cell[   10713] = 32'h0;  // 32'h6739431d;
    ram_cell[   10714] = 32'h0;  // 32'h129b6ba9;
    ram_cell[   10715] = 32'h0;  // 32'hf4002173;
    ram_cell[   10716] = 32'h0;  // 32'hc09cf1d0;
    ram_cell[   10717] = 32'h0;  // 32'hdbd8c879;
    ram_cell[   10718] = 32'h0;  // 32'hb4ce6769;
    ram_cell[   10719] = 32'h0;  // 32'h9e24eb5f;
    ram_cell[   10720] = 32'h0;  // 32'h6c287782;
    ram_cell[   10721] = 32'h0;  // 32'h6ce4a299;
    ram_cell[   10722] = 32'h0;  // 32'h5731fa06;
    ram_cell[   10723] = 32'h0;  // 32'he2523de5;
    ram_cell[   10724] = 32'h0;  // 32'h14f0d980;
    ram_cell[   10725] = 32'h0;  // 32'h48b6827f;
    ram_cell[   10726] = 32'h0;  // 32'hac5d4927;
    ram_cell[   10727] = 32'h0;  // 32'hfcffd196;
    ram_cell[   10728] = 32'h0;  // 32'he578c58a;
    ram_cell[   10729] = 32'h0;  // 32'h876013bd;
    ram_cell[   10730] = 32'h0;  // 32'h6e9d5916;
    ram_cell[   10731] = 32'h0;  // 32'hdb4aa777;
    ram_cell[   10732] = 32'h0;  // 32'hdebb7da6;
    ram_cell[   10733] = 32'h0;  // 32'h0b672875;
    ram_cell[   10734] = 32'h0;  // 32'h5c538871;
    ram_cell[   10735] = 32'h0;  // 32'hc98d77d0;
    ram_cell[   10736] = 32'h0;  // 32'h6c513af1;
    ram_cell[   10737] = 32'h0;  // 32'hd137565d;
    ram_cell[   10738] = 32'h0;  // 32'h2516b71b;
    ram_cell[   10739] = 32'h0;  // 32'h1a0997ff;
    ram_cell[   10740] = 32'h0;  // 32'hf6872214;
    ram_cell[   10741] = 32'h0;  // 32'h209ae850;
    ram_cell[   10742] = 32'h0;  // 32'hcfdaf471;
    ram_cell[   10743] = 32'h0;  // 32'h1f533432;
    ram_cell[   10744] = 32'h0;  // 32'hb7c599d4;
    ram_cell[   10745] = 32'h0;  // 32'h99f31a37;
    ram_cell[   10746] = 32'h0;  // 32'ha6f13683;
    ram_cell[   10747] = 32'h0;  // 32'hb108cebd;
    ram_cell[   10748] = 32'h0;  // 32'hdff854f4;
    ram_cell[   10749] = 32'h0;  // 32'hee72a85c;
    ram_cell[   10750] = 32'h0;  // 32'h2fa97b3d;
    ram_cell[   10751] = 32'h0;  // 32'he0502e22;
    ram_cell[   10752] = 32'h0;  // 32'h506db97b;
    ram_cell[   10753] = 32'h0;  // 32'h70510d99;
    ram_cell[   10754] = 32'h0;  // 32'hbb166f63;
    ram_cell[   10755] = 32'h0;  // 32'h099a3afe;
    ram_cell[   10756] = 32'h0;  // 32'h1c271f54;
    ram_cell[   10757] = 32'h0;  // 32'h9088a048;
    ram_cell[   10758] = 32'h0;  // 32'h3ef3d629;
    ram_cell[   10759] = 32'h0;  // 32'h9590a81e;
    ram_cell[   10760] = 32'h0;  // 32'hb732bd65;
    ram_cell[   10761] = 32'h0;  // 32'h9ec86b3b;
    ram_cell[   10762] = 32'h0;  // 32'heca21245;
    ram_cell[   10763] = 32'h0;  // 32'hcc470ccd;
    ram_cell[   10764] = 32'h0;  // 32'h59770d5a;
    ram_cell[   10765] = 32'h0;  // 32'h5963de94;
    ram_cell[   10766] = 32'h0;  // 32'hc8e9370c;
    ram_cell[   10767] = 32'h0;  // 32'h137f144b;
    ram_cell[   10768] = 32'h0;  // 32'hcec21762;
    ram_cell[   10769] = 32'h0;  // 32'hd2b704bb;
    ram_cell[   10770] = 32'h0;  // 32'h660d62d1;
    ram_cell[   10771] = 32'h0;  // 32'h52835844;
    ram_cell[   10772] = 32'h0;  // 32'ha0906e43;
    ram_cell[   10773] = 32'h0;  // 32'h7a5cc86c;
    ram_cell[   10774] = 32'h0;  // 32'he8985fb2;
    ram_cell[   10775] = 32'h0;  // 32'ha8845aef;
    ram_cell[   10776] = 32'h0;  // 32'hadcd9696;
    ram_cell[   10777] = 32'h0;  // 32'hd6c796f1;
    ram_cell[   10778] = 32'h0;  // 32'he913b217;
    ram_cell[   10779] = 32'h0;  // 32'h61c1ad50;
    ram_cell[   10780] = 32'h0;  // 32'hb3bb57b8;
    ram_cell[   10781] = 32'h0;  // 32'h3d011da8;
    ram_cell[   10782] = 32'h0;  // 32'h7249b38e;
    ram_cell[   10783] = 32'h0;  // 32'h0f3db386;
    ram_cell[   10784] = 32'h0;  // 32'ha60d9baa;
    ram_cell[   10785] = 32'h0;  // 32'hcf4acaab;
    ram_cell[   10786] = 32'h0;  // 32'ha067593a;
    ram_cell[   10787] = 32'h0;  // 32'hec65f758;
    ram_cell[   10788] = 32'h0;  // 32'hec57ef7a;
    ram_cell[   10789] = 32'h0;  // 32'heb0b15d9;
    ram_cell[   10790] = 32'h0;  // 32'h7a468616;
    ram_cell[   10791] = 32'h0;  // 32'hce58bcf1;
    ram_cell[   10792] = 32'h0;  // 32'h6569ab9b;
    ram_cell[   10793] = 32'h0;  // 32'h0a804c28;
    ram_cell[   10794] = 32'h0;  // 32'hc2244edf;
    ram_cell[   10795] = 32'h0;  // 32'h888d1e07;
    ram_cell[   10796] = 32'h0;  // 32'ha1c8ae5f;
    ram_cell[   10797] = 32'h0;  // 32'hba5f811f;
    ram_cell[   10798] = 32'h0;  // 32'h1b077686;
    ram_cell[   10799] = 32'h0;  // 32'h05143673;
    ram_cell[   10800] = 32'h0;  // 32'hb368d309;
    ram_cell[   10801] = 32'h0;  // 32'h49227b06;
    ram_cell[   10802] = 32'h0;  // 32'h4c663957;
    ram_cell[   10803] = 32'h0;  // 32'hf91bfc0f;
    ram_cell[   10804] = 32'h0;  // 32'hd76990e6;
    ram_cell[   10805] = 32'h0;  // 32'he04eee20;
    ram_cell[   10806] = 32'h0;  // 32'ha08ac76f;
    ram_cell[   10807] = 32'h0;  // 32'h6eed64cd;
    ram_cell[   10808] = 32'h0;  // 32'hac71b81b;
    ram_cell[   10809] = 32'h0;  // 32'h29a3e6fc;
    ram_cell[   10810] = 32'h0;  // 32'hab5f1556;
    ram_cell[   10811] = 32'h0;  // 32'h82aa9f4d;
    ram_cell[   10812] = 32'h0;  // 32'h10d21d30;
    ram_cell[   10813] = 32'h0;  // 32'hda4ccf23;
    ram_cell[   10814] = 32'h0;  // 32'hdacf59ff;
    ram_cell[   10815] = 32'h0;  // 32'h373ec718;
    ram_cell[   10816] = 32'h0;  // 32'hdb33e0a7;
    ram_cell[   10817] = 32'h0;  // 32'hd68ee30f;
    ram_cell[   10818] = 32'h0;  // 32'h9c454176;
    ram_cell[   10819] = 32'h0;  // 32'hcd92e035;
    ram_cell[   10820] = 32'h0;  // 32'h235e562e;
    ram_cell[   10821] = 32'h0;  // 32'he32bd73b;
    ram_cell[   10822] = 32'h0;  // 32'ha0bfc2d6;
    ram_cell[   10823] = 32'h0;  // 32'h8fb6eacd;
    ram_cell[   10824] = 32'h0;  // 32'h79a807b0;
    ram_cell[   10825] = 32'h0;  // 32'hca583469;
    ram_cell[   10826] = 32'h0;  // 32'hf1a835ef;
    ram_cell[   10827] = 32'h0;  // 32'hc47bf776;
    ram_cell[   10828] = 32'h0;  // 32'h0ad2b72a;
    ram_cell[   10829] = 32'h0;  // 32'h591e07de;
    ram_cell[   10830] = 32'h0;  // 32'h819840c2;
    ram_cell[   10831] = 32'h0;  // 32'h37f745e2;
    ram_cell[   10832] = 32'h0;  // 32'h1fae0a98;
    ram_cell[   10833] = 32'h0;  // 32'h21740009;
    ram_cell[   10834] = 32'h0;  // 32'he807cf92;
    ram_cell[   10835] = 32'h0;  // 32'h38c25299;
    ram_cell[   10836] = 32'h0;  // 32'h2e687206;
    ram_cell[   10837] = 32'h0;  // 32'h5fdd2504;
    ram_cell[   10838] = 32'h0;  // 32'hd1ac3c86;
    ram_cell[   10839] = 32'h0;  // 32'h29324c39;
    ram_cell[   10840] = 32'h0;  // 32'h9129ad76;
    ram_cell[   10841] = 32'h0;  // 32'h6061e88d;
    ram_cell[   10842] = 32'h0;  // 32'h7b2bf124;
    ram_cell[   10843] = 32'h0;  // 32'h00eb9609;
    ram_cell[   10844] = 32'h0;  // 32'h9bbb90e4;
    ram_cell[   10845] = 32'h0;  // 32'h4624eb77;
    ram_cell[   10846] = 32'h0;  // 32'hd3004f83;
    ram_cell[   10847] = 32'h0;  // 32'h444594e4;
    ram_cell[   10848] = 32'h0;  // 32'hb28ea6fd;
    ram_cell[   10849] = 32'h0;  // 32'hd17340df;
    ram_cell[   10850] = 32'h0;  // 32'h87b632f6;
    ram_cell[   10851] = 32'h0;  // 32'h8b72b0c7;
    ram_cell[   10852] = 32'h0;  // 32'hb445ca20;
    ram_cell[   10853] = 32'h0;  // 32'h491545e3;
    ram_cell[   10854] = 32'h0;  // 32'hf70cb005;
    ram_cell[   10855] = 32'h0;  // 32'h2861beef;
    ram_cell[   10856] = 32'h0;  // 32'h4549d12b;
    ram_cell[   10857] = 32'h0;  // 32'he777ccff;
    ram_cell[   10858] = 32'h0;  // 32'hdd285911;
    ram_cell[   10859] = 32'h0;  // 32'hfb99c0b1;
    ram_cell[   10860] = 32'h0;  // 32'h8248cc38;
    ram_cell[   10861] = 32'h0;  // 32'h209da4fa;
    ram_cell[   10862] = 32'h0;  // 32'hb0cb5764;
    ram_cell[   10863] = 32'h0;  // 32'h9fbd2b66;
    ram_cell[   10864] = 32'h0;  // 32'h859b3cf5;
    ram_cell[   10865] = 32'h0;  // 32'hcc812a07;
    ram_cell[   10866] = 32'h0;  // 32'hb1a6fd80;
    ram_cell[   10867] = 32'h0;  // 32'hdce2ec8c;
    ram_cell[   10868] = 32'h0;  // 32'hbd28a29a;
    ram_cell[   10869] = 32'h0;  // 32'h2613ee07;
    ram_cell[   10870] = 32'h0;  // 32'hc5272c6d;
    ram_cell[   10871] = 32'h0;  // 32'h45f169ee;
    ram_cell[   10872] = 32'h0;  // 32'hae2a90a4;
    ram_cell[   10873] = 32'h0;  // 32'hbb081494;
    ram_cell[   10874] = 32'h0;  // 32'h6cac0732;
    ram_cell[   10875] = 32'h0;  // 32'h431e6163;
    ram_cell[   10876] = 32'h0;  // 32'hdf27be9a;
    ram_cell[   10877] = 32'h0;  // 32'h7187c5d1;
    ram_cell[   10878] = 32'h0;  // 32'h7fd6d553;
    ram_cell[   10879] = 32'h0;  // 32'h281efe65;
    ram_cell[   10880] = 32'h0;  // 32'hf886d906;
    ram_cell[   10881] = 32'h0;  // 32'h96d705a7;
    ram_cell[   10882] = 32'h0;  // 32'hd6c304ff;
    ram_cell[   10883] = 32'h0;  // 32'h2c79648b;
    ram_cell[   10884] = 32'h0;  // 32'hb029b816;
    ram_cell[   10885] = 32'h0;  // 32'ha03ea8b1;
    ram_cell[   10886] = 32'h0;  // 32'he8ebdde7;
    ram_cell[   10887] = 32'h0;  // 32'hb9d16e40;
    ram_cell[   10888] = 32'h0;  // 32'he70c5179;
    ram_cell[   10889] = 32'h0;  // 32'ha0f1096a;
    ram_cell[   10890] = 32'h0;  // 32'hc9320f24;
    ram_cell[   10891] = 32'h0;  // 32'hc3328bde;
    ram_cell[   10892] = 32'h0;  // 32'hb8730634;
    ram_cell[   10893] = 32'h0;  // 32'ha7400572;
    ram_cell[   10894] = 32'h0;  // 32'h3ea13020;
    ram_cell[   10895] = 32'h0;  // 32'h9f2a80e0;
    ram_cell[   10896] = 32'h0;  // 32'h7d992b78;
    ram_cell[   10897] = 32'h0;  // 32'h95237f71;
    ram_cell[   10898] = 32'h0;  // 32'hc7103fd3;
    ram_cell[   10899] = 32'h0;  // 32'h4dd06b11;
    ram_cell[   10900] = 32'h0;  // 32'h7f772d47;
    ram_cell[   10901] = 32'h0;  // 32'hfb96e07a;
    ram_cell[   10902] = 32'h0;  // 32'h4c6b1773;
    ram_cell[   10903] = 32'h0;  // 32'h6b1b9200;
    ram_cell[   10904] = 32'h0;  // 32'h186c9a70;
    ram_cell[   10905] = 32'h0;  // 32'ha3382705;
    ram_cell[   10906] = 32'h0;  // 32'h63ede97f;
    ram_cell[   10907] = 32'h0;  // 32'hdb4c6cf0;
    ram_cell[   10908] = 32'h0;  // 32'hdefe2994;
    ram_cell[   10909] = 32'h0;  // 32'hb5221edd;
    ram_cell[   10910] = 32'h0;  // 32'h0045472f;
    ram_cell[   10911] = 32'h0;  // 32'h74826ced;
    ram_cell[   10912] = 32'h0;  // 32'h317b909f;
    ram_cell[   10913] = 32'h0;  // 32'hc85a4815;
    ram_cell[   10914] = 32'h0;  // 32'hd66c7b8c;
    ram_cell[   10915] = 32'h0;  // 32'h8840ae39;
    ram_cell[   10916] = 32'h0;  // 32'hba21b451;
    ram_cell[   10917] = 32'h0;  // 32'he6604074;
    ram_cell[   10918] = 32'h0;  // 32'had6bfad3;
    ram_cell[   10919] = 32'h0;  // 32'h54946a25;
    ram_cell[   10920] = 32'h0;  // 32'h04a67120;
    ram_cell[   10921] = 32'h0;  // 32'he834a4de;
    ram_cell[   10922] = 32'h0;  // 32'h6af3d2e9;
    ram_cell[   10923] = 32'h0;  // 32'hab37cbe4;
    ram_cell[   10924] = 32'h0;  // 32'h03aa3347;
    ram_cell[   10925] = 32'h0;  // 32'he662bf9f;
    ram_cell[   10926] = 32'h0;  // 32'h916e84a8;
    ram_cell[   10927] = 32'h0;  // 32'h8a7c649d;
    ram_cell[   10928] = 32'h0;  // 32'h200dc276;
    ram_cell[   10929] = 32'h0;  // 32'h53915b30;
    ram_cell[   10930] = 32'h0;  // 32'hc8850185;
    ram_cell[   10931] = 32'h0;  // 32'h87e296df;
    ram_cell[   10932] = 32'h0;  // 32'h68ed4d42;
    ram_cell[   10933] = 32'h0;  // 32'hc2ed2937;
    ram_cell[   10934] = 32'h0;  // 32'h24bf8e4f;
    ram_cell[   10935] = 32'h0;  // 32'h26d56611;
    ram_cell[   10936] = 32'h0;  // 32'hfe3e8c19;
    ram_cell[   10937] = 32'h0;  // 32'h0c75b0db;
    ram_cell[   10938] = 32'h0;  // 32'h9ab6aef3;
    ram_cell[   10939] = 32'h0;  // 32'hc7e71936;
    ram_cell[   10940] = 32'h0;  // 32'h1e41872c;
    ram_cell[   10941] = 32'h0;  // 32'ha7258ae3;
    ram_cell[   10942] = 32'h0;  // 32'h21557ce6;
    ram_cell[   10943] = 32'h0;  // 32'h09a82f90;
    ram_cell[   10944] = 32'h0;  // 32'hb29bfdce;
    ram_cell[   10945] = 32'h0;  // 32'hab0e5aeb;
    ram_cell[   10946] = 32'h0;  // 32'hb859ea46;
    ram_cell[   10947] = 32'h0;  // 32'h17b7bf73;
    ram_cell[   10948] = 32'h0;  // 32'ha9cddfc7;
    ram_cell[   10949] = 32'h0;  // 32'hf6a5f669;
    ram_cell[   10950] = 32'h0;  // 32'hc841a559;
    ram_cell[   10951] = 32'h0;  // 32'h7657e80a;
    ram_cell[   10952] = 32'h0;  // 32'h1a5095ab;
    ram_cell[   10953] = 32'h0;  // 32'h0a83eeb8;
    ram_cell[   10954] = 32'h0;  // 32'h39709af1;
    ram_cell[   10955] = 32'h0;  // 32'ha0a2c032;
    ram_cell[   10956] = 32'h0;  // 32'ha14e0a34;
    ram_cell[   10957] = 32'h0;  // 32'hf38de9fe;
    ram_cell[   10958] = 32'h0;  // 32'hf64b511b;
    ram_cell[   10959] = 32'h0;  // 32'h3a594b01;
    ram_cell[   10960] = 32'h0;  // 32'hc7662d8e;
    ram_cell[   10961] = 32'h0;  // 32'hcb6a8141;
    ram_cell[   10962] = 32'h0;  // 32'hcddfc8d0;
    ram_cell[   10963] = 32'h0;  // 32'h0f044374;
    ram_cell[   10964] = 32'h0;  // 32'h922e65bc;
    ram_cell[   10965] = 32'h0;  // 32'hddf89d60;
    ram_cell[   10966] = 32'h0;  // 32'h5c7e93c6;
    ram_cell[   10967] = 32'h0;  // 32'hf0cd19af;
    ram_cell[   10968] = 32'h0;  // 32'hed6d9eb3;
    ram_cell[   10969] = 32'h0;  // 32'h52943f8b;
    ram_cell[   10970] = 32'h0;  // 32'hb8e94363;
    ram_cell[   10971] = 32'h0;  // 32'hc899d5ae;
    ram_cell[   10972] = 32'h0;  // 32'hbe226802;
    ram_cell[   10973] = 32'h0;  // 32'hdb30b261;
    ram_cell[   10974] = 32'h0;  // 32'h7e4a8cf3;
    ram_cell[   10975] = 32'h0;  // 32'he35a67c6;
    ram_cell[   10976] = 32'h0;  // 32'h0194e771;
    ram_cell[   10977] = 32'h0;  // 32'hf6516b6d;
    ram_cell[   10978] = 32'h0;  // 32'h414f6d8b;
    ram_cell[   10979] = 32'h0;  // 32'h6f74bc26;
    ram_cell[   10980] = 32'h0;  // 32'h5d0d7b27;
    ram_cell[   10981] = 32'h0;  // 32'hbe4cd1ef;
    ram_cell[   10982] = 32'h0;  // 32'h2554f8c9;
    ram_cell[   10983] = 32'h0;  // 32'hd97ced1c;
    ram_cell[   10984] = 32'h0;  // 32'h889cc81f;
    ram_cell[   10985] = 32'h0;  // 32'h7b1032b3;
    ram_cell[   10986] = 32'h0;  // 32'hb15cb991;
    ram_cell[   10987] = 32'h0;  // 32'hd3914e9d;
    ram_cell[   10988] = 32'h0;  // 32'h15ed9d31;
    ram_cell[   10989] = 32'h0;  // 32'hbbd3b3ed;
    ram_cell[   10990] = 32'h0;  // 32'h27aec544;
    ram_cell[   10991] = 32'h0;  // 32'hb37ea13d;
    ram_cell[   10992] = 32'h0;  // 32'ha2272f8e;
    ram_cell[   10993] = 32'h0;  // 32'h3f15697a;
    ram_cell[   10994] = 32'h0;  // 32'hc55044e9;
    ram_cell[   10995] = 32'h0;  // 32'h69f8bd04;
    ram_cell[   10996] = 32'h0;  // 32'h5e299a4d;
    ram_cell[   10997] = 32'h0;  // 32'h55c2e12c;
    ram_cell[   10998] = 32'h0;  // 32'hf15c7f83;
    ram_cell[   10999] = 32'h0;  // 32'h8e51cc63;
    ram_cell[   11000] = 32'h0;  // 32'h8a30b0b0;
    ram_cell[   11001] = 32'h0;  // 32'h0526e19c;
    ram_cell[   11002] = 32'h0;  // 32'hfc3fe039;
    ram_cell[   11003] = 32'h0;  // 32'h84d90e29;
    ram_cell[   11004] = 32'h0;  // 32'hb1636c2f;
    ram_cell[   11005] = 32'h0;  // 32'h157a9e41;
    ram_cell[   11006] = 32'h0;  // 32'h7d5f3e13;
    ram_cell[   11007] = 32'h0;  // 32'hf5e54123;
    ram_cell[   11008] = 32'h0;  // 32'hb4fac5c2;
    ram_cell[   11009] = 32'h0;  // 32'h32211c96;
    ram_cell[   11010] = 32'h0;  // 32'he3965063;
    ram_cell[   11011] = 32'h0;  // 32'heff73e2d;
    ram_cell[   11012] = 32'h0;  // 32'hd9b962d5;
    ram_cell[   11013] = 32'h0;  // 32'h6216a07c;
    ram_cell[   11014] = 32'h0;  // 32'hfa036b6f;
    ram_cell[   11015] = 32'h0;  // 32'h397eabf8;
    ram_cell[   11016] = 32'h0;  // 32'h8dad0531;
    ram_cell[   11017] = 32'h0;  // 32'ha2dfee88;
    ram_cell[   11018] = 32'h0;  // 32'hf2f3fd48;
    ram_cell[   11019] = 32'h0;  // 32'h7a183700;
    ram_cell[   11020] = 32'h0;  // 32'h33cedcaa;
    ram_cell[   11021] = 32'h0;  // 32'h7648216e;
    ram_cell[   11022] = 32'h0;  // 32'h42d51665;
    ram_cell[   11023] = 32'h0;  // 32'h82d7eb4d;
    ram_cell[   11024] = 32'h0;  // 32'h5593a5ea;
    ram_cell[   11025] = 32'h0;  // 32'hf2fe5bb4;
    ram_cell[   11026] = 32'h0;  // 32'h3b4b482e;
    ram_cell[   11027] = 32'h0;  // 32'h0c1ea96b;
    ram_cell[   11028] = 32'h0;  // 32'h000c8bf1;
    ram_cell[   11029] = 32'h0;  // 32'h320cafbf;
    ram_cell[   11030] = 32'h0;  // 32'h48ac4e7b;
    ram_cell[   11031] = 32'h0;  // 32'h31ac2144;
    ram_cell[   11032] = 32'h0;  // 32'h114d1852;
    ram_cell[   11033] = 32'h0;  // 32'hf6b24b17;
    ram_cell[   11034] = 32'h0;  // 32'h462d92a7;
    ram_cell[   11035] = 32'h0;  // 32'he7f92ba7;
    ram_cell[   11036] = 32'h0;  // 32'h66c9f6d5;
    ram_cell[   11037] = 32'h0;  // 32'he2609b36;
    ram_cell[   11038] = 32'h0;  // 32'hd7b770ce;
    ram_cell[   11039] = 32'h0;  // 32'h20aeb6cb;
    ram_cell[   11040] = 32'h0;  // 32'h77c4392f;
    ram_cell[   11041] = 32'h0;  // 32'h0148d619;
    ram_cell[   11042] = 32'h0;  // 32'h8d297757;
    ram_cell[   11043] = 32'h0;  // 32'h9b588824;
    ram_cell[   11044] = 32'h0;  // 32'h39bc6771;
    ram_cell[   11045] = 32'h0;  // 32'hfa57fc80;
    ram_cell[   11046] = 32'h0;  // 32'h8d34a4dc;
    ram_cell[   11047] = 32'h0;  // 32'he2e981c3;
    ram_cell[   11048] = 32'h0;  // 32'h431c4239;
    ram_cell[   11049] = 32'h0;  // 32'h170d666b;
    ram_cell[   11050] = 32'h0;  // 32'h2ebea573;
    ram_cell[   11051] = 32'h0;  // 32'h3b2b9ff0;
    ram_cell[   11052] = 32'h0;  // 32'hc4f9ad16;
    ram_cell[   11053] = 32'h0;  // 32'h10dc21a8;
    ram_cell[   11054] = 32'h0;  // 32'he3ae2fef;
    ram_cell[   11055] = 32'h0;  // 32'h4c7c2b55;
    ram_cell[   11056] = 32'h0;  // 32'had229f03;
    ram_cell[   11057] = 32'h0;  // 32'h97cd2830;
    ram_cell[   11058] = 32'h0;  // 32'he03e7b0a;
    ram_cell[   11059] = 32'h0;  // 32'h672df604;
    ram_cell[   11060] = 32'h0;  // 32'hfc19c4bf;
    ram_cell[   11061] = 32'h0;  // 32'hfeb63ef5;
    ram_cell[   11062] = 32'h0;  // 32'h9d47d263;
    ram_cell[   11063] = 32'h0;  // 32'h2e581dd6;
    ram_cell[   11064] = 32'h0;  // 32'h5ead4f49;
    ram_cell[   11065] = 32'h0;  // 32'h1996e27a;
    ram_cell[   11066] = 32'h0;  // 32'h17b9637d;
    ram_cell[   11067] = 32'h0;  // 32'ha9c33467;
    ram_cell[   11068] = 32'h0;  // 32'h0181eb30;
    ram_cell[   11069] = 32'h0;  // 32'h31d96627;
    ram_cell[   11070] = 32'h0;  // 32'h40d5f459;
    ram_cell[   11071] = 32'h0;  // 32'h6312cb2f;
    ram_cell[   11072] = 32'h0;  // 32'hca49b41b;
    ram_cell[   11073] = 32'h0;  // 32'ha44fd2ce;
    ram_cell[   11074] = 32'h0;  // 32'h30960df1;
    ram_cell[   11075] = 32'h0;  // 32'hb5a03871;
    ram_cell[   11076] = 32'h0;  // 32'he380750e;
    ram_cell[   11077] = 32'h0;  // 32'hea4ead8b;
    ram_cell[   11078] = 32'h0;  // 32'h789b379c;
    ram_cell[   11079] = 32'h0;  // 32'h3832ba3f;
    ram_cell[   11080] = 32'h0;  // 32'hb3c08ede;
    ram_cell[   11081] = 32'h0;  // 32'h7aeb3421;
    ram_cell[   11082] = 32'h0;  // 32'h140a87b4;
    ram_cell[   11083] = 32'h0;  // 32'h9afef0e6;
    ram_cell[   11084] = 32'h0;  // 32'hdd973e24;
    ram_cell[   11085] = 32'h0;  // 32'h287ff2bd;
    ram_cell[   11086] = 32'h0;  // 32'he936db0a;
    ram_cell[   11087] = 32'h0;  // 32'h82e327c3;
    ram_cell[   11088] = 32'h0;  // 32'h127e1ac7;
    ram_cell[   11089] = 32'h0;  // 32'hb859abfd;
    ram_cell[   11090] = 32'h0;  // 32'h3475197d;
    ram_cell[   11091] = 32'h0;  // 32'hdaea3d5d;
    ram_cell[   11092] = 32'h0;  // 32'hf2a6fd3c;
    ram_cell[   11093] = 32'h0;  // 32'hcef48e75;
    ram_cell[   11094] = 32'h0;  // 32'hdd8e35c1;
    ram_cell[   11095] = 32'h0;  // 32'hd7aacdfe;
    ram_cell[   11096] = 32'h0;  // 32'h77c70dec;
    ram_cell[   11097] = 32'h0;  // 32'h944cdc70;
    ram_cell[   11098] = 32'h0;  // 32'h381b5a22;
    ram_cell[   11099] = 32'h0;  // 32'hb371e0a2;
    ram_cell[   11100] = 32'h0;  // 32'h1cbe09fc;
    ram_cell[   11101] = 32'h0;  // 32'hb0ffefe4;
    ram_cell[   11102] = 32'h0;  // 32'h57731893;
    ram_cell[   11103] = 32'h0;  // 32'h928cbf03;
    ram_cell[   11104] = 32'h0;  // 32'hdd8cec00;
    ram_cell[   11105] = 32'h0;  // 32'h1be358bc;
    ram_cell[   11106] = 32'h0;  // 32'h5be66513;
    ram_cell[   11107] = 32'h0;  // 32'hf60c4f62;
    ram_cell[   11108] = 32'h0;  // 32'h2b2dfa33;
    ram_cell[   11109] = 32'h0;  // 32'ha9759e76;
    ram_cell[   11110] = 32'h0;  // 32'hf2f5a530;
    ram_cell[   11111] = 32'h0;  // 32'h1707b329;
    ram_cell[   11112] = 32'h0;  // 32'h7539db7c;
    ram_cell[   11113] = 32'h0;  // 32'hb568ed46;
    ram_cell[   11114] = 32'h0;  // 32'h202722ef;
    ram_cell[   11115] = 32'h0;  // 32'h7e4ea1d6;
    ram_cell[   11116] = 32'h0;  // 32'hb52d5b23;
    ram_cell[   11117] = 32'h0;  // 32'h6be56b8d;
    ram_cell[   11118] = 32'h0;  // 32'hf99e3717;
    ram_cell[   11119] = 32'h0;  // 32'h2e9c91b2;
    ram_cell[   11120] = 32'h0;  // 32'h4455a818;
    ram_cell[   11121] = 32'h0;  // 32'he80a9b15;
    ram_cell[   11122] = 32'h0;  // 32'h04665449;
    ram_cell[   11123] = 32'h0;  // 32'hfe11f234;
    ram_cell[   11124] = 32'h0;  // 32'h5089fcb3;
    ram_cell[   11125] = 32'h0;  // 32'h1bc02c67;
    ram_cell[   11126] = 32'h0;  // 32'he5690c65;
    ram_cell[   11127] = 32'h0;  // 32'hdd720728;
    ram_cell[   11128] = 32'h0;  // 32'h7e550d56;
    ram_cell[   11129] = 32'h0;  // 32'h892944bc;
    ram_cell[   11130] = 32'h0;  // 32'hd5ebcea5;
    ram_cell[   11131] = 32'h0;  // 32'h8200ece1;
    ram_cell[   11132] = 32'h0;  // 32'hc14cdc38;
    ram_cell[   11133] = 32'h0;  // 32'hdddd097f;
    ram_cell[   11134] = 32'h0;  // 32'h99612e03;
    ram_cell[   11135] = 32'h0;  // 32'hd19ddde7;
    ram_cell[   11136] = 32'h0;  // 32'h28ab7ce1;
    ram_cell[   11137] = 32'h0;  // 32'h95759d56;
    ram_cell[   11138] = 32'h0;  // 32'hb68ed5c7;
    ram_cell[   11139] = 32'h0;  // 32'h68eb0b93;
    ram_cell[   11140] = 32'h0;  // 32'h4cfce0a4;
    ram_cell[   11141] = 32'h0;  // 32'ha2854803;
    ram_cell[   11142] = 32'h0;  // 32'hc54ebb65;
    ram_cell[   11143] = 32'h0;  // 32'hefbcb908;
    ram_cell[   11144] = 32'h0;  // 32'h67032396;
    ram_cell[   11145] = 32'h0;  // 32'h150f19af;
    ram_cell[   11146] = 32'h0;  // 32'h295c9e94;
    ram_cell[   11147] = 32'h0;  // 32'hf87ea237;
    ram_cell[   11148] = 32'h0;  // 32'hbc7060ab;
    ram_cell[   11149] = 32'h0;  // 32'h468eff2f;
    ram_cell[   11150] = 32'h0;  // 32'h887ac5b5;
    ram_cell[   11151] = 32'h0;  // 32'h5d60d906;
    ram_cell[   11152] = 32'h0;  // 32'h63e476a4;
    ram_cell[   11153] = 32'h0;  // 32'h01145b8e;
    ram_cell[   11154] = 32'h0;  // 32'h519e34a4;
    ram_cell[   11155] = 32'h0;  // 32'h9e241095;
    ram_cell[   11156] = 32'h0;  // 32'h8af0ded0;
    ram_cell[   11157] = 32'h0;  // 32'h57b08395;
    ram_cell[   11158] = 32'h0;  // 32'hc16e70d0;
    ram_cell[   11159] = 32'h0;  // 32'hb02c05c3;
    ram_cell[   11160] = 32'h0;  // 32'hb523e31e;
    ram_cell[   11161] = 32'h0;  // 32'h087be128;
    ram_cell[   11162] = 32'h0;  // 32'h3b2c9203;
    ram_cell[   11163] = 32'h0;  // 32'hac5d3c63;
    ram_cell[   11164] = 32'h0;  // 32'ha5035df8;
    ram_cell[   11165] = 32'h0;  // 32'h621c30c2;
    ram_cell[   11166] = 32'h0;  // 32'h22956e93;
    ram_cell[   11167] = 32'h0;  // 32'h54cbbeb3;
    ram_cell[   11168] = 32'h0;  // 32'he67ed240;
    ram_cell[   11169] = 32'h0;  // 32'hb6c1342b;
    ram_cell[   11170] = 32'h0;  // 32'hc3df62fd;
    ram_cell[   11171] = 32'h0;  // 32'h98ea4bb2;
    ram_cell[   11172] = 32'h0;  // 32'hb464ae65;
    ram_cell[   11173] = 32'h0;  // 32'heed0bb20;
    ram_cell[   11174] = 32'h0;  // 32'ha8e0be82;
    ram_cell[   11175] = 32'h0;  // 32'h169b59fa;
    ram_cell[   11176] = 32'h0;  // 32'h121eb265;
    ram_cell[   11177] = 32'h0;  // 32'hb66f5bdb;
    ram_cell[   11178] = 32'h0;  // 32'h9fffe324;
    ram_cell[   11179] = 32'h0;  // 32'hcfccb342;
    ram_cell[   11180] = 32'h0;  // 32'h016f0d51;
    ram_cell[   11181] = 32'h0;  // 32'hf4f9df0d;
    ram_cell[   11182] = 32'h0;  // 32'h601dd5a6;
    ram_cell[   11183] = 32'h0;  // 32'hd38ee49a;
    ram_cell[   11184] = 32'h0;  // 32'hee14ce4e;
    ram_cell[   11185] = 32'h0;  // 32'h100b2ea5;
    ram_cell[   11186] = 32'h0;  // 32'hebb81afd;
    ram_cell[   11187] = 32'h0;  // 32'h886ed76a;
    ram_cell[   11188] = 32'h0;  // 32'h11418b70;
    ram_cell[   11189] = 32'h0;  // 32'h05305615;
    ram_cell[   11190] = 32'h0;  // 32'he2f3fd6f;
    ram_cell[   11191] = 32'h0;  // 32'h8694bf9b;
    ram_cell[   11192] = 32'h0;  // 32'h74240c05;
    ram_cell[   11193] = 32'h0;  // 32'hce3d8ec9;
    ram_cell[   11194] = 32'h0;  // 32'h81cae2db;
    ram_cell[   11195] = 32'h0;  // 32'h4be977cf;
    ram_cell[   11196] = 32'h0;  // 32'h625cc68c;
    ram_cell[   11197] = 32'h0;  // 32'h6bbfee2b;
    ram_cell[   11198] = 32'h0;  // 32'h62689d65;
    ram_cell[   11199] = 32'h0;  // 32'h234a7a3c;
    ram_cell[   11200] = 32'h0;  // 32'ha4dc0b32;
    ram_cell[   11201] = 32'h0;  // 32'h97832793;
    ram_cell[   11202] = 32'h0;  // 32'hc618ddcc;
    ram_cell[   11203] = 32'h0;  // 32'h3dbc8d26;
    ram_cell[   11204] = 32'h0;  // 32'h2247ace0;
    ram_cell[   11205] = 32'h0;  // 32'hbb028cd0;
    ram_cell[   11206] = 32'h0;  // 32'h43e9101e;
    ram_cell[   11207] = 32'h0;  // 32'hf5239895;
    ram_cell[   11208] = 32'h0;  // 32'h4f7a4380;
    ram_cell[   11209] = 32'h0;  // 32'h742be9b9;
    ram_cell[   11210] = 32'h0;  // 32'h147fc445;
    ram_cell[   11211] = 32'h0;  // 32'h710eccdf;
    ram_cell[   11212] = 32'h0;  // 32'h11e09f66;
    ram_cell[   11213] = 32'h0;  // 32'hd11215ed;
    ram_cell[   11214] = 32'h0;  // 32'hc9087cc5;
    ram_cell[   11215] = 32'h0;  // 32'h1f2ec0be;
    ram_cell[   11216] = 32'h0;  // 32'h573e6ec9;
    ram_cell[   11217] = 32'h0;  // 32'h21e38fab;
    ram_cell[   11218] = 32'h0;  // 32'h8cefdd45;
    ram_cell[   11219] = 32'h0;  // 32'h022c8dda;
    ram_cell[   11220] = 32'h0;  // 32'h1f5794ee;
    ram_cell[   11221] = 32'h0;  // 32'h4beb6d92;
    ram_cell[   11222] = 32'h0;  // 32'h201ae7ba;
    ram_cell[   11223] = 32'h0;  // 32'h1a77adc6;
    ram_cell[   11224] = 32'h0;  // 32'h2a596ed9;
    ram_cell[   11225] = 32'h0;  // 32'h78cf59ef;
    ram_cell[   11226] = 32'h0;  // 32'h16b2011c;
    ram_cell[   11227] = 32'h0;  // 32'ha8720563;
    ram_cell[   11228] = 32'h0;  // 32'head118c8;
    ram_cell[   11229] = 32'h0;  // 32'he931abe0;
    ram_cell[   11230] = 32'h0;  // 32'hdbccb3f5;
    ram_cell[   11231] = 32'h0;  // 32'hcd12978f;
    ram_cell[   11232] = 32'h0;  // 32'h291f756b;
    ram_cell[   11233] = 32'h0;  // 32'h6a2bc6c8;
    ram_cell[   11234] = 32'h0;  // 32'h25c05c74;
    ram_cell[   11235] = 32'h0;  // 32'h88e60d39;
    ram_cell[   11236] = 32'h0;  // 32'h53a8e226;
    ram_cell[   11237] = 32'h0;  // 32'hd93bf389;
    ram_cell[   11238] = 32'h0;  // 32'ha349045b;
    ram_cell[   11239] = 32'h0;  // 32'h8da43549;
    ram_cell[   11240] = 32'h0;  // 32'h4ab46a0c;
    ram_cell[   11241] = 32'h0;  // 32'hd910df52;
    ram_cell[   11242] = 32'h0;  // 32'he9ccea32;
    ram_cell[   11243] = 32'h0;  // 32'hd3df486e;
    ram_cell[   11244] = 32'h0;  // 32'h96d30eea;
    ram_cell[   11245] = 32'h0;  // 32'hd4675ea4;
    ram_cell[   11246] = 32'h0;  // 32'h7162c1b7;
    ram_cell[   11247] = 32'h0;  // 32'hf9a3f9fb;
    ram_cell[   11248] = 32'h0;  // 32'h970fabdc;
    ram_cell[   11249] = 32'h0;  // 32'hb7857f4e;
    ram_cell[   11250] = 32'h0;  // 32'hff5a6d19;
    ram_cell[   11251] = 32'h0;  // 32'h561b4af8;
    ram_cell[   11252] = 32'h0;  // 32'hceeae348;
    ram_cell[   11253] = 32'h0;  // 32'hf4d60909;
    ram_cell[   11254] = 32'h0;  // 32'h0ea3fb52;
    ram_cell[   11255] = 32'h0;  // 32'h2a444332;
    ram_cell[   11256] = 32'h0;  // 32'hf0221d81;
    ram_cell[   11257] = 32'h0;  // 32'h6bfa1533;
    ram_cell[   11258] = 32'h0;  // 32'h22103706;
    ram_cell[   11259] = 32'h0;  // 32'hc5475b10;
    ram_cell[   11260] = 32'h0;  // 32'h17c84e13;
    ram_cell[   11261] = 32'h0;  // 32'h919112bb;
    ram_cell[   11262] = 32'h0;  // 32'h26fd70a5;
    ram_cell[   11263] = 32'h0;  // 32'h8c13ed21;
    ram_cell[   11264] = 32'h0;  // 32'h4b494556;
    ram_cell[   11265] = 32'h0;  // 32'he6219123;
    ram_cell[   11266] = 32'h0;  // 32'hbb8497c5;
    ram_cell[   11267] = 32'h0;  // 32'h2033df30;
    ram_cell[   11268] = 32'h0;  // 32'h4dd69aa9;
    ram_cell[   11269] = 32'h0;  // 32'ha377f8a2;
    ram_cell[   11270] = 32'h0;  // 32'h7636b963;
    ram_cell[   11271] = 32'h0;  // 32'h93a938ed;
    ram_cell[   11272] = 32'h0;  // 32'hfb72096d;
    ram_cell[   11273] = 32'h0;  // 32'hec3130f5;
    ram_cell[   11274] = 32'h0;  // 32'h613db067;
    ram_cell[   11275] = 32'h0;  // 32'h731350f8;
    ram_cell[   11276] = 32'h0;  // 32'h3e4c3653;
    ram_cell[   11277] = 32'h0;  // 32'h021ae30c;
    ram_cell[   11278] = 32'h0;  // 32'h59aebc9b;
    ram_cell[   11279] = 32'h0;  // 32'h1592202f;
    ram_cell[   11280] = 32'h0;  // 32'h4edb917a;
    ram_cell[   11281] = 32'h0;  // 32'hd0ba9333;
    ram_cell[   11282] = 32'h0;  // 32'h2d7f9c51;
    ram_cell[   11283] = 32'h0;  // 32'hf193d848;
    ram_cell[   11284] = 32'h0;  // 32'h42bafe2c;
    ram_cell[   11285] = 32'h0;  // 32'h5637cda3;
    ram_cell[   11286] = 32'h0;  // 32'h93dc6bc4;
    ram_cell[   11287] = 32'h0;  // 32'h3c00bb19;
    ram_cell[   11288] = 32'h0;  // 32'h3773ced5;
    ram_cell[   11289] = 32'h0;  // 32'h6a6387d7;
    ram_cell[   11290] = 32'h0;  // 32'h90b0b95d;
    ram_cell[   11291] = 32'h0;  // 32'hd8a060c6;
    ram_cell[   11292] = 32'h0;  // 32'hd5e3fcca;
    ram_cell[   11293] = 32'h0;  // 32'h9404e35d;
    ram_cell[   11294] = 32'h0;  // 32'h2df5e7f6;
    ram_cell[   11295] = 32'h0;  // 32'h06d63ca5;
    ram_cell[   11296] = 32'h0;  // 32'h6498dd1b;
    ram_cell[   11297] = 32'h0;  // 32'ha0079750;
    ram_cell[   11298] = 32'h0;  // 32'ha15b2cad;
    ram_cell[   11299] = 32'h0;  // 32'h0b994ef3;
    ram_cell[   11300] = 32'h0;  // 32'h4e2ae253;
    ram_cell[   11301] = 32'h0;  // 32'h74960d40;
    ram_cell[   11302] = 32'h0;  // 32'hf90ef2bb;
    ram_cell[   11303] = 32'h0;  // 32'h13e303e0;
    ram_cell[   11304] = 32'h0;  // 32'h3f031a55;
    ram_cell[   11305] = 32'h0;  // 32'hbd15819b;
    ram_cell[   11306] = 32'h0;  // 32'h732a4c53;
    ram_cell[   11307] = 32'h0;  // 32'hfd46b7c2;
    ram_cell[   11308] = 32'h0;  // 32'hce8d5ee2;
    ram_cell[   11309] = 32'h0;  // 32'h545a3538;
    ram_cell[   11310] = 32'h0;  // 32'h7af11b3f;
    ram_cell[   11311] = 32'h0;  // 32'hbefbd9a0;
    ram_cell[   11312] = 32'h0;  // 32'h2e4f0d3d;
    ram_cell[   11313] = 32'h0;  // 32'hf7f9f256;
    ram_cell[   11314] = 32'h0;  // 32'h23bc8dae;
    ram_cell[   11315] = 32'h0;  // 32'hcf7bd6ac;
    ram_cell[   11316] = 32'h0;  // 32'h9a61c8e9;
    ram_cell[   11317] = 32'h0;  // 32'hb0cf5c2c;
    ram_cell[   11318] = 32'h0;  // 32'h64931afd;
    ram_cell[   11319] = 32'h0;  // 32'h54169148;
    ram_cell[   11320] = 32'h0;  // 32'h6c2ac235;
    ram_cell[   11321] = 32'h0;  // 32'h74c9360f;
    ram_cell[   11322] = 32'h0;  // 32'hecf291ba;
    ram_cell[   11323] = 32'h0;  // 32'h992f362c;
    ram_cell[   11324] = 32'h0;  // 32'h10399fde;
    ram_cell[   11325] = 32'h0;  // 32'hd534e82f;
    ram_cell[   11326] = 32'h0;  // 32'h0e5176e6;
    ram_cell[   11327] = 32'h0;  // 32'h30f67e47;
    ram_cell[   11328] = 32'h0;  // 32'h5631d484;
    ram_cell[   11329] = 32'h0;  // 32'h0ccdcdaa;
    ram_cell[   11330] = 32'h0;  // 32'hc9631a06;
    ram_cell[   11331] = 32'h0;  // 32'h227264da;
    ram_cell[   11332] = 32'h0;  // 32'h32ec8ff7;
    ram_cell[   11333] = 32'h0;  // 32'h74802992;
    ram_cell[   11334] = 32'h0;  // 32'h985a457b;
    ram_cell[   11335] = 32'h0;  // 32'h19c35abf;
    ram_cell[   11336] = 32'h0;  // 32'h3cfade1d;
    ram_cell[   11337] = 32'h0;  // 32'hdbcc2dd5;
    ram_cell[   11338] = 32'h0;  // 32'hcbd8a699;
    ram_cell[   11339] = 32'h0;  // 32'hf316c4de;
    ram_cell[   11340] = 32'h0;  // 32'h08c8e4e9;
    ram_cell[   11341] = 32'h0;  // 32'ha59eb686;
    ram_cell[   11342] = 32'h0;  // 32'h066db447;
    ram_cell[   11343] = 32'h0;  // 32'h7ef1eff2;
    ram_cell[   11344] = 32'h0;  // 32'hc3479fc8;
    ram_cell[   11345] = 32'h0;  // 32'h34014b2f;
    ram_cell[   11346] = 32'h0;  // 32'h37e93cae;
    ram_cell[   11347] = 32'h0;  // 32'hf01e1b4b;
    ram_cell[   11348] = 32'h0;  // 32'h86b70d5b;
    ram_cell[   11349] = 32'h0;  // 32'h8d428d75;
    ram_cell[   11350] = 32'h0;  // 32'h23fe4af2;
    ram_cell[   11351] = 32'h0;  // 32'h53e52d06;
    ram_cell[   11352] = 32'h0;  // 32'ha7c4c23a;
    ram_cell[   11353] = 32'h0;  // 32'h9bbddeb4;
    ram_cell[   11354] = 32'h0;  // 32'h37e5e576;
    ram_cell[   11355] = 32'h0;  // 32'hb6b37160;
    ram_cell[   11356] = 32'h0;  // 32'h271b4ef1;
    ram_cell[   11357] = 32'h0;  // 32'h70fc38eb;
    ram_cell[   11358] = 32'h0;  // 32'hfbef54eb;
    ram_cell[   11359] = 32'h0;  // 32'h8addde70;
    ram_cell[   11360] = 32'h0;  // 32'hd3591635;
    ram_cell[   11361] = 32'h0;  // 32'hb1b1115e;
    ram_cell[   11362] = 32'h0;  // 32'h1cba9589;
    ram_cell[   11363] = 32'h0;  // 32'h741fbd04;
    ram_cell[   11364] = 32'h0;  // 32'h815898da;
    ram_cell[   11365] = 32'h0;  // 32'h0dba3aa5;
    ram_cell[   11366] = 32'h0;  // 32'h6d9b7d03;
    ram_cell[   11367] = 32'h0;  // 32'h76172489;
    ram_cell[   11368] = 32'h0;  // 32'h26d4ddf7;
    ram_cell[   11369] = 32'h0;  // 32'h04cd7d47;
    ram_cell[   11370] = 32'h0;  // 32'h647561a8;
    ram_cell[   11371] = 32'h0;  // 32'h523739c9;
    ram_cell[   11372] = 32'h0;  // 32'h823c4803;
    ram_cell[   11373] = 32'h0;  // 32'hedb69ca6;
    ram_cell[   11374] = 32'h0;  // 32'h06f85ab3;
    ram_cell[   11375] = 32'h0;  // 32'h15dc13d7;
    ram_cell[   11376] = 32'h0;  // 32'h675c1f86;
    ram_cell[   11377] = 32'h0;  // 32'h1d576799;
    ram_cell[   11378] = 32'h0;  // 32'h830fdd37;
    ram_cell[   11379] = 32'h0;  // 32'hc647bad8;
    ram_cell[   11380] = 32'h0;  // 32'hd1a388c8;
    ram_cell[   11381] = 32'h0;  // 32'h7add2c71;
    ram_cell[   11382] = 32'h0;  // 32'h9a2b090a;
    ram_cell[   11383] = 32'h0;  // 32'h16d332a9;
    ram_cell[   11384] = 32'h0;  // 32'h7d800234;
    ram_cell[   11385] = 32'h0;  // 32'h27ee084d;
    ram_cell[   11386] = 32'h0;  // 32'he6156456;
    ram_cell[   11387] = 32'h0;  // 32'h10ffd8f0;
    ram_cell[   11388] = 32'h0;  // 32'hd53e3a9e;
    ram_cell[   11389] = 32'h0;  // 32'h25817a04;
    ram_cell[   11390] = 32'h0;  // 32'ha1b64905;
    ram_cell[   11391] = 32'h0;  // 32'hc2f7159f;
    ram_cell[   11392] = 32'h0;  // 32'h002eb609;
    ram_cell[   11393] = 32'h0;  // 32'hf974f13d;
    ram_cell[   11394] = 32'h0;  // 32'hebf36d52;
    ram_cell[   11395] = 32'h0;  // 32'hc1e9054f;
    ram_cell[   11396] = 32'h0;  // 32'hc8d5087d;
    ram_cell[   11397] = 32'h0;  // 32'h3db6c42c;
    ram_cell[   11398] = 32'h0;  // 32'h34c83a34;
    ram_cell[   11399] = 32'h0;  // 32'hf938572e;
    ram_cell[   11400] = 32'h0;  // 32'h8e92870a;
    ram_cell[   11401] = 32'h0;  // 32'h1469c3a2;
    ram_cell[   11402] = 32'h0;  // 32'h44c4287c;
    ram_cell[   11403] = 32'h0;  // 32'h05d01625;
    ram_cell[   11404] = 32'h0;  // 32'h909a3bd4;
    ram_cell[   11405] = 32'h0;  // 32'h8d83c824;
    ram_cell[   11406] = 32'h0;  // 32'h13c3a642;
    ram_cell[   11407] = 32'h0;  // 32'h255d0b25;
    ram_cell[   11408] = 32'h0;  // 32'hb1cba93b;
    ram_cell[   11409] = 32'h0;  // 32'h74de09f9;
    ram_cell[   11410] = 32'h0;  // 32'hb39ffbe5;
    ram_cell[   11411] = 32'h0;  // 32'hd080ad51;
    ram_cell[   11412] = 32'h0;  // 32'hb3afcf47;
    ram_cell[   11413] = 32'h0;  // 32'h28c841e1;
    ram_cell[   11414] = 32'h0;  // 32'h8103fd4b;
    ram_cell[   11415] = 32'h0;  // 32'hb7fc3648;
    ram_cell[   11416] = 32'h0;  // 32'hb5f6ea44;
    ram_cell[   11417] = 32'h0;  // 32'h41468641;
    ram_cell[   11418] = 32'h0;  // 32'h19d6b64b;
    ram_cell[   11419] = 32'h0;  // 32'h54e481b1;
    ram_cell[   11420] = 32'h0;  // 32'h8f944292;
    ram_cell[   11421] = 32'h0;  // 32'hba4bf058;
    ram_cell[   11422] = 32'h0;  // 32'h347df4a1;
    ram_cell[   11423] = 32'h0;  // 32'h11dcec49;
    ram_cell[   11424] = 32'h0;  // 32'h267b8659;
    ram_cell[   11425] = 32'h0;  // 32'h4418eaa0;
    ram_cell[   11426] = 32'h0;  // 32'hcf8fbcd6;
    ram_cell[   11427] = 32'h0;  // 32'h8bf70411;
    ram_cell[   11428] = 32'h0;  // 32'h9d1b9820;
    ram_cell[   11429] = 32'h0;  // 32'h7ee42367;
    ram_cell[   11430] = 32'h0;  // 32'hf39fcd81;
    ram_cell[   11431] = 32'h0;  // 32'h8d5a877c;
    ram_cell[   11432] = 32'h0;  // 32'h2863acf8;
    ram_cell[   11433] = 32'h0;  // 32'h1812b750;
    ram_cell[   11434] = 32'h0;  // 32'h67145e25;
    ram_cell[   11435] = 32'h0;  // 32'hf159099d;
    ram_cell[   11436] = 32'h0;  // 32'hde0c86ad;
    ram_cell[   11437] = 32'h0;  // 32'h268585e9;
    ram_cell[   11438] = 32'h0;  // 32'h48a223b1;
    ram_cell[   11439] = 32'h0;  // 32'h9c50e2ab;
    ram_cell[   11440] = 32'h0;  // 32'hf08af699;
    ram_cell[   11441] = 32'h0;  // 32'hae8ce46e;
    ram_cell[   11442] = 32'h0;  // 32'h7e0d3d4c;
    ram_cell[   11443] = 32'h0;  // 32'h1d21754f;
    ram_cell[   11444] = 32'h0;  // 32'h23e7c8f7;
    ram_cell[   11445] = 32'h0;  // 32'hd151d923;
    ram_cell[   11446] = 32'h0;  // 32'hdda17b49;
    ram_cell[   11447] = 32'h0;  // 32'h62148260;
    ram_cell[   11448] = 32'h0;  // 32'h430727aa;
    ram_cell[   11449] = 32'h0;  // 32'hd08d10eb;
    ram_cell[   11450] = 32'h0;  // 32'h0a390f20;
    ram_cell[   11451] = 32'h0;  // 32'h434b9b13;
    ram_cell[   11452] = 32'h0;  // 32'hb0d8c4f4;
    ram_cell[   11453] = 32'h0;  // 32'h9e138dc5;
    ram_cell[   11454] = 32'h0;  // 32'h61987192;
    ram_cell[   11455] = 32'h0;  // 32'h7a2b50c3;
    ram_cell[   11456] = 32'h0;  // 32'h3bcad10f;
    ram_cell[   11457] = 32'h0;  // 32'hca110cf7;
    ram_cell[   11458] = 32'h0;  // 32'h281c2858;
    ram_cell[   11459] = 32'h0;  // 32'h5fa24a4f;
    ram_cell[   11460] = 32'h0;  // 32'h4d43ebd5;
    ram_cell[   11461] = 32'h0;  // 32'h64ed8f43;
    ram_cell[   11462] = 32'h0;  // 32'ha3c865b4;
    ram_cell[   11463] = 32'h0;  // 32'hd4d8d369;
    ram_cell[   11464] = 32'h0;  // 32'h4f0874a4;
    ram_cell[   11465] = 32'h0;  // 32'h8de8d4a0;
    ram_cell[   11466] = 32'h0;  // 32'he48d68e1;
    ram_cell[   11467] = 32'h0;  // 32'h1879e26d;
    ram_cell[   11468] = 32'h0;  // 32'h9e4b5d11;
    ram_cell[   11469] = 32'h0;  // 32'he233efc3;
    ram_cell[   11470] = 32'h0;  // 32'h4a1c86bd;
    ram_cell[   11471] = 32'h0;  // 32'hc69e8427;
    ram_cell[   11472] = 32'h0;  // 32'h1fc2f1b9;
    ram_cell[   11473] = 32'h0;  // 32'h30b99c4a;
    ram_cell[   11474] = 32'h0;  // 32'h1f7aa4ca;
    ram_cell[   11475] = 32'h0;  // 32'h3efb89c6;
    ram_cell[   11476] = 32'h0;  // 32'h0dc6cd91;
    ram_cell[   11477] = 32'h0;  // 32'h15e20521;
    ram_cell[   11478] = 32'h0;  // 32'h6075a1ca;
    ram_cell[   11479] = 32'h0;  // 32'h2b8485e1;
    ram_cell[   11480] = 32'h0;  // 32'hd9a3b3ba;
    ram_cell[   11481] = 32'h0;  // 32'h53029cfe;
    ram_cell[   11482] = 32'h0;  // 32'h4bd554d4;
    ram_cell[   11483] = 32'h0;  // 32'h8e30869a;
    ram_cell[   11484] = 32'h0;  // 32'hf64c30e4;
    ram_cell[   11485] = 32'h0;  // 32'h525997c8;
    ram_cell[   11486] = 32'h0;  // 32'h6f286214;
    ram_cell[   11487] = 32'h0;  // 32'h1f387769;
    ram_cell[   11488] = 32'h0;  // 32'h19e719a6;
    ram_cell[   11489] = 32'h0;  // 32'hd9402aef;
    ram_cell[   11490] = 32'h0;  // 32'h39f7ef43;
    ram_cell[   11491] = 32'h0;  // 32'had3e9b34;
    ram_cell[   11492] = 32'h0;  // 32'h4f53698b;
    ram_cell[   11493] = 32'h0;  // 32'h9e62e17c;
    ram_cell[   11494] = 32'h0;  // 32'h78e95e68;
    ram_cell[   11495] = 32'h0;  // 32'hd6b38d27;
    ram_cell[   11496] = 32'h0;  // 32'h4b6c7d62;
    ram_cell[   11497] = 32'h0;  // 32'ha8f43df6;
    ram_cell[   11498] = 32'h0;  // 32'hc7fe4a49;
    ram_cell[   11499] = 32'h0;  // 32'h7771935e;
    ram_cell[   11500] = 32'h0;  // 32'hc264589a;
    ram_cell[   11501] = 32'h0;  // 32'h3c548aac;
    ram_cell[   11502] = 32'h0;  // 32'h1c52e3db;
    ram_cell[   11503] = 32'h0;  // 32'hd2aba53c;
    ram_cell[   11504] = 32'h0;  // 32'h4a6ab517;
    ram_cell[   11505] = 32'h0;  // 32'hed3223ad;
    ram_cell[   11506] = 32'h0;  // 32'hf693ef18;
    ram_cell[   11507] = 32'h0;  // 32'h3c7a3005;
    ram_cell[   11508] = 32'h0;  // 32'hf8878082;
    ram_cell[   11509] = 32'h0;  // 32'hc87b6b64;
    ram_cell[   11510] = 32'h0;  // 32'h5869a46a;
    ram_cell[   11511] = 32'h0;  // 32'hf58ab258;
    ram_cell[   11512] = 32'h0;  // 32'hf9adc438;
    ram_cell[   11513] = 32'h0;  // 32'he229d8ff;
    ram_cell[   11514] = 32'h0;  // 32'h20243b26;
    ram_cell[   11515] = 32'h0;  // 32'h43cb3989;
    ram_cell[   11516] = 32'h0;  // 32'ha7316be2;
    ram_cell[   11517] = 32'h0;  // 32'h26ac80bc;
    ram_cell[   11518] = 32'h0;  // 32'hd4cce5bd;
    ram_cell[   11519] = 32'h0;  // 32'h8979e098;
    ram_cell[   11520] = 32'h0;  // 32'hed0bb4e0;
    ram_cell[   11521] = 32'h0;  // 32'he2fc91bf;
    ram_cell[   11522] = 32'h0;  // 32'h1347cafe;
    ram_cell[   11523] = 32'h0;  // 32'h18589677;
    ram_cell[   11524] = 32'h0;  // 32'h1bb3527e;
    ram_cell[   11525] = 32'h0;  // 32'h2e4dd752;
    ram_cell[   11526] = 32'h0;  // 32'hc47a857a;
    ram_cell[   11527] = 32'h0;  // 32'h46d309b1;
    ram_cell[   11528] = 32'h0;  // 32'ha97d26f6;
    ram_cell[   11529] = 32'h0;  // 32'h7815b525;
    ram_cell[   11530] = 32'h0;  // 32'hf6b0060d;
    ram_cell[   11531] = 32'h0;  // 32'hffac66fc;
    ram_cell[   11532] = 32'h0;  // 32'h25b22d36;
    ram_cell[   11533] = 32'h0;  // 32'h82778353;
    ram_cell[   11534] = 32'h0;  // 32'hcd2b6b1a;
    ram_cell[   11535] = 32'h0;  // 32'h6d748088;
    ram_cell[   11536] = 32'h0;  // 32'h67f54ee9;
    ram_cell[   11537] = 32'h0;  // 32'habaadf3e;
    ram_cell[   11538] = 32'h0;  // 32'h5fd2a69d;
    ram_cell[   11539] = 32'h0;  // 32'he28dbc11;
    ram_cell[   11540] = 32'h0;  // 32'h7602eb9b;
    ram_cell[   11541] = 32'h0;  // 32'h3a190ca5;
    ram_cell[   11542] = 32'h0;  // 32'h143cec6d;
    ram_cell[   11543] = 32'h0;  // 32'h285403ab;
    ram_cell[   11544] = 32'h0;  // 32'h6c4826b1;
    ram_cell[   11545] = 32'h0;  // 32'h1e64a8bc;
    ram_cell[   11546] = 32'h0;  // 32'h8f90d4e6;
    ram_cell[   11547] = 32'h0;  // 32'h0dc72c9b;
    ram_cell[   11548] = 32'h0;  // 32'h38a5ae33;
    ram_cell[   11549] = 32'h0;  // 32'h620b2d69;
    ram_cell[   11550] = 32'h0;  // 32'hc3bad39d;
    ram_cell[   11551] = 32'h0;  // 32'h2fdff96d;
    ram_cell[   11552] = 32'h0;  // 32'h995da319;
    ram_cell[   11553] = 32'h0;  // 32'h8e7d24e6;
    ram_cell[   11554] = 32'h0;  // 32'ha33349f7;
    ram_cell[   11555] = 32'h0;  // 32'hb4f874c8;
    ram_cell[   11556] = 32'h0;  // 32'hfed44de9;
    ram_cell[   11557] = 32'h0;  // 32'ha08076db;
    ram_cell[   11558] = 32'h0;  // 32'hadc6888e;
    ram_cell[   11559] = 32'h0;  // 32'h2d6cff03;
    ram_cell[   11560] = 32'h0;  // 32'he8820652;
    ram_cell[   11561] = 32'h0;  // 32'h8abc7743;
    ram_cell[   11562] = 32'h0;  // 32'h9ef40bb9;
    ram_cell[   11563] = 32'h0;  // 32'h5001c3d1;
    ram_cell[   11564] = 32'h0;  // 32'h6e0df928;
    ram_cell[   11565] = 32'h0;  // 32'he072f200;
    ram_cell[   11566] = 32'h0;  // 32'hd5669361;
    ram_cell[   11567] = 32'h0;  // 32'h42811159;
    ram_cell[   11568] = 32'h0;  // 32'h723feb53;
    ram_cell[   11569] = 32'h0;  // 32'h695228d7;
    ram_cell[   11570] = 32'h0;  // 32'h2592b2e8;
    ram_cell[   11571] = 32'h0;  // 32'hd198f9ca;
    ram_cell[   11572] = 32'h0;  // 32'hc35f4822;
    ram_cell[   11573] = 32'h0;  // 32'hf8d13d6e;
    ram_cell[   11574] = 32'h0;  // 32'h6f969376;
    ram_cell[   11575] = 32'h0;  // 32'hc62d85f3;
    ram_cell[   11576] = 32'h0;  // 32'hcf2f4cff;
    ram_cell[   11577] = 32'h0;  // 32'h6385089e;
    ram_cell[   11578] = 32'h0;  // 32'hb9d5c3b8;
    ram_cell[   11579] = 32'h0;  // 32'hd5e89f07;
    ram_cell[   11580] = 32'h0;  // 32'hc9cd9ad8;
    ram_cell[   11581] = 32'h0;  // 32'he54c1198;
    ram_cell[   11582] = 32'h0;  // 32'h0a705e1a;
    ram_cell[   11583] = 32'h0;  // 32'hec5c1c63;
    ram_cell[   11584] = 32'h0;  // 32'h678579a1;
    ram_cell[   11585] = 32'h0;  // 32'he55d1c68;
    ram_cell[   11586] = 32'h0;  // 32'he385509e;
    ram_cell[   11587] = 32'h0;  // 32'h53950ffa;
    ram_cell[   11588] = 32'h0;  // 32'hf6be8edd;
    ram_cell[   11589] = 32'h0;  // 32'hbebe9d92;
    ram_cell[   11590] = 32'h0;  // 32'h4aed87e2;
    ram_cell[   11591] = 32'h0;  // 32'h8fd504bc;
    ram_cell[   11592] = 32'h0;  // 32'h9091b90e;
    ram_cell[   11593] = 32'h0;  // 32'h75095768;
    ram_cell[   11594] = 32'h0;  // 32'h6035579f;
    ram_cell[   11595] = 32'h0;  // 32'h8ce41d07;
    ram_cell[   11596] = 32'h0;  // 32'h55ccf114;
    ram_cell[   11597] = 32'h0;  // 32'he86e48f4;
    ram_cell[   11598] = 32'h0;  // 32'h29317a4a;
    ram_cell[   11599] = 32'h0;  // 32'hd07a35c7;
    ram_cell[   11600] = 32'h0;  // 32'h6701bb4d;
    ram_cell[   11601] = 32'h0;  // 32'he2912169;
    ram_cell[   11602] = 32'h0;  // 32'h518ecf47;
    ram_cell[   11603] = 32'h0;  // 32'h6fc17b6d;
    ram_cell[   11604] = 32'h0;  // 32'hf1751f84;
    ram_cell[   11605] = 32'h0;  // 32'hd1bf1e58;
    ram_cell[   11606] = 32'h0;  // 32'h207c5161;
    ram_cell[   11607] = 32'h0;  // 32'h057d013d;
    ram_cell[   11608] = 32'h0;  // 32'h403af051;
    ram_cell[   11609] = 32'h0;  // 32'h2f9d6653;
    ram_cell[   11610] = 32'h0;  // 32'h1068b910;
    ram_cell[   11611] = 32'h0;  // 32'h9c62ec14;
    ram_cell[   11612] = 32'h0;  // 32'hd502482f;
    ram_cell[   11613] = 32'h0;  // 32'h62ed2774;
    ram_cell[   11614] = 32'h0;  // 32'hcb63a32e;
    ram_cell[   11615] = 32'h0;  // 32'h5d20dc67;
    ram_cell[   11616] = 32'h0;  // 32'hb4e09086;
    ram_cell[   11617] = 32'h0;  // 32'hb9b71e07;
    ram_cell[   11618] = 32'h0;  // 32'h07d1d5b3;
    ram_cell[   11619] = 32'h0;  // 32'h8af5fb49;
    ram_cell[   11620] = 32'h0;  // 32'h2dafff4b;
    ram_cell[   11621] = 32'h0;  // 32'h82b8e957;
    ram_cell[   11622] = 32'h0;  // 32'h29a81e40;
    ram_cell[   11623] = 32'h0;  // 32'hbeac33a3;
    ram_cell[   11624] = 32'h0;  // 32'hcec32217;
    ram_cell[   11625] = 32'h0;  // 32'hb3dc4483;
    ram_cell[   11626] = 32'h0;  // 32'hd07d479c;
    ram_cell[   11627] = 32'h0;  // 32'h7ea6c2e3;
    ram_cell[   11628] = 32'h0;  // 32'h8460bfa6;
    ram_cell[   11629] = 32'h0;  // 32'h477b93b1;
    ram_cell[   11630] = 32'h0;  // 32'hf1cb155a;
    ram_cell[   11631] = 32'h0;  // 32'hd921873d;
    ram_cell[   11632] = 32'h0;  // 32'h7e75d2b4;
    ram_cell[   11633] = 32'h0;  // 32'h1f543776;
    ram_cell[   11634] = 32'h0;  // 32'he172e598;
    ram_cell[   11635] = 32'h0;  // 32'h5722b412;
    ram_cell[   11636] = 32'h0;  // 32'h761eea9c;
    ram_cell[   11637] = 32'h0;  // 32'hdeb01089;
    ram_cell[   11638] = 32'h0;  // 32'h4f1fc5b6;
    ram_cell[   11639] = 32'h0;  // 32'ha9bda269;
    ram_cell[   11640] = 32'h0;  // 32'hc10b4785;
    ram_cell[   11641] = 32'h0;  // 32'hda016788;
    ram_cell[   11642] = 32'h0;  // 32'h4d5712eb;
    ram_cell[   11643] = 32'h0;  // 32'h605ab59d;
    ram_cell[   11644] = 32'h0;  // 32'hcda126db;
    ram_cell[   11645] = 32'h0;  // 32'hb5efcc79;
    ram_cell[   11646] = 32'h0;  // 32'h95de1973;
    ram_cell[   11647] = 32'h0;  // 32'h5816afe8;
    ram_cell[   11648] = 32'h0;  // 32'h1e3ab4b4;
    ram_cell[   11649] = 32'h0;  // 32'h64f814e0;
    ram_cell[   11650] = 32'h0;  // 32'hb0a71255;
    ram_cell[   11651] = 32'h0;  // 32'hf4bd54f4;
    ram_cell[   11652] = 32'h0;  // 32'h259749e7;
    ram_cell[   11653] = 32'h0;  // 32'h3f2fd575;
    ram_cell[   11654] = 32'h0;  // 32'hf495c413;
    ram_cell[   11655] = 32'h0;  // 32'ha5fa9ad9;
    ram_cell[   11656] = 32'h0;  // 32'h197dea38;
    ram_cell[   11657] = 32'h0;  // 32'h1a5de848;
    ram_cell[   11658] = 32'h0;  // 32'h46c18265;
    ram_cell[   11659] = 32'h0;  // 32'h769aa67c;
    ram_cell[   11660] = 32'h0;  // 32'hf9e01eaf;
    ram_cell[   11661] = 32'h0;  // 32'hb743a046;
    ram_cell[   11662] = 32'h0;  // 32'h61048c5b;
    ram_cell[   11663] = 32'h0;  // 32'h863a77ff;
    ram_cell[   11664] = 32'h0;  // 32'h849b20c5;
    ram_cell[   11665] = 32'h0;  // 32'h41c5beb8;
    ram_cell[   11666] = 32'h0;  // 32'hddce1423;
    ram_cell[   11667] = 32'h0;  // 32'ha0ff1f18;
    ram_cell[   11668] = 32'h0;  // 32'h40f96a11;
    ram_cell[   11669] = 32'h0;  // 32'h16cc630c;
    ram_cell[   11670] = 32'h0;  // 32'hdfe24f98;
    ram_cell[   11671] = 32'h0;  // 32'heb27ec38;
    ram_cell[   11672] = 32'h0;  // 32'he58031f0;
    ram_cell[   11673] = 32'h0;  // 32'h51fd260a;
    ram_cell[   11674] = 32'h0;  // 32'h8e462702;
    ram_cell[   11675] = 32'h0;  // 32'h77fb3445;
    ram_cell[   11676] = 32'h0;  // 32'h17d19174;
    ram_cell[   11677] = 32'h0;  // 32'hfaa45eba;
    ram_cell[   11678] = 32'h0;  // 32'hba17624c;
    ram_cell[   11679] = 32'h0;  // 32'h5a4b3600;
    ram_cell[   11680] = 32'h0;  // 32'hcb7ebe94;
    ram_cell[   11681] = 32'h0;  // 32'h02985da6;
    ram_cell[   11682] = 32'h0;  // 32'h2264a2d4;
    ram_cell[   11683] = 32'h0;  // 32'h0cc9106f;
    ram_cell[   11684] = 32'h0;  // 32'h0738dacc;
    ram_cell[   11685] = 32'h0;  // 32'h4f2779af;
    ram_cell[   11686] = 32'h0;  // 32'h9e3ad9dd;
    ram_cell[   11687] = 32'h0;  // 32'h83f52553;
    ram_cell[   11688] = 32'h0;  // 32'hd10a8035;
    ram_cell[   11689] = 32'h0;  // 32'h021af608;
    ram_cell[   11690] = 32'h0;  // 32'h46b5d20b;
    ram_cell[   11691] = 32'h0;  // 32'h46b83756;
    ram_cell[   11692] = 32'h0;  // 32'h986ccf08;
    ram_cell[   11693] = 32'h0;  // 32'hf5a71782;
    ram_cell[   11694] = 32'h0;  // 32'h2221908f;
    ram_cell[   11695] = 32'h0;  // 32'hded3077f;
    ram_cell[   11696] = 32'h0;  // 32'h11b7c53d;
    ram_cell[   11697] = 32'h0;  // 32'h9794c467;
    ram_cell[   11698] = 32'h0;  // 32'ha0acc5e1;
    ram_cell[   11699] = 32'h0;  // 32'h3f3ccfd1;
    ram_cell[   11700] = 32'h0;  // 32'h59717ab9;
    ram_cell[   11701] = 32'h0;  // 32'h3a5d572d;
    ram_cell[   11702] = 32'h0;  // 32'hdb33dfb8;
    ram_cell[   11703] = 32'h0;  // 32'h692e99cb;
    ram_cell[   11704] = 32'h0;  // 32'h4d25dd43;
    ram_cell[   11705] = 32'h0;  // 32'h19460391;
    ram_cell[   11706] = 32'h0;  // 32'hef795a44;
    ram_cell[   11707] = 32'h0;  // 32'he0343fe8;
    ram_cell[   11708] = 32'h0;  // 32'h6934bbfd;
    ram_cell[   11709] = 32'h0;  // 32'h1bb42c2e;
    ram_cell[   11710] = 32'h0;  // 32'h93eadb0b;
    ram_cell[   11711] = 32'h0;  // 32'h58c63b48;
    ram_cell[   11712] = 32'h0;  // 32'ha8dda77a;
    ram_cell[   11713] = 32'h0;  // 32'h221b9500;
    ram_cell[   11714] = 32'h0;  // 32'h7b47f485;
    ram_cell[   11715] = 32'h0;  // 32'h75d08e47;
    ram_cell[   11716] = 32'h0;  // 32'hf47bcadc;
    ram_cell[   11717] = 32'h0;  // 32'h56ea8326;
    ram_cell[   11718] = 32'h0;  // 32'hb4ceaefb;
    ram_cell[   11719] = 32'h0;  // 32'h485298d8;
    ram_cell[   11720] = 32'h0;  // 32'h3418b4ae;
    ram_cell[   11721] = 32'h0;  // 32'ha3dd38fe;
    ram_cell[   11722] = 32'h0;  // 32'ha3499879;
    ram_cell[   11723] = 32'h0;  // 32'haa69ae55;
    ram_cell[   11724] = 32'h0;  // 32'he8f72054;
    ram_cell[   11725] = 32'h0;  // 32'h625f7f4a;
    ram_cell[   11726] = 32'h0;  // 32'hd78cbd08;
    ram_cell[   11727] = 32'h0;  // 32'hb27ffeb6;
    ram_cell[   11728] = 32'h0;  // 32'hfe6d4d2f;
    ram_cell[   11729] = 32'h0;  // 32'hbee4a52f;
    ram_cell[   11730] = 32'h0;  // 32'hd056ee4a;
    ram_cell[   11731] = 32'h0;  // 32'hfb8634c9;
    ram_cell[   11732] = 32'h0;  // 32'h15851939;
    ram_cell[   11733] = 32'h0;  // 32'h93cadeed;
    ram_cell[   11734] = 32'h0;  // 32'hc196208d;
    ram_cell[   11735] = 32'h0;  // 32'h75dbd321;
    ram_cell[   11736] = 32'h0;  // 32'hb09ced7b;
    ram_cell[   11737] = 32'h0;  // 32'h8a51d13e;
    ram_cell[   11738] = 32'h0;  // 32'hddd7ca5b;
    ram_cell[   11739] = 32'h0;  // 32'h6bd477d9;
    ram_cell[   11740] = 32'h0;  // 32'h2d2bb77d;
    ram_cell[   11741] = 32'h0;  // 32'h66e56920;
    ram_cell[   11742] = 32'h0;  // 32'h94c57dec;
    ram_cell[   11743] = 32'h0;  // 32'haebd237e;
    ram_cell[   11744] = 32'h0;  // 32'h763a6e7b;
    ram_cell[   11745] = 32'h0;  // 32'h13145bdb;
    ram_cell[   11746] = 32'h0;  // 32'ha5c80ff5;
    ram_cell[   11747] = 32'h0;  // 32'h2c64b9e1;
    ram_cell[   11748] = 32'h0;  // 32'hb5bf85ec;
    ram_cell[   11749] = 32'h0;  // 32'hbf150edf;
    ram_cell[   11750] = 32'h0;  // 32'h76621fee;
    ram_cell[   11751] = 32'h0;  // 32'h4b2512ee;
    ram_cell[   11752] = 32'h0;  // 32'hbe85a0fd;
    ram_cell[   11753] = 32'h0;  // 32'h85026535;
    ram_cell[   11754] = 32'h0;  // 32'hee00f4bf;
    ram_cell[   11755] = 32'h0;  // 32'hf171352b;
    ram_cell[   11756] = 32'h0;  // 32'h84ba8f80;
    ram_cell[   11757] = 32'h0;  // 32'h34f17b92;
    ram_cell[   11758] = 32'h0;  // 32'h0808ac35;
    ram_cell[   11759] = 32'h0;  // 32'h670c8170;
    ram_cell[   11760] = 32'h0;  // 32'h8c24b418;
    ram_cell[   11761] = 32'h0;  // 32'hbef0dc31;
    ram_cell[   11762] = 32'h0;  // 32'h5c4be2c7;
    ram_cell[   11763] = 32'h0;  // 32'h20ffb82e;
    ram_cell[   11764] = 32'h0;  // 32'ha7213d6b;
    ram_cell[   11765] = 32'h0;  // 32'h7c35419e;
    ram_cell[   11766] = 32'h0;  // 32'h36c964cf;
    ram_cell[   11767] = 32'h0;  // 32'hf79508fe;
    ram_cell[   11768] = 32'h0;  // 32'h4b429a64;
    ram_cell[   11769] = 32'h0;  // 32'hca7e8e6c;
    ram_cell[   11770] = 32'h0;  // 32'h090b61ed;
    ram_cell[   11771] = 32'h0;  // 32'hdd245826;
    ram_cell[   11772] = 32'h0;  // 32'h968e24a7;
    ram_cell[   11773] = 32'h0;  // 32'h1eb4d083;
    ram_cell[   11774] = 32'h0;  // 32'h429a97d4;
    ram_cell[   11775] = 32'h0;  // 32'ha1a8a3b3;
    ram_cell[   11776] = 32'h0;  // 32'h87d49801;
    ram_cell[   11777] = 32'h0;  // 32'h9d48a562;
    ram_cell[   11778] = 32'h0;  // 32'h942725cf;
    ram_cell[   11779] = 32'h0;  // 32'h5d08321a;
    ram_cell[   11780] = 32'h0;  // 32'hefafa233;
    ram_cell[   11781] = 32'h0;  // 32'hf9dab0b4;
    ram_cell[   11782] = 32'h0;  // 32'h0baf6913;
    ram_cell[   11783] = 32'h0;  // 32'h4093001d;
    ram_cell[   11784] = 32'h0;  // 32'ha327a029;
    ram_cell[   11785] = 32'h0;  // 32'he95c646f;
    ram_cell[   11786] = 32'h0;  // 32'h5a8932af;
    ram_cell[   11787] = 32'h0;  // 32'h013c6fa0;
    ram_cell[   11788] = 32'h0;  // 32'h3f5d29a5;
    ram_cell[   11789] = 32'h0;  // 32'hd89d4725;
    ram_cell[   11790] = 32'h0;  // 32'h8849a720;
    ram_cell[   11791] = 32'h0;  // 32'hdcc84d95;
    ram_cell[   11792] = 32'h0;  // 32'he842efbb;
    ram_cell[   11793] = 32'h0;  // 32'h06327a44;
    ram_cell[   11794] = 32'h0;  // 32'h4fbe07ea;
    ram_cell[   11795] = 32'h0;  // 32'hb65561e3;
    ram_cell[   11796] = 32'h0;  // 32'ha0945f3e;
    ram_cell[   11797] = 32'h0;  // 32'h6efd19f3;
    ram_cell[   11798] = 32'h0;  // 32'h11e95206;
    ram_cell[   11799] = 32'h0;  // 32'h44412f18;
    ram_cell[   11800] = 32'h0;  // 32'hec3677f9;
    ram_cell[   11801] = 32'h0;  // 32'h49d63171;
    ram_cell[   11802] = 32'h0;  // 32'hb44c5dec;
    ram_cell[   11803] = 32'h0;  // 32'ha0413eae;
    ram_cell[   11804] = 32'h0;  // 32'hc389f422;
    ram_cell[   11805] = 32'h0;  // 32'h699691f2;
    ram_cell[   11806] = 32'h0;  // 32'h9bf784c9;
    ram_cell[   11807] = 32'h0;  // 32'h2edd2166;
    ram_cell[   11808] = 32'h0;  // 32'hd4330864;
    ram_cell[   11809] = 32'h0;  // 32'h31446be1;
    ram_cell[   11810] = 32'h0;  // 32'h02e88963;
    ram_cell[   11811] = 32'h0;  // 32'hfde61187;
    ram_cell[   11812] = 32'h0;  // 32'hcfbfa537;
    ram_cell[   11813] = 32'h0;  // 32'h4ed6a0ca;
    ram_cell[   11814] = 32'h0;  // 32'ha6eb862d;
    ram_cell[   11815] = 32'h0;  // 32'h96e4554c;
    ram_cell[   11816] = 32'h0;  // 32'h5c40d69f;
    ram_cell[   11817] = 32'h0;  // 32'hc53ff886;
    ram_cell[   11818] = 32'h0;  // 32'h4d622a86;
    ram_cell[   11819] = 32'h0;  // 32'h5199c819;
    ram_cell[   11820] = 32'h0;  // 32'hde2111e4;
    ram_cell[   11821] = 32'h0;  // 32'h8bd1bacd;
    ram_cell[   11822] = 32'h0;  // 32'hd797915e;
    ram_cell[   11823] = 32'h0;  // 32'h203075a8;
    ram_cell[   11824] = 32'h0;  // 32'h12b7d2df;
    ram_cell[   11825] = 32'h0;  // 32'h51526739;
    ram_cell[   11826] = 32'h0;  // 32'h4e0c8a71;
    ram_cell[   11827] = 32'h0;  // 32'h1e38215e;
    ram_cell[   11828] = 32'h0;  // 32'hc9d47d3b;
    ram_cell[   11829] = 32'h0;  // 32'h9ee42978;
    ram_cell[   11830] = 32'h0;  // 32'ha6ead116;
    ram_cell[   11831] = 32'h0;  // 32'h74c24941;
    ram_cell[   11832] = 32'h0;  // 32'h23d60f5a;
    ram_cell[   11833] = 32'h0;  // 32'h5ec67fe9;
    ram_cell[   11834] = 32'h0;  // 32'hf6dd5ffd;
    ram_cell[   11835] = 32'h0;  // 32'h851921fe;
    ram_cell[   11836] = 32'h0;  // 32'h620c03db;
    ram_cell[   11837] = 32'h0;  // 32'h8b49c713;
    ram_cell[   11838] = 32'h0;  // 32'h493debff;
    ram_cell[   11839] = 32'h0;  // 32'h09e8d4c1;
    ram_cell[   11840] = 32'h0;  // 32'hd76b2dbf;
    ram_cell[   11841] = 32'h0;  // 32'h026892e3;
    ram_cell[   11842] = 32'h0;  // 32'h39566d6f;
    ram_cell[   11843] = 32'h0;  // 32'ha37fe55f;
    ram_cell[   11844] = 32'h0;  // 32'h78d36694;
    ram_cell[   11845] = 32'h0;  // 32'hb28a7ecc;
    ram_cell[   11846] = 32'h0;  // 32'heb728087;
    ram_cell[   11847] = 32'h0;  // 32'h7cbbbb69;
    ram_cell[   11848] = 32'h0;  // 32'he8b9176f;
    ram_cell[   11849] = 32'h0;  // 32'hdee76aea;
    ram_cell[   11850] = 32'h0;  // 32'hdf2a2b1c;
    ram_cell[   11851] = 32'h0;  // 32'h0749bf88;
    ram_cell[   11852] = 32'h0;  // 32'hfe01c41c;
    ram_cell[   11853] = 32'h0;  // 32'hce2c44a1;
    ram_cell[   11854] = 32'h0;  // 32'h61e04139;
    ram_cell[   11855] = 32'h0;  // 32'h2334895c;
    ram_cell[   11856] = 32'h0;  // 32'h6f1298db;
    ram_cell[   11857] = 32'h0;  // 32'h83831cb9;
    ram_cell[   11858] = 32'h0;  // 32'h9335cb38;
    ram_cell[   11859] = 32'h0;  // 32'h8ba89f94;
    ram_cell[   11860] = 32'h0;  // 32'h818f34e1;
    ram_cell[   11861] = 32'h0;  // 32'hcecc54a8;
    ram_cell[   11862] = 32'h0;  // 32'h1ab599d2;
    ram_cell[   11863] = 32'h0;  // 32'hd0b77d35;
    ram_cell[   11864] = 32'h0;  // 32'h605ccc06;
    ram_cell[   11865] = 32'h0;  // 32'h66b5d7d2;
    ram_cell[   11866] = 32'h0;  // 32'hea0fe4d9;
    ram_cell[   11867] = 32'h0;  // 32'he0ab40fa;
    ram_cell[   11868] = 32'h0;  // 32'ha566ce95;
    ram_cell[   11869] = 32'h0;  // 32'h0db2c3d4;
    ram_cell[   11870] = 32'h0;  // 32'h2116e6c3;
    ram_cell[   11871] = 32'h0;  // 32'h8ec6ee22;
    ram_cell[   11872] = 32'h0;  // 32'h3efc80e4;
    ram_cell[   11873] = 32'h0;  // 32'h31be1bfa;
    ram_cell[   11874] = 32'h0;  // 32'h77f729e6;
    ram_cell[   11875] = 32'h0;  // 32'h3948ed35;
    ram_cell[   11876] = 32'h0;  // 32'h119c2d26;
    ram_cell[   11877] = 32'h0;  // 32'h83284837;
    ram_cell[   11878] = 32'h0;  // 32'h8688b9c4;
    ram_cell[   11879] = 32'h0;  // 32'h07257655;
    ram_cell[   11880] = 32'h0;  // 32'hd839ae26;
    ram_cell[   11881] = 32'h0;  // 32'h8b89fc22;
    ram_cell[   11882] = 32'h0;  // 32'h91cb27ff;
    ram_cell[   11883] = 32'h0;  // 32'h3d2db861;
    ram_cell[   11884] = 32'h0;  // 32'h1117ca75;
    ram_cell[   11885] = 32'h0;  // 32'hbbeeab2a;
    ram_cell[   11886] = 32'h0;  // 32'hae91d647;
    ram_cell[   11887] = 32'h0;  // 32'h57f51ef5;
    ram_cell[   11888] = 32'h0;  // 32'h741be55a;
    ram_cell[   11889] = 32'h0;  // 32'h1d8529b6;
    ram_cell[   11890] = 32'h0;  // 32'hecf6563a;
    ram_cell[   11891] = 32'h0;  // 32'hba83cb32;
    ram_cell[   11892] = 32'h0;  // 32'he496843f;
    ram_cell[   11893] = 32'h0;  // 32'hbf8d614e;
    ram_cell[   11894] = 32'h0;  // 32'hf49cf6ce;
    ram_cell[   11895] = 32'h0;  // 32'h0ad3a6f4;
    ram_cell[   11896] = 32'h0;  // 32'hef5bd94d;
    ram_cell[   11897] = 32'h0;  // 32'he2001c86;
    ram_cell[   11898] = 32'h0;  // 32'hbd3e1929;
    ram_cell[   11899] = 32'h0;  // 32'hff645747;
    ram_cell[   11900] = 32'h0;  // 32'h127bf14c;
    ram_cell[   11901] = 32'h0;  // 32'hb4ed9148;
    ram_cell[   11902] = 32'h0;  // 32'haef8e64e;
    ram_cell[   11903] = 32'h0;  // 32'h5c32e166;
    ram_cell[   11904] = 32'h0;  // 32'hac9ada6c;
    ram_cell[   11905] = 32'h0;  // 32'h61c348af;
    ram_cell[   11906] = 32'h0;  // 32'h623af3bf;
    ram_cell[   11907] = 32'h0;  // 32'ha16c4283;
    ram_cell[   11908] = 32'h0;  // 32'h3a849eb6;
    ram_cell[   11909] = 32'h0;  // 32'h6c1dd749;
    ram_cell[   11910] = 32'h0;  // 32'hed1b3fe7;
    ram_cell[   11911] = 32'h0;  // 32'h61bc7e85;
    ram_cell[   11912] = 32'h0;  // 32'h828e2f23;
    ram_cell[   11913] = 32'h0;  // 32'h06db1031;
    ram_cell[   11914] = 32'h0;  // 32'h45986117;
    ram_cell[   11915] = 32'h0;  // 32'h470576d8;
    ram_cell[   11916] = 32'h0;  // 32'hf551f62f;
    ram_cell[   11917] = 32'h0;  // 32'hc3997683;
    ram_cell[   11918] = 32'h0;  // 32'h25570bc7;
    ram_cell[   11919] = 32'h0;  // 32'h629c5e1b;
    ram_cell[   11920] = 32'h0;  // 32'hbcf0c4b7;
    ram_cell[   11921] = 32'h0;  // 32'hd92c6865;
    ram_cell[   11922] = 32'h0;  // 32'h7518aad4;
    ram_cell[   11923] = 32'h0;  // 32'h8a0091c7;
    ram_cell[   11924] = 32'h0;  // 32'h1f6090ca;
    ram_cell[   11925] = 32'h0;  // 32'he92b28f3;
    ram_cell[   11926] = 32'h0;  // 32'h25354335;
    ram_cell[   11927] = 32'h0;  // 32'h542a94c7;
    ram_cell[   11928] = 32'h0;  // 32'h31053af0;
    ram_cell[   11929] = 32'h0;  // 32'h62fe7906;
    ram_cell[   11930] = 32'h0;  // 32'h064cb7c1;
    ram_cell[   11931] = 32'h0;  // 32'h8b9cbf3f;
    ram_cell[   11932] = 32'h0;  // 32'h657c9980;
    ram_cell[   11933] = 32'h0;  // 32'hbd1d761b;
    ram_cell[   11934] = 32'h0;  // 32'hb7432569;
    ram_cell[   11935] = 32'h0;  // 32'hfacf83b1;
    ram_cell[   11936] = 32'h0;  // 32'h48347b9c;
    ram_cell[   11937] = 32'h0;  // 32'h7f31304e;
    ram_cell[   11938] = 32'h0;  // 32'h506b5b8f;
    ram_cell[   11939] = 32'h0;  // 32'h65b5e4dc;
    ram_cell[   11940] = 32'h0;  // 32'h8151f8b5;
    ram_cell[   11941] = 32'h0;  // 32'hf9cd198b;
    ram_cell[   11942] = 32'h0;  // 32'h075b9019;
    ram_cell[   11943] = 32'h0;  // 32'ha7272221;
    ram_cell[   11944] = 32'h0;  // 32'h56e420e0;
    ram_cell[   11945] = 32'h0;  // 32'h6a9d27ba;
    ram_cell[   11946] = 32'h0;  // 32'h4842895f;
    ram_cell[   11947] = 32'h0;  // 32'h8dc9e6c4;
    ram_cell[   11948] = 32'h0;  // 32'hca15b478;
    ram_cell[   11949] = 32'h0;  // 32'hde6ab190;
    ram_cell[   11950] = 32'h0;  // 32'hecedf5ba;
    ram_cell[   11951] = 32'h0;  // 32'ha811da39;
    ram_cell[   11952] = 32'h0;  // 32'h425da3f8;
    ram_cell[   11953] = 32'h0;  // 32'hf7925ae9;
    ram_cell[   11954] = 32'h0;  // 32'hc8743c8a;
    ram_cell[   11955] = 32'h0;  // 32'h09f0d49e;
    ram_cell[   11956] = 32'h0;  // 32'h2ea8c710;
    ram_cell[   11957] = 32'h0;  // 32'h09549d8d;
    ram_cell[   11958] = 32'h0;  // 32'hb7aeeca3;
    ram_cell[   11959] = 32'h0;  // 32'h34e13d87;
    ram_cell[   11960] = 32'h0;  // 32'hb18f1363;
    ram_cell[   11961] = 32'h0;  // 32'h6a568b39;
    ram_cell[   11962] = 32'h0;  // 32'h4edc7eaa;
    ram_cell[   11963] = 32'h0;  // 32'h219e3b56;
    ram_cell[   11964] = 32'h0;  // 32'hf96cbf42;
    ram_cell[   11965] = 32'h0;  // 32'h42f14287;
    ram_cell[   11966] = 32'h0;  // 32'ha362b8c4;
    ram_cell[   11967] = 32'h0;  // 32'h73ddee19;
    ram_cell[   11968] = 32'h0;  // 32'hf223e08a;
    ram_cell[   11969] = 32'h0;  // 32'ha74fed08;
    ram_cell[   11970] = 32'h0;  // 32'hfe83b27c;
    ram_cell[   11971] = 32'h0;  // 32'hdb284a8b;
    ram_cell[   11972] = 32'h0;  // 32'hcc848085;
    ram_cell[   11973] = 32'h0;  // 32'hf7115a1a;
    ram_cell[   11974] = 32'h0;  // 32'hff99aa21;
    ram_cell[   11975] = 32'h0;  // 32'h82b8ad98;
    ram_cell[   11976] = 32'h0;  // 32'he8044420;
    ram_cell[   11977] = 32'h0;  // 32'h8bdf01ae;
    ram_cell[   11978] = 32'h0;  // 32'he67f06c9;
    ram_cell[   11979] = 32'h0;  // 32'hb0ce5b25;
    ram_cell[   11980] = 32'h0;  // 32'ha0958677;
    ram_cell[   11981] = 32'h0;  // 32'hf315c7d6;
    ram_cell[   11982] = 32'h0;  // 32'h88ccf833;
    ram_cell[   11983] = 32'h0;  // 32'h49bc987c;
    ram_cell[   11984] = 32'h0;  // 32'h5b400849;
    ram_cell[   11985] = 32'h0;  // 32'hc6edded8;
    ram_cell[   11986] = 32'h0;  // 32'hbf111131;
    ram_cell[   11987] = 32'h0;  // 32'ha0cf503f;
    ram_cell[   11988] = 32'h0;  // 32'h33a00ef0;
    ram_cell[   11989] = 32'h0;  // 32'hb964b267;
    ram_cell[   11990] = 32'h0;  // 32'h69f6883e;
    ram_cell[   11991] = 32'h0;  // 32'hd1c082cb;
    ram_cell[   11992] = 32'h0;  // 32'h8f5b90c3;
    ram_cell[   11993] = 32'h0;  // 32'h113f4139;
    ram_cell[   11994] = 32'h0;  // 32'h29482d36;
    ram_cell[   11995] = 32'h0;  // 32'h9f9dc64e;
    ram_cell[   11996] = 32'h0;  // 32'h259e720f;
    ram_cell[   11997] = 32'h0;  // 32'hed8043cc;
    ram_cell[   11998] = 32'h0;  // 32'h61cf5976;
    ram_cell[   11999] = 32'h0;  // 32'h37b79809;
    ram_cell[   12000] = 32'h0;  // 32'hf31d03ac;
    ram_cell[   12001] = 32'h0;  // 32'h2920a372;
    ram_cell[   12002] = 32'h0;  // 32'hbd8a91be;
    ram_cell[   12003] = 32'h0;  // 32'h8071e6b7;
    ram_cell[   12004] = 32'h0;  // 32'hf0ac190b;
    ram_cell[   12005] = 32'h0;  // 32'h2556a2e7;
    ram_cell[   12006] = 32'h0;  // 32'h9dced300;
    ram_cell[   12007] = 32'h0;  // 32'hcc96d19e;
    ram_cell[   12008] = 32'h0;  // 32'hf659a0df;
    ram_cell[   12009] = 32'h0;  // 32'ha140a773;
    ram_cell[   12010] = 32'h0;  // 32'hc564c22d;
    ram_cell[   12011] = 32'h0;  // 32'h68e231c4;
    ram_cell[   12012] = 32'h0;  // 32'ha1cae321;
    ram_cell[   12013] = 32'h0;  // 32'h1a1f6a17;
    ram_cell[   12014] = 32'h0;  // 32'hbd4c41aa;
    ram_cell[   12015] = 32'h0;  // 32'h39c99f84;
    ram_cell[   12016] = 32'h0;  // 32'hec589548;
    ram_cell[   12017] = 32'h0;  // 32'hef88b61e;
    ram_cell[   12018] = 32'h0;  // 32'h87ecb4fc;
    ram_cell[   12019] = 32'h0;  // 32'had192028;
    ram_cell[   12020] = 32'h0;  // 32'hd32cac72;
    ram_cell[   12021] = 32'h0;  // 32'h95f003ef;
    ram_cell[   12022] = 32'h0;  // 32'h8d2580b6;
    ram_cell[   12023] = 32'h0;  // 32'h58ae3350;
    ram_cell[   12024] = 32'h0;  // 32'h6fbec5c0;
    ram_cell[   12025] = 32'h0;  // 32'heb47315d;
    ram_cell[   12026] = 32'h0;  // 32'hf01f85ca;
    ram_cell[   12027] = 32'h0;  // 32'hc3d47ad6;
    ram_cell[   12028] = 32'h0;  // 32'h9536f35d;
    ram_cell[   12029] = 32'h0;  // 32'h7817dc69;
    ram_cell[   12030] = 32'h0;  // 32'h020167b2;
    ram_cell[   12031] = 32'h0;  // 32'ha2b63a63;
    ram_cell[   12032] = 32'h0;  // 32'h3c81d534;
    ram_cell[   12033] = 32'h0;  // 32'hc99a0969;
    ram_cell[   12034] = 32'h0;  // 32'hf4606c18;
    ram_cell[   12035] = 32'h0;  // 32'h4f5d817e;
    ram_cell[   12036] = 32'h0;  // 32'hda54f5d5;
    ram_cell[   12037] = 32'h0;  // 32'haa5216bb;
    ram_cell[   12038] = 32'h0;  // 32'h0caf9719;
    ram_cell[   12039] = 32'h0;  // 32'h447a6d82;
    ram_cell[   12040] = 32'h0;  // 32'h693bd505;
    ram_cell[   12041] = 32'h0;  // 32'haace9976;
    ram_cell[   12042] = 32'h0;  // 32'h3e440fca;
    ram_cell[   12043] = 32'h0;  // 32'h11f1b88d;
    ram_cell[   12044] = 32'h0;  // 32'he5b906a9;
    ram_cell[   12045] = 32'h0;  // 32'hf82bf9ef;
    ram_cell[   12046] = 32'h0;  // 32'h27b1fa34;
    ram_cell[   12047] = 32'h0;  // 32'h7976d7aa;
    ram_cell[   12048] = 32'h0;  // 32'h53a2dcdb;
    ram_cell[   12049] = 32'h0;  // 32'he36c8738;
    ram_cell[   12050] = 32'h0;  // 32'he2be50c8;
    ram_cell[   12051] = 32'h0;  // 32'h577238a4;
    ram_cell[   12052] = 32'h0;  // 32'h6a7a425d;
    ram_cell[   12053] = 32'h0;  // 32'hf312a87a;
    ram_cell[   12054] = 32'h0;  // 32'h281fb26f;
    ram_cell[   12055] = 32'h0;  // 32'h7c14c2d6;
    ram_cell[   12056] = 32'h0;  // 32'h8c8f4418;
    ram_cell[   12057] = 32'h0;  // 32'hf4cd9c41;
    ram_cell[   12058] = 32'h0;  // 32'h0e80ae10;
    ram_cell[   12059] = 32'h0;  // 32'h42ae1061;
    ram_cell[   12060] = 32'h0;  // 32'h9a6c7f5a;
    ram_cell[   12061] = 32'h0;  // 32'h16241345;
    ram_cell[   12062] = 32'h0;  // 32'h1ef92a9b;
    ram_cell[   12063] = 32'h0;  // 32'h60b7af13;
    ram_cell[   12064] = 32'h0;  // 32'h50527bd6;
    ram_cell[   12065] = 32'h0;  // 32'h9a6e5b69;
    ram_cell[   12066] = 32'h0;  // 32'hfc192fd0;
    ram_cell[   12067] = 32'h0;  // 32'h89ba744d;
    ram_cell[   12068] = 32'h0;  // 32'h60e83fc0;
    ram_cell[   12069] = 32'h0;  // 32'h7145daaa;
    ram_cell[   12070] = 32'h0;  // 32'h847be43b;
    ram_cell[   12071] = 32'h0;  // 32'h7bcc56d5;
    ram_cell[   12072] = 32'h0;  // 32'h56e9da9c;
    ram_cell[   12073] = 32'h0;  // 32'h4375a918;
    ram_cell[   12074] = 32'h0;  // 32'h0d64ef76;
    ram_cell[   12075] = 32'h0;  // 32'hd01b6b93;
    ram_cell[   12076] = 32'h0;  // 32'ha3b0bc37;
    ram_cell[   12077] = 32'h0;  // 32'h5b8a64f8;
    ram_cell[   12078] = 32'h0;  // 32'h3f80a654;
    ram_cell[   12079] = 32'h0;  // 32'h1f75d84e;
    ram_cell[   12080] = 32'h0;  // 32'hcef6a791;
    ram_cell[   12081] = 32'h0;  // 32'hc7966582;
    ram_cell[   12082] = 32'h0;  // 32'h3b566905;
    ram_cell[   12083] = 32'h0;  // 32'hf203358b;
    ram_cell[   12084] = 32'h0;  // 32'h3e3e9e8b;
    ram_cell[   12085] = 32'h0;  // 32'hb98118db;
    ram_cell[   12086] = 32'h0;  // 32'h955ab9ef;
    ram_cell[   12087] = 32'h0;  // 32'h6aa86ce1;
    ram_cell[   12088] = 32'h0;  // 32'hf5e04d51;
    ram_cell[   12089] = 32'h0;  // 32'h316ea88e;
    ram_cell[   12090] = 32'h0;  // 32'h7507c8e8;
    ram_cell[   12091] = 32'h0;  // 32'hc9c5ff2c;
    ram_cell[   12092] = 32'h0;  // 32'h74e335a6;
    ram_cell[   12093] = 32'h0;  // 32'hc23580ef;
    ram_cell[   12094] = 32'h0;  // 32'hbb6cad20;
    ram_cell[   12095] = 32'h0;  // 32'h006ee623;
    ram_cell[   12096] = 32'h0;  // 32'h0918b10e;
    ram_cell[   12097] = 32'h0;  // 32'hb1472f60;
    ram_cell[   12098] = 32'h0;  // 32'h64cce9bf;
    ram_cell[   12099] = 32'h0;  // 32'hf8107bb7;
    ram_cell[   12100] = 32'h0;  // 32'h1f9d2760;
    ram_cell[   12101] = 32'h0;  // 32'h4cae98e0;
    ram_cell[   12102] = 32'h0;  // 32'h1f129b0f;
    ram_cell[   12103] = 32'h0;  // 32'hea6fadf3;
    ram_cell[   12104] = 32'h0;  // 32'h8056a108;
    ram_cell[   12105] = 32'h0;  // 32'h7ba29640;
    ram_cell[   12106] = 32'h0;  // 32'h0f67b833;
    ram_cell[   12107] = 32'h0;  // 32'hee760b59;
    ram_cell[   12108] = 32'h0;  // 32'h8fde92d9;
    ram_cell[   12109] = 32'h0;  // 32'hd5abd19d;
    ram_cell[   12110] = 32'h0;  // 32'hd1cedddd;
    ram_cell[   12111] = 32'h0;  // 32'h68ef8cf0;
    ram_cell[   12112] = 32'h0;  // 32'haa62e831;
    ram_cell[   12113] = 32'h0;  // 32'h44f619b0;
    ram_cell[   12114] = 32'h0;  // 32'hb4facc8a;
    ram_cell[   12115] = 32'h0;  // 32'hfc50f3f1;
    ram_cell[   12116] = 32'h0;  // 32'h0fd29b05;
    ram_cell[   12117] = 32'h0;  // 32'h2ad6410a;
    ram_cell[   12118] = 32'h0;  // 32'hdbedfad0;
    ram_cell[   12119] = 32'h0;  // 32'hdc468890;
    ram_cell[   12120] = 32'h0;  // 32'h086154c9;
    ram_cell[   12121] = 32'h0;  // 32'h22d8cce8;
    ram_cell[   12122] = 32'h0;  // 32'hd1badc78;
    ram_cell[   12123] = 32'h0;  // 32'h922e17de;
    ram_cell[   12124] = 32'h0;  // 32'hfcf5eff5;
    ram_cell[   12125] = 32'h0;  // 32'hc2667268;
    ram_cell[   12126] = 32'h0;  // 32'hbef34d85;
    ram_cell[   12127] = 32'h0;  // 32'hca04cbbb;
    ram_cell[   12128] = 32'h0;  // 32'hac2c18e1;
    ram_cell[   12129] = 32'h0;  // 32'h50171817;
    ram_cell[   12130] = 32'h0;  // 32'hf5bab7b0;
    ram_cell[   12131] = 32'h0;  // 32'h6e78f854;
    ram_cell[   12132] = 32'h0;  // 32'h0c9ae2f7;
    ram_cell[   12133] = 32'h0;  // 32'h9bab8738;
    ram_cell[   12134] = 32'h0;  // 32'h5352e783;
    ram_cell[   12135] = 32'h0;  // 32'h82216774;
    ram_cell[   12136] = 32'h0;  // 32'h6854e0bd;
    ram_cell[   12137] = 32'h0;  // 32'hb20f485a;
    ram_cell[   12138] = 32'h0;  // 32'h3fc2dcc8;
    ram_cell[   12139] = 32'h0;  // 32'h6db97b47;
    ram_cell[   12140] = 32'h0;  // 32'hf38aba63;
    ram_cell[   12141] = 32'h0;  // 32'he82ad0aa;
    ram_cell[   12142] = 32'h0;  // 32'h5fcee872;
    ram_cell[   12143] = 32'h0;  // 32'h7ce4996b;
    ram_cell[   12144] = 32'h0;  // 32'hf837f277;
    ram_cell[   12145] = 32'h0;  // 32'h212d3d3d;
    ram_cell[   12146] = 32'h0;  // 32'h22d18204;
    ram_cell[   12147] = 32'h0;  // 32'h31689d72;
    ram_cell[   12148] = 32'h0;  // 32'h1ede370d;
    ram_cell[   12149] = 32'h0;  // 32'h32d10db1;
    ram_cell[   12150] = 32'h0;  // 32'hbbdc5cf7;
    ram_cell[   12151] = 32'h0;  // 32'h376db554;
    ram_cell[   12152] = 32'h0;  // 32'hd16f1879;
    ram_cell[   12153] = 32'h0;  // 32'h1fff2dfa;
    ram_cell[   12154] = 32'h0;  // 32'h1bd1624e;
    ram_cell[   12155] = 32'h0;  // 32'h5c19f599;
    ram_cell[   12156] = 32'h0;  // 32'h7568b0a0;
    ram_cell[   12157] = 32'h0;  // 32'h49a4d977;
    ram_cell[   12158] = 32'h0;  // 32'h0d033a94;
    ram_cell[   12159] = 32'h0;  // 32'h18da1b50;
    ram_cell[   12160] = 32'h0;  // 32'h4d0cb27a;
    ram_cell[   12161] = 32'h0;  // 32'h9236a3d1;
    ram_cell[   12162] = 32'h0;  // 32'haf221922;
    ram_cell[   12163] = 32'h0;  // 32'hd0f7f8f8;
    ram_cell[   12164] = 32'h0;  // 32'haa1c6c74;
    ram_cell[   12165] = 32'h0;  // 32'hf76871a9;
    ram_cell[   12166] = 32'h0;  // 32'ha7a0f54d;
    ram_cell[   12167] = 32'h0;  // 32'h38c2ce22;
    ram_cell[   12168] = 32'h0;  // 32'hf4646c93;
    ram_cell[   12169] = 32'h0;  // 32'hd6a0fc18;
    ram_cell[   12170] = 32'h0;  // 32'hd52e7db4;
    ram_cell[   12171] = 32'h0;  // 32'hd0419aaf;
    ram_cell[   12172] = 32'h0;  // 32'h460e8c46;
    ram_cell[   12173] = 32'h0;  // 32'h5dc32d9f;
    ram_cell[   12174] = 32'h0;  // 32'h6536a891;
    ram_cell[   12175] = 32'h0;  // 32'h7bf06ca3;
    ram_cell[   12176] = 32'h0;  // 32'h0ae01697;
    ram_cell[   12177] = 32'h0;  // 32'he3bb9922;
    ram_cell[   12178] = 32'h0;  // 32'he8976e03;
    ram_cell[   12179] = 32'h0;  // 32'h746d6c9f;
    ram_cell[   12180] = 32'h0;  // 32'h9d55a64c;
    ram_cell[   12181] = 32'h0;  // 32'h1fd3dad7;
    ram_cell[   12182] = 32'h0;  // 32'h50a08634;
    ram_cell[   12183] = 32'h0;  // 32'h97845224;
    ram_cell[   12184] = 32'h0;  // 32'hac04e709;
    ram_cell[   12185] = 32'h0;  // 32'h4295f74d;
    ram_cell[   12186] = 32'h0;  // 32'hfe9dfde8;
    ram_cell[   12187] = 32'h0;  // 32'h573fb125;
    ram_cell[   12188] = 32'h0;  // 32'hcd5d101e;
    ram_cell[   12189] = 32'h0;  // 32'h1b97f3d4;
    ram_cell[   12190] = 32'h0;  // 32'h781a4d19;
    ram_cell[   12191] = 32'h0;  // 32'h14deaa49;
    ram_cell[   12192] = 32'h0;  // 32'h635e5121;
    ram_cell[   12193] = 32'h0;  // 32'h7a85bda8;
    ram_cell[   12194] = 32'h0;  // 32'h0b297a5f;
    ram_cell[   12195] = 32'h0;  // 32'hf96dfc2f;
    ram_cell[   12196] = 32'h0;  // 32'ha15ddd9e;
    ram_cell[   12197] = 32'h0;  // 32'hae620f92;
    ram_cell[   12198] = 32'h0;  // 32'h83342ead;
    ram_cell[   12199] = 32'h0;  // 32'hbabda127;
    ram_cell[   12200] = 32'h0;  // 32'h0ed412cc;
    ram_cell[   12201] = 32'h0;  // 32'h6dca72fc;
    ram_cell[   12202] = 32'h0;  // 32'h19cc07b8;
    ram_cell[   12203] = 32'h0;  // 32'ha02ba2b9;
    ram_cell[   12204] = 32'h0;  // 32'h4f6a8177;
    ram_cell[   12205] = 32'h0;  // 32'h8201318d;
    ram_cell[   12206] = 32'h0;  // 32'h1e205821;
    ram_cell[   12207] = 32'h0;  // 32'h1dd7b67f;
    ram_cell[   12208] = 32'h0;  // 32'hdf831772;
    ram_cell[   12209] = 32'h0;  // 32'he4df8fc1;
    ram_cell[   12210] = 32'h0;  // 32'h76cab64e;
    ram_cell[   12211] = 32'h0;  // 32'hc6f7a1fe;
    ram_cell[   12212] = 32'h0;  // 32'hf7642938;
    ram_cell[   12213] = 32'h0;  // 32'h10688442;
    ram_cell[   12214] = 32'h0;  // 32'h1566c42d;
    ram_cell[   12215] = 32'h0;  // 32'h9d8b9eec;
    ram_cell[   12216] = 32'h0;  // 32'h89c51836;
    ram_cell[   12217] = 32'h0;  // 32'hc5520a78;
    ram_cell[   12218] = 32'h0;  // 32'h5141af46;
    ram_cell[   12219] = 32'h0;  // 32'h51342cfb;
    ram_cell[   12220] = 32'h0;  // 32'hfef8bd0c;
    ram_cell[   12221] = 32'h0;  // 32'hb565027d;
    ram_cell[   12222] = 32'h0;  // 32'h35a2bafb;
    ram_cell[   12223] = 32'h0;  // 32'hd9427856;
    ram_cell[   12224] = 32'h0;  // 32'hcba49ff7;
    ram_cell[   12225] = 32'h0;  // 32'hfc745019;
    ram_cell[   12226] = 32'h0;  // 32'h72a3c821;
    ram_cell[   12227] = 32'h0;  // 32'h3792c4fd;
    ram_cell[   12228] = 32'h0;  // 32'he5905afa;
    ram_cell[   12229] = 32'h0;  // 32'hb2fe6d71;
    ram_cell[   12230] = 32'h0;  // 32'hff60d728;
    ram_cell[   12231] = 32'h0;  // 32'he86112bd;
    ram_cell[   12232] = 32'h0;  // 32'ha5e0307a;
    ram_cell[   12233] = 32'h0;  // 32'h50831bd0;
    ram_cell[   12234] = 32'h0;  // 32'hbe4c9035;
    ram_cell[   12235] = 32'h0;  // 32'hf8b6367b;
    ram_cell[   12236] = 32'h0;  // 32'h277f2f0c;
    ram_cell[   12237] = 32'h0;  // 32'h3d7b866f;
    ram_cell[   12238] = 32'h0;  // 32'h9fe46648;
    ram_cell[   12239] = 32'h0;  // 32'hb00cf113;
    ram_cell[   12240] = 32'h0;  // 32'h926f4fde;
    ram_cell[   12241] = 32'h0;  // 32'h6ea6ee42;
    ram_cell[   12242] = 32'h0;  // 32'h2d8918cc;
    ram_cell[   12243] = 32'h0;  // 32'h591269d0;
    ram_cell[   12244] = 32'h0;  // 32'hac8dc1f9;
    ram_cell[   12245] = 32'h0;  // 32'hf73589e7;
    ram_cell[   12246] = 32'h0;  // 32'ha31d5921;
    ram_cell[   12247] = 32'h0;  // 32'h4781741e;
    ram_cell[   12248] = 32'h0;  // 32'hadddb74b;
    ram_cell[   12249] = 32'h0;  // 32'h1ce4463e;
    ram_cell[   12250] = 32'h0;  // 32'hf6737760;
    ram_cell[   12251] = 32'h0;  // 32'h4622eb39;
    ram_cell[   12252] = 32'h0;  // 32'h2785191d;
    ram_cell[   12253] = 32'h0;  // 32'h1c4fbe85;
    ram_cell[   12254] = 32'h0;  // 32'hce768e33;
    ram_cell[   12255] = 32'h0;  // 32'hfbe37f88;
    ram_cell[   12256] = 32'h0;  // 32'h467f4a39;
    ram_cell[   12257] = 32'h0;  // 32'h267cda6b;
    ram_cell[   12258] = 32'h0;  // 32'h0db44fd3;
    ram_cell[   12259] = 32'h0;  // 32'h9128a236;
    ram_cell[   12260] = 32'h0;  // 32'h28b674f2;
    ram_cell[   12261] = 32'h0;  // 32'h3b6db736;
    ram_cell[   12262] = 32'h0;  // 32'h1928476c;
    ram_cell[   12263] = 32'h0;  // 32'hdaa99d2f;
    ram_cell[   12264] = 32'h0;  // 32'h1f58c194;
    ram_cell[   12265] = 32'h0;  // 32'h6df0eca2;
    ram_cell[   12266] = 32'h0;  // 32'ha688119b;
    ram_cell[   12267] = 32'h0;  // 32'hfaee4763;
    ram_cell[   12268] = 32'h0;  // 32'h055bb2e9;
    ram_cell[   12269] = 32'h0;  // 32'hd55b21b5;
    ram_cell[   12270] = 32'h0;  // 32'h23ee8813;
    ram_cell[   12271] = 32'h0;  // 32'h5280b948;
    ram_cell[   12272] = 32'h0;  // 32'h683e8b72;
    ram_cell[   12273] = 32'h0;  // 32'h524999d8;
    ram_cell[   12274] = 32'h0;  // 32'ha5360314;
    ram_cell[   12275] = 32'h0;  // 32'h19de2e9f;
    ram_cell[   12276] = 32'h0;  // 32'hf241d5c1;
    ram_cell[   12277] = 32'h0;  // 32'hbe19af3b;
    ram_cell[   12278] = 32'h0;  // 32'hbd45cc05;
    ram_cell[   12279] = 32'h0;  // 32'hcf2a2df8;
    ram_cell[   12280] = 32'h0;  // 32'hb5f397c8;
    ram_cell[   12281] = 32'h0;  // 32'h71e20881;
    ram_cell[   12282] = 32'h0;  // 32'haa69f713;
    ram_cell[   12283] = 32'h0;  // 32'h6aca7767;
    ram_cell[   12284] = 32'h0;  // 32'hc12fc7bf;
    ram_cell[   12285] = 32'h0;  // 32'h70107888;
    ram_cell[   12286] = 32'h0;  // 32'hc312dcc3;
    ram_cell[   12287] = 32'h0;  // 32'hbd708e31;
    ram_cell[   12288] = 32'h0;  // 32'h92a3411e;
    ram_cell[   12289] = 32'h0;  // 32'h605c6b50;
    ram_cell[   12290] = 32'h0;  // 32'h2c82ff83;
    ram_cell[   12291] = 32'h0;  // 32'hbae1552c;
    ram_cell[   12292] = 32'h0;  // 32'hfc981fd1;
    ram_cell[   12293] = 32'h0;  // 32'h30df4ccf;
    ram_cell[   12294] = 32'h0;  // 32'h74e51a43;
    ram_cell[   12295] = 32'h0;  // 32'hafa1e36e;
    ram_cell[   12296] = 32'h0;  // 32'h7f12cce2;
    ram_cell[   12297] = 32'h0;  // 32'h2a152dbf;
    ram_cell[   12298] = 32'h0;  // 32'heff7a5bf;
    ram_cell[   12299] = 32'h0;  // 32'h5b33f617;
    ram_cell[   12300] = 32'h0;  // 32'hafc8c0b4;
    ram_cell[   12301] = 32'h0;  // 32'h2dbbfe01;
    ram_cell[   12302] = 32'h0;  // 32'he2e6f160;
    ram_cell[   12303] = 32'h0;  // 32'hb54c98a1;
    ram_cell[   12304] = 32'h0;  // 32'h69a730da;
    ram_cell[   12305] = 32'h0;  // 32'h5e02b538;
    ram_cell[   12306] = 32'h0;  // 32'h7c977f6a;
    ram_cell[   12307] = 32'h0;  // 32'hc490b07e;
    ram_cell[   12308] = 32'h0;  // 32'habc386be;
    ram_cell[   12309] = 32'h0;  // 32'hd221c99d;
    ram_cell[   12310] = 32'h0;  // 32'hc0c7b812;
    ram_cell[   12311] = 32'h0;  // 32'h0d79cf85;
    ram_cell[   12312] = 32'h0;  // 32'h4f59ee2b;
    ram_cell[   12313] = 32'h0;  // 32'hbe7d546c;
    ram_cell[   12314] = 32'h0;  // 32'hf0b3cbf7;
    ram_cell[   12315] = 32'h0;  // 32'h76df74af;
    ram_cell[   12316] = 32'h0;  // 32'h36b77d63;
    ram_cell[   12317] = 32'h0;  // 32'h9d6b7b98;
    ram_cell[   12318] = 32'h0;  // 32'habf43ab7;
    ram_cell[   12319] = 32'h0;  // 32'hc350e06b;
    ram_cell[   12320] = 32'h0;  // 32'hd2851f3b;
    ram_cell[   12321] = 32'h0;  // 32'hff0bf4a8;
    ram_cell[   12322] = 32'h0;  // 32'h5ab4efcd;
    ram_cell[   12323] = 32'h0;  // 32'h59162d1a;
    ram_cell[   12324] = 32'h0;  // 32'h0bdd1d9f;
    ram_cell[   12325] = 32'h0;  // 32'hfd799a1f;
    ram_cell[   12326] = 32'h0;  // 32'hd1971df6;
    ram_cell[   12327] = 32'h0;  // 32'h0f07fb85;
    ram_cell[   12328] = 32'h0;  // 32'hd0c30f5f;
    ram_cell[   12329] = 32'h0;  // 32'h5dc977ef;
    ram_cell[   12330] = 32'h0;  // 32'h3b216fa0;
    ram_cell[   12331] = 32'h0;  // 32'hbd2c0415;
    ram_cell[   12332] = 32'h0;  // 32'h4c152312;
    ram_cell[   12333] = 32'h0;  // 32'hd7115b91;
    ram_cell[   12334] = 32'h0;  // 32'hb38fcc36;
    ram_cell[   12335] = 32'h0;  // 32'he973dab5;
    ram_cell[   12336] = 32'h0;  // 32'h1c112f12;
    ram_cell[   12337] = 32'h0;  // 32'hdea5a85d;
    ram_cell[   12338] = 32'h0;  // 32'h6fb6d882;
    ram_cell[   12339] = 32'h0;  // 32'h130ed43e;
    ram_cell[   12340] = 32'h0;  // 32'h90328ba2;
    ram_cell[   12341] = 32'h0;  // 32'h34110614;
    ram_cell[   12342] = 32'h0;  // 32'h060fcca4;
    ram_cell[   12343] = 32'h0;  // 32'hea59aa0b;
    ram_cell[   12344] = 32'h0;  // 32'h20ab8f91;
    ram_cell[   12345] = 32'h0;  // 32'h067a81fe;
    ram_cell[   12346] = 32'h0;  // 32'h2313193d;
    ram_cell[   12347] = 32'h0;  // 32'h1789052b;
    ram_cell[   12348] = 32'h0;  // 32'he137b071;
    ram_cell[   12349] = 32'h0;  // 32'hcfb6a32c;
    ram_cell[   12350] = 32'h0;  // 32'h0a748963;
    ram_cell[   12351] = 32'h0;  // 32'h36b9cf4a;
    ram_cell[   12352] = 32'h0;  // 32'h6b4cdc47;
    ram_cell[   12353] = 32'h0;  // 32'hee642040;
    ram_cell[   12354] = 32'h0;  // 32'h8bee3d2f;
    ram_cell[   12355] = 32'h0;  // 32'hd5a01738;
    ram_cell[   12356] = 32'h0;  // 32'h7b74238d;
    ram_cell[   12357] = 32'h0;  // 32'h12bac260;
    ram_cell[   12358] = 32'h0;  // 32'h348c2723;
    ram_cell[   12359] = 32'h0;  // 32'hcda30c4a;
    ram_cell[   12360] = 32'h0;  // 32'h0aa86925;
    ram_cell[   12361] = 32'h0;  // 32'h5e85eb5c;
    ram_cell[   12362] = 32'h0;  // 32'ha4dc1bfa;
    ram_cell[   12363] = 32'h0;  // 32'h54181883;
    ram_cell[   12364] = 32'h0;  // 32'h894e8693;
    ram_cell[   12365] = 32'h0;  // 32'hac3c5994;
    ram_cell[   12366] = 32'h0;  // 32'h55314f59;
    ram_cell[   12367] = 32'h0;  // 32'h42b4e7da;
    ram_cell[   12368] = 32'h0;  // 32'hbc9cc43a;
    ram_cell[   12369] = 32'h0;  // 32'hd8a185ae;
    ram_cell[   12370] = 32'h0;  // 32'ha47ea940;
    ram_cell[   12371] = 32'h0;  // 32'hef46f8e1;
    ram_cell[   12372] = 32'h0;  // 32'he54873e8;
    ram_cell[   12373] = 32'h0;  // 32'hc99fcbf2;
    ram_cell[   12374] = 32'h0;  // 32'h130ba2d4;
    ram_cell[   12375] = 32'h0;  // 32'h93d7242e;
    ram_cell[   12376] = 32'h0;  // 32'h539f5ab5;
    ram_cell[   12377] = 32'h0;  // 32'ha2093588;
    ram_cell[   12378] = 32'h0;  // 32'h71b78171;
    ram_cell[   12379] = 32'h0;  // 32'hfc6ac08d;
    ram_cell[   12380] = 32'h0;  // 32'h21004f3d;
    ram_cell[   12381] = 32'h0;  // 32'ha0764843;
    ram_cell[   12382] = 32'h0;  // 32'ha9047405;
    ram_cell[   12383] = 32'h0;  // 32'h4190b040;
    ram_cell[   12384] = 32'h0;  // 32'habaa7d6c;
    ram_cell[   12385] = 32'h0;  // 32'h6d225a46;
    ram_cell[   12386] = 32'h0;  // 32'hf809ac20;
    ram_cell[   12387] = 32'h0;  // 32'h7ba167c9;
    ram_cell[   12388] = 32'h0;  // 32'h30ea30ae;
    ram_cell[   12389] = 32'h0;  // 32'h9bfb4167;
    ram_cell[   12390] = 32'h0;  // 32'head5767e;
    ram_cell[   12391] = 32'h0;  // 32'h50354334;
    ram_cell[   12392] = 32'h0;  // 32'h23289901;
    ram_cell[   12393] = 32'h0;  // 32'h2fbe8278;
    ram_cell[   12394] = 32'h0;  // 32'h82bf0a99;
    ram_cell[   12395] = 32'h0;  // 32'hf073d36b;
    ram_cell[   12396] = 32'h0;  // 32'h8d6ca631;
    ram_cell[   12397] = 32'h0;  // 32'h8074d7b2;
    ram_cell[   12398] = 32'h0;  // 32'h82a4ea5d;
    ram_cell[   12399] = 32'h0;  // 32'h4987ef8f;
    ram_cell[   12400] = 32'h0;  // 32'h638692c8;
    ram_cell[   12401] = 32'h0;  // 32'h2b40faee;
    ram_cell[   12402] = 32'h0;  // 32'hf9a1904a;
    ram_cell[   12403] = 32'h0;  // 32'h8077a2c7;
    ram_cell[   12404] = 32'h0;  // 32'h8a38caa6;
    ram_cell[   12405] = 32'h0;  // 32'hebb35141;
    ram_cell[   12406] = 32'h0;  // 32'h91ebe61c;
    ram_cell[   12407] = 32'h0;  // 32'ha135cb83;
    ram_cell[   12408] = 32'h0;  // 32'h260e24fe;
    ram_cell[   12409] = 32'h0;  // 32'h3dc234e4;
    ram_cell[   12410] = 32'h0;  // 32'hc0b9b82f;
    ram_cell[   12411] = 32'h0;  // 32'h053090f9;
    ram_cell[   12412] = 32'h0;  // 32'h2c681852;
    ram_cell[   12413] = 32'h0;  // 32'h4265d390;
    ram_cell[   12414] = 32'h0;  // 32'h57eecdf9;
    ram_cell[   12415] = 32'h0;  // 32'hc7f57d12;
    ram_cell[   12416] = 32'h0;  // 32'hd99cfca3;
    ram_cell[   12417] = 32'h0;  // 32'h2ac2ef81;
    ram_cell[   12418] = 32'h0;  // 32'h2fceb7e5;
    ram_cell[   12419] = 32'h0;  // 32'hf9df7dd4;
    ram_cell[   12420] = 32'h0;  // 32'h14dff360;
    ram_cell[   12421] = 32'h0;  // 32'h99d4251e;
    ram_cell[   12422] = 32'h0;  // 32'h25cb077d;
    ram_cell[   12423] = 32'h0;  // 32'h177da204;
    ram_cell[   12424] = 32'h0;  // 32'hacf093a7;
    ram_cell[   12425] = 32'h0;  // 32'h9c56959a;
    ram_cell[   12426] = 32'h0;  // 32'h4c891cbb;
    ram_cell[   12427] = 32'h0;  // 32'h8e5f50d0;
    ram_cell[   12428] = 32'h0;  // 32'hf3af436e;
    ram_cell[   12429] = 32'h0;  // 32'hae47111f;
    ram_cell[   12430] = 32'h0;  // 32'hb481c97c;
    ram_cell[   12431] = 32'h0;  // 32'h4d8836d2;
    ram_cell[   12432] = 32'h0;  // 32'h25cbcf6f;
    ram_cell[   12433] = 32'h0;  // 32'h9bd34ab5;
    ram_cell[   12434] = 32'h0;  // 32'h1e6b37b2;
    ram_cell[   12435] = 32'h0;  // 32'h38421153;
    ram_cell[   12436] = 32'h0;  // 32'h45ef4e2f;
    ram_cell[   12437] = 32'h0;  // 32'hd2c01b08;
    ram_cell[   12438] = 32'h0;  // 32'hc331c079;
    ram_cell[   12439] = 32'h0;  // 32'h67eddf07;
    ram_cell[   12440] = 32'h0;  // 32'hd5a23a57;
    ram_cell[   12441] = 32'h0;  // 32'h71c9f8e6;
    ram_cell[   12442] = 32'h0;  // 32'h99b4687d;
    ram_cell[   12443] = 32'h0;  // 32'h8f634b9b;
    ram_cell[   12444] = 32'h0;  // 32'h4e4d1126;
    ram_cell[   12445] = 32'h0;  // 32'h005c5c5b;
    ram_cell[   12446] = 32'h0;  // 32'hbbfc65ad;
    ram_cell[   12447] = 32'h0;  // 32'h7aac6eac;
    ram_cell[   12448] = 32'h0;  // 32'h66e4d824;
    ram_cell[   12449] = 32'h0;  // 32'h436f0bad;
    ram_cell[   12450] = 32'h0;  // 32'hf5037c93;
    ram_cell[   12451] = 32'h0;  // 32'h4d545c16;
    ram_cell[   12452] = 32'h0;  // 32'hab31ce8d;
    ram_cell[   12453] = 32'h0;  // 32'h00e6de31;
    ram_cell[   12454] = 32'h0;  // 32'h00170e71;
    ram_cell[   12455] = 32'h0;  // 32'hca209929;
    ram_cell[   12456] = 32'h0;  // 32'ha52ae023;
    ram_cell[   12457] = 32'h0;  // 32'h64fe6fd0;
    ram_cell[   12458] = 32'h0;  // 32'h9c17396d;
    ram_cell[   12459] = 32'h0;  // 32'hb88751a1;
    ram_cell[   12460] = 32'h0;  // 32'he51f5949;
    ram_cell[   12461] = 32'h0;  // 32'hc99493f9;
    ram_cell[   12462] = 32'h0;  // 32'hc1ead743;
    ram_cell[   12463] = 32'h0;  // 32'h61a598e5;
    ram_cell[   12464] = 32'h0;  // 32'h51a72117;
    ram_cell[   12465] = 32'h0;  // 32'h5506b0f2;
    ram_cell[   12466] = 32'h0;  // 32'h46a48da3;
    ram_cell[   12467] = 32'h0;  // 32'h41074c6e;
    ram_cell[   12468] = 32'h0;  // 32'he468a605;
    ram_cell[   12469] = 32'h0;  // 32'h0b23903d;
    ram_cell[   12470] = 32'h0;  // 32'hc9ce6457;
    ram_cell[   12471] = 32'h0;  // 32'hd16203fc;
    ram_cell[   12472] = 32'h0;  // 32'h73e3a059;
    ram_cell[   12473] = 32'h0;  // 32'he12b43c5;
    ram_cell[   12474] = 32'h0;  // 32'h45d9a992;
    ram_cell[   12475] = 32'h0;  // 32'h04b084e2;
    ram_cell[   12476] = 32'h0;  // 32'h3b201bff;
    ram_cell[   12477] = 32'h0;  // 32'ha3da349e;
    ram_cell[   12478] = 32'h0;  // 32'h95aed7d8;
    ram_cell[   12479] = 32'h0;  // 32'hc9dd387a;
    ram_cell[   12480] = 32'h0;  // 32'hffa6ab53;
    ram_cell[   12481] = 32'h0;  // 32'hfc12311e;
    ram_cell[   12482] = 32'h0;  // 32'h10a8a843;
    ram_cell[   12483] = 32'h0;  // 32'h12152887;
    ram_cell[   12484] = 32'h0;  // 32'h445c5436;
    ram_cell[   12485] = 32'h0;  // 32'h3c8ac202;
    ram_cell[   12486] = 32'h0;  // 32'h00e546e8;
    ram_cell[   12487] = 32'h0;  // 32'h227fb562;
    ram_cell[   12488] = 32'h0;  // 32'h254cc4ac;
    ram_cell[   12489] = 32'h0;  // 32'h797799b4;
    ram_cell[   12490] = 32'h0;  // 32'hd9e5b482;
    ram_cell[   12491] = 32'h0;  // 32'hbddcec26;
    ram_cell[   12492] = 32'h0;  // 32'haea6056f;
    ram_cell[   12493] = 32'h0;  // 32'ha194b0ab;
    ram_cell[   12494] = 32'h0;  // 32'hc8ef01ff;
    ram_cell[   12495] = 32'h0;  // 32'hec4dabb1;
    ram_cell[   12496] = 32'h0;  // 32'h4586b2ce;
    ram_cell[   12497] = 32'h0;  // 32'ha359471f;
    ram_cell[   12498] = 32'h0;  // 32'hd9844a0f;
    ram_cell[   12499] = 32'h0;  // 32'h8451ed96;
    ram_cell[   12500] = 32'h0;  // 32'hfef3e2b1;
    ram_cell[   12501] = 32'h0;  // 32'hd5053627;
    ram_cell[   12502] = 32'h0;  // 32'h45b298f5;
    ram_cell[   12503] = 32'h0;  // 32'h0df468ae;
    ram_cell[   12504] = 32'h0;  // 32'hc0457c42;
    ram_cell[   12505] = 32'h0;  // 32'h8a70b37c;
    ram_cell[   12506] = 32'h0;  // 32'hbcba027b;
    ram_cell[   12507] = 32'h0;  // 32'h456e05f0;
    ram_cell[   12508] = 32'h0;  // 32'hc1586fd5;
    ram_cell[   12509] = 32'h0;  // 32'h4cab2459;
    ram_cell[   12510] = 32'h0;  // 32'h371f8d9f;
    ram_cell[   12511] = 32'h0;  // 32'hd01fb917;
    ram_cell[   12512] = 32'h0;  // 32'h0f69aadc;
    ram_cell[   12513] = 32'h0;  // 32'h9b4874ec;
    ram_cell[   12514] = 32'h0;  // 32'h87777de5;
    ram_cell[   12515] = 32'h0;  // 32'h95fddd09;
    ram_cell[   12516] = 32'h0;  // 32'h9aead3bc;
    ram_cell[   12517] = 32'h0;  // 32'hb6ff3bc0;
    ram_cell[   12518] = 32'h0;  // 32'h2a9bc396;
    ram_cell[   12519] = 32'h0;  // 32'hb36d2bf4;
    ram_cell[   12520] = 32'h0;  // 32'h627d600c;
    ram_cell[   12521] = 32'h0;  // 32'h824e2e04;
    ram_cell[   12522] = 32'h0;  // 32'h4062fd28;
    ram_cell[   12523] = 32'h0;  // 32'h148ddc01;
    ram_cell[   12524] = 32'h0;  // 32'h61b57730;
    ram_cell[   12525] = 32'h0;  // 32'h1a6694ff;
    ram_cell[   12526] = 32'h0;  // 32'h4d3622b7;
    ram_cell[   12527] = 32'h0;  // 32'hb34de91b;
    ram_cell[   12528] = 32'h0;  // 32'h79897530;
    ram_cell[   12529] = 32'h0;  // 32'h08b8ff3f;
    ram_cell[   12530] = 32'h0;  // 32'hd565b63c;
    ram_cell[   12531] = 32'h0;  // 32'h4af1a1c0;
    ram_cell[   12532] = 32'h0;  // 32'h87e99773;
    ram_cell[   12533] = 32'h0;  // 32'hfdb4af7d;
    ram_cell[   12534] = 32'h0;  // 32'h42fd9c07;
    ram_cell[   12535] = 32'h0;  // 32'h613b1205;
    ram_cell[   12536] = 32'h0;  // 32'hacf2369c;
    ram_cell[   12537] = 32'h0;  // 32'h1ae67008;
    ram_cell[   12538] = 32'h0;  // 32'h5f5ca2ea;
    ram_cell[   12539] = 32'h0;  // 32'hf9dc0d5e;
    ram_cell[   12540] = 32'h0;  // 32'h6122bf86;
    ram_cell[   12541] = 32'h0;  // 32'h80744ec6;
    ram_cell[   12542] = 32'h0;  // 32'h7508bb33;
    ram_cell[   12543] = 32'h0;  // 32'h4762dcea;
    ram_cell[   12544] = 32'h0;  // 32'hc26053c9;
    ram_cell[   12545] = 32'h0;  // 32'hc6d6de43;
    ram_cell[   12546] = 32'h0;  // 32'h879ebb45;
    ram_cell[   12547] = 32'h0;  // 32'h9940a9b4;
    ram_cell[   12548] = 32'h0;  // 32'h842ab976;
    ram_cell[   12549] = 32'h0;  // 32'h51680b5d;
    ram_cell[   12550] = 32'h0;  // 32'h8083b778;
    ram_cell[   12551] = 32'h0;  // 32'h2a90277a;
    ram_cell[   12552] = 32'h0;  // 32'hdbeefa32;
    ram_cell[   12553] = 32'h0;  // 32'h30103c2e;
    ram_cell[   12554] = 32'h0;  // 32'hfac39ce3;
    ram_cell[   12555] = 32'h0;  // 32'hbb91ba7f;
    ram_cell[   12556] = 32'h0;  // 32'h1b156233;
    ram_cell[   12557] = 32'h0;  // 32'h74aaf247;
    ram_cell[   12558] = 32'h0;  // 32'h3dcbc994;
    ram_cell[   12559] = 32'h0;  // 32'h4eb56fbe;
    ram_cell[   12560] = 32'h0;  // 32'h18d45802;
    ram_cell[   12561] = 32'h0;  // 32'h23252c68;
    ram_cell[   12562] = 32'h0;  // 32'h0bd45e2f;
    ram_cell[   12563] = 32'h0;  // 32'h92324af4;
    ram_cell[   12564] = 32'h0;  // 32'hcdcd5e0c;
    ram_cell[   12565] = 32'h0;  // 32'hcce4444e;
    ram_cell[   12566] = 32'h0;  // 32'hc347145d;
    ram_cell[   12567] = 32'h0;  // 32'hd82080fc;
    ram_cell[   12568] = 32'h0;  // 32'hd8f57107;
    ram_cell[   12569] = 32'h0;  // 32'h3ebf0b12;
    ram_cell[   12570] = 32'h0;  // 32'he654fc8f;
    ram_cell[   12571] = 32'h0;  // 32'h6ae59ad5;
    ram_cell[   12572] = 32'h0;  // 32'h3a9262c6;
    ram_cell[   12573] = 32'h0;  // 32'heac23775;
    ram_cell[   12574] = 32'h0;  // 32'hb9cc768d;
    ram_cell[   12575] = 32'h0;  // 32'h9ec8427d;
    ram_cell[   12576] = 32'h0;  // 32'h5fb92eee;
    ram_cell[   12577] = 32'h0;  // 32'h953811a0;
    ram_cell[   12578] = 32'h0;  // 32'h09d4116e;
    ram_cell[   12579] = 32'h0;  // 32'h8132f0b4;
    ram_cell[   12580] = 32'h0;  // 32'h4f15d6e5;
    ram_cell[   12581] = 32'h0;  // 32'hce3cdeac;
    ram_cell[   12582] = 32'h0;  // 32'he929e206;
    ram_cell[   12583] = 32'h0;  // 32'h6c26da69;
    ram_cell[   12584] = 32'h0;  // 32'h0bedaf64;
    ram_cell[   12585] = 32'h0;  // 32'h2f064afe;
    ram_cell[   12586] = 32'h0;  // 32'hd4a6c3b9;
    ram_cell[   12587] = 32'h0;  // 32'h84696438;
    ram_cell[   12588] = 32'h0;  // 32'ha9ec3681;
    ram_cell[   12589] = 32'h0;  // 32'h4312ed7a;
    ram_cell[   12590] = 32'h0;  // 32'hfeee1986;
    ram_cell[   12591] = 32'h0;  // 32'h75d37859;
    ram_cell[   12592] = 32'h0;  // 32'h67eb6cc3;
    ram_cell[   12593] = 32'h0;  // 32'h7d257a5b;
    ram_cell[   12594] = 32'h0;  // 32'h7c25455f;
    ram_cell[   12595] = 32'h0;  // 32'h2b65e331;
    ram_cell[   12596] = 32'h0;  // 32'h6b69d5a7;
    ram_cell[   12597] = 32'h0;  // 32'h24b08590;
    ram_cell[   12598] = 32'h0;  // 32'h577eac43;
    ram_cell[   12599] = 32'h0;  // 32'hc3fe91dc;
    ram_cell[   12600] = 32'h0;  // 32'hb3ea768e;
    ram_cell[   12601] = 32'h0;  // 32'h6b5c585f;
    ram_cell[   12602] = 32'h0;  // 32'hfb472677;
    ram_cell[   12603] = 32'h0;  // 32'hcb29f87b;
    ram_cell[   12604] = 32'h0;  // 32'h99331b49;
    ram_cell[   12605] = 32'h0;  // 32'h01db4723;
    ram_cell[   12606] = 32'h0;  // 32'h79ef7515;
    ram_cell[   12607] = 32'h0;  // 32'h9248fba4;
    ram_cell[   12608] = 32'h0;  // 32'hf8793736;
    ram_cell[   12609] = 32'h0;  // 32'h360c8f2c;
    ram_cell[   12610] = 32'h0;  // 32'hf330a324;
    ram_cell[   12611] = 32'h0;  // 32'h1b7f8d91;
    ram_cell[   12612] = 32'h0;  // 32'h853825dc;
    ram_cell[   12613] = 32'h0;  // 32'he4d86b22;
    ram_cell[   12614] = 32'h0;  // 32'h90c72efa;
    ram_cell[   12615] = 32'h0;  // 32'he008f637;
    ram_cell[   12616] = 32'h0;  // 32'h67323f41;
    ram_cell[   12617] = 32'h0;  // 32'h8f7cf830;
    ram_cell[   12618] = 32'h0;  // 32'h6e8e597f;
    ram_cell[   12619] = 32'h0;  // 32'ha2541a5f;
    ram_cell[   12620] = 32'h0;  // 32'h52a0dd76;
    ram_cell[   12621] = 32'h0;  // 32'h945592f5;
    ram_cell[   12622] = 32'h0;  // 32'h404127bd;
    ram_cell[   12623] = 32'h0;  // 32'ha824e767;
    ram_cell[   12624] = 32'h0;  // 32'h03408bb3;
    ram_cell[   12625] = 32'h0;  // 32'hc877f5a5;
    ram_cell[   12626] = 32'h0;  // 32'hf0024a8d;
    ram_cell[   12627] = 32'h0;  // 32'h3c423e34;
    ram_cell[   12628] = 32'h0;  // 32'h5c08880b;
    ram_cell[   12629] = 32'h0;  // 32'h63d341a8;
    ram_cell[   12630] = 32'h0;  // 32'hd2a3e9fd;
    ram_cell[   12631] = 32'h0;  // 32'ha18d5384;
    ram_cell[   12632] = 32'h0;  // 32'h1778d4e8;
    ram_cell[   12633] = 32'h0;  // 32'h31471ed3;
    ram_cell[   12634] = 32'h0;  // 32'h4704e31c;
    ram_cell[   12635] = 32'h0;  // 32'h2c9df269;
    ram_cell[   12636] = 32'h0;  // 32'hc7d8998e;
    ram_cell[   12637] = 32'h0;  // 32'hcfc97927;
    ram_cell[   12638] = 32'h0;  // 32'hf760df90;
    ram_cell[   12639] = 32'h0;  // 32'h67cf8081;
    ram_cell[   12640] = 32'h0;  // 32'h0e14476f;
    ram_cell[   12641] = 32'h0;  // 32'h11fd991e;
    ram_cell[   12642] = 32'h0;  // 32'hdca98ba1;
    ram_cell[   12643] = 32'h0;  // 32'haed98c5a;
    ram_cell[   12644] = 32'h0;  // 32'hce40ab61;
    ram_cell[   12645] = 32'h0;  // 32'hdd49d796;
    ram_cell[   12646] = 32'h0;  // 32'h65d6f45c;
    ram_cell[   12647] = 32'h0;  // 32'h3d18fea7;
    ram_cell[   12648] = 32'h0;  // 32'h4558c4b9;
    ram_cell[   12649] = 32'h0;  // 32'hab005047;
    ram_cell[   12650] = 32'h0;  // 32'h513c3a88;
    ram_cell[   12651] = 32'h0;  // 32'h6509c105;
    ram_cell[   12652] = 32'h0;  // 32'h72e70884;
    ram_cell[   12653] = 32'h0;  // 32'he55c142a;
    ram_cell[   12654] = 32'h0;  // 32'h86161ba8;
    ram_cell[   12655] = 32'h0;  // 32'h387132fb;
    ram_cell[   12656] = 32'h0;  // 32'hbc000c2f;
    ram_cell[   12657] = 32'h0;  // 32'h1d1fbc25;
    ram_cell[   12658] = 32'h0;  // 32'h1c28bd2e;
    ram_cell[   12659] = 32'h0;  // 32'he1ddc271;
    ram_cell[   12660] = 32'h0;  // 32'h9bc31d9f;
    ram_cell[   12661] = 32'h0;  // 32'h36331b9c;
    ram_cell[   12662] = 32'h0;  // 32'h527c4869;
    ram_cell[   12663] = 32'h0;  // 32'haa788625;
    ram_cell[   12664] = 32'h0;  // 32'he2bc9ed1;
    ram_cell[   12665] = 32'h0;  // 32'h9d8f6030;
    ram_cell[   12666] = 32'h0;  // 32'h8d9da3d1;
    ram_cell[   12667] = 32'h0;  // 32'h5b2cc9fa;
    ram_cell[   12668] = 32'h0;  // 32'h019df223;
    ram_cell[   12669] = 32'h0;  // 32'h8d814ef9;
    ram_cell[   12670] = 32'h0;  // 32'hab3fafd0;
    ram_cell[   12671] = 32'h0;  // 32'h48373150;
    ram_cell[   12672] = 32'h0;  // 32'hd67ac38e;
    ram_cell[   12673] = 32'h0;  // 32'ha619e01b;
    ram_cell[   12674] = 32'h0;  // 32'hea5ec423;
    ram_cell[   12675] = 32'h0;  // 32'h446ec671;
    ram_cell[   12676] = 32'h0;  // 32'h212463c0;
    ram_cell[   12677] = 32'h0;  // 32'h370f41b0;
    ram_cell[   12678] = 32'h0;  // 32'h523825d9;
    ram_cell[   12679] = 32'h0;  // 32'h592ab2f2;
    ram_cell[   12680] = 32'h0;  // 32'h008ed0e2;
    ram_cell[   12681] = 32'h0;  // 32'h1dedcf0e;
    ram_cell[   12682] = 32'h0;  // 32'h250839ee;
    ram_cell[   12683] = 32'h0;  // 32'h8e83ea0b;
    ram_cell[   12684] = 32'h0;  // 32'h3fc34b9d;
    ram_cell[   12685] = 32'h0;  // 32'h9e4a4998;
    ram_cell[   12686] = 32'h0;  // 32'h7b4cd2bd;
    ram_cell[   12687] = 32'h0;  // 32'h354d974e;
    ram_cell[   12688] = 32'h0;  // 32'hab00c54f;
    ram_cell[   12689] = 32'h0;  // 32'ha7bcf466;
    ram_cell[   12690] = 32'h0;  // 32'h1d000da0;
    ram_cell[   12691] = 32'h0;  // 32'h8591da07;
    ram_cell[   12692] = 32'h0;  // 32'hbd38da8d;
    ram_cell[   12693] = 32'h0;  // 32'h48bf199a;
    ram_cell[   12694] = 32'h0;  // 32'h3a60884a;
    ram_cell[   12695] = 32'h0;  // 32'h10c32ecf;
    ram_cell[   12696] = 32'h0;  // 32'h4a4247fe;
    ram_cell[   12697] = 32'h0;  // 32'h03b0037f;
    ram_cell[   12698] = 32'h0;  // 32'hc264911f;
    ram_cell[   12699] = 32'h0;  // 32'h2cc87d9f;
    ram_cell[   12700] = 32'h0;  // 32'hcc2f6007;
    ram_cell[   12701] = 32'h0;  // 32'he01296d6;
    ram_cell[   12702] = 32'h0;  // 32'h6385f5e6;
    ram_cell[   12703] = 32'h0;  // 32'h3c8966f4;
    ram_cell[   12704] = 32'h0;  // 32'h530949c6;
    ram_cell[   12705] = 32'h0;  // 32'h881d674e;
    ram_cell[   12706] = 32'h0;  // 32'h1eb6620e;
    ram_cell[   12707] = 32'h0;  // 32'hbc19a225;
    ram_cell[   12708] = 32'h0;  // 32'h7c8ed3eb;
    ram_cell[   12709] = 32'h0;  // 32'h3e5be373;
    ram_cell[   12710] = 32'h0;  // 32'h16d2d98b;
    ram_cell[   12711] = 32'h0;  // 32'h7a5b36a8;
    ram_cell[   12712] = 32'h0;  // 32'h94aef0dc;
    ram_cell[   12713] = 32'h0;  // 32'ha3ea5873;
    ram_cell[   12714] = 32'h0;  // 32'h0183432c;
    ram_cell[   12715] = 32'h0;  // 32'he1160315;
    ram_cell[   12716] = 32'h0;  // 32'hd9b16c25;
    ram_cell[   12717] = 32'h0;  // 32'h0b8cd74d;
    ram_cell[   12718] = 32'h0;  // 32'h8601e7ad;
    ram_cell[   12719] = 32'h0;  // 32'hf8529c45;
    ram_cell[   12720] = 32'h0;  // 32'hf429597e;
    ram_cell[   12721] = 32'h0;  // 32'h52c50212;
    ram_cell[   12722] = 32'h0;  // 32'hf45f3008;
    ram_cell[   12723] = 32'h0;  // 32'h79f31733;
    ram_cell[   12724] = 32'h0;  // 32'hbad36c55;
    ram_cell[   12725] = 32'h0;  // 32'h2a9ffe4a;
    ram_cell[   12726] = 32'h0;  // 32'h2ac40dcd;
    ram_cell[   12727] = 32'h0;  // 32'ha80e9f67;
    ram_cell[   12728] = 32'h0;  // 32'h235c888d;
    ram_cell[   12729] = 32'h0;  // 32'h8f786167;
    ram_cell[   12730] = 32'h0;  // 32'hd9201617;
    ram_cell[   12731] = 32'h0;  // 32'he39db957;
    ram_cell[   12732] = 32'h0;  // 32'ha4b177d6;
    ram_cell[   12733] = 32'h0;  // 32'h8ee697d9;
    ram_cell[   12734] = 32'h0;  // 32'hea879b22;
    ram_cell[   12735] = 32'h0;  // 32'h93fab016;
    ram_cell[   12736] = 32'h0;  // 32'h830c239f;
    ram_cell[   12737] = 32'h0;  // 32'ha9ac828d;
    ram_cell[   12738] = 32'h0;  // 32'hcee185c4;
    ram_cell[   12739] = 32'h0;  // 32'h94a682d1;
    ram_cell[   12740] = 32'h0;  // 32'hac11f7c3;
    ram_cell[   12741] = 32'h0;  // 32'hd1c4f95e;
    ram_cell[   12742] = 32'h0;  // 32'h3ade4e6c;
    ram_cell[   12743] = 32'h0;  // 32'h7de457b6;
    ram_cell[   12744] = 32'h0;  // 32'h97c31917;
    ram_cell[   12745] = 32'h0;  // 32'hedb43c36;
    ram_cell[   12746] = 32'h0;  // 32'he87bd066;
    ram_cell[   12747] = 32'h0;  // 32'h0d4b5418;
    ram_cell[   12748] = 32'h0;  // 32'hbbe9cc56;
    ram_cell[   12749] = 32'h0;  // 32'h622e86d4;
    ram_cell[   12750] = 32'h0;  // 32'h68b057b9;
    ram_cell[   12751] = 32'h0;  // 32'he2889bb9;
    ram_cell[   12752] = 32'h0;  // 32'hbd06b8b4;
    ram_cell[   12753] = 32'h0;  // 32'h824baac5;
    ram_cell[   12754] = 32'h0;  // 32'h6e08b17b;
    ram_cell[   12755] = 32'h0;  // 32'h197bd49f;
    ram_cell[   12756] = 32'h0;  // 32'h7a5266bf;
    ram_cell[   12757] = 32'h0;  // 32'h7f44aaaf;
    ram_cell[   12758] = 32'h0;  // 32'hf8c87951;
    ram_cell[   12759] = 32'h0;  // 32'h69ff18de;
    ram_cell[   12760] = 32'h0;  // 32'hc942a31d;
    ram_cell[   12761] = 32'h0;  // 32'h50f91ef1;
    ram_cell[   12762] = 32'h0;  // 32'h5cbf010a;
    ram_cell[   12763] = 32'h0;  // 32'hffc51b70;
    ram_cell[   12764] = 32'h0;  // 32'he60c511a;
    ram_cell[   12765] = 32'h0;  // 32'h85e9c996;
    ram_cell[   12766] = 32'h0;  // 32'h65e0b7d8;
    ram_cell[   12767] = 32'h0;  // 32'h937fd02e;
    ram_cell[   12768] = 32'h0;  // 32'h03fff196;
    ram_cell[   12769] = 32'h0;  // 32'h1aa6cbe0;
    ram_cell[   12770] = 32'h0;  // 32'hc544d026;
    ram_cell[   12771] = 32'h0;  // 32'h35b8b017;
    ram_cell[   12772] = 32'h0;  // 32'h28e41fe3;
    ram_cell[   12773] = 32'h0;  // 32'h3f03320a;
    ram_cell[   12774] = 32'h0;  // 32'h545f1559;
    ram_cell[   12775] = 32'h0;  // 32'h1da8652f;
    ram_cell[   12776] = 32'h0;  // 32'h6ece90e5;
    ram_cell[   12777] = 32'h0;  // 32'hb93f6d9b;
    ram_cell[   12778] = 32'h0;  // 32'h01438640;
    ram_cell[   12779] = 32'h0;  // 32'hbbf41bef;
    ram_cell[   12780] = 32'h0;  // 32'h8775e625;
    ram_cell[   12781] = 32'h0;  // 32'h7470ea5f;
    ram_cell[   12782] = 32'h0;  // 32'h909104da;
    ram_cell[   12783] = 32'h0;  // 32'he2afff05;
    ram_cell[   12784] = 32'h0;  // 32'h23708879;
    ram_cell[   12785] = 32'h0;  // 32'h412da762;
    ram_cell[   12786] = 32'h0;  // 32'h33d20bb0;
    ram_cell[   12787] = 32'h0;  // 32'hae3968e7;
    ram_cell[   12788] = 32'h0;  // 32'hebbe18b8;
    ram_cell[   12789] = 32'h0;  // 32'hd5accda5;
    ram_cell[   12790] = 32'h0;  // 32'hb404ed36;
    ram_cell[   12791] = 32'h0;  // 32'hd375bf84;
    ram_cell[   12792] = 32'h0;  // 32'hc441543b;
    ram_cell[   12793] = 32'h0;  // 32'h54f5ed20;
    ram_cell[   12794] = 32'h0;  // 32'hc351aa0d;
    ram_cell[   12795] = 32'h0;  // 32'ha25434eb;
    ram_cell[   12796] = 32'h0;  // 32'hef129a86;
    ram_cell[   12797] = 32'h0;  // 32'hb06fa267;
    ram_cell[   12798] = 32'h0;  // 32'hf6219ede;
    ram_cell[   12799] = 32'h0;  // 32'h3f1f716e;
    ram_cell[   12800] = 32'h0;  // 32'h8e501568;
    ram_cell[   12801] = 32'h0;  // 32'ha5d2ffb4;
    ram_cell[   12802] = 32'h0;  // 32'hcf448509;
    ram_cell[   12803] = 32'h0;  // 32'h3173a7c3;
    ram_cell[   12804] = 32'h0;  // 32'h91812181;
    ram_cell[   12805] = 32'h0;  // 32'ha9a29969;
    ram_cell[   12806] = 32'h0;  // 32'habddc19d;
    ram_cell[   12807] = 32'h0;  // 32'h121be30f;
    ram_cell[   12808] = 32'h0;  // 32'h022897ab;
    ram_cell[   12809] = 32'h0;  // 32'h6a02fd83;
    ram_cell[   12810] = 32'h0;  // 32'h84733e2d;
    ram_cell[   12811] = 32'h0;  // 32'ha089d3b1;
    ram_cell[   12812] = 32'h0;  // 32'h643549fe;
    ram_cell[   12813] = 32'h0;  // 32'hb1e77cf0;
    ram_cell[   12814] = 32'h0;  // 32'h541a9c42;
    ram_cell[   12815] = 32'h0;  // 32'h65a6dc69;
    ram_cell[   12816] = 32'h0;  // 32'hc5b1f045;
    ram_cell[   12817] = 32'h0;  // 32'h3bf9056a;
    ram_cell[   12818] = 32'h0;  // 32'h2bc5edc8;
    ram_cell[   12819] = 32'h0;  // 32'hdfb20922;
    ram_cell[   12820] = 32'h0;  // 32'h49384cb6;
    ram_cell[   12821] = 32'h0;  // 32'h51db8c77;
    ram_cell[   12822] = 32'h0;  // 32'h0c5dcf52;
    ram_cell[   12823] = 32'h0;  // 32'hc406da8e;
    ram_cell[   12824] = 32'h0;  // 32'h35d11aea;
    ram_cell[   12825] = 32'h0;  // 32'h77d2586f;
    ram_cell[   12826] = 32'h0;  // 32'h8dbc0a78;
    ram_cell[   12827] = 32'h0;  // 32'h76c3fdba;
    ram_cell[   12828] = 32'h0;  // 32'hcf693b97;
    ram_cell[   12829] = 32'h0;  // 32'h0d123e63;
    ram_cell[   12830] = 32'h0;  // 32'hd68284cd;
    ram_cell[   12831] = 32'h0;  // 32'h71f81625;
    ram_cell[   12832] = 32'h0;  // 32'h6bf673d7;
    ram_cell[   12833] = 32'h0;  // 32'h3fed214e;
    ram_cell[   12834] = 32'h0;  // 32'ha742768b;
    ram_cell[   12835] = 32'h0;  // 32'h26ec458a;
    ram_cell[   12836] = 32'h0;  // 32'hf2e953fb;
    ram_cell[   12837] = 32'h0;  // 32'h3fa0535f;
    ram_cell[   12838] = 32'h0;  // 32'hecb44adf;
    ram_cell[   12839] = 32'h0;  // 32'ha67f269f;
    ram_cell[   12840] = 32'h0;  // 32'hca912a87;
    ram_cell[   12841] = 32'h0;  // 32'h5bc83288;
    ram_cell[   12842] = 32'h0;  // 32'h2eadb154;
    ram_cell[   12843] = 32'h0;  // 32'hcecff48b;
    ram_cell[   12844] = 32'h0;  // 32'h2187b7f8;
    ram_cell[   12845] = 32'h0;  // 32'h77b85f5a;
    ram_cell[   12846] = 32'h0;  // 32'hd09f4b21;
    ram_cell[   12847] = 32'h0;  // 32'h0f8900f4;
    ram_cell[   12848] = 32'h0;  // 32'ha1ca941f;
    ram_cell[   12849] = 32'h0;  // 32'h1a9d10ff;
    ram_cell[   12850] = 32'h0;  // 32'h1b4f0593;
    ram_cell[   12851] = 32'h0;  // 32'ha0d65fa7;
    ram_cell[   12852] = 32'h0;  // 32'hc7a81108;
    ram_cell[   12853] = 32'h0;  // 32'h9fdc3a68;
    ram_cell[   12854] = 32'h0;  // 32'h34e0e175;
    ram_cell[   12855] = 32'h0;  // 32'h783bfdb0;
    ram_cell[   12856] = 32'h0;  // 32'h4ccc697c;
    ram_cell[   12857] = 32'h0;  // 32'h19e1c4db;
    ram_cell[   12858] = 32'h0;  // 32'h533e37a7;
    ram_cell[   12859] = 32'h0;  // 32'hb92b1dd4;
    ram_cell[   12860] = 32'h0;  // 32'h6e227fb5;
    ram_cell[   12861] = 32'h0;  // 32'h97bba148;
    ram_cell[   12862] = 32'h0;  // 32'h6564dae3;
    ram_cell[   12863] = 32'h0;  // 32'he9d65e93;
    ram_cell[   12864] = 32'h0;  // 32'ha531cda5;
    ram_cell[   12865] = 32'h0;  // 32'h77dfb421;
    ram_cell[   12866] = 32'h0;  // 32'hc498cfa3;
    ram_cell[   12867] = 32'h0;  // 32'hd264e864;
    ram_cell[   12868] = 32'h0;  // 32'h652023d8;
    ram_cell[   12869] = 32'h0;  // 32'he48b2431;
    ram_cell[   12870] = 32'h0;  // 32'h2d73eb8a;
    ram_cell[   12871] = 32'h0;  // 32'hfd604f2b;
    ram_cell[   12872] = 32'h0;  // 32'h07046113;
    ram_cell[   12873] = 32'h0;  // 32'h7b488c3b;
    ram_cell[   12874] = 32'h0;  // 32'h4463dc39;
    ram_cell[   12875] = 32'h0;  // 32'h8bcf2eed;
    ram_cell[   12876] = 32'h0;  // 32'he3cef51f;
    ram_cell[   12877] = 32'h0;  // 32'h8ec822b9;
    ram_cell[   12878] = 32'h0;  // 32'h86e464fc;
    ram_cell[   12879] = 32'h0;  // 32'h828499fe;
    ram_cell[   12880] = 32'h0;  // 32'h0f32b09b;
    ram_cell[   12881] = 32'h0;  // 32'h454cb0e7;
    ram_cell[   12882] = 32'h0;  // 32'hd8e4a6b9;
    ram_cell[   12883] = 32'h0;  // 32'hb3bd4e97;
    ram_cell[   12884] = 32'h0;  // 32'hea197a6f;
    ram_cell[   12885] = 32'h0;  // 32'hd64bb51a;
    ram_cell[   12886] = 32'h0;  // 32'hc4370037;
    ram_cell[   12887] = 32'h0;  // 32'h360bdf3a;
    ram_cell[   12888] = 32'h0;  // 32'h5e2fa86d;
    ram_cell[   12889] = 32'h0;  // 32'h07f3467f;
    ram_cell[   12890] = 32'h0;  // 32'ha19b1b6d;
    ram_cell[   12891] = 32'h0;  // 32'h9d429794;
    ram_cell[   12892] = 32'h0;  // 32'h4794d1d5;
    ram_cell[   12893] = 32'h0;  // 32'h8cbe8c68;
    ram_cell[   12894] = 32'h0;  // 32'hd90eb5f5;
    ram_cell[   12895] = 32'h0;  // 32'heb02aae8;
    ram_cell[   12896] = 32'h0;  // 32'h1d8f97da;
    ram_cell[   12897] = 32'h0;  // 32'hc6fc0570;
    ram_cell[   12898] = 32'h0;  // 32'h6badf2a9;
    ram_cell[   12899] = 32'h0;  // 32'hb959af1d;
    ram_cell[   12900] = 32'h0;  // 32'h80419cef;
    ram_cell[   12901] = 32'h0;  // 32'h8d3ce2d1;
    ram_cell[   12902] = 32'h0;  // 32'h9d838ed6;
    ram_cell[   12903] = 32'h0;  // 32'hae43a850;
    ram_cell[   12904] = 32'h0;  // 32'hb5c8f787;
    ram_cell[   12905] = 32'h0;  // 32'h05231e43;
    ram_cell[   12906] = 32'h0;  // 32'hfc30bd34;
    ram_cell[   12907] = 32'h0;  // 32'h96d0e569;
    ram_cell[   12908] = 32'h0;  // 32'h89665a98;
    ram_cell[   12909] = 32'h0;  // 32'h96ffe6e1;
    ram_cell[   12910] = 32'h0;  // 32'h11176a06;
    ram_cell[   12911] = 32'h0;  // 32'h7679ac1e;
    ram_cell[   12912] = 32'h0;  // 32'hb0c0fd08;
    ram_cell[   12913] = 32'h0;  // 32'ha95c3e06;
    ram_cell[   12914] = 32'h0;  // 32'h2c072d6a;
    ram_cell[   12915] = 32'h0;  // 32'h9c6dcf6e;
    ram_cell[   12916] = 32'h0;  // 32'h0bec728b;
    ram_cell[   12917] = 32'h0;  // 32'h19b6d146;
    ram_cell[   12918] = 32'h0;  // 32'ha1d00bfd;
    ram_cell[   12919] = 32'h0;  // 32'h905ca570;
    ram_cell[   12920] = 32'h0;  // 32'h968d7084;
    ram_cell[   12921] = 32'h0;  // 32'hfc401cd6;
    ram_cell[   12922] = 32'h0;  // 32'h4c9a0742;
    ram_cell[   12923] = 32'h0;  // 32'h670260a8;
    ram_cell[   12924] = 32'h0;  // 32'h60c52a76;
    ram_cell[   12925] = 32'h0;  // 32'h3ba99aaf;
    ram_cell[   12926] = 32'h0;  // 32'hea9c698f;
    ram_cell[   12927] = 32'h0;  // 32'h73683352;
    ram_cell[   12928] = 32'h0;  // 32'h32f8166f;
    ram_cell[   12929] = 32'h0;  // 32'hce925bab;
    ram_cell[   12930] = 32'h0;  // 32'h8d54ba40;
    ram_cell[   12931] = 32'h0;  // 32'hb422e57d;
    ram_cell[   12932] = 32'h0;  // 32'h8f3f5e9f;
    ram_cell[   12933] = 32'h0;  // 32'ha847ac54;
    ram_cell[   12934] = 32'h0;  // 32'h29023e0c;
    ram_cell[   12935] = 32'h0;  // 32'h96d0ba78;
    ram_cell[   12936] = 32'h0;  // 32'hecbef729;
    ram_cell[   12937] = 32'h0;  // 32'h4e995976;
    ram_cell[   12938] = 32'h0;  // 32'h2f660ab3;
    ram_cell[   12939] = 32'h0;  // 32'h6f17f9a4;
    ram_cell[   12940] = 32'h0;  // 32'hb894f5fc;
    ram_cell[   12941] = 32'h0;  // 32'hb31e25aa;
    ram_cell[   12942] = 32'h0;  // 32'hce891d1b;
    ram_cell[   12943] = 32'h0;  // 32'hdf82bfcf;
    ram_cell[   12944] = 32'h0;  // 32'h73d0140c;
    ram_cell[   12945] = 32'h0;  // 32'he09f8e00;
    ram_cell[   12946] = 32'h0;  // 32'h5b935919;
    ram_cell[   12947] = 32'h0;  // 32'h787e8ad6;
    ram_cell[   12948] = 32'h0;  // 32'hb8e5904d;
    ram_cell[   12949] = 32'h0;  // 32'h1966618b;
    ram_cell[   12950] = 32'h0;  // 32'h2a4b86f4;
    ram_cell[   12951] = 32'h0;  // 32'h3ffa1a2d;
    ram_cell[   12952] = 32'h0;  // 32'h7ec21a88;
    ram_cell[   12953] = 32'h0;  // 32'hefb9a95d;
    ram_cell[   12954] = 32'h0;  // 32'h03583bee;
    ram_cell[   12955] = 32'h0;  // 32'h85efe7bc;
    ram_cell[   12956] = 32'h0;  // 32'hf51bedba;
    ram_cell[   12957] = 32'h0;  // 32'h888d7f55;
    ram_cell[   12958] = 32'h0;  // 32'hd3ce99bd;
    ram_cell[   12959] = 32'h0;  // 32'h7c17e200;
    ram_cell[   12960] = 32'h0;  // 32'h8e36d354;
    ram_cell[   12961] = 32'h0;  // 32'h7da43131;
    ram_cell[   12962] = 32'h0;  // 32'hff4fe274;
    ram_cell[   12963] = 32'h0;  // 32'h3237fb6f;
    ram_cell[   12964] = 32'h0;  // 32'hbe00854d;
    ram_cell[   12965] = 32'h0;  // 32'h4d0b85e9;
    ram_cell[   12966] = 32'h0;  // 32'h562bb007;
    ram_cell[   12967] = 32'h0;  // 32'h985f3cf4;
    ram_cell[   12968] = 32'h0;  // 32'h6b1f806c;
    ram_cell[   12969] = 32'h0;  // 32'h986eaad0;
    ram_cell[   12970] = 32'h0;  // 32'h146bef93;
    ram_cell[   12971] = 32'h0;  // 32'h2fbcaac6;
    ram_cell[   12972] = 32'h0;  // 32'hf8c66a89;
    ram_cell[   12973] = 32'h0;  // 32'hc339df24;
    ram_cell[   12974] = 32'h0;  // 32'h0da28a03;
    ram_cell[   12975] = 32'h0;  // 32'h0e07ef28;
    ram_cell[   12976] = 32'h0;  // 32'hedc40f00;
    ram_cell[   12977] = 32'h0;  // 32'ha35647f2;
    ram_cell[   12978] = 32'h0;  // 32'h32aee1e7;
    ram_cell[   12979] = 32'h0;  // 32'h92b45d3d;
    ram_cell[   12980] = 32'h0;  // 32'hccfbe31d;
    ram_cell[   12981] = 32'h0;  // 32'h53cbe691;
    ram_cell[   12982] = 32'h0;  // 32'h696d9f03;
    ram_cell[   12983] = 32'h0;  // 32'h2eaf82c0;
    ram_cell[   12984] = 32'h0;  // 32'h61adae87;
    ram_cell[   12985] = 32'h0;  // 32'h52efc559;
    ram_cell[   12986] = 32'h0;  // 32'h902a30a1;
    ram_cell[   12987] = 32'h0;  // 32'hdbcb283e;
    ram_cell[   12988] = 32'h0;  // 32'h0b313eeb;
    ram_cell[   12989] = 32'h0;  // 32'h76ea8c5f;
    ram_cell[   12990] = 32'h0;  // 32'h67237f19;
    ram_cell[   12991] = 32'h0;  // 32'hcbd827b4;
    ram_cell[   12992] = 32'h0;  // 32'h9af8f1c6;
    ram_cell[   12993] = 32'h0;  // 32'he43b7059;
    ram_cell[   12994] = 32'h0;  // 32'h30c26ed7;
    ram_cell[   12995] = 32'h0;  // 32'h513d8815;
    ram_cell[   12996] = 32'h0;  // 32'h302b4aa4;
    ram_cell[   12997] = 32'h0;  // 32'hae51f315;
    ram_cell[   12998] = 32'h0;  // 32'h27907670;
    ram_cell[   12999] = 32'h0;  // 32'h96848678;
    ram_cell[   13000] = 32'h0;  // 32'h837eafc2;
    ram_cell[   13001] = 32'h0;  // 32'h15462c78;
    ram_cell[   13002] = 32'h0;  // 32'h549f6569;
    ram_cell[   13003] = 32'h0;  // 32'hed519468;
    ram_cell[   13004] = 32'h0;  // 32'ha4040ca5;
    ram_cell[   13005] = 32'h0;  // 32'hd8478f6f;
    ram_cell[   13006] = 32'h0;  // 32'h720de181;
    ram_cell[   13007] = 32'h0;  // 32'h4799130b;
    ram_cell[   13008] = 32'h0;  // 32'hfac2e1ca;
    ram_cell[   13009] = 32'h0;  // 32'h7af66e65;
    ram_cell[   13010] = 32'h0;  // 32'h8d6d4f03;
    ram_cell[   13011] = 32'h0;  // 32'h1b0511d2;
    ram_cell[   13012] = 32'h0;  // 32'hc7cd90a5;
    ram_cell[   13013] = 32'h0;  // 32'heed069f0;
    ram_cell[   13014] = 32'h0;  // 32'hb0c4428d;
    ram_cell[   13015] = 32'h0;  // 32'h7ad3dab7;
    ram_cell[   13016] = 32'h0;  // 32'h405c13ec;
    ram_cell[   13017] = 32'h0;  // 32'hbd1d3956;
    ram_cell[   13018] = 32'h0;  // 32'h0811c63b;
    ram_cell[   13019] = 32'h0;  // 32'h882573c7;
    ram_cell[   13020] = 32'h0;  // 32'hff15bae5;
    ram_cell[   13021] = 32'h0;  // 32'ha9f3d6de;
    ram_cell[   13022] = 32'h0;  // 32'he7730aa6;
    ram_cell[   13023] = 32'h0;  // 32'hffa8fb58;
    ram_cell[   13024] = 32'h0;  // 32'h0cce2e4f;
    ram_cell[   13025] = 32'h0;  // 32'h1d94d131;
    ram_cell[   13026] = 32'h0;  // 32'hcad826c1;
    ram_cell[   13027] = 32'h0;  // 32'h46bc33cb;
    ram_cell[   13028] = 32'h0;  // 32'h5e155d1f;
    ram_cell[   13029] = 32'h0;  // 32'ha05f7556;
    ram_cell[   13030] = 32'h0;  // 32'hd4f683ae;
    ram_cell[   13031] = 32'h0;  // 32'heb1adfcd;
    ram_cell[   13032] = 32'h0;  // 32'h2cf79108;
    ram_cell[   13033] = 32'h0;  // 32'hc1518c1b;
    ram_cell[   13034] = 32'h0;  // 32'h1355b2f8;
    ram_cell[   13035] = 32'h0;  // 32'ha69c521f;
    ram_cell[   13036] = 32'h0;  // 32'h00b4f21e;
    ram_cell[   13037] = 32'h0;  // 32'h21c2dd65;
    ram_cell[   13038] = 32'h0;  // 32'h945b0633;
    ram_cell[   13039] = 32'h0;  // 32'he26d4c4a;
    ram_cell[   13040] = 32'h0;  // 32'h44935440;
    ram_cell[   13041] = 32'h0;  // 32'haab30290;
    ram_cell[   13042] = 32'h0;  // 32'h92af1088;
    ram_cell[   13043] = 32'h0;  // 32'h6017a3e3;
    ram_cell[   13044] = 32'h0;  // 32'h8739bd3d;
    ram_cell[   13045] = 32'h0;  // 32'h339d7337;
    ram_cell[   13046] = 32'h0;  // 32'h03bb7c24;
    ram_cell[   13047] = 32'h0;  // 32'hbab846b3;
    ram_cell[   13048] = 32'h0;  // 32'hc37c1991;
    ram_cell[   13049] = 32'h0;  // 32'h58dbecd6;
    ram_cell[   13050] = 32'h0;  // 32'h93ad42e6;
    ram_cell[   13051] = 32'h0;  // 32'hefd15100;
    ram_cell[   13052] = 32'h0;  // 32'h2703104a;
    ram_cell[   13053] = 32'h0;  // 32'h0690c2a5;
    ram_cell[   13054] = 32'h0;  // 32'h8c6b8b64;
    ram_cell[   13055] = 32'h0;  // 32'hdf15620b;
    ram_cell[   13056] = 32'h0;  // 32'hf5e5de5d;
    ram_cell[   13057] = 32'h0;  // 32'h32e5f8a2;
    ram_cell[   13058] = 32'h0;  // 32'hec20b369;
    ram_cell[   13059] = 32'h0;  // 32'h87429c6c;
    ram_cell[   13060] = 32'h0;  // 32'h1817c11f;
    ram_cell[   13061] = 32'h0;  // 32'h7caa051d;
    ram_cell[   13062] = 32'h0;  // 32'ha4f8d3eb;
    ram_cell[   13063] = 32'h0;  // 32'h88e9c773;
    ram_cell[   13064] = 32'h0;  // 32'hd8e1a590;
    ram_cell[   13065] = 32'h0;  // 32'h4a4a3ecc;
    ram_cell[   13066] = 32'h0;  // 32'h81c552d1;
    ram_cell[   13067] = 32'h0;  // 32'hbd018ffb;
    ram_cell[   13068] = 32'h0;  // 32'h67c38319;
    ram_cell[   13069] = 32'h0;  // 32'hd3866bcf;
    ram_cell[   13070] = 32'h0;  // 32'h8eca4213;
    ram_cell[   13071] = 32'h0;  // 32'hc78701c6;
    ram_cell[   13072] = 32'h0;  // 32'hc1062bb5;
    ram_cell[   13073] = 32'h0;  // 32'h1146cac9;
    ram_cell[   13074] = 32'h0;  // 32'hcfbd3169;
    ram_cell[   13075] = 32'h0;  // 32'hafc94210;
    ram_cell[   13076] = 32'h0;  // 32'haea86b07;
    ram_cell[   13077] = 32'h0;  // 32'h83a1676c;
    ram_cell[   13078] = 32'h0;  // 32'h45862da2;
    ram_cell[   13079] = 32'h0;  // 32'h6bd764cc;
    ram_cell[   13080] = 32'h0;  // 32'h1f1b9b08;
    ram_cell[   13081] = 32'h0;  // 32'h65863683;
    ram_cell[   13082] = 32'h0;  // 32'hc209c14c;
    ram_cell[   13083] = 32'h0;  // 32'h0b0b2547;
    ram_cell[   13084] = 32'h0;  // 32'h184f1e41;
    ram_cell[   13085] = 32'h0;  // 32'hea7deb5f;
    ram_cell[   13086] = 32'h0;  // 32'h6db9ec28;
    ram_cell[   13087] = 32'h0;  // 32'h00a2f3b2;
    ram_cell[   13088] = 32'h0;  // 32'h3abbdb81;
    ram_cell[   13089] = 32'h0;  // 32'hae60a79c;
    ram_cell[   13090] = 32'h0;  // 32'hffcb84fd;
    ram_cell[   13091] = 32'h0;  // 32'hbdcebca2;
    ram_cell[   13092] = 32'h0;  // 32'h081d0897;
    ram_cell[   13093] = 32'h0;  // 32'hd7202aef;
    ram_cell[   13094] = 32'h0;  // 32'h1adf25a9;
    ram_cell[   13095] = 32'h0;  // 32'h87ad218a;
    ram_cell[   13096] = 32'h0;  // 32'h0b3d4beb;
    ram_cell[   13097] = 32'h0;  // 32'hcbc1bb93;
    ram_cell[   13098] = 32'h0;  // 32'hf796a92d;
    ram_cell[   13099] = 32'h0;  // 32'hfa681805;
    ram_cell[   13100] = 32'h0;  // 32'hedcff6e8;
    ram_cell[   13101] = 32'h0;  // 32'hd2ae9670;
    ram_cell[   13102] = 32'h0;  // 32'hb332b8c1;
    ram_cell[   13103] = 32'h0;  // 32'h464397fa;
    ram_cell[   13104] = 32'h0;  // 32'h204818a4;
    ram_cell[   13105] = 32'h0;  // 32'h525d6c2d;
    ram_cell[   13106] = 32'h0;  // 32'h8e3067f5;
    ram_cell[   13107] = 32'h0;  // 32'h9cf358ad;
    ram_cell[   13108] = 32'h0;  // 32'h30a8409d;
    ram_cell[   13109] = 32'h0;  // 32'hf7116641;
    ram_cell[   13110] = 32'h0;  // 32'hf5782807;
    ram_cell[   13111] = 32'h0;  // 32'hba4b2310;
    ram_cell[   13112] = 32'h0;  // 32'hf3071f3d;
    ram_cell[   13113] = 32'h0;  // 32'hf10e5c22;
    ram_cell[   13114] = 32'h0;  // 32'h2bf55849;
    ram_cell[   13115] = 32'h0;  // 32'hdc1950fb;
    ram_cell[   13116] = 32'h0;  // 32'h52cd2a08;
    ram_cell[   13117] = 32'h0;  // 32'hfc74d7c5;
    ram_cell[   13118] = 32'h0;  // 32'hbed8d6e3;
    ram_cell[   13119] = 32'h0;  // 32'he696dc21;
    ram_cell[   13120] = 32'h0;  // 32'h66df24e2;
    ram_cell[   13121] = 32'h0;  // 32'h43ec3184;
    ram_cell[   13122] = 32'h0;  // 32'hf810f606;
    ram_cell[   13123] = 32'h0;  // 32'h91fdf0b5;
    ram_cell[   13124] = 32'h0;  // 32'hd01e7b09;
    ram_cell[   13125] = 32'h0;  // 32'hea02f51d;
    ram_cell[   13126] = 32'h0;  // 32'hc1de865c;
    ram_cell[   13127] = 32'h0;  // 32'h8bf2cdb7;
    ram_cell[   13128] = 32'h0;  // 32'h5d2fbab6;
    ram_cell[   13129] = 32'h0;  // 32'h41f9d0f3;
    ram_cell[   13130] = 32'h0;  // 32'h9d1bba18;
    ram_cell[   13131] = 32'h0;  // 32'h2d823bd1;
    ram_cell[   13132] = 32'h0;  // 32'h0ec04729;
    ram_cell[   13133] = 32'h0;  // 32'h3aa8a04b;
    ram_cell[   13134] = 32'h0;  // 32'h51d1386c;
    ram_cell[   13135] = 32'h0;  // 32'h474f5b25;
    ram_cell[   13136] = 32'h0;  // 32'h52f6bbc7;
    ram_cell[   13137] = 32'h0;  // 32'h4c62c62c;
    ram_cell[   13138] = 32'h0;  // 32'h98d6bc09;
    ram_cell[   13139] = 32'h0;  // 32'h5445b0c5;
    ram_cell[   13140] = 32'h0;  // 32'hff171978;
    ram_cell[   13141] = 32'h0;  // 32'h88dc7ba8;
    ram_cell[   13142] = 32'h0;  // 32'h9df95758;
    ram_cell[   13143] = 32'h0;  // 32'ha4bd30de;
    ram_cell[   13144] = 32'h0;  // 32'h974c8a3c;
    ram_cell[   13145] = 32'h0;  // 32'h77f2fc8b;
    ram_cell[   13146] = 32'h0;  // 32'h44521585;
    ram_cell[   13147] = 32'h0;  // 32'he039dc1a;
    ram_cell[   13148] = 32'h0;  // 32'h279000dc;
    ram_cell[   13149] = 32'h0;  // 32'he9e4fc5b;
    ram_cell[   13150] = 32'h0;  // 32'h3b8c4f3f;
    ram_cell[   13151] = 32'h0;  // 32'ha04fa28a;
    ram_cell[   13152] = 32'h0;  // 32'h4a9a2161;
    ram_cell[   13153] = 32'h0;  // 32'h41b08a2e;
    ram_cell[   13154] = 32'h0;  // 32'hca53858e;
    ram_cell[   13155] = 32'h0;  // 32'he19f6466;
    ram_cell[   13156] = 32'h0;  // 32'h8d87063e;
    ram_cell[   13157] = 32'h0;  // 32'h3cf2a0e0;
    ram_cell[   13158] = 32'h0;  // 32'hf0e7f7f1;
    ram_cell[   13159] = 32'h0;  // 32'h8526e585;
    ram_cell[   13160] = 32'h0;  // 32'hea9a64b4;
    ram_cell[   13161] = 32'h0;  // 32'hd2d1c4c7;
    ram_cell[   13162] = 32'h0;  // 32'h23901f3d;
    ram_cell[   13163] = 32'h0;  // 32'hc47692cf;
    ram_cell[   13164] = 32'h0;  // 32'he0e3c1f0;
    ram_cell[   13165] = 32'h0;  // 32'hc1ec1327;
    ram_cell[   13166] = 32'h0;  // 32'h9a7cf68e;
    ram_cell[   13167] = 32'h0;  // 32'h118c620f;
    ram_cell[   13168] = 32'h0;  // 32'h73edd288;
    ram_cell[   13169] = 32'h0;  // 32'h71d78b3f;
    ram_cell[   13170] = 32'h0;  // 32'h6e6ebc59;
    ram_cell[   13171] = 32'h0;  // 32'h21fcee39;
    ram_cell[   13172] = 32'h0;  // 32'h06d8acf4;
    ram_cell[   13173] = 32'h0;  // 32'h0aae9dc5;
    ram_cell[   13174] = 32'h0;  // 32'hbeb4c768;
    ram_cell[   13175] = 32'h0;  // 32'hdcbaf07e;
    ram_cell[   13176] = 32'h0;  // 32'h6cf1979b;
    ram_cell[   13177] = 32'h0;  // 32'h82f7163d;
    ram_cell[   13178] = 32'h0;  // 32'h6c6b2704;
    ram_cell[   13179] = 32'h0;  // 32'haddc959a;
    ram_cell[   13180] = 32'h0;  // 32'h4b570715;
    ram_cell[   13181] = 32'h0;  // 32'had33d1ba;
    ram_cell[   13182] = 32'h0;  // 32'h7f8d6890;
    ram_cell[   13183] = 32'h0;  // 32'h79d08a00;
    ram_cell[   13184] = 32'h0;  // 32'hf509246a;
    ram_cell[   13185] = 32'h0;  // 32'hc20dfb43;
    ram_cell[   13186] = 32'h0;  // 32'h95ae8d7c;
    ram_cell[   13187] = 32'h0;  // 32'h5ebb1a4e;
    ram_cell[   13188] = 32'h0;  // 32'hc5b30412;
    ram_cell[   13189] = 32'h0;  // 32'h594959c5;
    ram_cell[   13190] = 32'h0;  // 32'h695198e5;
    ram_cell[   13191] = 32'h0;  // 32'h82f94bb4;
    ram_cell[   13192] = 32'h0;  // 32'hd48fdd01;
    ram_cell[   13193] = 32'h0;  // 32'hd5275638;
    ram_cell[   13194] = 32'h0;  // 32'h20aec9de;
    ram_cell[   13195] = 32'h0;  // 32'he5871797;
    ram_cell[   13196] = 32'h0;  // 32'h1ce2fd44;
    ram_cell[   13197] = 32'h0;  // 32'hc97970b3;
    ram_cell[   13198] = 32'h0;  // 32'h6bd963da;
    ram_cell[   13199] = 32'h0;  // 32'h2330f853;
    ram_cell[   13200] = 32'h0;  // 32'he374e00b;
    ram_cell[   13201] = 32'h0;  // 32'hd4bde3e7;
    ram_cell[   13202] = 32'h0;  // 32'hbda2b19d;
    ram_cell[   13203] = 32'h0;  // 32'h91681f34;
    ram_cell[   13204] = 32'h0;  // 32'hd2a09292;
    ram_cell[   13205] = 32'h0;  // 32'h906c67a0;
    ram_cell[   13206] = 32'h0;  // 32'h1a766561;
    ram_cell[   13207] = 32'h0;  // 32'hcc33ba0c;
    ram_cell[   13208] = 32'h0;  // 32'h40522bf7;
    ram_cell[   13209] = 32'h0;  // 32'h21265ba7;
    ram_cell[   13210] = 32'h0;  // 32'he66d4433;
    ram_cell[   13211] = 32'h0;  // 32'h05837d53;
    ram_cell[   13212] = 32'h0;  // 32'hfc4ee2c0;
    ram_cell[   13213] = 32'h0;  // 32'h8f96e3bb;
    ram_cell[   13214] = 32'h0;  // 32'h283ff0b4;
    ram_cell[   13215] = 32'h0;  // 32'hb2c372c7;
    ram_cell[   13216] = 32'h0;  // 32'hb72a2aed;
    ram_cell[   13217] = 32'h0;  // 32'hc8216564;
    ram_cell[   13218] = 32'h0;  // 32'h618b5a07;
    ram_cell[   13219] = 32'h0;  // 32'h95f7d3f7;
    ram_cell[   13220] = 32'h0;  // 32'hb350eb12;
    ram_cell[   13221] = 32'h0;  // 32'h4c0f89ac;
    ram_cell[   13222] = 32'h0;  // 32'hd601de99;
    ram_cell[   13223] = 32'h0;  // 32'h7c532d51;
    ram_cell[   13224] = 32'h0;  // 32'hacf91e55;
    ram_cell[   13225] = 32'h0;  // 32'h3f1d1d45;
    ram_cell[   13226] = 32'h0;  // 32'hf3a903b2;
    ram_cell[   13227] = 32'h0;  // 32'h00a7084e;
    ram_cell[   13228] = 32'h0;  // 32'hf0d97b57;
    ram_cell[   13229] = 32'h0;  // 32'ha20942a0;
    ram_cell[   13230] = 32'h0;  // 32'h9d9bf3cc;
    ram_cell[   13231] = 32'h0;  // 32'h63d3e28b;
    ram_cell[   13232] = 32'h0;  // 32'h99233f5e;
    ram_cell[   13233] = 32'h0;  // 32'h71227417;
    ram_cell[   13234] = 32'h0;  // 32'h2fb3423a;
    ram_cell[   13235] = 32'h0;  // 32'hb126c92a;
    ram_cell[   13236] = 32'h0;  // 32'h58bd8da3;
    ram_cell[   13237] = 32'h0;  // 32'habde98f9;
    ram_cell[   13238] = 32'h0;  // 32'hadb13193;
    ram_cell[   13239] = 32'h0;  // 32'h90a4879c;
    ram_cell[   13240] = 32'h0;  // 32'h8b1c1f61;
    ram_cell[   13241] = 32'h0;  // 32'h8e20d87b;
    ram_cell[   13242] = 32'h0;  // 32'h4200cfc1;
    ram_cell[   13243] = 32'h0;  // 32'h28bc0565;
    ram_cell[   13244] = 32'h0;  // 32'hb5933fe1;
    ram_cell[   13245] = 32'h0;  // 32'h864cce2c;
    ram_cell[   13246] = 32'h0;  // 32'hf413c11a;
    ram_cell[   13247] = 32'h0;  // 32'h675b2aec;
    ram_cell[   13248] = 32'h0;  // 32'hfa63128e;
    ram_cell[   13249] = 32'h0;  // 32'h683fa978;
    ram_cell[   13250] = 32'h0;  // 32'hd9f00e00;
    ram_cell[   13251] = 32'h0;  // 32'h647a3cf9;
    ram_cell[   13252] = 32'h0;  // 32'hb52edd8d;
    ram_cell[   13253] = 32'h0;  // 32'h4ef73f35;
    ram_cell[   13254] = 32'h0;  // 32'h29cf3b81;
    ram_cell[   13255] = 32'h0;  // 32'hbda081e4;
    ram_cell[   13256] = 32'h0;  // 32'ha3e465db;
    ram_cell[   13257] = 32'h0;  // 32'hc42c7f2c;
    ram_cell[   13258] = 32'h0;  // 32'had4cfb82;
    ram_cell[   13259] = 32'h0;  // 32'hc53729d4;
    ram_cell[   13260] = 32'h0;  // 32'h3a15833b;
    ram_cell[   13261] = 32'h0;  // 32'h9d7f0269;
    ram_cell[   13262] = 32'h0;  // 32'h5d858e64;
    ram_cell[   13263] = 32'h0;  // 32'heefe69fb;
    ram_cell[   13264] = 32'h0;  // 32'h97b99e8e;
    ram_cell[   13265] = 32'h0;  // 32'h2925dcc6;
    ram_cell[   13266] = 32'h0;  // 32'hd92585c5;
    ram_cell[   13267] = 32'h0;  // 32'h9e2beafb;
    ram_cell[   13268] = 32'h0;  // 32'hd85c93ad;
    ram_cell[   13269] = 32'h0;  // 32'h35998d90;
    ram_cell[   13270] = 32'h0;  // 32'h563dd331;
    ram_cell[   13271] = 32'h0;  // 32'h6a8e2788;
    ram_cell[   13272] = 32'h0;  // 32'h28fce454;
    ram_cell[   13273] = 32'h0;  // 32'h36c4aac5;
    ram_cell[   13274] = 32'h0;  // 32'ha561bfac;
    ram_cell[   13275] = 32'h0;  // 32'h90419c83;
    ram_cell[   13276] = 32'h0;  // 32'h1d22aca4;
    ram_cell[   13277] = 32'h0;  // 32'h10d5df65;
    ram_cell[   13278] = 32'h0;  // 32'hcb4a4f5a;
    ram_cell[   13279] = 32'h0;  // 32'h466d457e;
    ram_cell[   13280] = 32'h0;  // 32'h597ec995;
    ram_cell[   13281] = 32'h0;  // 32'hbcad51d3;
    ram_cell[   13282] = 32'h0;  // 32'he9afa236;
    ram_cell[   13283] = 32'h0;  // 32'h37e816e8;
    ram_cell[   13284] = 32'h0;  // 32'h39b4354f;
    ram_cell[   13285] = 32'h0;  // 32'h66be5682;
    ram_cell[   13286] = 32'h0;  // 32'ha958ac39;
    ram_cell[   13287] = 32'h0;  // 32'h47e4e84e;
    ram_cell[   13288] = 32'h0;  // 32'h29fccbf6;
    ram_cell[   13289] = 32'h0;  // 32'h30bc488d;
    ram_cell[   13290] = 32'h0;  // 32'h2db172e5;
    ram_cell[   13291] = 32'h0;  // 32'he8547650;
    ram_cell[   13292] = 32'h0;  // 32'hee729372;
    ram_cell[   13293] = 32'h0;  // 32'hb5007993;
    ram_cell[   13294] = 32'h0;  // 32'h8defa5b7;
    ram_cell[   13295] = 32'h0;  // 32'h89807bd2;
    ram_cell[   13296] = 32'h0;  // 32'h05615f8e;
    ram_cell[   13297] = 32'h0;  // 32'hd8a7046f;
    ram_cell[   13298] = 32'h0;  // 32'h4e802fc8;
    ram_cell[   13299] = 32'h0;  // 32'h71209f1d;
    ram_cell[   13300] = 32'h0;  // 32'h91c71a76;
    ram_cell[   13301] = 32'h0;  // 32'h7b90662e;
    ram_cell[   13302] = 32'h0;  // 32'h286edfa4;
    ram_cell[   13303] = 32'h0;  // 32'haa0f9680;
    ram_cell[   13304] = 32'h0;  // 32'h2a7c18f6;
    ram_cell[   13305] = 32'h0;  // 32'hc708af67;
    ram_cell[   13306] = 32'h0;  // 32'hccc9abd0;
    ram_cell[   13307] = 32'h0;  // 32'hc9fa19a1;
    ram_cell[   13308] = 32'h0;  // 32'h9482e1e7;
    ram_cell[   13309] = 32'h0;  // 32'h63fed14a;
    ram_cell[   13310] = 32'h0;  // 32'haed5e647;
    ram_cell[   13311] = 32'h0;  // 32'ha4e0e540;
    ram_cell[   13312] = 32'h0;  // 32'h4fb74d67;
    ram_cell[   13313] = 32'h0;  // 32'h76286994;
    ram_cell[   13314] = 32'h0;  // 32'h78a22b13;
    ram_cell[   13315] = 32'h0;  // 32'h459df7df;
    ram_cell[   13316] = 32'h0;  // 32'hbe47d116;
    ram_cell[   13317] = 32'h0;  // 32'h565c66c3;
    ram_cell[   13318] = 32'h0;  // 32'h07fcbefa;
    ram_cell[   13319] = 32'h0;  // 32'hde110982;
    ram_cell[   13320] = 32'h0;  // 32'h0c122cfc;
    ram_cell[   13321] = 32'h0;  // 32'h9b23e43a;
    ram_cell[   13322] = 32'h0;  // 32'hb3a14217;
    ram_cell[   13323] = 32'h0;  // 32'hff49e7dc;
    ram_cell[   13324] = 32'h0;  // 32'hd13e2195;
    ram_cell[   13325] = 32'h0;  // 32'h0d06dec6;
    ram_cell[   13326] = 32'h0;  // 32'h38e05a66;
    ram_cell[   13327] = 32'h0;  // 32'h695ded47;
    ram_cell[   13328] = 32'h0;  // 32'h3d8693b1;
    ram_cell[   13329] = 32'h0;  // 32'h5e02ba3f;
    ram_cell[   13330] = 32'h0;  // 32'h6a062581;
    ram_cell[   13331] = 32'h0;  // 32'h10f362bd;
    ram_cell[   13332] = 32'h0;  // 32'h54a46264;
    ram_cell[   13333] = 32'h0;  // 32'ha2deff0a;
    ram_cell[   13334] = 32'h0;  // 32'hc0db31a0;
    ram_cell[   13335] = 32'h0;  // 32'h59601cb1;
    ram_cell[   13336] = 32'h0;  // 32'h18837c69;
    ram_cell[   13337] = 32'h0;  // 32'ha2354d96;
    ram_cell[   13338] = 32'h0;  // 32'h2d816b93;
    ram_cell[   13339] = 32'h0;  // 32'hf4de1382;
    ram_cell[   13340] = 32'h0;  // 32'h46808605;
    ram_cell[   13341] = 32'h0;  // 32'hc0fbaf5b;
    ram_cell[   13342] = 32'h0;  // 32'h71d57d3e;
    ram_cell[   13343] = 32'h0;  // 32'hc782d327;
    ram_cell[   13344] = 32'h0;  // 32'h021bee04;
    ram_cell[   13345] = 32'h0;  // 32'hd1a9ea3f;
    ram_cell[   13346] = 32'h0;  // 32'h194e7993;
    ram_cell[   13347] = 32'h0;  // 32'hbcf5ec6b;
    ram_cell[   13348] = 32'h0;  // 32'h704a5198;
    ram_cell[   13349] = 32'h0;  // 32'hdf810f5b;
    ram_cell[   13350] = 32'h0;  // 32'h6e08178c;
    ram_cell[   13351] = 32'h0;  // 32'hbd821848;
    ram_cell[   13352] = 32'h0;  // 32'hde51c320;
    ram_cell[   13353] = 32'h0;  // 32'h317cd032;
    ram_cell[   13354] = 32'h0;  // 32'h14ad2306;
    ram_cell[   13355] = 32'h0;  // 32'h20c803a1;
    ram_cell[   13356] = 32'h0;  // 32'hd0e627fd;
    ram_cell[   13357] = 32'h0;  // 32'h73f6a591;
    ram_cell[   13358] = 32'h0;  // 32'hc3dab858;
    ram_cell[   13359] = 32'h0;  // 32'h546a541d;
    ram_cell[   13360] = 32'h0;  // 32'hbc2f189b;
    ram_cell[   13361] = 32'h0;  // 32'h8100ff1a;
    ram_cell[   13362] = 32'h0;  // 32'hcb4592ac;
    ram_cell[   13363] = 32'h0;  // 32'he73d902e;
    ram_cell[   13364] = 32'h0;  // 32'h4e2063ce;
    ram_cell[   13365] = 32'h0;  // 32'h49b108e2;
    ram_cell[   13366] = 32'h0;  // 32'h483f47a9;
    ram_cell[   13367] = 32'h0;  // 32'hc17d9cbb;
    ram_cell[   13368] = 32'h0;  // 32'hb5994836;
    ram_cell[   13369] = 32'h0;  // 32'hd3055a7d;
    ram_cell[   13370] = 32'h0;  // 32'h0d18a29e;
    ram_cell[   13371] = 32'h0;  // 32'h5909a6c4;
    ram_cell[   13372] = 32'h0;  // 32'he8edf5f3;
    ram_cell[   13373] = 32'h0;  // 32'h0e9b2af7;
    ram_cell[   13374] = 32'h0;  // 32'hd21f973f;
    ram_cell[   13375] = 32'h0;  // 32'hef7b020b;
    ram_cell[   13376] = 32'h0;  // 32'h4b7e75aa;
    ram_cell[   13377] = 32'h0;  // 32'h4419a183;
    ram_cell[   13378] = 32'h0;  // 32'h6ce92e44;
    ram_cell[   13379] = 32'h0;  // 32'hf888a573;
    ram_cell[   13380] = 32'h0;  // 32'hdffb6357;
    ram_cell[   13381] = 32'h0;  // 32'h2c00b508;
    ram_cell[   13382] = 32'h0;  // 32'hbdd86bcd;
    ram_cell[   13383] = 32'h0;  // 32'h4d14ece3;
    ram_cell[   13384] = 32'h0;  // 32'h63d4f060;
    ram_cell[   13385] = 32'h0;  // 32'h738f4c88;
    ram_cell[   13386] = 32'h0;  // 32'hb1d6c8fd;
    ram_cell[   13387] = 32'h0;  // 32'hbb8085a0;
    ram_cell[   13388] = 32'h0;  // 32'h6d581f7e;
    ram_cell[   13389] = 32'h0;  // 32'h753d982f;
    ram_cell[   13390] = 32'h0;  // 32'he0d55bd2;
    ram_cell[   13391] = 32'h0;  // 32'h75e9b8db;
    ram_cell[   13392] = 32'h0;  // 32'h2e6e2ece;
    ram_cell[   13393] = 32'h0;  // 32'he870da8b;
    ram_cell[   13394] = 32'h0;  // 32'ha31988ff;
    ram_cell[   13395] = 32'h0;  // 32'h760e26eb;
    ram_cell[   13396] = 32'h0;  // 32'h982eeb9f;
    ram_cell[   13397] = 32'h0;  // 32'h3f898018;
    ram_cell[   13398] = 32'h0;  // 32'h0ffc7f45;
    ram_cell[   13399] = 32'h0;  // 32'h18d4d206;
    ram_cell[   13400] = 32'h0;  // 32'h8feef1d8;
    ram_cell[   13401] = 32'h0;  // 32'h9316ed3f;
    ram_cell[   13402] = 32'h0;  // 32'hce5752cb;
    ram_cell[   13403] = 32'h0;  // 32'h019a5c4f;
    ram_cell[   13404] = 32'h0;  // 32'hd7c19e21;
    ram_cell[   13405] = 32'h0;  // 32'h5b41260b;
    ram_cell[   13406] = 32'h0;  // 32'h359a941e;
    ram_cell[   13407] = 32'h0;  // 32'h3a558c6d;
    ram_cell[   13408] = 32'h0;  // 32'hc3254378;
    ram_cell[   13409] = 32'h0;  // 32'hd42d80be;
    ram_cell[   13410] = 32'h0;  // 32'h1fc5b45e;
    ram_cell[   13411] = 32'h0;  // 32'h0c810949;
    ram_cell[   13412] = 32'h0;  // 32'hb347fa90;
    ram_cell[   13413] = 32'h0;  // 32'h3c40e9a2;
    ram_cell[   13414] = 32'h0;  // 32'h8b3f989a;
    ram_cell[   13415] = 32'h0;  // 32'h5037b0e8;
    ram_cell[   13416] = 32'h0;  // 32'hc50322e2;
    ram_cell[   13417] = 32'h0;  // 32'hdc52c672;
    ram_cell[   13418] = 32'h0;  // 32'h8891c4c0;
    ram_cell[   13419] = 32'h0;  // 32'hd90a3efb;
    ram_cell[   13420] = 32'h0;  // 32'h1db96e3b;
    ram_cell[   13421] = 32'h0;  // 32'h5e1426f2;
    ram_cell[   13422] = 32'h0;  // 32'h15bbf426;
    ram_cell[   13423] = 32'h0;  // 32'h30927141;
    ram_cell[   13424] = 32'h0;  // 32'h4d3902a5;
    ram_cell[   13425] = 32'h0;  // 32'hbae79b68;
    ram_cell[   13426] = 32'h0;  // 32'h60b9d9c8;
    ram_cell[   13427] = 32'h0;  // 32'h11d1b6e0;
    ram_cell[   13428] = 32'h0;  // 32'h26e55cf2;
    ram_cell[   13429] = 32'h0;  // 32'h737dc45a;
    ram_cell[   13430] = 32'h0;  // 32'h2b9e27ba;
    ram_cell[   13431] = 32'h0;  // 32'h50473b0a;
    ram_cell[   13432] = 32'h0;  // 32'he692f41e;
    ram_cell[   13433] = 32'h0;  // 32'haf82758c;
    ram_cell[   13434] = 32'h0;  // 32'h5f3e883f;
    ram_cell[   13435] = 32'h0;  // 32'h89d447b0;
    ram_cell[   13436] = 32'h0;  // 32'hae52079f;
    ram_cell[   13437] = 32'h0;  // 32'hec57ea30;
    ram_cell[   13438] = 32'h0;  // 32'h480070f4;
    ram_cell[   13439] = 32'h0;  // 32'h4bec2e62;
    ram_cell[   13440] = 32'h0;  // 32'h2e031128;
    ram_cell[   13441] = 32'h0;  // 32'habc6fb4e;
    ram_cell[   13442] = 32'h0;  // 32'h9dd29c93;
    ram_cell[   13443] = 32'h0;  // 32'h06f8522b;
    ram_cell[   13444] = 32'h0;  // 32'h9fd20ce0;
    ram_cell[   13445] = 32'h0;  // 32'h17ba231c;
    ram_cell[   13446] = 32'h0;  // 32'h19771ecd;
    ram_cell[   13447] = 32'h0;  // 32'h62d129f6;
    ram_cell[   13448] = 32'h0;  // 32'h7933a7d6;
    ram_cell[   13449] = 32'h0;  // 32'h3ca5b86e;
    ram_cell[   13450] = 32'h0;  // 32'hdc127a45;
    ram_cell[   13451] = 32'h0;  // 32'h97632738;
    ram_cell[   13452] = 32'h0;  // 32'hd33e0188;
    ram_cell[   13453] = 32'h0;  // 32'h61e300a7;
    ram_cell[   13454] = 32'h0;  // 32'h37f18d29;
    ram_cell[   13455] = 32'h0;  // 32'he9826d9e;
    ram_cell[   13456] = 32'h0;  // 32'h80aa8651;
    ram_cell[   13457] = 32'h0;  // 32'h5b08abc6;
    ram_cell[   13458] = 32'h0;  // 32'haed52454;
    ram_cell[   13459] = 32'h0;  // 32'h2552056d;
    ram_cell[   13460] = 32'h0;  // 32'hed6154b0;
    ram_cell[   13461] = 32'h0;  // 32'hea034f51;
    ram_cell[   13462] = 32'h0;  // 32'he69f9b74;
    ram_cell[   13463] = 32'h0;  // 32'h8af90a77;
    ram_cell[   13464] = 32'h0;  // 32'hb0e39949;
    ram_cell[   13465] = 32'h0;  // 32'hf5f51199;
    ram_cell[   13466] = 32'h0;  // 32'h0e1cf341;
    ram_cell[   13467] = 32'h0;  // 32'hd8973c9e;
    ram_cell[   13468] = 32'h0;  // 32'h203db4e4;
    ram_cell[   13469] = 32'h0;  // 32'h5ebbac97;
    ram_cell[   13470] = 32'h0;  // 32'h8b4e49e8;
    ram_cell[   13471] = 32'h0;  // 32'h85568bb7;
    ram_cell[   13472] = 32'h0;  // 32'h5813b9c5;
    ram_cell[   13473] = 32'h0;  // 32'h010ebd37;
    ram_cell[   13474] = 32'h0;  // 32'h747f3b16;
    ram_cell[   13475] = 32'h0;  // 32'h85892175;
    ram_cell[   13476] = 32'h0;  // 32'h81f65a67;
    ram_cell[   13477] = 32'h0;  // 32'hc05f1184;
    ram_cell[   13478] = 32'h0;  // 32'h233a9e6f;
    ram_cell[   13479] = 32'h0;  // 32'hd8cea61c;
    ram_cell[   13480] = 32'h0;  // 32'h496bfb08;
    ram_cell[   13481] = 32'h0;  // 32'h784f3935;
    ram_cell[   13482] = 32'h0;  // 32'h069fc305;
    ram_cell[   13483] = 32'h0;  // 32'h8ff2400c;
    ram_cell[   13484] = 32'h0;  // 32'h5b90bb63;
    ram_cell[   13485] = 32'h0;  // 32'hc70db577;
    ram_cell[   13486] = 32'h0;  // 32'ha01bbfce;
    ram_cell[   13487] = 32'h0;  // 32'hbd03298c;
    ram_cell[   13488] = 32'h0;  // 32'hadcac17c;
    ram_cell[   13489] = 32'h0;  // 32'hc63cb218;
    ram_cell[   13490] = 32'h0;  // 32'h62890a28;
    ram_cell[   13491] = 32'h0;  // 32'he3d014b1;
    ram_cell[   13492] = 32'h0;  // 32'h3a22c79e;
    ram_cell[   13493] = 32'h0;  // 32'h954b979e;
    ram_cell[   13494] = 32'h0;  // 32'h10a6f279;
    ram_cell[   13495] = 32'h0;  // 32'hb956029d;
    ram_cell[   13496] = 32'h0;  // 32'ha7ba4118;
    ram_cell[   13497] = 32'h0;  // 32'h77c1e8b0;
    ram_cell[   13498] = 32'h0;  // 32'h8aebd9a8;
    ram_cell[   13499] = 32'h0;  // 32'hda701db7;
    ram_cell[   13500] = 32'h0;  // 32'h4dad6850;
    ram_cell[   13501] = 32'h0;  // 32'h0a6bf296;
    ram_cell[   13502] = 32'h0;  // 32'hdec81123;
    ram_cell[   13503] = 32'h0;  // 32'hbffabdb1;
    ram_cell[   13504] = 32'h0;  // 32'h5ade79ef;
    ram_cell[   13505] = 32'h0;  // 32'h09111d2a;
    ram_cell[   13506] = 32'h0;  // 32'h7a91e05c;
    ram_cell[   13507] = 32'h0;  // 32'haaf1a547;
    ram_cell[   13508] = 32'h0;  // 32'h3eec4939;
    ram_cell[   13509] = 32'h0;  // 32'h86f6072a;
    ram_cell[   13510] = 32'h0;  // 32'h36b13944;
    ram_cell[   13511] = 32'h0;  // 32'h787cb5d7;
    ram_cell[   13512] = 32'h0;  // 32'he9a3d01f;
    ram_cell[   13513] = 32'h0;  // 32'h76187684;
    ram_cell[   13514] = 32'h0;  // 32'h6e2fcce8;
    ram_cell[   13515] = 32'h0;  // 32'h4dbf03d1;
    ram_cell[   13516] = 32'h0;  // 32'h2d56ca10;
    ram_cell[   13517] = 32'h0;  // 32'h4e7b788a;
    ram_cell[   13518] = 32'h0;  // 32'h26a8cacf;
    ram_cell[   13519] = 32'h0;  // 32'h229894b4;
    ram_cell[   13520] = 32'h0;  // 32'h1019163b;
    ram_cell[   13521] = 32'h0;  // 32'hff1bfceb;
    ram_cell[   13522] = 32'h0;  // 32'hef42e970;
    ram_cell[   13523] = 32'h0;  // 32'he2801365;
    ram_cell[   13524] = 32'h0;  // 32'h45f3c7a9;
    ram_cell[   13525] = 32'h0;  // 32'hf84d641c;
    ram_cell[   13526] = 32'h0;  // 32'h6d95b830;
    ram_cell[   13527] = 32'h0;  // 32'h101c2181;
    ram_cell[   13528] = 32'h0;  // 32'h03378c12;
    ram_cell[   13529] = 32'h0;  // 32'h789ed872;
    ram_cell[   13530] = 32'h0;  // 32'hbee77564;
    ram_cell[   13531] = 32'h0;  // 32'he851d45c;
    ram_cell[   13532] = 32'h0;  // 32'hb3ab778d;
    ram_cell[   13533] = 32'h0;  // 32'h1592bf28;
    ram_cell[   13534] = 32'h0;  // 32'h4d504989;
    ram_cell[   13535] = 32'h0;  // 32'h54f7331d;
    ram_cell[   13536] = 32'h0;  // 32'h79e5a0fe;
    ram_cell[   13537] = 32'h0;  // 32'ha28b249b;
    ram_cell[   13538] = 32'h0;  // 32'h1686d029;
    ram_cell[   13539] = 32'h0;  // 32'h82e63ae3;
    ram_cell[   13540] = 32'h0;  // 32'h2d962cea;
    ram_cell[   13541] = 32'h0;  // 32'hefaddd24;
    ram_cell[   13542] = 32'h0;  // 32'h1efa8640;
    ram_cell[   13543] = 32'h0;  // 32'h036cbe9c;
    ram_cell[   13544] = 32'h0;  // 32'hd1741280;
    ram_cell[   13545] = 32'h0;  // 32'hfb4f76a1;
    ram_cell[   13546] = 32'h0;  // 32'hb65fdf83;
    ram_cell[   13547] = 32'h0;  // 32'heaa44674;
    ram_cell[   13548] = 32'h0;  // 32'h54b92dd0;
    ram_cell[   13549] = 32'h0;  // 32'h2d339694;
    ram_cell[   13550] = 32'h0;  // 32'h3b932b87;
    ram_cell[   13551] = 32'h0;  // 32'h672e5eba;
    ram_cell[   13552] = 32'h0;  // 32'h88b729c1;
    ram_cell[   13553] = 32'h0;  // 32'h770aeb53;
    ram_cell[   13554] = 32'h0;  // 32'h50b2dd97;
    ram_cell[   13555] = 32'h0;  // 32'ha79212f7;
    ram_cell[   13556] = 32'h0;  // 32'h9477122e;
    ram_cell[   13557] = 32'h0;  // 32'hcac15a35;
    ram_cell[   13558] = 32'h0;  // 32'h1160b2d8;
    ram_cell[   13559] = 32'h0;  // 32'h1dd7c6f3;
    ram_cell[   13560] = 32'h0;  // 32'hcae416d7;
    ram_cell[   13561] = 32'h0;  // 32'h3cae3859;
    ram_cell[   13562] = 32'h0;  // 32'h49b27365;
    ram_cell[   13563] = 32'h0;  // 32'hccc952ad;
    ram_cell[   13564] = 32'h0;  // 32'hb3f7b826;
    ram_cell[   13565] = 32'h0;  // 32'h3060b99d;
    ram_cell[   13566] = 32'h0;  // 32'h060d311a;
    ram_cell[   13567] = 32'h0;  // 32'ha88bffb7;
    ram_cell[   13568] = 32'h0;  // 32'hbbc0723d;
    ram_cell[   13569] = 32'h0;  // 32'h95590a4c;
    ram_cell[   13570] = 32'h0;  // 32'h1f549915;
    ram_cell[   13571] = 32'h0;  // 32'hcbae9d3e;
    ram_cell[   13572] = 32'h0;  // 32'h148f3e09;
    ram_cell[   13573] = 32'h0;  // 32'h1aacdaae;
    ram_cell[   13574] = 32'h0;  // 32'hecf0729c;
    ram_cell[   13575] = 32'h0;  // 32'hdc9bf958;
    ram_cell[   13576] = 32'h0;  // 32'hf7b896b4;
    ram_cell[   13577] = 32'h0;  // 32'h5f6eedcd;
    ram_cell[   13578] = 32'h0;  // 32'h52d42f36;
    ram_cell[   13579] = 32'h0;  // 32'h0fb72e3d;
    ram_cell[   13580] = 32'h0;  // 32'h7cd9f495;
    ram_cell[   13581] = 32'h0;  // 32'he8ca95a5;
    ram_cell[   13582] = 32'h0;  // 32'h3315d78c;
    ram_cell[   13583] = 32'h0;  // 32'hba4456ee;
    ram_cell[   13584] = 32'h0;  // 32'h9f67b203;
    ram_cell[   13585] = 32'h0;  // 32'h718d19b8;
    ram_cell[   13586] = 32'h0;  // 32'hd3a9b7e2;
    ram_cell[   13587] = 32'h0;  // 32'h037037d6;
    ram_cell[   13588] = 32'h0;  // 32'h7ec8b68a;
    ram_cell[   13589] = 32'h0;  // 32'hf89047c9;
    ram_cell[   13590] = 32'h0;  // 32'h558d3ae1;
    ram_cell[   13591] = 32'h0;  // 32'h476601fc;
    ram_cell[   13592] = 32'h0;  // 32'hccad5832;
    ram_cell[   13593] = 32'h0;  // 32'h23618914;
    ram_cell[   13594] = 32'h0;  // 32'h8f970cc6;
    ram_cell[   13595] = 32'h0;  // 32'hb8118ca9;
    ram_cell[   13596] = 32'h0;  // 32'h25447c86;
    ram_cell[   13597] = 32'h0;  // 32'h9af3e907;
    ram_cell[   13598] = 32'h0;  // 32'h87060033;
    ram_cell[   13599] = 32'h0;  // 32'h3d869f62;
    ram_cell[   13600] = 32'h0;  // 32'h800b76b7;
    ram_cell[   13601] = 32'h0;  // 32'h55b7ba1e;
    ram_cell[   13602] = 32'h0;  // 32'h07e1328c;
    ram_cell[   13603] = 32'h0;  // 32'h4f956463;
    ram_cell[   13604] = 32'h0;  // 32'hbe1acd3b;
    ram_cell[   13605] = 32'h0;  // 32'h5db9511d;
    ram_cell[   13606] = 32'h0;  // 32'h8582089d;
    ram_cell[   13607] = 32'h0;  // 32'h507a1177;
    ram_cell[   13608] = 32'h0;  // 32'h5969f46f;
    ram_cell[   13609] = 32'h0;  // 32'h690a5035;
    ram_cell[   13610] = 32'h0;  // 32'h65ffa2ae;
    ram_cell[   13611] = 32'h0;  // 32'ha5b700ce;
    ram_cell[   13612] = 32'h0;  // 32'h68e8584d;
    ram_cell[   13613] = 32'h0;  // 32'h46c1212a;
    ram_cell[   13614] = 32'h0;  // 32'h0a3f3482;
    ram_cell[   13615] = 32'h0;  // 32'h539a8ee7;
    ram_cell[   13616] = 32'h0;  // 32'h1b523973;
    ram_cell[   13617] = 32'h0;  // 32'hb2f4f517;
    ram_cell[   13618] = 32'h0;  // 32'h883c88a9;
    ram_cell[   13619] = 32'h0;  // 32'hf486a762;
    ram_cell[   13620] = 32'h0;  // 32'h2103a9d6;
    ram_cell[   13621] = 32'h0;  // 32'h62b34d7f;
    ram_cell[   13622] = 32'h0;  // 32'h62fd88a8;
    ram_cell[   13623] = 32'h0;  // 32'h57ad1f8a;
    ram_cell[   13624] = 32'h0;  // 32'h45177509;
    ram_cell[   13625] = 32'h0;  // 32'h0b270b07;
    ram_cell[   13626] = 32'h0;  // 32'h6e65a14b;
    ram_cell[   13627] = 32'h0;  // 32'h025731a5;
    ram_cell[   13628] = 32'h0;  // 32'h21d7e6ca;
    ram_cell[   13629] = 32'h0;  // 32'hc04690b3;
    ram_cell[   13630] = 32'h0;  // 32'h4c3b9579;
    ram_cell[   13631] = 32'h0;  // 32'h0aa45e66;
    ram_cell[   13632] = 32'h0;  // 32'h78307eee;
    ram_cell[   13633] = 32'h0;  // 32'h4a56d237;
    ram_cell[   13634] = 32'h0;  // 32'heff17571;
    ram_cell[   13635] = 32'h0;  // 32'hc8d12d91;
    ram_cell[   13636] = 32'h0;  // 32'hc522ad73;
    ram_cell[   13637] = 32'h0;  // 32'h6da57705;
    ram_cell[   13638] = 32'h0;  // 32'h5aedab34;
    ram_cell[   13639] = 32'h0;  // 32'hb4599bb9;
    ram_cell[   13640] = 32'h0;  // 32'h5aac1aa8;
    ram_cell[   13641] = 32'h0;  // 32'h66608665;
    ram_cell[   13642] = 32'h0;  // 32'hea6b3675;
    ram_cell[   13643] = 32'h0;  // 32'h7cac336f;
    ram_cell[   13644] = 32'h0;  // 32'h35338eac;
    ram_cell[   13645] = 32'h0;  // 32'h92383658;
    ram_cell[   13646] = 32'h0;  // 32'ha30d3b2e;
    ram_cell[   13647] = 32'h0;  // 32'h82f21963;
    ram_cell[   13648] = 32'h0;  // 32'h2025ffab;
    ram_cell[   13649] = 32'h0;  // 32'h3078c25d;
    ram_cell[   13650] = 32'h0;  // 32'h2a3d5d22;
    ram_cell[   13651] = 32'h0;  // 32'h8ed13723;
    ram_cell[   13652] = 32'h0;  // 32'hac4b0105;
    ram_cell[   13653] = 32'h0;  // 32'he6e2fd7b;
    ram_cell[   13654] = 32'h0;  // 32'h849488ea;
    ram_cell[   13655] = 32'h0;  // 32'hb05b110f;
    ram_cell[   13656] = 32'h0;  // 32'ha56ba017;
    ram_cell[   13657] = 32'h0;  // 32'h6d871c81;
    ram_cell[   13658] = 32'h0;  // 32'h5f54ec1f;
    ram_cell[   13659] = 32'h0;  // 32'ha4899ebd;
    ram_cell[   13660] = 32'h0;  // 32'ha37f7d97;
    ram_cell[   13661] = 32'h0;  // 32'h76f9d765;
    ram_cell[   13662] = 32'h0;  // 32'h440ccf63;
    ram_cell[   13663] = 32'h0;  // 32'h9bd2c741;
    ram_cell[   13664] = 32'h0;  // 32'hc5105ded;
    ram_cell[   13665] = 32'h0;  // 32'he51b39ee;
    ram_cell[   13666] = 32'h0;  // 32'hc4d399b5;
    ram_cell[   13667] = 32'h0;  // 32'hee3c584e;
    ram_cell[   13668] = 32'h0;  // 32'he242c455;
    ram_cell[   13669] = 32'h0;  // 32'h09b57ecf;
    ram_cell[   13670] = 32'h0;  // 32'h6c3a699e;
    ram_cell[   13671] = 32'h0;  // 32'hc04ba54d;
    ram_cell[   13672] = 32'h0;  // 32'hb59f734b;
    ram_cell[   13673] = 32'h0;  // 32'h03c32fba;
    ram_cell[   13674] = 32'h0;  // 32'hc55b8040;
    ram_cell[   13675] = 32'h0;  // 32'ha54a39c6;
    ram_cell[   13676] = 32'h0;  // 32'hb6dbc845;
    ram_cell[   13677] = 32'h0;  // 32'hcaddc39e;
    ram_cell[   13678] = 32'h0;  // 32'h033df875;
    ram_cell[   13679] = 32'h0;  // 32'h83dc97cb;
    ram_cell[   13680] = 32'h0;  // 32'ha7cd08cb;
    ram_cell[   13681] = 32'h0;  // 32'h86f48cde;
    ram_cell[   13682] = 32'h0;  // 32'h2f259ce6;
    ram_cell[   13683] = 32'h0;  // 32'h229466bf;
    ram_cell[   13684] = 32'h0;  // 32'hd17c7e74;
    ram_cell[   13685] = 32'h0;  // 32'h2adf4fd0;
    ram_cell[   13686] = 32'h0;  // 32'he6dfa2dc;
    ram_cell[   13687] = 32'h0;  // 32'hdc3236ac;
    ram_cell[   13688] = 32'h0;  // 32'h750b0c90;
    ram_cell[   13689] = 32'h0;  // 32'h26cb91d0;
    ram_cell[   13690] = 32'h0;  // 32'h8b124a90;
    ram_cell[   13691] = 32'h0;  // 32'he4f5d553;
    ram_cell[   13692] = 32'h0;  // 32'h8b04fb97;
    ram_cell[   13693] = 32'h0;  // 32'hb69b7f94;
    ram_cell[   13694] = 32'h0;  // 32'h08befa75;
    ram_cell[   13695] = 32'h0;  // 32'h46e551f5;
    ram_cell[   13696] = 32'h0;  // 32'h535f85fe;
    ram_cell[   13697] = 32'h0;  // 32'h43705ee6;
    ram_cell[   13698] = 32'h0;  // 32'hf47a0f1f;
    ram_cell[   13699] = 32'h0;  // 32'h40de0882;
    ram_cell[   13700] = 32'h0;  // 32'h1949ea83;
    ram_cell[   13701] = 32'h0;  // 32'hd191b47a;
    ram_cell[   13702] = 32'h0;  // 32'h378ce1b3;
    ram_cell[   13703] = 32'h0;  // 32'hdf7e351b;
    ram_cell[   13704] = 32'h0;  // 32'h6d5ef67b;
    ram_cell[   13705] = 32'h0;  // 32'he97ad3cb;
    ram_cell[   13706] = 32'h0;  // 32'h19a742b5;
    ram_cell[   13707] = 32'h0;  // 32'hd1085761;
    ram_cell[   13708] = 32'h0;  // 32'hb3085bc5;
    ram_cell[   13709] = 32'h0;  // 32'ha521a6bd;
    ram_cell[   13710] = 32'h0;  // 32'hf7fe7c1a;
    ram_cell[   13711] = 32'h0;  // 32'h26822461;
    ram_cell[   13712] = 32'h0;  // 32'ha93900c7;
    ram_cell[   13713] = 32'h0;  // 32'h8ae5e457;
    ram_cell[   13714] = 32'h0;  // 32'h4994aea7;
    ram_cell[   13715] = 32'h0;  // 32'hc7827bf6;
    ram_cell[   13716] = 32'h0;  // 32'h0de6dcd3;
    ram_cell[   13717] = 32'h0;  // 32'hf13a220f;
    ram_cell[   13718] = 32'h0;  // 32'h498068ec;
    ram_cell[   13719] = 32'h0;  // 32'h80830afc;
    ram_cell[   13720] = 32'h0;  // 32'h20fc0e25;
    ram_cell[   13721] = 32'h0;  // 32'h5dbed792;
    ram_cell[   13722] = 32'h0;  // 32'h122b90f2;
    ram_cell[   13723] = 32'h0;  // 32'h5712b74b;
    ram_cell[   13724] = 32'h0;  // 32'h15ab2c0c;
    ram_cell[   13725] = 32'h0;  // 32'h56fc9732;
    ram_cell[   13726] = 32'h0;  // 32'h9fe1f0d3;
    ram_cell[   13727] = 32'h0;  // 32'hf406f3a6;
    ram_cell[   13728] = 32'h0;  // 32'h47980da1;
    ram_cell[   13729] = 32'h0;  // 32'h4364534e;
    ram_cell[   13730] = 32'h0;  // 32'h1847a748;
    ram_cell[   13731] = 32'h0;  // 32'h3a5d823b;
    ram_cell[   13732] = 32'h0;  // 32'ha8c0f26b;
    ram_cell[   13733] = 32'h0;  // 32'he3fb7c5e;
    ram_cell[   13734] = 32'h0;  // 32'hf1e50859;
    ram_cell[   13735] = 32'h0;  // 32'h29f2cb34;
    ram_cell[   13736] = 32'h0;  // 32'hade1b8a9;
    ram_cell[   13737] = 32'h0;  // 32'h0f2a14eb;
    ram_cell[   13738] = 32'h0;  // 32'h10b0931b;
    ram_cell[   13739] = 32'h0;  // 32'h7482d076;
    ram_cell[   13740] = 32'h0;  // 32'h13236110;
    ram_cell[   13741] = 32'h0;  // 32'h128f3db1;
    ram_cell[   13742] = 32'h0;  // 32'ha2344e4f;
    ram_cell[   13743] = 32'h0;  // 32'h5145a5c7;
    ram_cell[   13744] = 32'h0;  // 32'h405b5561;
    ram_cell[   13745] = 32'h0;  // 32'haa515d88;
    ram_cell[   13746] = 32'h0;  // 32'h32c4bb7e;
    ram_cell[   13747] = 32'h0;  // 32'hea946091;
    ram_cell[   13748] = 32'h0;  // 32'h5baa2c5c;
    ram_cell[   13749] = 32'h0;  // 32'he38b756f;
    ram_cell[   13750] = 32'h0;  // 32'h78a21884;
    ram_cell[   13751] = 32'h0;  // 32'h0f95cef0;
    ram_cell[   13752] = 32'h0;  // 32'h67947d02;
    ram_cell[   13753] = 32'h0;  // 32'h6fcc189d;
    ram_cell[   13754] = 32'h0;  // 32'hc8854640;
    ram_cell[   13755] = 32'h0;  // 32'h85ca5068;
    ram_cell[   13756] = 32'h0;  // 32'h791fc138;
    ram_cell[   13757] = 32'h0;  // 32'hd9674d2e;
    ram_cell[   13758] = 32'h0;  // 32'h8c5af9d0;
    ram_cell[   13759] = 32'h0;  // 32'hc5a5201a;
    ram_cell[   13760] = 32'h0;  // 32'h626563bc;
    ram_cell[   13761] = 32'h0;  // 32'hd82da0de;
    ram_cell[   13762] = 32'h0;  // 32'h8204fc1e;
    ram_cell[   13763] = 32'h0;  // 32'h11d74499;
    ram_cell[   13764] = 32'h0;  // 32'hb40eb881;
    ram_cell[   13765] = 32'h0;  // 32'hcefe91ea;
    ram_cell[   13766] = 32'h0;  // 32'hb53a2f4f;
    ram_cell[   13767] = 32'h0;  // 32'h283db3bd;
    ram_cell[   13768] = 32'h0;  // 32'h19cf7dfa;
    ram_cell[   13769] = 32'h0;  // 32'hd574ad73;
    ram_cell[   13770] = 32'h0;  // 32'hcb62313b;
    ram_cell[   13771] = 32'h0;  // 32'hc92131c9;
    ram_cell[   13772] = 32'h0;  // 32'h9645ec40;
    ram_cell[   13773] = 32'h0;  // 32'hc007c09c;
    ram_cell[   13774] = 32'h0;  // 32'ha0f9890b;
    ram_cell[   13775] = 32'h0;  // 32'h324dbe29;
    ram_cell[   13776] = 32'h0;  // 32'heba8995e;
    ram_cell[   13777] = 32'h0;  // 32'hd40230db;
    ram_cell[   13778] = 32'h0;  // 32'h2b4d0e50;
    ram_cell[   13779] = 32'h0;  // 32'he8107d75;
    ram_cell[   13780] = 32'h0;  // 32'h7bf4bb50;
    ram_cell[   13781] = 32'h0;  // 32'heb5c4271;
    ram_cell[   13782] = 32'h0;  // 32'h227b5b78;
    ram_cell[   13783] = 32'h0;  // 32'hed4b6134;
    ram_cell[   13784] = 32'h0;  // 32'h9f5cfaf5;
    ram_cell[   13785] = 32'h0;  // 32'h24123547;
    ram_cell[   13786] = 32'h0;  // 32'ha75ebbad;
    ram_cell[   13787] = 32'h0;  // 32'h95895014;
    ram_cell[   13788] = 32'h0;  // 32'h897c71b2;
    ram_cell[   13789] = 32'h0;  // 32'hf3cf8120;
    ram_cell[   13790] = 32'h0;  // 32'he13a02a4;
    ram_cell[   13791] = 32'h0;  // 32'hc1c156f0;
    ram_cell[   13792] = 32'h0;  // 32'h6043f57e;
    ram_cell[   13793] = 32'h0;  // 32'hf46107c5;
    ram_cell[   13794] = 32'h0;  // 32'ha9982c34;
    ram_cell[   13795] = 32'h0;  // 32'hb0613e93;
    ram_cell[   13796] = 32'h0;  // 32'h83e06a5e;
    ram_cell[   13797] = 32'h0;  // 32'h815c216c;
    ram_cell[   13798] = 32'h0;  // 32'h65363ee9;
    ram_cell[   13799] = 32'h0;  // 32'hd6398557;
    ram_cell[   13800] = 32'h0;  // 32'h27278a1c;
    ram_cell[   13801] = 32'h0;  // 32'hf252447d;
    ram_cell[   13802] = 32'h0;  // 32'hf67cd4b3;
    ram_cell[   13803] = 32'h0;  // 32'h3f828d92;
    ram_cell[   13804] = 32'h0;  // 32'hcf42bd13;
    ram_cell[   13805] = 32'h0;  // 32'h79807050;
    ram_cell[   13806] = 32'h0;  // 32'h5273d073;
    ram_cell[   13807] = 32'h0;  // 32'h6259be5a;
    ram_cell[   13808] = 32'h0;  // 32'h7ac38a99;
    ram_cell[   13809] = 32'h0;  // 32'hde90ebf1;
    ram_cell[   13810] = 32'h0;  // 32'hb727f653;
    ram_cell[   13811] = 32'h0;  // 32'h05d9e89e;
    ram_cell[   13812] = 32'h0;  // 32'hd1322779;
    ram_cell[   13813] = 32'h0;  // 32'he12a341f;
    ram_cell[   13814] = 32'h0;  // 32'hb2b0f1db;
    ram_cell[   13815] = 32'h0;  // 32'ha2a5d175;
    ram_cell[   13816] = 32'h0;  // 32'h5ca1a490;
    ram_cell[   13817] = 32'h0;  // 32'h87a8b21e;
    ram_cell[   13818] = 32'h0;  // 32'h5760d92b;
    ram_cell[   13819] = 32'h0;  // 32'h6a9de057;
    ram_cell[   13820] = 32'h0;  // 32'h90e4332c;
    ram_cell[   13821] = 32'h0;  // 32'h74e1c584;
    ram_cell[   13822] = 32'h0;  // 32'h9644509c;
    ram_cell[   13823] = 32'h0;  // 32'hd585b563;
    ram_cell[   13824] = 32'h0;  // 32'h811aa342;
    ram_cell[   13825] = 32'h0;  // 32'hdd44c87f;
    ram_cell[   13826] = 32'h0;  // 32'h22ddeef2;
    ram_cell[   13827] = 32'h0;  // 32'ha705c263;
    ram_cell[   13828] = 32'h0;  // 32'hee5866ce;
    ram_cell[   13829] = 32'h0;  // 32'he3e1c8ef;
    ram_cell[   13830] = 32'h0;  // 32'h324513fc;
    ram_cell[   13831] = 32'h0;  // 32'h72531cb1;
    ram_cell[   13832] = 32'h0;  // 32'h2816e0c3;
    ram_cell[   13833] = 32'h0;  // 32'h9115f990;
    ram_cell[   13834] = 32'h0;  // 32'hca52dabd;
    ram_cell[   13835] = 32'h0;  // 32'hc1dcf8ed;
    ram_cell[   13836] = 32'h0;  // 32'h148a08a8;
    ram_cell[   13837] = 32'h0;  // 32'h017de5b4;
    ram_cell[   13838] = 32'h0;  // 32'he71748c5;
    ram_cell[   13839] = 32'h0;  // 32'h63544104;
    ram_cell[   13840] = 32'h0;  // 32'h77b1fe36;
    ram_cell[   13841] = 32'h0;  // 32'h2615c9eb;
    ram_cell[   13842] = 32'h0;  // 32'hc3bd76bf;
    ram_cell[   13843] = 32'h0;  // 32'h679b9659;
    ram_cell[   13844] = 32'h0;  // 32'h199b883c;
    ram_cell[   13845] = 32'h0;  // 32'h712ea15e;
    ram_cell[   13846] = 32'h0;  // 32'hab4c5b85;
    ram_cell[   13847] = 32'h0;  // 32'h79a0134d;
    ram_cell[   13848] = 32'h0;  // 32'h81b5b1f1;
    ram_cell[   13849] = 32'h0;  // 32'ha5720454;
    ram_cell[   13850] = 32'h0;  // 32'he333efcc;
    ram_cell[   13851] = 32'h0;  // 32'h26b90594;
    ram_cell[   13852] = 32'h0;  // 32'h5184a6ed;
    ram_cell[   13853] = 32'h0;  // 32'h66a4ff96;
    ram_cell[   13854] = 32'h0;  // 32'hea825d8a;
    ram_cell[   13855] = 32'h0;  // 32'hf192872e;
    ram_cell[   13856] = 32'h0;  // 32'h7113a7f6;
    ram_cell[   13857] = 32'h0;  // 32'h82ede44d;
    ram_cell[   13858] = 32'h0;  // 32'h6d3318dd;
    ram_cell[   13859] = 32'h0;  // 32'he3075411;
    ram_cell[   13860] = 32'h0;  // 32'h20d9a700;
    ram_cell[   13861] = 32'h0;  // 32'ha24e9530;
    ram_cell[   13862] = 32'h0;  // 32'h0119c931;
    ram_cell[   13863] = 32'h0;  // 32'hbfe833a5;
    ram_cell[   13864] = 32'h0;  // 32'ha4d83f37;
    ram_cell[   13865] = 32'h0;  // 32'h8d2bda6b;
    ram_cell[   13866] = 32'h0;  // 32'h1e8ddb51;
    ram_cell[   13867] = 32'h0;  // 32'h2161010f;
    ram_cell[   13868] = 32'h0;  // 32'hc5e4c19f;
    ram_cell[   13869] = 32'h0;  // 32'h32735944;
    ram_cell[   13870] = 32'h0;  // 32'he1ceead4;
    ram_cell[   13871] = 32'h0;  // 32'heeaefe92;
    ram_cell[   13872] = 32'h0;  // 32'he34cacd9;
    ram_cell[   13873] = 32'h0;  // 32'h3094e964;
    ram_cell[   13874] = 32'h0;  // 32'h319cf4cd;
    ram_cell[   13875] = 32'h0;  // 32'h6bbcd332;
    ram_cell[   13876] = 32'h0;  // 32'hef321cb8;
    ram_cell[   13877] = 32'h0;  // 32'h906fe85d;
    ram_cell[   13878] = 32'h0;  // 32'h2f7ff9ea;
    ram_cell[   13879] = 32'h0;  // 32'hf178127b;
    ram_cell[   13880] = 32'h0;  // 32'heb0bb696;
    ram_cell[   13881] = 32'h0;  // 32'h3ef62079;
    ram_cell[   13882] = 32'h0;  // 32'h5569f3af;
    ram_cell[   13883] = 32'h0;  // 32'h852e4ac3;
    ram_cell[   13884] = 32'h0;  // 32'he1dd77a4;
    ram_cell[   13885] = 32'h0;  // 32'he18ca36d;
    ram_cell[   13886] = 32'h0;  // 32'h8454c3b0;
    ram_cell[   13887] = 32'h0;  // 32'hd4b3cc8e;
    ram_cell[   13888] = 32'h0;  // 32'haeb931d1;
    ram_cell[   13889] = 32'h0;  // 32'hbdbc3e93;
    ram_cell[   13890] = 32'h0;  // 32'h46e629df;
    ram_cell[   13891] = 32'h0;  // 32'hd7591dc6;
    ram_cell[   13892] = 32'h0;  // 32'h9abd1cd2;
    ram_cell[   13893] = 32'h0;  // 32'h723a2c95;
    ram_cell[   13894] = 32'h0;  // 32'h2c36e728;
    ram_cell[   13895] = 32'h0;  // 32'ha136de90;
    ram_cell[   13896] = 32'h0;  // 32'h94cdb1f1;
    ram_cell[   13897] = 32'h0;  // 32'h56772910;
    ram_cell[   13898] = 32'h0;  // 32'h4b1e7729;
    ram_cell[   13899] = 32'h0;  // 32'h1f0006f6;
    ram_cell[   13900] = 32'h0;  // 32'h5ec07431;
    ram_cell[   13901] = 32'h0;  // 32'hb2d8188c;
    ram_cell[   13902] = 32'h0;  // 32'h5575e49b;
    ram_cell[   13903] = 32'h0;  // 32'h57f00b9a;
    ram_cell[   13904] = 32'h0;  // 32'hc5e9fccb;
    ram_cell[   13905] = 32'h0;  // 32'h43b5939a;
    ram_cell[   13906] = 32'h0;  // 32'h45cc597a;
    ram_cell[   13907] = 32'h0;  // 32'ha2d0fa5f;
    ram_cell[   13908] = 32'h0;  // 32'h23b9b0ca;
    ram_cell[   13909] = 32'h0;  // 32'h6bcf38e5;
    ram_cell[   13910] = 32'h0;  // 32'h96ce6282;
    ram_cell[   13911] = 32'h0;  // 32'h0071e1ab;
    ram_cell[   13912] = 32'h0;  // 32'h20fef192;
    ram_cell[   13913] = 32'h0;  // 32'h6f2f5424;
    ram_cell[   13914] = 32'h0;  // 32'h16ab6acc;
    ram_cell[   13915] = 32'h0;  // 32'hf2807951;
    ram_cell[   13916] = 32'h0;  // 32'h2ea1af1a;
    ram_cell[   13917] = 32'h0;  // 32'h8fa61453;
    ram_cell[   13918] = 32'h0;  // 32'hd767030a;
    ram_cell[   13919] = 32'h0;  // 32'h6cf92ffa;
    ram_cell[   13920] = 32'h0;  // 32'hdd60adfe;
    ram_cell[   13921] = 32'h0;  // 32'hed1729c3;
    ram_cell[   13922] = 32'h0;  // 32'hb6471881;
    ram_cell[   13923] = 32'h0;  // 32'h7aa4bc35;
    ram_cell[   13924] = 32'h0;  // 32'hd80d5688;
    ram_cell[   13925] = 32'h0;  // 32'hd9e9569b;
    ram_cell[   13926] = 32'h0;  // 32'hb35287b7;
    ram_cell[   13927] = 32'h0;  // 32'h3c694a29;
    ram_cell[   13928] = 32'h0;  // 32'hfb55ec04;
    ram_cell[   13929] = 32'h0;  // 32'h033335e7;
    ram_cell[   13930] = 32'h0;  // 32'h7aa1b957;
    ram_cell[   13931] = 32'h0;  // 32'hce9eb573;
    ram_cell[   13932] = 32'h0;  // 32'hae9f2efe;
    ram_cell[   13933] = 32'h0;  // 32'hb9bd420c;
    ram_cell[   13934] = 32'h0;  // 32'h67a7653b;
    ram_cell[   13935] = 32'h0;  // 32'hf8f0a3af;
    ram_cell[   13936] = 32'h0;  // 32'h28fac9da;
    ram_cell[   13937] = 32'h0;  // 32'hbfbed640;
    ram_cell[   13938] = 32'h0;  // 32'h58e3560b;
    ram_cell[   13939] = 32'h0;  // 32'haaedbbe2;
    ram_cell[   13940] = 32'h0;  // 32'h88ae4dbb;
    ram_cell[   13941] = 32'h0;  // 32'h20b76e38;
    ram_cell[   13942] = 32'h0;  // 32'hb3784a0e;
    ram_cell[   13943] = 32'h0;  // 32'h8c517ffd;
    ram_cell[   13944] = 32'h0;  // 32'h2fb38631;
    ram_cell[   13945] = 32'h0;  // 32'h78525dce;
    ram_cell[   13946] = 32'h0;  // 32'h272da7df;
    ram_cell[   13947] = 32'h0;  // 32'h4e156986;
    ram_cell[   13948] = 32'h0;  // 32'he852619e;
    ram_cell[   13949] = 32'h0;  // 32'h8a4729c8;
    ram_cell[   13950] = 32'h0;  // 32'h47588a3d;
    ram_cell[   13951] = 32'h0;  // 32'hda4a4659;
    ram_cell[   13952] = 32'h0;  // 32'hd021b26e;
    ram_cell[   13953] = 32'h0;  // 32'hb88ff851;
    ram_cell[   13954] = 32'h0;  // 32'he8722028;
    ram_cell[   13955] = 32'h0;  // 32'h79a5c3d0;
    ram_cell[   13956] = 32'h0;  // 32'hb7717990;
    ram_cell[   13957] = 32'h0;  // 32'h54393b97;
    ram_cell[   13958] = 32'h0;  // 32'h0cfb083d;
    ram_cell[   13959] = 32'h0;  // 32'hedad595a;
    ram_cell[   13960] = 32'h0;  // 32'h425ce727;
    ram_cell[   13961] = 32'h0;  // 32'hdbbad502;
    ram_cell[   13962] = 32'h0;  // 32'h55782459;
    ram_cell[   13963] = 32'h0;  // 32'hdfb5d36a;
    ram_cell[   13964] = 32'h0;  // 32'h55cb1db3;
    ram_cell[   13965] = 32'h0;  // 32'hd1c7dc3f;
    ram_cell[   13966] = 32'h0;  // 32'h4f84905c;
    ram_cell[   13967] = 32'h0;  // 32'h91b7015b;
    ram_cell[   13968] = 32'h0;  // 32'h7f256917;
    ram_cell[   13969] = 32'h0;  // 32'hf6bdd095;
    ram_cell[   13970] = 32'h0;  // 32'h8dbf257e;
    ram_cell[   13971] = 32'h0;  // 32'h6e7c3fad;
    ram_cell[   13972] = 32'h0;  // 32'hcb269fe7;
    ram_cell[   13973] = 32'h0;  // 32'h79166146;
    ram_cell[   13974] = 32'h0;  // 32'h862107a0;
    ram_cell[   13975] = 32'h0;  // 32'h77b4d3c6;
    ram_cell[   13976] = 32'h0;  // 32'hf16edecb;
    ram_cell[   13977] = 32'h0;  // 32'h4c6e3650;
    ram_cell[   13978] = 32'h0;  // 32'h3407240d;
    ram_cell[   13979] = 32'h0;  // 32'h5e3ad54e;
    ram_cell[   13980] = 32'h0;  // 32'h0448e73e;
    ram_cell[   13981] = 32'h0;  // 32'hd5e7da99;
    ram_cell[   13982] = 32'h0;  // 32'hc93a850c;
    ram_cell[   13983] = 32'h0;  // 32'h7180bc72;
    ram_cell[   13984] = 32'h0;  // 32'h054cd278;
    ram_cell[   13985] = 32'h0;  // 32'hfbf2a4ad;
    ram_cell[   13986] = 32'h0;  // 32'h48f0184a;
    ram_cell[   13987] = 32'h0;  // 32'ha236ebe4;
    ram_cell[   13988] = 32'h0;  // 32'h552b1332;
    ram_cell[   13989] = 32'h0;  // 32'h25b5001e;
    ram_cell[   13990] = 32'h0;  // 32'h1c9d0024;
    ram_cell[   13991] = 32'h0;  // 32'hfb955966;
    ram_cell[   13992] = 32'h0;  // 32'h15b4a574;
    ram_cell[   13993] = 32'h0;  // 32'h5ad7e5ab;
    ram_cell[   13994] = 32'h0;  // 32'hdfaaeacb;
    ram_cell[   13995] = 32'h0;  // 32'hc135c8ab;
    ram_cell[   13996] = 32'h0;  // 32'ha9e2d8dd;
    ram_cell[   13997] = 32'h0;  // 32'h47ba78b7;
    ram_cell[   13998] = 32'h0;  // 32'hcf349379;
    ram_cell[   13999] = 32'h0;  // 32'hc2219747;
    ram_cell[   14000] = 32'h0;  // 32'hc76d6ccd;
    ram_cell[   14001] = 32'h0;  // 32'hebcaf287;
    ram_cell[   14002] = 32'h0;  // 32'h5c3ce6a5;
    ram_cell[   14003] = 32'h0;  // 32'h32f08440;
    ram_cell[   14004] = 32'h0;  // 32'h145636ce;
    ram_cell[   14005] = 32'h0;  // 32'ha2d671d9;
    ram_cell[   14006] = 32'h0;  // 32'h4f371504;
    ram_cell[   14007] = 32'h0;  // 32'hf2d03218;
    ram_cell[   14008] = 32'h0;  // 32'h162e1c71;
    ram_cell[   14009] = 32'h0;  // 32'h5d94fdb2;
    ram_cell[   14010] = 32'h0;  // 32'hed5e0e4f;
    ram_cell[   14011] = 32'h0;  // 32'h307c84e6;
    ram_cell[   14012] = 32'h0;  // 32'h3f6cb439;
    ram_cell[   14013] = 32'h0;  // 32'h379f8053;
    ram_cell[   14014] = 32'h0;  // 32'h749540f6;
    ram_cell[   14015] = 32'h0;  // 32'h85701fb5;
    ram_cell[   14016] = 32'h0;  // 32'h4511ebce;
    ram_cell[   14017] = 32'h0;  // 32'h96b99754;
    ram_cell[   14018] = 32'h0;  // 32'h6fae1e10;
    ram_cell[   14019] = 32'h0;  // 32'hf736880f;
    ram_cell[   14020] = 32'h0;  // 32'h6b67c876;
    ram_cell[   14021] = 32'h0;  // 32'h2c881ed2;
    ram_cell[   14022] = 32'h0;  // 32'h363de5af;
    ram_cell[   14023] = 32'h0;  // 32'hd87523ee;
    ram_cell[   14024] = 32'h0;  // 32'h21292474;
    ram_cell[   14025] = 32'h0;  // 32'ha7ee391e;
    ram_cell[   14026] = 32'h0;  // 32'h6217cccc;
    ram_cell[   14027] = 32'h0;  // 32'h1f3a407c;
    ram_cell[   14028] = 32'h0;  // 32'h32f06f87;
    ram_cell[   14029] = 32'h0;  // 32'h8b978176;
    ram_cell[   14030] = 32'h0;  // 32'h9ffc7c57;
    ram_cell[   14031] = 32'h0;  // 32'hdc100c9e;
    ram_cell[   14032] = 32'h0;  // 32'h379949b5;
    ram_cell[   14033] = 32'h0;  // 32'he79092cc;
    ram_cell[   14034] = 32'h0;  // 32'haf6052b3;
    ram_cell[   14035] = 32'h0;  // 32'h64a11dab;
    ram_cell[   14036] = 32'h0;  // 32'h0273d128;
    ram_cell[   14037] = 32'h0;  // 32'h3259b172;
    ram_cell[   14038] = 32'h0;  // 32'hd0df9940;
    ram_cell[   14039] = 32'h0;  // 32'h14994162;
    ram_cell[   14040] = 32'h0;  // 32'h23dc1419;
    ram_cell[   14041] = 32'h0;  // 32'h2afa0793;
    ram_cell[   14042] = 32'h0;  // 32'h0ef46ad8;
    ram_cell[   14043] = 32'h0;  // 32'h53649684;
    ram_cell[   14044] = 32'h0;  // 32'h6f661100;
    ram_cell[   14045] = 32'h0;  // 32'h83646b8a;
    ram_cell[   14046] = 32'h0;  // 32'h0e1f94e1;
    ram_cell[   14047] = 32'h0;  // 32'h3f7b1f1a;
    ram_cell[   14048] = 32'h0;  // 32'h32d0393f;
    ram_cell[   14049] = 32'h0;  // 32'h77c9537e;
    ram_cell[   14050] = 32'h0;  // 32'had1f9827;
    ram_cell[   14051] = 32'h0;  // 32'h8f49e3d7;
    ram_cell[   14052] = 32'h0;  // 32'hedd4ba29;
    ram_cell[   14053] = 32'h0;  // 32'hd948734a;
    ram_cell[   14054] = 32'h0;  // 32'h2fb628b5;
    ram_cell[   14055] = 32'h0;  // 32'hd1e124f5;
    ram_cell[   14056] = 32'h0;  // 32'hda57a6d0;
    ram_cell[   14057] = 32'h0;  // 32'hdf4e9c85;
    ram_cell[   14058] = 32'h0;  // 32'hc1871915;
    ram_cell[   14059] = 32'h0;  // 32'he2c1a9eb;
    ram_cell[   14060] = 32'h0;  // 32'h5874965b;
    ram_cell[   14061] = 32'h0;  // 32'haaf862f9;
    ram_cell[   14062] = 32'h0;  // 32'hd0b84680;
    ram_cell[   14063] = 32'h0;  // 32'h7f6f73c7;
    ram_cell[   14064] = 32'h0;  // 32'h7e8b9d97;
    ram_cell[   14065] = 32'h0;  // 32'h0320c128;
    ram_cell[   14066] = 32'h0;  // 32'heee9275f;
    ram_cell[   14067] = 32'h0;  // 32'h31e4779b;
    ram_cell[   14068] = 32'h0;  // 32'h537e8598;
    ram_cell[   14069] = 32'h0;  // 32'h1665d90c;
    ram_cell[   14070] = 32'h0;  // 32'h38fb8703;
    ram_cell[   14071] = 32'h0;  // 32'had84c701;
    ram_cell[   14072] = 32'h0;  // 32'hde143069;
    ram_cell[   14073] = 32'h0;  // 32'h3e12de3a;
    ram_cell[   14074] = 32'h0;  // 32'h6f88490e;
    ram_cell[   14075] = 32'h0;  // 32'h6e4d1c39;
    ram_cell[   14076] = 32'h0;  // 32'hb1a7942e;
    ram_cell[   14077] = 32'h0;  // 32'h0794ec59;
    ram_cell[   14078] = 32'h0;  // 32'h5bef6369;
    ram_cell[   14079] = 32'h0;  // 32'h3e1a2b96;
    ram_cell[   14080] = 32'h0;  // 32'h38f8802e;
    ram_cell[   14081] = 32'h0;  // 32'ha88269cb;
    ram_cell[   14082] = 32'h0;  // 32'h29a66aec;
    ram_cell[   14083] = 32'h0;  // 32'h44ebe7f9;
    ram_cell[   14084] = 32'h0;  // 32'h2d7052fb;
    ram_cell[   14085] = 32'h0;  // 32'h28334b58;
    ram_cell[   14086] = 32'h0;  // 32'he622f563;
    ram_cell[   14087] = 32'h0;  // 32'hce8a129e;
    ram_cell[   14088] = 32'h0;  // 32'hf5eb680e;
    ram_cell[   14089] = 32'h0;  // 32'hbb2a0467;
    ram_cell[   14090] = 32'h0;  // 32'h3f349319;
    ram_cell[   14091] = 32'h0;  // 32'h70a2c1e6;
    ram_cell[   14092] = 32'h0;  // 32'h2a570ad8;
    ram_cell[   14093] = 32'h0;  // 32'hdd0846fd;
    ram_cell[   14094] = 32'h0;  // 32'h0fa5cf1c;
    ram_cell[   14095] = 32'h0;  // 32'h79f6c3ba;
    ram_cell[   14096] = 32'h0;  // 32'hacc8ff89;
    ram_cell[   14097] = 32'h0;  // 32'h4a1d04dd;
    ram_cell[   14098] = 32'h0;  // 32'hb94e90c1;
    ram_cell[   14099] = 32'h0;  // 32'hafb07ead;
    ram_cell[   14100] = 32'h0;  // 32'h4f65dbd9;
    ram_cell[   14101] = 32'h0;  // 32'h37559b2f;
    ram_cell[   14102] = 32'h0;  // 32'h8d534ece;
    ram_cell[   14103] = 32'h0;  // 32'h678333f1;
    ram_cell[   14104] = 32'h0;  // 32'h4e34627f;
    ram_cell[   14105] = 32'h0;  // 32'he44c4f94;
    ram_cell[   14106] = 32'h0;  // 32'h4b162c2e;
    ram_cell[   14107] = 32'h0;  // 32'h70453723;
    ram_cell[   14108] = 32'h0;  // 32'h642e5531;
    ram_cell[   14109] = 32'h0;  // 32'h290f1587;
    ram_cell[   14110] = 32'h0;  // 32'h09380020;
    ram_cell[   14111] = 32'h0;  // 32'ha91302ba;
    ram_cell[   14112] = 32'h0;  // 32'hf8e50f27;
    ram_cell[   14113] = 32'h0;  // 32'h4f478561;
    ram_cell[   14114] = 32'h0;  // 32'h8748f452;
    ram_cell[   14115] = 32'h0;  // 32'h7575a70d;
    ram_cell[   14116] = 32'h0;  // 32'h4ce0c156;
    ram_cell[   14117] = 32'h0;  // 32'h3adef7d2;
    ram_cell[   14118] = 32'h0;  // 32'hef6b6941;
    ram_cell[   14119] = 32'h0;  // 32'hd3a0e7bf;
    ram_cell[   14120] = 32'h0;  // 32'h9f7b273d;
    ram_cell[   14121] = 32'h0;  // 32'ha950d102;
    ram_cell[   14122] = 32'h0;  // 32'h58bbcbcb;
    ram_cell[   14123] = 32'h0;  // 32'h25f0559d;
    ram_cell[   14124] = 32'h0;  // 32'hb1129460;
    ram_cell[   14125] = 32'h0;  // 32'h9238537f;
    ram_cell[   14126] = 32'h0;  // 32'h7fd84ed7;
    ram_cell[   14127] = 32'h0;  // 32'h8bbcee48;
    ram_cell[   14128] = 32'h0;  // 32'h98ffce29;
    ram_cell[   14129] = 32'h0;  // 32'hba9016d1;
    ram_cell[   14130] = 32'h0;  // 32'h4d62445a;
    ram_cell[   14131] = 32'h0;  // 32'h48725b6a;
    ram_cell[   14132] = 32'h0;  // 32'h2501ddae;
    ram_cell[   14133] = 32'h0;  // 32'h37e7eac6;
    ram_cell[   14134] = 32'h0;  // 32'h8f315a97;
    ram_cell[   14135] = 32'h0;  // 32'hef1a0207;
    ram_cell[   14136] = 32'h0;  // 32'hf288d562;
    ram_cell[   14137] = 32'h0;  // 32'h6a449343;
    ram_cell[   14138] = 32'h0;  // 32'h4de7f7d2;
    ram_cell[   14139] = 32'h0;  // 32'h9149f480;
    ram_cell[   14140] = 32'h0;  // 32'hea38f947;
    ram_cell[   14141] = 32'h0;  // 32'h3f0800a6;
    ram_cell[   14142] = 32'h0;  // 32'hb9093234;
    ram_cell[   14143] = 32'h0;  // 32'h93c60b3d;
    ram_cell[   14144] = 32'h0;  // 32'h35d10182;
    ram_cell[   14145] = 32'h0;  // 32'hc2acb9cd;
    ram_cell[   14146] = 32'h0;  // 32'hddac238c;
    ram_cell[   14147] = 32'h0;  // 32'hf54b168a;
    ram_cell[   14148] = 32'h0;  // 32'h570c99ea;
    ram_cell[   14149] = 32'h0;  // 32'h7bb0a775;
    ram_cell[   14150] = 32'h0;  // 32'h337a3e6d;
    ram_cell[   14151] = 32'h0;  // 32'he36c88ab;
    ram_cell[   14152] = 32'h0;  // 32'h951804dd;
    ram_cell[   14153] = 32'h0;  // 32'h3dbf4ce1;
    ram_cell[   14154] = 32'h0;  // 32'h7ed71494;
    ram_cell[   14155] = 32'h0;  // 32'h1770d46a;
    ram_cell[   14156] = 32'h0;  // 32'h2a2cd1f7;
    ram_cell[   14157] = 32'h0;  // 32'hbb179a68;
    ram_cell[   14158] = 32'h0;  // 32'h5e7318b4;
    ram_cell[   14159] = 32'h0;  // 32'h86bee93e;
    ram_cell[   14160] = 32'h0;  // 32'hc106a422;
    ram_cell[   14161] = 32'h0;  // 32'h816d62b5;
    ram_cell[   14162] = 32'h0;  // 32'ha21beead;
    ram_cell[   14163] = 32'h0;  // 32'hd6c19161;
    ram_cell[   14164] = 32'h0;  // 32'h7c87053c;
    ram_cell[   14165] = 32'h0;  // 32'hc16a04a3;
    ram_cell[   14166] = 32'h0;  // 32'h9f3db49c;
    ram_cell[   14167] = 32'h0;  // 32'habcbd13d;
    ram_cell[   14168] = 32'h0;  // 32'hdc46da0a;
    ram_cell[   14169] = 32'h0;  // 32'h48c3daee;
    ram_cell[   14170] = 32'h0;  // 32'h76eca872;
    ram_cell[   14171] = 32'h0;  // 32'h5acac588;
    ram_cell[   14172] = 32'h0;  // 32'h22b317bc;
    ram_cell[   14173] = 32'h0;  // 32'he13ee553;
    ram_cell[   14174] = 32'h0;  // 32'ha92759b4;
    ram_cell[   14175] = 32'h0;  // 32'hc5c358e2;
    ram_cell[   14176] = 32'h0;  // 32'hb8b0e82c;
    ram_cell[   14177] = 32'h0;  // 32'hf7612063;
    ram_cell[   14178] = 32'h0;  // 32'hda4e7ec3;
    ram_cell[   14179] = 32'h0;  // 32'h43eacb42;
    ram_cell[   14180] = 32'h0;  // 32'h9c33b026;
    ram_cell[   14181] = 32'h0;  // 32'h9f7936cc;
    ram_cell[   14182] = 32'h0;  // 32'hf902de67;
    ram_cell[   14183] = 32'h0;  // 32'ha85c7288;
    ram_cell[   14184] = 32'h0;  // 32'h9e56d888;
    ram_cell[   14185] = 32'h0;  // 32'h2a81ea13;
    ram_cell[   14186] = 32'h0;  // 32'h68b04695;
    ram_cell[   14187] = 32'h0;  // 32'h0e11bbd8;
    ram_cell[   14188] = 32'h0;  // 32'hae2efa96;
    ram_cell[   14189] = 32'h0;  // 32'he1ed566e;
    ram_cell[   14190] = 32'h0;  // 32'h50d6f362;
    ram_cell[   14191] = 32'h0;  // 32'h71f26df3;
    ram_cell[   14192] = 32'h0;  // 32'h5e0a5631;
    ram_cell[   14193] = 32'h0;  // 32'h0356f3b1;
    ram_cell[   14194] = 32'h0;  // 32'hd1f709fe;
    ram_cell[   14195] = 32'h0;  // 32'h56af9334;
    ram_cell[   14196] = 32'h0;  // 32'h4becd581;
    ram_cell[   14197] = 32'h0;  // 32'h5100b824;
    ram_cell[   14198] = 32'h0;  // 32'h6dbddbfa;
    ram_cell[   14199] = 32'h0;  // 32'h9de1b2dc;
    ram_cell[   14200] = 32'h0;  // 32'ha5781607;
    ram_cell[   14201] = 32'h0;  // 32'h65f1f8f4;
    ram_cell[   14202] = 32'h0;  // 32'habfe2a2c;
    ram_cell[   14203] = 32'h0;  // 32'h0e9f3b68;
    ram_cell[   14204] = 32'h0;  // 32'hd5e1fa6d;
    ram_cell[   14205] = 32'h0;  // 32'hcf7fe7a4;
    ram_cell[   14206] = 32'h0;  // 32'hfc6c0170;
    ram_cell[   14207] = 32'h0;  // 32'h4fb58985;
    ram_cell[   14208] = 32'h0;  // 32'h9de706bf;
    ram_cell[   14209] = 32'h0;  // 32'h84d43d79;
    ram_cell[   14210] = 32'h0;  // 32'h12a6f19e;
    ram_cell[   14211] = 32'h0;  // 32'h22a544d7;
    ram_cell[   14212] = 32'h0;  // 32'h982635fd;
    ram_cell[   14213] = 32'h0;  // 32'h988df9df;
    ram_cell[   14214] = 32'h0;  // 32'hbde6f721;
    ram_cell[   14215] = 32'h0;  // 32'h2d7fd185;
    ram_cell[   14216] = 32'h0;  // 32'h48a2cf25;
    ram_cell[   14217] = 32'h0;  // 32'h2db513c0;
    ram_cell[   14218] = 32'h0;  // 32'h87b793fa;
    ram_cell[   14219] = 32'h0;  // 32'h42290a6c;
    ram_cell[   14220] = 32'h0;  // 32'hcbe506c0;
    ram_cell[   14221] = 32'h0;  // 32'hbb2c011a;
    ram_cell[   14222] = 32'h0;  // 32'he7ac7b25;
    ram_cell[   14223] = 32'h0;  // 32'hc2d36d66;
    ram_cell[   14224] = 32'h0;  // 32'h76a5681e;
    ram_cell[   14225] = 32'h0;  // 32'hca92181f;
    ram_cell[   14226] = 32'h0;  // 32'h967236c3;
    ram_cell[   14227] = 32'h0;  // 32'h16af68fe;
    ram_cell[   14228] = 32'h0;  // 32'h317c1fd7;
    ram_cell[   14229] = 32'h0;  // 32'h2fa7c798;
    ram_cell[   14230] = 32'h0;  // 32'h0a6f834c;
    ram_cell[   14231] = 32'h0;  // 32'hce86bdf1;
    ram_cell[   14232] = 32'h0;  // 32'h3072b2ab;
    ram_cell[   14233] = 32'h0;  // 32'h8cef0bf7;
    ram_cell[   14234] = 32'h0;  // 32'hbca57ce1;
    ram_cell[   14235] = 32'h0;  // 32'hf1023e2d;
    ram_cell[   14236] = 32'h0;  // 32'h40d681a9;
    ram_cell[   14237] = 32'h0;  // 32'hb62e757a;
    ram_cell[   14238] = 32'h0;  // 32'h870e5f9d;
    ram_cell[   14239] = 32'h0;  // 32'h752d9ba9;
    ram_cell[   14240] = 32'h0;  // 32'h577bfaba;
    ram_cell[   14241] = 32'h0;  // 32'h9d8d45d8;
    ram_cell[   14242] = 32'h0;  // 32'h457c4495;
    ram_cell[   14243] = 32'h0;  // 32'h2cd2e1f0;
    ram_cell[   14244] = 32'h0;  // 32'h6f9f1d5c;
    ram_cell[   14245] = 32'h0;  // 32'hde4bc125;
    ram_cell[   14246] = 32'h0;  // 32'hbfdd10cf;
    ram_cell[   14247] = 32'h0;  // 32'h00682b93;
    ram_cell[   14248] = 32'h0;  // 32'hfa001d6f;
    ram_cell[   14249] = 32'h0;  // 32'h274c5854;
    ram_cell[   14250] = 32'h0;  // 32'h0799f3ff;
    ram_cell[   14251] = 32'h0;  // 32'hce99cfef;
    ram_cell[   14252] = 32'h0;  // 32'h1a56eb31;
    ram_cell[   14253] = 32'h0;  // 32'h72f18b30;
    ram_cell[   14254] = 32'h0;  // 32'h734bc934;
    ram_cell[   14255] = 32'h0;  // 32'h472b800a;
    ram_cell[   14256] = 32'h0;  // 32'hcea5b21d;
    ram_cell[   14257] = 32'h0;  // 32'hc0577567;
    ram_cell[   14258] = 32'h0;  // 32'hd6a4d194;
    ram_cell[   14259] = 32'h0;  // 32'h767d3dfb;
    ram_cell[   14260] = 32'h0;  // 32'hc0703640;
    ram_cell[   14261] = 32'h0;  // 32'hdef9f701;
    ram_cell[   14262] = 32'h0;  // 32'h38720300;
    ram_cell[   14263] = 32'h0;  // 32'hb88f761e;
    ram_cell[   14264] = 32'h0;  // 32'h28c0a383;
    ram_cell[   14265] = 32'h0;  // 32'h34e45d17;
    ram_cell[   14266] = 32'h0;  // 32'h647c2fbd;
    ram_cell[   14267] = 32'h0;  // 32'hec4b28b3;
    ram_cell[   14268] = 32'h0;  // 32'ha56b85aa;
    ram_cell[   14269] = 32'h0;  // 32'hac671c66;
    ram_cell[   14270] = 32'h0;  // 32'hfdbe5ebb;
    ram_cell[   14271] = 32'h0;  // 32'h6e39a7fb;
    ram_cell[   14272] = 32'h0;  // 32'hb868f984;
    ram_cell[   14273] = 32'h0;  // 32'h713624f4;
    ram_cell[   14274] = 32'h0;  // 32'h444efec2;
    ram_cell[   14275] = 32'h0;  // 32'h83794466;
    ram_cell[   14276] = 32'h0;  // 32'h8885bb60;
    ram_cell[   14277] = 32'h0;  // 32'h3095ac83;
    ram_cell[   14278] = 32'h0;  // 32'h164dcbee;
    ram_cell[   14279] = 32'h0;  // 32'h0198a01f;
    ram_cell[   14280] = 32'h0;  // 32'hcf9f4cdd;
    ram_cell[   14281] = 32'h0;  // 32'h95f5b18b;
    ram_cell[   14282] = 32'h0;  // 32'h0046934d;
    ram_cell[   14283] = 32'h0;  // 32'he0b3766d;
    ram_cell[   14284] = 32'h0;  // 32'hb4e094a6;
    ram_cell[   14285] = 32'h0;  // 32'hf88cc40e;
    ram_cell[   14286] = 32'h0;  // 32'h7b6cca72;
    ram_cell[   14287] = 32'h0;  // 32'h2d9b97ca;
    ram_cell[   14288] = 32'h0;  // 32'hd7d5e112;
    ram_cell[   14289] = 32'h0;  // 32'h013568ff;
    ram_cell[   14290] = 32'h0;  // 32'h5df972c0;
    ram_cell[   14291] = 32'h0;  // 32'h89434668;
    ram_cell[   14292] = 32'h0;  // 32'h661988b6;
    ram_cell[   14293] = 32'h0;  // 32'h991c4a23;
    ram_cell[   14294] = 32'h0;  // 32'h0bfdcc2d;
    ram_cell[   14295] = 32'h0;  // 32'h0d7caeca;
    ram_cell[   14296] = 32'h0;  // 32'h13942452;
    ram_cell[   14297] = 32'h0;  // 32'h45521f09;
    ram_cell[   14298] = 32'h0;  // 32'h7631a48e;
    ram_cell[   14299] = 32'h0;  // 32'h5ebd6fe7;
    ram_cell[   14300] = 32'h0;  // 32'h1766a662;
    ram_cell[   14301] = 32'h0;  // 32'h4fb46589;
    ram_cell[   14302] = 32'h0;  // 32'h62f96555;
    ram_cell[   14303] = 32'h0;  // 32'h1d1dd652;
    ram_cell[   14304] = 32'h0;  // 32'hf9525207;
    ram_cell[   14305] = 32'h0;  // 32'h457d2f7d;
    ram_cell[   14306] = 32'h0;  // 32'hb138a282;
    ram_cell[   14307] = 32'h0;  // 32'h3ce859d3;
    ram_cell[   14308] = 32'h0;  // 32'hfe237b35;
    ram_cell[   14309] = 32'h0;  // 32'h78219c75;
    ram_cell[   14310] = 32'h0;  // 32'h13bc29f0;
    ram_cell[   14311] = 32'h0;  // 32'hb442c22a;
    ram_cell[   14312] = 32'h0;  // 32'h9d3dcbb0;
    ram_cell[   14313] = 32'h0;  // 32'h3a9846ba;
    ram_cell[   14314] = 32'h0;  // 32'h39c7f172;
    ram_cell[   14315] = 32'h0;  // 32'hd7f596c9;
    ram_cell[   14316] = 32'h0;  // 32'hac651cbf;
    ram_cell[   14317] = 32'h0;  // 32'hfed53e01;
    ram_cell[   14318] = 32'h0;  // 32'hb7e5a0e9;
    ram_cell[   14319] = 32'h0;  // 32'h643e4ee6;
    ram_cell[   14320] = 32'h0;  // 32'h7878c99a;
    ram_cell[   14321] = 32'h0;  // 32'hd786c13d;
    ram_cell[   14322] = 32'h0;  // 32'h902d92b1;
    ram_cell[   14323] = 32'h0;  // 32'h499ccbea;
    ram_cell[   14324] = 32'h0;  // 32'hc60e6019;
    ram_cell[   14325] = 32'h0;  // 32'hcd9fba82;
    ram_cell[   14326] = 32'h0;  // 32'h9c60a251;
    ram_cell[   14327] = 32'h0;  // 32'h7e4ccd20;
    ram_cell[   14328] = 32'h0;  // 32'h7f23ec47;
    ram_cell[   14329] = 32'h0;  // 32'hd7e2814f;
    ram_cell[   14330] = 32'h0;  // 32'hb8246462;
    ram_cell[   14331] = 32'h0;  // 32'h5ab970af;
    ram_cell[   14332] = 32'h0;  // 32'h6bd07df5;
    ram_cell[   14333] = 32'h0;  // 32'h72e8f1b1;
    ram_cell[   14334] = 32'h0;  // 32'h036d3853;
    ram_cell[   14335] = 32'h0;  // 32'h9d713c60;
    ram_cell[   14336] = 32'h0;  // 32'h852323be;
    ram_cell[   14337] = 32'h0;  // 32'he749b7e8;
    ram_cell[   14338] = 32'h0;  // 32'h40cb42f6;
    ram_cell[   14339] = 32'h0;  // 32'hc75e9d0d;
    ram_cell[   14340] = 32'h0;  // 32'hf3131781;
    ram_cell[   14341] = 32'h0;  // 32'h1238adf4;
    ram_cell[   14342] = 32'h0;  // 32'ha0026021;
    ram_cell[   14343] = 32'h0;  // 32'h6a6b9b94;
    ram_cell[   14344] = 32'h0;  // 32'hf1de139d;
    ram_cell[   14345] = 32'h0;  // 32'hcfef232f;
    ram_cell[   14346] = 32'h0;  // 32'h5c789b7e;
    ram_cell[   14347] = 32'h0;  // 32'h60e935c3;
    ram_cell[   14348] = 32'h0;  // 32'h52219e81;
    ram_cell[   14349] = 32'h0;  // 32'hf61a0a31;
    ram_cell[   14350] = 32'h0;  // 32'h3ddbf090;
    ram_cell[   14351] = 32'h0;  // 32'h5b54b9d0;
    ram_cell[   14352] = 32'h0;  // 32'h43b25d40;
    ram_cell[   14353] = 32'h0;  // 32'h7ad30cf9;
    ram_cell[   14354] = 32'h0;  // 32'hd9bd5e03;
    ram_cell[   14355] = 32'h0;  // 32'h82070245;
    ram_cell[   14356] = 32'h0;  // 32'h1a293a83;
    ram_cell[   14357] = 32'h0;  // 32'hc599b994;
    ram_cell[   14358] = 32'h0;  // 32'hc201fcc1;
    ram_cell[   14359] = 32'h0;  // 32'ha4ea5a1c;
    ram_cell[   14360] = 32'h0;  // 32'h92b01ddc;
    ram_cell[   14361] = 32'h0;  // 32'hba71bd72;
    ram_cell[   14362] = 32'h0;  // 32'h886e7a64;
    ram_cell[   14363] = 32'h0;  // 32'h801fe22a;
    ram_cell[   14364] = 32'h0;  // 32'haf654237;
    ram_cell[   14365] = 32'h0;  // 32'hcdb612f2;
    ram_cell[   14366] = 32'h0;  // 32'h0a605ff8;
    ram_cell[   14367] = 32'h0;  // 32'hc6622e50;
    ram_cell[   14368] = 32'h0;  // 32'h58de6418;
    ram_cell[   14369] = 32'h0;  // 32'h64afa3ab;
    ram_cell[   14370] = 32'h0;  // 32'hfc5fd790;
    ram_cell[   14371] = 32'h0;  // 32'h90360d67;
    ram_cell[   14372] = 32'h0;  // 32'h92441c25;
    ram_cell[   14373] = 32'h0;  // 32'hcdadc098;
    ram_cell[   14374] = 32'h0;  // 32'h1f4511c5;
    ram_cell[   14375] = 32'h0;  // 32'h68dcfbcc;
    ram_cell[   14376] = 32'h0;  // 32'h8360c22b;
    ram_cell[   14377] = 32'h0;  // 32'h3320360e;
    ram_cell[   14378] = 32'h0;  // 32'hc7459794;
    ram_cell[   14379] = 32'h0;  // 32'hfdade721;
    ram_cell[   14380] = 32'h0;  // 32'h813b8765;
    ram_cell[   14381] = 32'h0;  // 32'hf425c6f7;
    ram_cell[   14382] = 32'h0;  // 32'hfc22c53a;
    ram_cell[   14383] = 32'h0;  // 32'hc8635172;
    ram_cell[   14384] = 32'h0;  // 32'hfc719cba;
    ram_cell[   14385] = 32'h0;  // 32'h742b9c91;
    ram_cell[   14386] = 32'h0;  // 32'h13370a90;
    ram_cell[   14387] = 32'h0;  // 32'hd59cf7c2;
    ram_cell[   14388] = 32'h0;  // 32'ha47c6728;
    ram_cell[   14389] = 32'h0;  // 32'hb936c642;
    ram_cell[   14390] = 32'h0;  // 32'h35dd2893;
    ram_cell[   14391] = 32'h0;  // 32'h306c7340;
    ram_cell[   14392] = 32'h0;  // 32'h21cb4e34;
    ram_cell[   14393] = 32'h0;  // 32'hf3d4f795;
    ram_cell[   14394] = 32'h0;  // 32'hb3a472b6;
    ram_cell[   14395] = 32'h0;  // 32'h012bccde;
    ram_cell[   14396] = 32'h0;  // 32'ha860f618;
    ram_cell[   14397] = 32'h0;  // 32'h7cfe85e5;
    ram_cell[   14398] = 32'h0;  // 32'h36cc6885;
    ram_cell[   14399] = 32'h0;  // 32'hbfc08cae;
    ram_cell[   14400] = 32'h0;  // 32'hd2a64559;
    ram_cell[   14401] = 32'h0;  // 32'h5ca4643a;
    ram_cell[   14402] = 32'h0;  // 32'h4d91bcca;
    ram_cell[   14403] = 32'h0;  // 32'hff83d92e;
    ram_cell[   14404] = 32'h0;  // 32'hedfd1180;
    ram_cell[   14405] = 32'h0;  // 32'hb5052580;
    ram_cell[   14406] = 32'h0;  // 32'hfd5ba466;
    ram_cell[   14407] = 32'h0;  // 32'hb7ab44a4;
    ram_cell[   14408] = 32'h0;  // 32'h6646c168;
    ram_cell[   14409] = 32'h0;  // 32'hd5323383;
    ram_cell[   14410] = 32'h0;  // 32'h7469a615;
    ram_cell[   14411] = 32'h0;  // 32'hcce8f493;
    ram_cell[   14412] = 32'h0;  // 32'h8afa7469;
    ram_cell[   14413] = 32'h0;  // 32'h4ab92e49;
    ram_cell[   14414] = 32'h0;  // 32'haa492e76;
    ram_cell[   14415] = 32'h0;  // 32'h82e08eeb;
    ram_cell[   14416] = 32'h0;  // 32'hce612957;
    ram_cell[   14417] = 32'h0;  // 32'h2aca917d;
    ram_cell[   14418] = 32'h0;  // 32'hf5146ed7;
    ram_cell[   14419] = 32'h0;  // 32'h0686d425;
    ram_cell[   14420] = 32'h0;  // 32'he3d311a5;
    ram_cell[   14421] = 32'h0;  // 32'h4080335c;
    ram_cell[   14422] = 32'h0;  // 32'h6b532ba6;
    ram_cell[   14423] = 32'h0;  // 32'h16239506;
    ram_cell[   14424] = 32'h0;  // 32'h6b5421bb;
    ram_cell[   14425] = 32'h0;  // 32'h6ed548c3;
    ram_cell[   14426] = 32'h0;  // 32'h6f231edb;
    ram_cell[   14427] = 32'h0;  // 32'h7c634667;
    ram_cell[   14428] = 32'h0;  // 32'he1d2feb3;
    ram_cell[   14429] = 32'h0;  // 32'hf4d643c2;
    ram_cell[   14430] = 32'h0;  // 32'h8dac28b4;
    ram_cell[   14431] = 32'h0;  // 32'hd1813d0f;
    ram_cell[   14432] = 32'h0;  // 32'h4e2b93db;
    ram_cell[   14433] = 32'h0;  // 32'he5601df3;
    ram_cell[   14434] = 32'h0;  // 32'hd0404b00;
    ram_cell[   14435] = 32'h0;  // 32'h0a2fe662;
    ram_cell[   14436] = 32'h0;  // 32'hbddf9fce;
    ram_cell[   14437] = 32'h0;  // 32'h9dba6b76;
    ram_cell[   14438] = 32'h0;  // 32'hb6178c82;
    ram_cell[   14439] = 32'h0;  // 32'hd7043972;
    ram_cell[   14440] = 32'h0;  // 32'hbb938df4;
    ram_cell[   14441] = 32'h0;  // 32'hf9b86d73;
    ram_cell[   14442] = 32'h0;  // 32'hb34f6c31;
    ram_cell[   14443] = 32'h0;  // 32'h64a49df8;
    ram_cell[   14444] = 32'h0;  // 32'hf03517da;
    ram_cell[   14445] = 32'h0;  // 32'hf3646943;
    ram_cell[   14446] = 32'h0;  // 32'hd25c45da;
    ram_cell[   14447] = 32'h0;  // 32'h6b9d5656;
    ram_cell[   14448] = 32'h0;  // 32'h9f098fab;
    ram_cell[   14449] = 32'h0;  // 32'h7636c3ab;
    ram_cell[   14450] = 32'h0;  // 32'h36f55de6;
    ram_cell[   14451] = 32'h0;  // 32'hfb5c634c;
    ram_cell[   14452] = 32'h0;  // 32'h96198653;
    ram_cell[   14453] = 32'h0;  // 32'h75857cbb;
    ram_cell[   14454] = 32'h0;  // 32'h2d7e2bf1;
    ram_cell[   14455] = 32'h0;  // 32'hcf32dbbe;
    ram_cell[   14456] = 32'h0;  // 32'he21f7925;
    ram_cell[   14457] = 32'h0;  // 32'h2bea2ee9;
    ram_cell[   14458] = 32'h0;  // 32'he344156f;
    ram_cell[   14459] = 32'h0;  // 32'h24c8eb2c;
    ram_cell[   14460] = 32'h0;  // 32'h13d151af;
    ram_cell[   14461] = 32'h0;  // 32'h91af653e;
    ram_cell[   14462] = 32'h0;  // 32'h5a973bf2;
    ram_cell[   14463] = 32'h0;  // 32'h1170cfb8;
    ram_cell[   14464] = 32'h0;  // 32'he081be48;
    ram_cell[   14465] = 32'h0;  // 32'h26e69e5f;
    ram_cell[   14466] = 32'h0;  // 32'h5e6eb068;
    ram_cell[   14467] = 32'h0;  // 32'h1c7d36b6;
    ram_cell[   14468] = 32'h0;  // 32'h8890fe6c;
    ram_cell[   14469] = 32'h0;  // 32'h35041ea6;
    ram_cell[   14470] = 32'h0;  // 32'h4c57d1a2;
    ram_cell[   14471] = 32'h0;  // 32'haeba915e;
    ram_cell[   14472] = 32'h0;  // 32'hc79e38bd;
    ram_cell[   14473] = 32'h0;  // 32'h5b1f5b45;
    ram_cell[   14474] = 32'h0;  // 32'he9a9e1e4;
    ram_cell[   14475] = 32'h0;  // 32'hcb6c1927;
    ram_cell[   14476] = 32'h0;  // 32'hcd63578f;
    ram_cell[   14477] = 32'h0;  // 32'h1bcdc12f;
    ram_cell[   14478] = 32'h0;  // 32'hc12438a5;
    ram_cell[   14479] = 32'h0;  // 32'h5ee85dfc;
    ram_cell[   14480] = 32'h0;  // 32'h7c217759;
    ram_cell[   14481] = 32'h0;  // 32'hd2c0143b;
    ram_cell[   14482] = 32'h0;  // 32'hcd6ed76a;
    ram_cell[   14483] = 32'h0;  // 32'h8ff73323;
    ram_cell[   14484] = 32'h0;  // 32'hbf1eef7c;
    ram_cell[   14485] = 32'h0;  // 32'h67f5d9b2;
    ram_cell[   14486] = 32'h0;  // 32'h655c780d;
    ram_cell[   14487] = 32'h0;  // 32'heb0956c8;
    ram_cell[   14488] = 32'h0;  // 32'hcefcb6a4;
    ram_cell[   14489] = 32'h0;  // 32'hd705bed4;
    ram_cell[   14490] = 32'h0;  // 32'he4aeaaa6;
    ram_cell[   14491] = 32'h0;  // 32'hcf8eb1ec;
    ram_cell[   14492] = 32'h0;  // 32'hbed47cfc;
    ram_cell[   14493] = 32'h0;  // 32'h7a764830;
    ram_cell[   14494] = 32'h0;  // 32'h99600f46;
    ram_cell[   14495] = 32'h0;  // 32'h49d3d06f;
    ram_cell[   14496] = 32'h0;  // 32'h53dca3e0;
    ram_cell[   14497] = 32'h0;  // 32'h6e4513d9;
    ram_cell[   14498] = 32'h0;  // 32'hf6fe56b4;
    ram_cell[   14499] = 32'h0;  // 32'h226f7d7a;
    ram_cell[   14500] = 32'h0;  // 32'hd926de6e;
    ram_cell[   14501] = 32'h0;  // 32'h9e50f229;
    ram_cell[   14502] = 32'h0;  // 32'h2251ec9c;
    ram_cell[   14503] = 32'h0;  // 32'hec212b33;
    ram_cell[   14504] = 32'h0;  // 32'h82f97677;
    ram_cell[   14505] = 32'h0;  // 32'haa6b57d0;
    ram_cell[   14506] = 32'h0;  // 32'hc7e3a0f5;
    ram_cell[   14507] = 32'h0;  // 32'h33148224;
    ram_cell[   14508] = 32'h0;  // 32'h2b723a21;
    ram_cell[   14509] = 32'h0;  // 32'hc36c8846;
    ram_cell[   14510] = 32'h0;  // 32'hb2fb8c97;
    ram_cell[   14511] = 32'h0;  // 32'hc85e9834;
    ram_cell[   14512] = 32'h0;  // 32'h1d78af6e;
    ram_cell[   14513] = 32'h0;  // 32'h4768d2e8;
    ram_cell[   14514] = 32'h0;  // 32'h8c25abf4;
    ram_cell[   14515] = 32'h0;  // 32'h36bd13d6;
    ram_cell[   14516] = 32'h0;  // 32'h1ab397a7;
    ram_cell[   14517] = 32'h0;  // 32'hb1cb449d;
    ram_cell[   14518] = 32'h0;  // 32'h20ab408e;
    ram_cell[   14519] = 32'h0;  // 32'hbe2089fc;
    ram_cell[   14520] = 32'h0;  // 32'hd4edbe30;
    ram_cell[   14521] = 32'h0;  // 32'h4fa309c1;
    ram_cell[   14522] = 32'h0;  // 32'h8d33c5d0;
    ram_cell[   14523] = 32'h0;  // 32'he52faf9d;
    ram_cell[   14524] = 32'h0;  // 32'h01e578d8;
    ram_cell[   14525] = 32'h0;  // 32'h0d55f2a7;
    ram_cell[   14526] = 32'h0;  // 32'h015a40f0;
    ram_cell[   14527] = 32'h0;  // 32'hee6f0eb0;
    ram_cell[   14528] = 32'h0;  // 32'hd5b797cc;
    ram_cell[   14529] = 32'h0;  // 32'h9081abf8;
    ram_cell[   14530] = 32'h0;  // 32'hc04a4b0f;
    ram_cell[   14531] = 32'h0;  // 32'hf76c3787;
    ram_cell[   14532] = 32'h0;  // 32'hcb2ef96e;
    ram_cell[   14533] = 32'h0;  // 32'hcedd2adc;
    ram_cell[   14534] = 32'h0;  // 32'hf98e49c3;
    ram_cell[   14535] = 32'h0;  // 32'hf15d4789;
    ram_cell[   14536] = 32'h0;  // 32'hae47befc;
    ram_cell[   14537] = 32'h0;  // 32'h83553182;
    ram_cell[   14538] = 32'h0;  // 32'h00dd1aba;
    ram_cell[   14539] = 32'h0;  // 32'h0186531f;
    ram_cell[   14540] = 32'h0;  // 32'h005954bc;
    ram_cell[   14541] = 32'h0;  // 32'h8e9df025;
    ram_cell[   14542] = 32'h0;  // 32'h34c2eb4a;
    ram_cell[   14543] = 32'h0;  // 32'h242dec81;
    ram_cell[   14544] = 32'h0;  // 32'h4a9462f7;
    ram_cell[   14545] = 32'h0;  // 32'h8e4e3c1d;
    ram_cell[   14546] = 32'h0;  // 32'h77b1a94c;
    ram_cell[   14547] = 32'h0;  // 32'h6b845df8;
    ram_cell[   14548] = 32'h0;  // 32'h6861ee40;
    ram_cell[   14549] = 32'h0;  // 32'h0174f70b;
    ram_cell[   14550] = 32'h0;  // 32'h29fcf124;
    ram_cell[   14551] = 32'h0;  // 32'hce99caf5;
    ram_cell[   14552] = 32'h0;  // 32'h18cbebcb;
    ram_cell[   14553] = 32'h0;  // 32'h47cc53b6;
    ram_cell[   14554] = 32'h0;  // 32'hc21b4f9b;
    ram_cell[   14555] = 32'h0;  // 32'hda933667;
    ram_cell[   14556] = 32'h0;  // 32'h17239457;
    ram_cell[   14557] = 32'h0;  // 32'he3229416;
    ram_cell[   14558] = 32'h0;  // 32'h8954fa04;
    ram_cell[   14559] = 32'h0;  // 32'hab73188a;
    ram_cell[   14560] = 32'h0;  // 32'hb4455213;
    ram_cell[   14561] = 32'h0;  // 32'h349d63e3;
    ram_cell[   14562] = 32'h0;  // 32'h5bfa925d;
    ram_cell[   14563] = 32'h0;  // 32'h8508f69a;
    ram_cell[   14564] = 32'h0;  // 32'h5f8ac74f;
    ram_cell[   14565] = 32'h0;  // 32'h41dded5c;
    ram_cell[   14566] = 32'h0;  // 32'h8d6e1147;
    ram_cell[   14567] = 32'h0;  // 32'ha07f0b85;
    ram_cell[   14568] = 32'h0;  // 32'hda6b3bc0;
    ram_cell[   14569] = 32'h0;  // 32'h2b798c8c;
    ram_cell[   14570] = 32'h0;  // 32'h6e63816a;
    ram_cell[   14571] = 32'h0;  // 32'h6a12c657;
    ram_cell[   14572] = 32'h0;  // 32'h1c721ff3;
    ram_cell[   14573] = 32'h0;  // 32'h37985622;
    ram_cell[   14574] = 32'h0;  // 32'h5d66792c;
    ram_cell[   14575] = 32'h0;  // 32'hb68a3783;
    ram_cell[   14576] = 32'h0;  // 32'h9473d917;
    ram_cell[   14577] = 32'h0;  // 32'h1ff7cf82;
    ram_cell[   14578] = 32'h0;  // 32'ha5133628;
    ram_cell[   14579] = 32'h0;  // 32'h8e8de321;
    ram_cell[   14580] = 32'h0;  // 32'h3c8a744e;
    ram_cell[   14581] = 32'h0;  // 32'h3c2b8c17;
    ram_cell[   14582] = 32'h0;  // 32'hfc77f129;
    ram_cell[   14583] = 32'h0;  // 32'h19ba0396;
    ram_cell[   14584] = 32'h0;  // 32'h49e91ec5;
    ram_cell[   14585] = 32'h0;  // 32'h3b30ea41;
    ram_cell[   14586] = 32'h0;  // 32'h3e1668b1;
    ram_cell[   14587] = 32'h0;  // 32'h0b8b58ff;
    ram_cell[   14588] = 32'h0;  // 32'ha73e648f;
    ram_cell[   14589] = 32'h0;  // 32'hefff86c7;
    ram_cell[   14590] = 32'h0;  // 32'h22471ef2;
    ram_cell[   14591] = 32'h0;  // 32'h2c34058a;
    ram_cell[   14592] = 32'h0;  // 32'hf90f1e6a;
    ram_cell[   14593] = 32'h0;  // 32'h98f1cf4f;
    ram_cell[   14594] = 32'h0;  // 32'h6a3f3956;
    ram_cell[   14595] = 32'h0;  // 32'h8c58f82c;
    ram_cell[   14596] = 32'h0;  // 32'h845e48fb;
    ram_cell[   14597] = 32'h0;  // 32'h02e4618d;
    ram_cell[   14598] = 32'h0;  // 32'h48c021ee;
    ram_cell[   14599] = 32'h0;  // 32'h4439f643;
    ram_cell[   14600] = 32'h0;  // 32'ha8f35b20;
    ram_cell[   14601] = 32'h0;  // 32'h47ec668c;
    ram_cell[   14602] = 32'h0;  // 32'h8f149aa2;
    ram_cell[   14603] = 32'h0;  // 32'hfdc96330;
    ram_cell[   14604] = 32'h0;  // 32'h35b4a218;
    ram_cell[   14605] = 32'h0;  // 32'hf4c06f94;
    ram_cell[   14606] = 32'h0;  // 32'h8a29890a;
    ram_cell[   14607] = 32'h0;  // 32'h460080ba;
    ram_cell[   14608] = 32'h0;  // 32'hb6013366;
    ram_cell[   14609] = 32'h0;  // 32'hc2edb4cc;
    ram_cell[   14610] = 32'h0;  // 32'h6ef849b5;
    ram_cell[   14611] = 32'h0;  // 32'h07798576;
    ram_cell[   14612] = 32'h0;  // 32'h1ac86283;
    ram_cell[   14613] = 32'h0;  // 32'h508da891;
    ram_cell[   14614] = 32'h0;  // 32'h52a045a7;
    ram_cell[   14615] = 32'h0;  // 32'hb607f4f1;
    ram_cell[   14616] = 32'h0;  // 32'h92a624dc;
    ram_cell[   14617] = 32'h0;  // 32'h3cd8fbfc;
    ram_cell[   14618] = 32'h0;  // 32'h3e46d65c;
    ram_cell[   14619] = 32'h0;  // 32'h3781b9cf;
    ram_cell[   14620] = 32'h0;  // 32'h4761f904;
    ram_cell[   14621] = 32'h0;  // 32'h83bae326;
    ram_cell[   14622] = 32'h0;  // 32'h36d31ec0;
    ram_cell[   14623] = 32'h0;  // 32'h31f123b9;
    ram_cell[   14624] = 32'h0;  // 32'h92c7adf0;
    ram_cell[   14625] = 32'h0;  // 32'hdbe060a6;
    ram_cell[   14626] = 32'h0;  // 32'h0d3a93b8;
    ram_cell[   14627] = 32'h0;  // 32'h310e401b;
    ram_cell[   14628] = 32'h0;  // 32'h46f08b66;
    ram_cell[   14629] = 32'h0;  // 32'h84390429;
    ram_cell[   14630] = 32'h0;  // 32'h31e388e8;
    ram_cell[   14631] = 32'h0;  // 32'h3d7eb4bd;
    ram_cell[   14632] = 32'h0;  // 32'he986a109;
    ram_cell[   14633] = 32'h0;  // 32'ha37a8e93;
    ram_cell[   14634] = 32'h0;  // 32'h5c590d6a;
    ram_cell[   14635] = 32'h0;  // 32'hec2b17ad;
    ram_cell[   14636] = 32'h0;  // 32'h9a65eff4;
    ram_cell[   14637] = 32'h0;  // 32'h1fe90cc2;
    ram_cell[   14638] = 32'h0;  // 32'hef809102;
    ram_cell[   14639] = 32'h0;  // 32'hcf81ead6;
    ram_cell[   14640] = 32'h0;  // 32'hac72ed64;
    ram_cell[   14641] = 32'h0;  // 32'he8df0950;
    ram_cell[   14642] = 32'h0;  // 32'hb7aee07b;
    ram_cell[   14643] = 32'h0;  // 32'h4f828250;
    ram_cell[   14644] = 32'h0;  // 32'hff251f47;
    ram_cell[   14645] = 32'h0;  // 32'h749e6783;
    ram_cell[   14646] = 32'h0;  // 32'h4e3d66b7;
    ram_cell[   14647] = 32'h0;  // 32'hd951f0d5;
    ram_cell[   14648] = 32'h0;  // 32'h1165739f;
    ram_cell[   14649] = 32'h0;  // 32'h5ac838b8;
    ram_cell[   14650] = 32'h0;  // 32'hc9a793f3;
    ram_cell[   14651] = 32'h0;  // 32'hf56ab600;
    ram_cell[   14652] = 32'h0;  // 32'h8b0b80ce;
    ram_cell[   14653] = 32'h0;  // 32'haa782cc8;
    ram_cell[   14654] = 32'h0;  // 32'h03adc1af;
    ram_cell[   14655] = 32'h0;  // 32'h8f554d1b;
    ram_cell[   14656] = 32'h0;  // 32'hb7c4cfd5;
    ram_cell[   14657] = 32'h0;  // 32'hd0c3437e;
    ram_cell[   14658] = 32'h0;  // 32'h3116c0b6;
    ram_cell[   14659] = 32'h0;  // 32'hb28f8512;
    ram_cell[   14660] = 32'h0;  // 32'had4d9892;
    ram_cell[   14661] = 32'h0;  // 32'hf73ebd25;
    ram_cell[   14662] = 32'h0;  // 32'h6fca83ca;
    ram_cell[   14663] = 32'h0;  // 32'hb7ff0837;
    ram_cell[   14664] = 32'h0;  // 32'h01cd210c;
    ram_cell[   14665] = 32'h0;  // 32'h202176d9;
    ram_cell[   14666] = 32'h0;  // 32'hf1dcbb61;
    ram_cell[   14667] = 32'h0;  // 32'h3f89d69c;
    ram_cell[   14668] = 32'h0;  // 32'h24442b23;
    ram_cell[   14669] = 32'h0;  // 32'h83bf93f7;
    ram_cell[   14670] = 32'h0;  // 32'h93326a00;
    ram_cell[   14671] = 32'h0;  // 32'h4d48330f;
    ram_cell[   14672] = 32'h0;  // 32'hbbe4f811;
    ram_cell[   14673] = 32'h0;  // 32'h8fdef724;
    ram_cell[   14674] = 32'h0;  // 32'hc36a2e72;
    ram_cell[   14675] = 32'h0;  // 32'h50946621;
    ram_cell[   14676] = 32'h0;  // 32'hdfebc5b7;
    ram_cell[   14677] = 32'h0;  // 32'h0da15581;
    ram_cell[   14678] = 32'h0;  // 32'hc78efb8a;
    ram_cell[   14679] = 32'h0;  // 32'h3bfa4bcb;
    ram_cell[   14680] = 32'h0;  // 32'h4f198edc;
    ram_cell[   14681] = 32'h0;  // 32'h40c45a7b;
    ram_cell[   14682] = 32'h0;  // 32'h781f0de5;
    ram_cell[   14683] = 32'h0;  // 32'h615f70b1;
    ram_cell[   14684] = 32'h0;  // 32'ha5019435;
    ram_cell[   14685] = 32'h0;  // 32'hd5e2d64c;
    ram_cell[   14686] = 32'h0;  // 32'h6c09663d;
    ram_cell[   14687] = 32'h0;  // 32'h0377e818;
    ram_cell[   14688] = 32'h0;  // 32'hb3fb854e;
    ram_cell[   14689] = 32'h0;  // 32'h8059e70a;
    ram_cell[   14690] = 32'h0;  // 32'h3b5e70d3;
    ram_cell[   14691] = 32'h0;  // 32'h34248858;
    ram_cell[   14692] = 32'h0;  // 32'hd0448ca0;
    ram_cell[   14693] = 32'h0;  // 32'hdb8a66c8;
    ram_cell[   14694] = 32'h0;  // 32'hcb932fbc;
    ram_cell[   14695] = 32'h0;  // 32'he3b7575c;
    ram_cell[   14696] = 32'h0;  // 32'h91837f7c;
    ram_cell[   14697] = 32'h0;  // 32'h3cb077a8;
    ram_cell[   14698] = 32'h0;  // 32'h49e9e328;
    ram_cell[   14699] = 32'h0;  // 32'hccbc6000;
    ram_cell[   14700] = 32'h0;  // 32'h20116f5f;
    ram_cell[   14701] = 32'h0;  // 32'h809a6651;
    ram_cell[   14702] = 32'h0;  // 32'h79a6f4c6;
    ram_cell[   14703] = 32'h0;  // 32'h8540fcd0;
    ram_cell[   14704] = 32'h0;  // 32'h409bd2f1;
    ram_cell[   14705] = 32'h0;  // 32'h9acf4adc;
    ram_cell[   14706] = 32'h0;  // 32'h866ee3a4;
    ram_cell[   14707] = 32'h0;  // 32'h50307619;
    ram_cell[   14708] = 32'h0;  // 32'hed059462;
    ram_cell[   14709] = 32'h0;  // 32'hdb2177f3;
    ram_cell[   14710] = 32'h0;  // 32'had3a43a4;
    ram_cell[   14711] = 32'h0;  // 32'h712a3197;
    ram_cell[   14712] = 32'h0;  // 32'hfc72082e;
    ram_cell[   14713] = 32'h0;  // 32'h8783dd3a;
    ram_cell[   14714] = 32'h0;  // 32'h592aca4d;
    ram_cell[   14715] = 32'h0;  // 32'ha0383f95;
    ram_cell[   14716] = 32'h0;  // 32'h4732dcb9;
    ram_cell[   14717] = 32'h0;  // 32'h1036ef05;
    ram_cell[   14718] = 32'h0;  // 32'hfdc499a0;
    ram_cell[   14719] = 32'h0;  // 32'h61fd97fb;
    ram_cell[   14720] = 32'h0;  // 32'h086024c2;
    ram_cell[   14721] = 32'h0;  // 32'h2ce4531b;
    ram_cell[   14722] = 32'h0;  // 32'hc2696d8e;
    ram_cell[   14723] = 32'h0;  // 32'hc09a3d17;
    ram_cell[   14724] = 32'h0;  // 32'hf670ea05;
    ram_cell[   14725] = 32'h0;  // 32'h4302acab;
    ram_cell[   14726] = 32'h0;  // 32'h42f9e16c;
    ram_cell[   14727] = 32'h0;  // 32'h9f3a3fdd;
    ram_cell[   14728] = 32'h0;  // 32'hb51dd215;
    ram_cell[   14729] = 32'h0;  // 32'habb8495e;
    ram_cell[   14730] = 32'h0;  // 32'hf63422bd;
    ram_cell[   14731] = 32'h0;  // 32'hbaf7b861;
    ram_cell[   14732] = 32'h0;  // 32'h5967d92f;
    ram_cell[   14733] = 32'h0;  // 32'hec9c6236;
    ram_cell[   14734] = 32'h0;  // 32'hd57b2f7b;
    ram_cell[   14735] = 32'h0;  // 32'hcc534bab;
    ram_cell[   14736] = 32'h0;  // 32'h60ce47a2;
    ram_cell[   14737] = 32'h0;  // 32'he9b15d95;
    ram_cell[   14738] = 32'h0;  // 32'h8beb98c3;
    ram_cell[   14739] = 32'h0;  // 32'h864dcbdb;
    ram_cell[   14740] = 32'h0;  // 32'hd9465ad8;
    ram_cell[   14741] = 32'h0;  // 32'h28c98fc8;
    ram_cell[   14742] = 32'h0;  // 32'h231305db;
    ram_cell[   14743] = 32'h0;  // 32'h2ed2d73c;
    ram_cell[   14744] = 32'h0;  // 32'hdbe1f5dd;
    ram_cell[   14745] = 32'h0;  // 32'h4e9bba9d;
    ram_cell[   14746] = 32'h0;  // 32'hc6e4d284;
    ram_cell[   14747] = 32'h0;  // 32'h4971ce17;
    ram_cell[   14748] = 32'h0;  // 32'hfe4fa1d1;
    ram_cell[   14749] = 32'h0;  // 32'h0f6c55bd;
    ram_cell[   14750] = 32'h0;  // 32'hd1ec9458;
    ram_cell[   14751] = 32'h0;  // 32'h1e16da10;
    ram_cell[   14752] = 32'h0;  // 32'h4826ad4a;
    ram_cell[   14753] = 32'h0;  // 32'hd48b2bbc;
    ram_cell[   14754] = 32'h0;  // 32'h49479734;
    ram_cell[   14755] = 32'h0;  // 32'h105b68e2;
    ram_cell[   14756] = 32'h0;  // 32'h2bcc0ef8;
    ram_cell[   14757] = 32'h0;  // 32'h57c83968;
    ram_cell[   14758] = 32'h0;  // 32'h9bd92faf;
    ram_cell[   14759] = 32'h0;  // 32'h75a5b2cc;
    ram_cell[   14760] = 32'h0;  // 32'h8d0e76de;
    ram_cell[   14761] = 32'h0;  // 32'hf1ab2caa;
    ram_cell[   14762] = 32'h0;  // 32'h309f6ea2;
    ram_cell[   14763] = 32'h0;  // 32'h12df3e6d;
    ram_cell[   14764] = 32'h0;  // 32'h46e12c94;
    ram_cell[   14765] = 32'h0;  // 32'ha9c93dc0;
    ram_cell[   14766] = 32'h0;  // 32'h9ca7be6a;
    ram_cell[   14767] = 32'h0;  // 32'he5e1e089;
    ram_cell[   14768] = 32'h0;  // 32'h51bdda26;
    ram_cell[   14769] = 32'h0;  // 32'h528a4ab8;
    ram_cell[   14770] = 32'h0;  // 32'h023ad5ac;
    ram_cell[   14771] = 32'h0;  // 32'hd11dd6fc;
    ram_cell[   14772] = 32'h0;  // 32'hb5e807de;
    ram_cell[   14773] = 32'h0;  // 32'ha3f38119;
    ram_cell[   14774] = 32'h0;  // 32'h90fb3ea2;
    ram_cell[   14775] = 32'h0;  // 32'h48106364;
    ram_cell[   14776] = 32'h0;  // 32'hd263b0d8;
    ram_cell[   14777] = 32'h0;  // 32'h3b54ef97;
    ram_cell[   14778] = 32'h0;  // 32'hb6fa02f5;
    ram_cell[   14779] = 32'h0;  // 32'hff8b4d04;
    ram_cell[   14780] = 32'h0;  // 32'ha8d0b9e3;
    ram_cell[   14781] = 32'h0;  // 32'hcc6643aa;
    ram_cell[   14782] = 32'h0;  // 32'h57b11d21;
    ram_cell[   14783] = 32'h0;  // 32'h3a6c9943;
    ram_cell[   14784] = 32'h0;  // 32'h8dd38a88;
    ram_cell[   14785] = 32'h0;  // 32'haf3fd7c2;
    ram_cell[   14786] = 32'h0;  // 32'h0076c2c5;
    ram_cell[   14787] = 32'h0;  // 32'hd454f3dc;
    ram_cell[   14788] = 32'h0;  // 32'h3c2ee139;
    ram_cell[   14789] = 32'h0;  // 32'hb7ba04d6;
    ram_cell[   14790] = 32'h0;  // 32'h68861b06;
    ram_cell[   14791] = 32'h0;  // 32'h051534aa;
    ram_cell[   14792] = 32'h0;  // 32'hfc7fef30;
    ram_cell[   14793] = 32'h0;  // 32'h103148d7;
    ram_cell[   14794] = 32'h0;  // 32'h76735b6a;
    ram_cell[   14795] = 32'h0;  // 32'hc86491a7;
    ram_cell[   14796] = 32'h0;  // 32'h34245e0d;
    ram_cell[   14797] = 32'h0;  // 32'h280afd98;
    ram_cell[   14798] = 32'h0;  // 32'h4f124ed9;
    ram_cell[   14799] = 32'h0;  // 32'h4791761e;
    ram_cell[   14800] = 32'h0;  // 32'h01cb0a24;
    ram_cell[   14801] = 32'h0;  // 32'hf37848de;
    ram_cell[   14802] = 32'h0;  // 32'h7cea30fb;
    ram_cell[   14803] = 32'h0;  // 32'h2de2bb06;
    ram_cell[   14804] = 32'h0;  // 32'hbfdff095;
    ram_cell[   14805] = 32'h0;  // 32'h4611cefd;
    ram_cell[   14806] = 32'h0;  // 32'h64afac32;
    ram_cell[   14807] = 32'h0;  // 32'hb0fd1aa4;
    ram_cell[   14808] = 32'h0;  // 32'hd8d35db2;
    ram_cell[   14809] = 32'h0;  // 32'h8e398976;
    ram_cell[   14810] = 32'h0;  // 32'hf4d462fd;
    ram_cell[   14811] = 32'h0;  // 32'h8dff21ed;
    ram_cell[   14812] = 32'h0;  // 32'h1801cf1e;
    ram_cell[   14813] = 32'h0;  // 32'hd6d35798;
    ram_cell[   14814] = 32'h0;  // 32'h55bf7a15;
    ram_cell[   14815] = 32'h0;  // 32'h03150b61;
    ram_cell[   14816] = 32'h0;  // 32'hf5b5277c;
    ram_cell[   14817] = 32'h0;  // 32'hb8001cd5;
    ram_cell[   14818] = 32'h0;  // 32'h78222f24;
    ram_cell[   14819] = 32'h0;  // 32'h3aae945d;
    ram_cell[   14820] = 32'h0;  // 32'h4ba1dc95;
    ram_cell[   14821] = 32'h0;  // 32'h085b7cc5;
    ram_cell[   14822] = 32'h0;  // 32'h16a839c7;
    ram_cell[   14823] = 32'h0;  // 32'hc79ea645;
    ram_cell[   14824] = 32'h0;  // 32'ha7790645;
    ram_cell[   14825] = 32'h0;  // 32'hdc9ac753;
    ram_cell[   14826] = 32'h0;  // 32'hd9674c42;
    ram_cell[   14827] = 32'h0;  // 32'ha059e639;
    ram_cell[   14828] = 32'h0;  // 32'he78de8a2;
    ram_cell[   14829] = 32'h0;  // 32'he3c6bf8d;
    ram_cell[   14830] = 32'h0;  // 32'hbe678967;
    ram_cell[   14831] = 32'h0;  // 32'h9b43636b;
    ram_cell[   14832] = 32'h0;  // 32'hbec2c033;
    ram_cell[   14833] = 32'h0;  // 32'h0a61ec26;
    ram_cell[   14834] = 32'h0;  // 32'hda247e8c;
    ram_cell[   14835] = 32'h0;  // 32'hf987d04a;
    ram_cell[   14836] = 32'h0;  // 32'hf2f303cd;
    ram_cell[   14837] = 32'h0;  // 32'hd9b17754;
    ram_cell[   14838] = 32'h0;  // 32'had9be4cf;
    ram_cell[   14839] = 32'h0;  // 32'h09a0c99e;
    ram_cell[   14840] = 32'h0;  // 32'h92c85e0b;
    ram_cell[   14841] = 32'h0;  // 32'h8c375a3e;
    ram_cell[   14842] = 32'h0;  // 32'h45b6ef69;
    ram_cell[   14843] = 32'h0;  // 32'h401f5244;
    ram_cell[   14844] = 32'h0;  // 32'h8a4ec6d3;
    ram_cell[   14845] = 32'h0;  // 32'h581e9291;
    ram_cell[   14846] = 32'h0;  // 32'hc65a79fa;
    ram_cell[   14847] = 32'h0;  // 32'h4fd5d115;
    ram_cell[   14848] = 32'h0;  // 32'h29ea6e63;
    ram_cell[   14849] = 32'h0;  // 32'heb63dc47;
    ram_cell[   14850] = 32'h0;  // 32'h29306e70;
    ram_cell[   14851] = 32'h0;  // 32'hb5a3c3e4;
    ram_cell[   14852] = 32'h0;  // 32'hb165503b;
    ram_cell[   14853] = 32'h0;  // 32'he52dfcb7;
    ram_cell[   14854] = 32'h0;  // 32'hc3b0f81b;
    ram_cell[   14855] = 32'h0;  // 32'h3fc06abb;
    ram_cell[   14856] = 32'h0;  // 32'he6ec1939;
    ram_cell[   14857] = 32'h0;  // 32'h666f65d0;
    ram_cell[   14858] = 32'h0;  // 32'h1c307e32;
    ram_cell[   14859] = 32'h0;  // 32'h664c1c98;
    ram_cell[   14860] = 32'h0;  // 32'h9467a8ba;
    ram_cell[   14861] = 32'h0;  // 32'h498c4b5d;
    ram_cell[   14862] = 32'h0;  // 32'he79bd435;
    ram_cell[   14863] = 32'h0;  // 32'ha473e56f;
    ram_cell[   14864] = 32'h0;  // 32'h7ed86d4a;
    ram_cell[   14865] = 32'h0;  // 32'hcf766f16;
    ram_cell[   14866] = 32'h0;  // 32'h25d48ac1;
    ram_cell[   14867] = 32'h0;  // 32'h6c950d0d;
    ram_cell[   14868] = 32'h0;  // 32'h2a80f538;
    ram_cell[   14869] = 32'h0;  // 32'hdc475896;
    ram_cell[   14870] = 32'h0;  // 32'h8489c4a1;
    ram_cell[   14871] = 32'h0;  // 32'hb5f55496;
    ram_cell[   14872] = 32'h0;  // 32'h7d5a8768;
    ram_cell[   14873] = 32'h0;  // 32'h4584700b;
    ram_cell[   14874] = 32'h0;  // 32'hd706a9d2;
    ram_cell[   14875] = 32'h0;  // 32'h7fe35536;
    ram_cell[   14876] = 32'h0;  // 32'h7195ebeb;
    ram_cell[   14877] = 32'h0;  // 32'h2e2afb73;
    ram_cell[   14878] = 32'h0;  // 32'h0b409143;
    ram_cell[   14879] = 32'h0;  // 32'h5b032a4a;
    ram_cell[   14880] = 32'h0;  // 32'h1757ebd7;
    ram_cell[   14881] = 32'h0;  // 32'hd8eb5723;
    ram_cell[   14882] = 32'h0;  // 32'h632f8eaf;
    ram_cell[   14883] = 32'h0;  // 32'h3a166bbb;
    ram_cell[   14884] = 32'h0;  // 32'hf79f94e1;
    ram_cell[   14885] = 32'h0;  // 32'h1669417d;
    ram_cell[   14886] = 32'h0;  // 32'h163578d0;
    ram_cell[   14887] = 32'h0;  // 32'h77cca1be;
    ram_cell[   14888] = 32'h0;  // 32'h3e4b0da0;
    ram_cell[   14889] = 32'h0;  // 32'h80a76ea2;
    ram_cell[   14890] = 32'h0;  // 32'haabd0369;
    ram_cell[   14891] = 32'h0;  // 32'h16eceac9;
    ram_cell[   14892] = 32'h0;  // 32'h9a856fa7;
    ram_cell[   14893] = 32'h0;  // 32'hef454719;
    ram_cell[   14894] = 32'h0;  // 32'h964558d6;
    ram_cell[   14895] = 32'h0;  // 32'h792e36d0;
    ram_cell[   14896] = 32'h0;  // 32'h671d1e93;
    ram_cell[   14897] = 32'h0;  // 32'ha761e7d3;
    ram_cell[   14898] = 32'h0;  // 32'hd091ed9f;
    ram_cell[   14899] = 32'h0;  // 32'h7e74f585;
    ram_cell[   14900] = 32'h0;  // 32'h460f1594;
    ram_cell[   14901] = 32'h0;  // 32'h496e803b;
    ram_cell[   14902] = 32'h0;  // 32'he04ca269;
    ram_cell[   14903] = 32'h0;  // 32'h5248ca8a;
    ram_cell[   14904] = 32'h0;  // 32'h3b46f55b;
    ram_cell[   14905] = 32'h0;  // 32'h2f2e94da;
    ram_cell[   14906] = 32'h0;  // 32'h7bc9a3fb;
    ram_cell[   14907] = 32'h0;  // 32'h1023f725;
    ram_cell[   14908] = 32'h0;  // 32'h5bd47296;
    ram_cell[   14909] = 32'h0;  // 32'hb4eaec4f;
    ram_cell[   14910] = 32'h0;  // 32'h99d4094f;
    ram_cell[   14911] = 32'h0;  // 32'hfbceafa4;
    ram_cell[   14912] = 32'h0;  // 32'h9745167b;
    ram_cell[   14913] = 32'h0;  // 32'hba8f7f04;
    ram_cell[   14914] = 32'h0;  // 32'ha6cceeca;
    ram_cell[   14915] = 32'h0;  // 32'h372878fb;
    ram_cell[   14916] = 32'h0;  // 32'h339fa1f0;
    ram_cell[   14917] = 32'h0;  // 32'he9fb67d9;
    ram_cell[   14918] = 32'h0;  // 32'h9f70db4e;
    ram_cell[   14919] = 32'h0;  // 32'h35e1ca61;
    ram_cell[   14920] = 32'h0;  // 32'heec54d5d;
    ram_cell[   14921] = 32'h0;  // 32'h40b9664a;
    ram_cell[   14922] = 32'h0;  // 32'he564a3ff;
    ram_cell[   14923] = 32'h0;  // 32'hb1141ca8;
    ram_cell[   14924] = 32'h0;  // 32'h572d07af;
    ram_cell[   14925] = 32'h0;  // 32'hfb415b65;
    ram_cell[   14926] = 32'h0;  // 32'h7596d24b;
    ram_cell[   14927] = 32'h0;  // 32'hf18c61b3;
    ram_cell[   14928] = 32'h0;  // 32'h36e730f8;
    ram_cell[   14929] = 32'h0;  // 32'hfe602941;
    ram_cell[   14930] = 32'h0;  // 32'h502af6c2;
    ram_cell[   14931] = 32'h0;  // 32'h49abfec6;
    ram_cell[   14932] = 32'h0;  // 32'h1e413f46;
    ram_cell[   14933] = 32'h0;  // 32'h17e5eea7;
    ram_cell[   14934] = 32'h0;  // 32'h9991efb6;
    ram_cell[   14935] = 32'h0;  // 32'he1e8b212;
    ram_cell[   14936] = 32'h0;  // 32'h00184672;
    ram_cell[   14937] = 32'h0;  // 32'h3f2be17b;
    ram_cell[   14938] = 32'h0;  // 32'hcd8ce92b;
    ram_cell[   14939] = 32'h0;  // 32'h0c9dad55;
    ram_cell[   14940] = 32'h0;  // 32'h90125a19;
    ram_cell[   14941] = 32'h0;  // 32'h31da0acf;
    ram_cell[   14942] = 32'h0;  // 32'h4c385b72;
    ram_cell[   14943] = 32'h0;  // 32'he57de6a2;
    ram_cell[   14944] = 32'h0;  // 32'hb4e5cd24;
    ram_cell[   14945] = 32'h0;  // 32'h50fd1900;
    ram_cell[   14946] = 32'h0;  // 32'he5b8657d;
    ram_cell[   14947] = 32'h0;  // 32'h006d7763;
    ram_cell[   14948] = 32'h0;  // 32'hb6d5f2ea;
    ram_cell[   14949] = 32'h0;  // 32'hcb102369;
    ram_cell[   14950] = 32'h0;  // 32'hd3f14e46;
    ram_cell[   14951] = 32'h0;  // 32'hf24d4329;
    ram_cell[   14952] = 32'h0;  // 32'h1f1cbf0a;
    ram_cell[   14953] = 32'h0;  // 32'h000e3fa1;
    ram_cell[   14954] = 32'h0;  // 32'h8d6df35f;
    ram_cell[   14955] = 32'h0;  // 32'hd43d194b;
    ram_cell[   14956] = 32'h0;  // 32'h5c99a61d;
    ram_cell[   14957] = 32'h0;  // 32'h2773e39c;
    ram_cell[   14958] = 32'h0;  // 32'h3946facc;
    ram_cell[   14959] = 32'h0;  // 32'h5d0c243b;
    ram_cell[   14960] = 32'h0;  // 32'h7f41c512;
    ram_cell[   14961] = 32'h0;  // 32'hb2131c8d;
    ram_cell[   14962] = 32'h0;  // 32'h83958a43;
    ram_cell[   14963] = 32'h0;  // 32'h392ac7bd;
    ram_cell[   14964] = 32'h0;  // 32'h10455621;
    ram_cell[   14965] = 32'h0;  // 32'hb1c21dec;
    ram_cell[   14966] = 32'h0;  // 32'h8919b880;
    ram_cell[   14967] = 32'h0;  // 32'hf07c463a;
    ram_cell[   14968] = 32'h0;  // 32'h9db781e0;
    ram_cell[   14969] = 32'h0;  // 32'h2bb77c44;
    ram_cell[   14970] = 32'h0;  // 32'ha036ffec;
    ram_cell[   14971] = 32'h0;  // 32'hf1a85568;
    ram_cell[   14972] = 32'h0;  // 32'h8417b2f3;
    ram_cell[   14973] = 32'h0;  // 32'h92e64ee5;
    ram_cell[   14974] = 32'h0;  // 32'h8dc3dc43;
    ram_cell[   14975] = 32'h0;  // 32'ha2c950db;
    ram_cell[   14976] = 32'h0;  // 32'h36648cd6;
    ram_cell[   14977] = 32'h0;  // 32'h45df3df6;
    ram_cell[   14978] = 32'h0;  // 32'h95b2ec6c;
    ram_cell[   14979] = 32'h0;  // 32'h6884c52d;
    ram_cell[   14980] = 32'h0;  // 32'h0838f7ed;
    ram_cell[   14981] = 32'h0;  // 32'hc7bccf7c;
    ram_cell[   14982] = 32'h0;  // 32'h452cb364;
    ram_cell[   14983] = 32'h0;  // 32'h592482e4;
    ram_cell[   14984] = 32'h0;  // 32'h028a1e31;
    ram_cell[   14985] = 32'h0;  // 32'ha08c7e83;
    ram_cell[   14986] = 32'h0;  // 32'h606d13a4;
    ram_cell[   14987] = 32'h0;  // 32'h13c5c979;
    ram_cell[   14988] = 32'h0;  // 32'hb8be92ba;
    ram_cell[   14989] = 32'h0;  // 32'h0f1cb97d;
    ram_cell[   14990] = 32'h0;  // 32'h6f847f90;
    ram_cell[   14991] = 32'h0;  // 32'had310def;
    ram_cell[   14992] = 32'h0;  // 32'h944b39dc;
    ram_cell[   14993] = 32'h0;  // 32'habc31ae8;
    ram_cell[   14994] = 32'h0;  // 32'h5eeac796;
    ram_cell[   14995] = 32'h0;  // 32'h9f8978bd;
    ram_cell[   14996] = 32'h0;  // 32'h30face53;
    ram_cell[   14997] = 32'h0;  // 32'h952bb6f4;
    ram_cell[   14998] = 32'h0;  // 32'h288b1eb0;
    ram_cell[   14999] = 32'h0;  // 32'hb55f0999;
    ram_cell[   15000] = 32'h0;  // 32'h2d0270fe;
    ram_cell[   15001] = 32'h0;  // 32'h2d208b9e;
    ram_cell[   15002] = 32'h0;  // 32'h1bb36e2b;
    ram_cell[   15003] = 32'h0;  // 32'hd0ed7360;
    ram_cell[   15004] = 32'h0;  // 32'h3c9c4a87;
    ram_cell[   15005] = 32'h0;  // 32'hc09e0d3b;
    ram_cell[   15006] = 32'h0;  // 32'hcd0f543e;
    ram_cell[   15007] = 32'h0;  // 32'hc6ccad81;
    ram_cell[   15008] = 32'h0;  // 32'h13ac7de0;
    ram_cell[   15009] = 32'h0;  // 32'h03e10ba1;
    ram_cell[   15010] = 32'h0;  // 32'hf3e4474f;
    ram_cell[   15011] = 32'h0;  // 32'hb68377a2;
    ram_cell[   15012] = 32'h0;  // 32'he8541273;
    ram_cell[   15013] = 32'h0;  // 32'hbe85713c;
    ram_cell[   15014] = 32'h0;  // 32'h6ac9102f;
    ram_cell[   15015] = 32'h0;  // 32'he8e8a6ab;
    ram_cell[   15016] = 32'h0;  // 32'ha9037543;
    ram_cell[   15017] = 32'h0;  // 32'h30377d12;
    ram_cell[   15018] = 32'h0;  // 32'h2c40927f;
    ram_cell[   15019] = 32'h0;  // 32'hb04519fd;
    ram_cell[   15020] = 32'h0;  // 32'hc9f3fc09;
    ram_cell[   15021] = 32'h0;  // 32'h4c47a39f;
    ram_cell[   15022] = 32'h0;  // 32'h2a72afff;
    ram_cell[   15023] = 32'h0;  // 32'hb8f1d5c0;
    ram_cell[   15024] = 32'h0;  // 32'h38d768fc;
    ram_cell[   15025] = 32'h0;  // 32'ha4b7cf8c;
    ram_cell[   15026] = 32'h0;  // 32'h8ca95061;
    ram_cell[   15027] = 32'h0;  // 32'h5f5491f3;
    ram_cell[   15028] = 32'h0;  // 32'h12391ca1;
    ram_cell[   15029] = 32'h0;  // 32'h7f6c61e8;
    ram_cell[   15030] = 32'h0;  // 32'h4d6192e0;
    ram_cell[   15031] = 32'h0;  // 32'h2cf1a52e;
    ram_cell[   15032] = 32'h0;  // 32'h9509a476;
    ram_cell[   15033] = 32'h0;  // 32'h7edf54d1;
    ram_cell[   15034] = 32'h0;  // 32'hbe4afdbc;
    ram_cell[   15035] = 32'h0;  // 32'h57122139;
    ram_cell[   15036] = 32'h0;  // 32'hb67ae4f0;
    ram_cell[   15037] = 32'h0;  // 32'h1dbc8cba;
    ram_cell[   15038] = 32'h0;  // 32'h0ceb0a5d;
    ram_cell[   15039] = 32'h0;  // 32'h69e37ad8;
    ram_cell[   15040] = 32'h0;  // 32'h76bf31d8;
    ram_cell[   15041] = 32'h0;  // 32'h77aa1791;
    ram_cell[   15042] = 32'h0;  // 32'h90c7b0b9;
    ram_cell[   15043] = 32'h0;  // 32'h4770ce2f;
    ram_cell[   15044] = 32'h0;  // 32'h10ba9d80;
    ram_cell[   15045] = 32'h0;  // 32'hb017ae6c;
    ram_cell[   15046] = 32'h0;  // 32'h5a2f123b;
    ram_cell[   15047] = 32'h0;  // 32'h85dfc4dc;
    ram_cell[   15048] = 32'h0;  // 32'h5a3864e1;
    ram_cell[   15049] = 32'h0;  // 32'h5ab78578;
    ram_cell[   15050] = 32'h0;  // 32'hbd515e0d;
    ram_cell[   15051] = 32'h0;  // 32'h4ea18aff;
    ram_cell[   15052] = 32'h0;  // 32'h671d381f;
    ram_cell[   15053] = 32'h0;  // 32'h0ed49cd2;
    ram_cell[   15054] = 32'h0;  // 32'hac68b938;
    ram_cell[   15055] = 32'h0;  // 32'h52491073;
    ram_cell[   15056] = 32'h0;  // 32'he105b5d2;
    ram_cell[   15057] = 32'h0;  // 32'hc485a6ad;
    ram_cell[   15058] = 32'h0;  // 32'hc8d5db10;
    ram_cell[   15059] = 32'h0;  // 32'h6a81620f;
    ram_cell[   15060] = 32'h0;  // 32'h55c0723f;
    ram_cell[   15061] = 32'h0;  // 32'hceefc203;
    ram_cell[   15062] = 32'h0;  // 32'h5e41a7ef;
    ram_cell[   15063] = 32'h0;  // 32'hf79a7114;
    ram_cell[   15064] = 32'h0;  // 32'hbae58dc7;
    ram_cell[   15065] = 32'h0;  // 32'hddab53e7;
    ram_cell[   15066] = 32'h0;  // 32'h414d403b;
    ram_cell[   15067] = 32'h0;  // 32'h7ee25799;
    ram_cell[   15068] = 32'h0;  // 32'h6a398fc9;
    ram_cell[   15069] = 32'h0;  // 32'hafe6f76a;
    ram_cell[   15070] = 32'h0;  // 32'h2ec08775;
    ram_cell[   15071] = 32'h0;  // 32'hd4e8377d;
    ram_cell[   15072] = 32'h0;  // 32'h7e9f9270;
    ram_cell[   15073] = 32'h0;  // 32'he18a0370;
    ram_cell[   15074] = 32'h0;  // 32'hf6c5538a;
    ram_cell[   15075] = 32'h0;  // 32'hbd3924bc;
    ram_cell[   15076] = 32'h0;  // 32'hb93e1f11;
    ram_cell[   15077] = 32'h0;  // 32'h347eafcf;
    ram_cell[   15078] = 32'h0;  // 32'hdfd2ca80;
    ram_cell[   15079] = 32'h0;  // 32'hcbfb3a85;
    ram_cell[   15080] = 32'h0;  // 32'hff98ef08;
    ram_cell[   15081] = 32'h0;  // 32'h292a1dd5;
    ram_cell[   15082] = 32'h0;  // 32'h22fc949d;
    ram_cell[   15083] = 32'h0;  // 32'h9be9704d;
    ram_cell[   15084] = 32'h0;  // 32'h8a66855e;
    ram_cell[   15085] = 32'h0;  // 32'h427c989d;
    ram_cell[   15086] = 32'h0;  // 32'hc3a29cff;
    ram_cell[   15087] = 32'h0;  // 32'h6e62dfac;
    ram_cell[   15088] = 32'h0;  // 32'h60f8b788;
    ram_cell[   15089] = 32'h0;  // 32'hc302ff0d;
    ram_cell[   15090] = 32'h0;  // 32'h669b003f;
    ram_cell[   15091] = 32'h0;  // 32'h655b5b51;
    ram_cell[   15092] = 32'h0;  // 32'h503bdebe;
    ram_cell[   15093] = 32'h0;  // 32'h4a5453db;
    ram_cell[   15094] = 32'h0;  // 32'h2c42f776;
    ram_cell[   15095] = 32'h0;  // 32'h91f90e1d;
    ram_cell[   15096] = 32'h0;  // 32'h48321fc5;
    ram_cell[   15097] = 32'h0;  // 32'h7b57865f;
    ram_cell[   15098] = 32'h0;  // 32'h6492dd53;
    ram_cell[   15099] = 32'h0;  // 32'h3df6cf39;
    ram_cell[   15100] = 32'h0;  // 32'h9c4b505c;
    ram_cell[   15101] = 32'h0;  // 32'hc5ee4ab3;
    ram_cell[   15102] = 32'h0;  // 32'hb5d2da14;
    ram_cell[   15103] = 32'h0;  // 32'h9c2d8311;
    ram_cell[   15104] = 32'h0;  // 32'h09cb888f;
    ram_cell[   15105] = 32'h0;  // 32'h8b97dcf5;
    ram_cell[   15106] = 32'h0;  // 32'h1a617793;
    ram_cell[   15107] = 32'h0;  // 32'ha86facd0;
    ram_cell[   15108] = 32'h0;  // 32'h0a68c173;
    ram_cell[   15109] = 32'h0;  // 32'hbbba3633;
    ram_cell[   15110] = 32'h0;  // 32'h82de51f9;
    ram_cell[   15111] = 32'h0;  // 32'h04727b24;
    ram_cell[   15112] = 32'h0;  // 32'h1a1185dc;
    ram_cell[   15113] = 32'h0;  // 32'hbd709b3c;
    ram_cell[   15114] = 32'h0;  // 32'hdf2209f8;
    ram_cell[   15115] = 32'h0;  // 32'h3f6fd2c8;
    ram_cell[   15116] = 32'h0;  // 32'hd045faca;
    ram_cell[   15117] = 32'h0;  // 32'haf140bfa;
    ram_cell[   15118] = 32'h0;  // 32'h953ea803;
    ram_cell[   15119] = 32'h0;  // 32'h8b80a8eb;
    ram_cell[   15120] = 32'h0;  // 32'h465d3f9d;
    ram_cell[   15121] = 32'h0;  // 32'h247c09d8;
    ram_cell[   15122] = 32'h0;  // 32'h4a6db14b;
    ram_cell[   15123] = 32'h0;  // 32'hf4a75d71;
    ram_cell[   15124] = 32'h0;  // 32'hf44ed655;
    ram_cell[   15125] = 32'h0;  // 32'ha5b4c5ad;
    ram_cell[   15126] = 32'h0;  // 32'h4eafaf61;
    ram_cell[   15127] = 32'h0;  // 32'h6a2fcdc6;
    ram_cell[   15128] = 32'h0;  // 32'h2591522f;
    ram_cell[   15129] = 32'h0;  // 32'h14ef0846;
    ram_cell[   15130] = 32'h0;  // 32'haeb2d31d;
    ram_cell[   15131] = 32'h0;  // 32'hbfa26098;
    ram_cell[   15132] = 32'h0;  // 32'hbd3c61c0;
    ram_cell[   15133] = 32'h0;  // 32'h19352a0e;
    ram_cell[   15134] = 32'h0;  // 32'hd34c95be;
    ram_cell[   15135] = 32'h0;  // 32'h627e1c47;
    ram_cell[   15136] = 32'h0;  // 32'h8bea722c;
    ram_cell[   15137] = 32'h0;  // 32'h8c37e5ac;
    ram_cell[   15138] = 32'h0;  // 32'h9dc0015a;
    ram_cell[   15139] = 32'h0;  // 32'h8068e8c3;
    ram_cell[   15140] = 32'h0;  // 32'hb736fb19;
    ram_cell[   15141] = 32'h0;  // 32'hbf33a2cc;
    ram_cell[   15142] = 32'h0;  // 32'h30be1072;
    ram_cell[   15143] = 32'h0;  // 32'h4eb4b8f4;
    ram_cell[   15144] = 32'h0;  // 32'he3be986f;
    ram_cell[   15145] = 32'h0;  // 32'he0435381;
    ram_cell[   15146] = 32'h0;  // 32'h60ed6cd9;
    ram_cell[   15147] = 32'h0;  // 32'hca3ffceb;
    ram_cell[   15148] = 32'h0;  // 32'h2d2ffcd9;
    ram_cell[   15149] = 32'h0;  // 32'hc78ace66;
    ram_cell[   15150] = 32'h0;  // 32'h509af9b3;
    ram_cell[   15151] = 32'h0;  // 32'had162df9;
    ram_cell[   15152] = 32'h0;  // 32'h2fbdfb57;
    ram_cell[   15153] = 32'h0;  // 32'h0fcb050d;
    ram_cell[   15154] = 32'h0;  // 32'ha1e4c4f5;
    ram_cell[   15155] = 32'h0;  // 32'h38332f1d;
    ram_cell[   15156] = 32'h0;  // 32'h19d0aa45;
    ram_cell[   15157] = 32'h0;  // 32'h988a45b7;
    ram_cell[   15158] = 32'h0;  // 32'h025fef1d;
    ram_cell[   15159] = 32'h0;  // 32'h6f85c8bf;
    ram_cell[   15160] = 32'h0;  // 32'h3f7dbe47;
    ram_cell[   15161] = 32'h0;  // 32'h79fc476d;
    ram_cell[   15162] = 32'h0;  // 32'hafeeccb3;
    ram_cell[   15163] = 32'h0;  // 32'hd6ed920c;
    ram_cell[   15164] = 32'h0;  // 32'hae19f2de;
    ram_cell[   15165] = 32'h0;  // 32'h892d7428;
    ram_cell[   15166] = 32'h0;  // 32'h28812b16;
    ram_cell[   15167] = 32'h0;  // 32'heea985a0;
    ram_cell[   15168] = 32'h0;  // 32'h32632cd3;
    ram_cell[   15169] = 32'h0;  // 32'hcdbdf1e8;
    ram_cell[   15170] = 32'h0;  // 32'h22209d8a;
    ram_cell[   15171] = 32'h0;  // 32'hb1497260;
    ram_cell[   15172] = 32'h0;  // 32'h6ff5dd59;
    ram_cell[   15173] = 32'h0;  // 32'h8cd93240;
    ram_cell[   15174] = 32'h0;  // 32'h9e980ff5;
    ram_cell[   15175] = 32'h0;  // 32'ha4b83f5f;
    ram_cell[   15176] = 32'h0;  // 32'h1cabc09a;
    ram_cell[   15177] = 32'h0;  // 32'hd3e83bb7;
    ram_cell[   15178] = 32'h0;  // 32'h90be345c;
    ram_cell[   15179] = 32'h0;  // 32'hc84ba976;
    ram_cell[   15180] = 32'h0;  // 32'hef533950;
    ram_cell[   15181] = 32'h0;  // 32'h4b9537d3;
    ram_cell[   15182] = 32'h0;  // 32'h8071e506;
    ram_cell[   15183] = 32'h0;  // 32'h25560297;
    ram_cell[   15184] = 32'h0;  // 32'h84d9212c;
    ram_cell[   15185] = 32'h0;  // 32'hb1d3c9b4;
    ram_cell[   15186] = 32'h0;  // 32'hcde64024;
    ram_cell[   15187] = 32'h0;  // 32'h5fa1df38;
    ram_cell[   15188] = 32'h0;  // 32'h56e1515d;
    ram_cell[   15189] = 32'h0;  // 32'h01a87100;
    ram_cell[   15190] = 32'h0;  // 32'hc7291fe6;
    ram_cell[   15191] = 32'h0;  // 32'h20d90e82;
    ram_cell[   15192] = 32'h0;  // 32'h322f6b57;
    ram_cell[   15193] = 32'h0;  // 32'h6215eb1b;
    ram_cell[   15194] = 32'h0;  // 32'h7a75bb68;
    ram_cell[   15195] = 32'h0;  // 32'h287f73b7;
    ram_cell[   15196] = 32'h0;  // 32'h664525a8;
    ram_cell[   15197] = 32'h0;  // 32'ha3632407;
    ram_cell[   15198] = 32'h0;  // 32'h656e1b84;
    ram_cell[   15199] = 32'h0;  // 32'h0b35b2a5;
    ram_cell[   15200] = 32'h0;  // 32'hbfa801c4;
    ram_cell[   15201] = 32'h0;  // 32'hdcbb376c;
    ram_cell[   15202] = 32'h0;  // 32'h0601a4f4;
    ram_cell[   15203] = 32'h0;  // 32'hef86bcc9;
    ram_cell[   15204] = 32'h0;  // 32'h0e69270c;
    ram_cell[   15205] = 32'h0;  // 32'hf20a1837;
    ram_cell[   15206] = 32'h0;  // 32'h25e4d120;
    ram_cell[   15207] = 32'h0;  // 32'h72a98a12;
    ram_cell[   15208] = 32'h0;  // 32'h03fdca49;
    ram_cell[   15209] = 32'h0;  // 32'hdac5c277;
    ram_cell[   15210] = 32'h0;  // 32'h8ab2f198;
    ram_cell[   15211] = 32'h0;  // 32'hf0b03b97;
    ram_cell[   15212] = 32'h0;  // 32'h47e9f336;
    ram_cell[   15213] = 32'h0;  // 32'h5fdf72c4;
    ram_cell[   15214] = 32'h0;  // 32'h98ee3f10;
    ram_cell[   15215] = 32'h0;  // 32'hb5bd8211;
    ram_cell[   15216] = 32'h0;  // 32'h0ece667b;
    ram_cell[   15217] = 32'h0;  // 32'h88cf1cec;
    ram_cell[   15218] = 32'h0;  // 32'h07af893e;
    ram_cell[   15219] = 32'h0;  // 32'h608c05e0;
    ram_cell[   15220] = 32'h0;  // 32'hee8be006;
    ram_cell[   15221] = 32'h0;  // 32'h53400fc9;
    ram_cell[   15222] = 32'h0;  // 32'h5bca23d4;
    ram_cell[   15223] = 32'h0;  // 32'h49a911d7;
    ram_cell[   15224] = 32'h0;  // 32'h14a3dab7;
    ram_cell[   15225] = 32'h0;  // 32'he2ad3487;
    ram_cell[   15226] = 32'h0;  // 32'h94821169;
    ram_cell[   15227] = 32'h0;  // 32'hd4a15acd;
    ram_cell[   15228] = 32'h0;  // 32'h4ce3e9e7;
    ram_cell[   15229] = 32'h0;  // 32'h41a4fdcc;
    ram_cell[   15230] = 32'h0;  // 32'hed773cbc;
    ram_cell[   15231] = 32'h0;  // 32'h8a2b7e92;
    ram_cell[   15232] = 32'h0;  // 32'h53efcc6c;
    ram_cell[   15233] = 32'h0;  // 32'hac28f7a4;
    ram_cell[   15234] = 32'h0;  // 32'h4d8b2469;
    ram_cell[   15235] = 32'h0;  // 32'h2c5ad598;
    ram_cell[   15236] = 32'h0;  // 32'h80d050da;
    ram_cell[   15237] = 32'h0;  // 32'h40e41b1c;
    ram_cell[   15238] = 32'h0;  // 32'hd69a41e2;
    ram_cell[   15239] = 32'h0;  // 32'h79ae4f3e;
    ram_cell[   15240] = 32'h0;  // 32'h14f21d45;
    ram_cell[   15241] = 32'h0;  // 32'h716e9e80;
    ram_cell[   15242] = 32'h0;  // 32'h46f5f6a4;
    ram_cell[   15243] = 32'h0;  // 32'h7e9ccd43;
    ram_cell[   15244] = 32'h0;  // 32'hd8b6326b;
    ram_cell[   15245] = 32'h0;  // 32'heccb6c86;
    ram_cell[   15246] = 32'h0;  // 32'haf153d2e;
    ram_cell[   15247] = 32'h0;  // 32'h6bb2a8ba;
    ram_cell[   15248] = 32'h0;  // 32'h5f191cbb;
    ram_cell[   15249] = 32'h0;  // 32'h2cc2cc48;
    ram_cell[   15250] = 32'h0;  // 32'h6a1fd06d;
    ram_cell[   15251] = 32'h0;  // 32'ha59c9e33;
    ram_cell[   15252] = 32'h0;  // 32'h2834e806;
    ram_cell[   15253] = 32'h0;  // 32'hae92e7d4;
    ram_cell[   15254] = 32'h0;  // 32'h7241ad8d;
    ram_cell[   15255] = 32'h0;  // 32'hb04d3a0f;
    ram_cell[   15256] = 32'h0;  // 32'h06d15daf;
    ram_cell[   15257] = 32'h0;  // 32'hdefa0ff3;
    ram_cell[   15258] = 32'h0;  // 32'hb729d87a;
    ram_cell[   15259] = 32'h0;  // 32'h27a9abbc;
    ram_cell[   15260] = 32'h0;  // 32'h7bfaba75;
    ram_cell[   15261] = 32'h0;  // 32'hf4b06bcd;
    ram_cell[   15262] = 32'h0;  // 32'h6ffd0e45;
    ram_cell[   15263] = 32'h0;  // 32'h320f4cce;
    ram_cell[   15264] = 32'h0;  // 32'h15d24202;
    ram_cell[   15265] = 32'h0;  // 32'h143bc3c5;
    ram_cell[   15266] = 32'h0;  // 32'h9be680a0;
    ram_cell[   15267] = 32'h0;  // 32'h2adf17f2;
    ram_cell[   15268] = 32'h0;  // 32'hc054f7f5;
    ram_cell[   15269] = 32'h0;  // 32'h4784a52f;
    ram_cell[   15270] = 32'h0;  // 32'h631ff3b1;
    ram_cell[   15271] = 32'h0;  // 32'h25199138;
    ram_cell[   15272] = 32'h0;  // 32'h8b96b670;
    ram_cell[   15273] = 32'h0;  // 32'h2123ab7d;
    ram_cell[   15274] = 32'h0;  // 32'h0be2d9ab;
    ram_cell[   15275] = 32'h0;  // 32'haec5108c;
    ram_cell[   15276] = 32'h0;  // 32'h4935cddb;
    ram_cell[   15277] = 32'h0;  // 32'hd013e3d5;
    ram_cell[   15278] = 32'h0;  // 32'hd10c2bcd;
    ram_cell[   15279] = 32'h0;  // 32'h4f62e4b4;
    ram_cell[   15280] = 32'h0;  // 32'h00f17b48;
    ram_cell[   15281] = 32'h0;  // 32'h82126043;
    ram_cell[   15282] = 32'h0;  // 32'h559eab12;
    ram_cell[   15283] = 32'h0;  // 32'hf0576b63;
    ram_cell[   15284] = 32'h0;  // 32'h410c21e7;
    ram_cell[   15285] = 32'h0;  // 32'h559141c9;
    ram_cell[   15286] = 32'h0;  // 32'h8fc2f04e;
    ram_cell[   15287] = 32'h0;  // 32'h3b8e2dcd;
    ram_cell[   15288] = 32'h0;  // 32'h66d46f9c;
    ram_cell[   15289] = 32'h0;  // 32'h2ba9cbde;
    ram_cell[   15290] = 32'h0;  // 32'h9ba442b6;
    ram_cell[   15291] = 32'h0;  // 32'h25cecd1f;
    ram_cell[   15292] = 32'h0;  // 32'h693f466c;
    ram_cell[   15293] = 32'h0;  // 32'hb0452d8b;
    ram_cell[   15294] = 32'h0;  // 32'h1cbd62ef;
    ram_cell[   15295] = 32'h0;  // 32'hebad49eb;
    ram_cell[   15296] = 32'h0;  // 32'he0d26600;
    ram_cell[   15297] = 32'h0;  // 32'h73f397bf;
    ram_cell[   15298] = 32'h0;  // 32'hb2005adb;
    ram_cell[   15299] = 32'h0;  // 32'h1caf8440;
    ram_cell[   15300] = 32'h0;  // 32'h0f9d867a;
    ram_cell[   15301] = 32'h0;  // 32'h33854aa5;
    ram_cell[   15302] = 32'h0;  // 32'h3cd46d23;
    ram_cell[   15303] = 32'h0;  // 32'hab81c039;
    ram_cell[   15304] = 32'h0;  // 32'he5f8b84b;
    ram_cell[   15305] = 32'h0;  // 32'h26b50d62;
    ram_cell[   15306] = 32'h0;  // 32'h76a932a8;
    ram_cell[   15307] = 32'h0;  // 32'h609c018f;
    ram_cell[   15308] = 32'h0;  // 32'h9bee8314;
    ram_cell[   15309] = 32'h0;  // 32'h761717da;
    ram_cell[   15310] = 32'h0;  // 32'h2d2e0f59;
    ram_cell[   15311] = 32'h0;  // 32'h847a7243;
    ram_cell[   15312] = 32'h0;  // 32'h6f5d7286;
    ram_cell[   15313] = 32'h0;  // 32'h160926ea;
    ram_cell[   15314] = 32'h0;  // 32'h4ee7cf4c;
    ram_cell[   15315] = 32'h0;  // 32'h52410135;
    ram_cell[   15316] = 32'h0;  // 32'h70228f23;
    ram_cell[   15317] = 32'h0;  // 32'h52b2a486;
    ram_cell[   15318] = 32'h0;  // 32'hd1f6fffb;
    ram_cell[   15319] = 32'h0;  // 32'h98939421;
    ram_cell[   15320] = 32'h0;  // 32'hd5f7aed1;
    ram_cell[   15321] = 32'h0;  // 32'h032bc396;
    ram_cell[   15322] = 32'h0;  // 32'h28ac5135;
    ram_cell[   15323] = 32'h0;  // 32'h970f4687;
    ram_cell[   15324] = 32'h0;  // 32'hc7209d41;
    ram_cell[   15325] = 32'h0;  // 32'h064c300d;
    ram_cell[   15326] = 32'h0;  // 32'h195b12f4;
    ram_cell[   15327] = 32'h0;  // 32'h2cd948e1;
    ram_cell[   15328] = 32'h0;  // 32'h77957d32;
    ram_cell[   15329] = 32'h0;  // 32'hb353bea7;
    ram_cell[   15330] = 32'h0;  // 32'h8298984f;
    ram_cell[   15331] = 32'h0;  // 32'h5f1d3963;
    ram_cell[   15332] = 32'h0;  // 32'hdbc8896e;
    ram_cell[   15333] = 32'h0;  // 32'hcabda25e;
    ram_cell[   15334] = 32'h0;  // 32'h14c4cb7c;
    ram_cell[   15335] = 32'h0;  // 32'h36ce2ef5;
    ram_cell[   15336] = 32'h0;  // 32'h58eaa756;
    ram_cell[   15337] = 32'h0;  // 32'h8704d7df;
    ram_cell[   15338] = 32'h0;  // 32'h263d6bc9;
    ram_cell[   15339] = 32'h0;  // 32'he1368c9d;
    ram_cell[   15340] = 32'h0;  // 32'h543f63d8;
    ram_cell[   15341] = 32'h0;  // 32'h66acd870;
    ram_cell[   15342] = 32'h0;  // 32'h2e9f149a;
    ram_cell[   15343] = 32'h0;  // 32'h2bd80a90;
    ram_cell[   15344] = 32'h0;  // 32'h33afcb03;
    ram_cell[   15345] = 32'h0;  // 32'h6e8159df;
    ram_cell[   15346] = 32'h0;  // 32'h7a6da6d7;
    ram_cell[   15347] = 32'h0;  // 32'had3c69a4;
    ram_cell[   15348] = 32'h0;  // 32'h76140785;
    ram_cell[   15349] = 32'h0;  // 32'hdfb19350;
    ram_cell[   15350] = 32'h0;  // 32'h53fd7774;
    ram_cell[   15351] = 32'h0;  // 32'hf0adc52e;
    ram_cell[   15352] = 32'h0;  // 32'he318fed8;
    ram_cell[   15353] = 32'h0;  // 32'h3cba3a88;
    ram_cell[   15354] = 32'h0;  // 32'h8d40b7a8;
    ram_cell[   15355] = 32'h0;  // 32'h54e3e79c;
    ram_cell[   15356] = 32'h0;  // 32'h8af155b4;
    ram_cell[   15357] = 32'h0;  // 32'h6dd7197a;
    ram_cell[   15358] = 32'h0;  // 32'h0b74df55;
    ram_cell[   15359] = 32'h0;  // 32'hba0668db;
    ram_cell[   15360] = 32'h0;  // 32'h14ea4100;
    ram_cell[   15361] = 32'h0;  // 32'hc000065b;
    ram_cell[   15362] = 32'h0;  // 32'h91b5d707;
    ram_cell[   15363] = 32'h0;  // 32'hc41f359c;
    ram_cell[   15364] = 32'h0;  // 32'h6142fc32;
    ram_cell[   15365] = 32'h0;  // 32'h3dbdb8de;
    ram_cell[   15366] = 32'h0;  // 32'hc7c6b307;
    ram_cell[   15367] = 32'h0;  // 32'hf1be2602;
    ram_cell[   15368] = 32'h0;  // 32'hf2e7ab98;
    ram_cell[   15369] = 32'h0;  // 32'he869310d;
    ram_cell[   15370] = 32'h0;  // 32'h9e015c50;
    ram_cell[   15371] = 32'h0;  // 32'hd03e50a9;
    ram_cell[   15372] = 32'h0;  // 32'h1889c2eb;
    ram_cell[   15373] = 32'h0;  // 32'h67d2aa71;
    ram_cell[   15374] = 32'h0;  // 32'h0157eed8;
    ram_cell[   15375] = 32'h0;  // 32'ha2ff1249;
    ram_cell[   15376] = 32'h0;  // 32'hd5a6f43b;
    ram_cell[   15377] = 32'h0;  // 32'h372d8d87;
    ram_cell[   15378] = 32'h0;  // 32'h9075e521;
    ram_cell[   15379] = 32'h0;  // 32'hb76af0d0;
    ram_cell[   15380] = 32'h0;  // 32'h489d715d;
    ram_cell[   15381] = 32'h0;  // 32'hbbb4a20b;
    ram_cell[   15382] = 32'h0;  // 32'h308020f3;
    ram_cell[   15383] = 32'h0;  // 32'haeca4550;
    ram_cell[   15384] = 32'h0;  // 32'h338e8fe4;
    ram_cell[   15385] = 32'h0;  // 32'h12840c21;
    ram_cell[   15386] = 32'h0;  // 32'hf6beaf23;
    ram_cell[   15387] = 32'h0;  // 32'h53ccc05b;
    ram_cell[   15388] = 32'h0;  // 32'h4e3bf660;
    ram_cell[   15389] = 32'h0;  // 32'h524a391d;
    ram_cell[   15390] = 32'h0;  // 32'h6657cde3;
    ram_cell[   15391] = 32'h0;  // 32'h4c7e6ce4;
    ram_cell[   15392] = 32'h0;  // 32'hd2e99954;
    ram_cell[   15393] = 32'h0;  // 32'hf693e4e0;
    ram_cell[   15394] = 32'h0;  // 32'hdaaa6b44;
    ram_cell[   15395] = 32'h0;  // 32'hb24f277c;
    ram_cell[   15396] = 32'h0;  // 32'h95ed2bf1;
    ram_cell[   15397] = 32'h0;  // 32'h27f33531;
    ram_cell[   15398] = 32'h0;  // 32'h73cb34e5;
    ram_cell[   15399] = 32'h0;  // 32'h3c2f196c;
    ram_cell[   15400] = 32'h0;  // 32'h2f1daf6a;
    ram_cell[   15401] = 32'h0;  // 32'h26c69476;
    ram_cell[   15402] = 32'h0;  // 32'heb96f619;
    ram_cell[   15403] = 32'h0;  // 32'hc8cbade1;
    ram_cell[   15404] = 32'h0;  // 32'h890f240b;
    ram_cell[   15405] = 32'h0;  // 32'hbfccc479;
    ram_cell[   15406] = 32'h0;  // 32'h209376f0;
    ram_cell[   15407] = 32'h0;  // 32'h039c4441;
    ram_cell[   15408] = 32'h0;  // 32'he049f7f0;
    ram_cell[   15409] = 32'h0;  // 32'h6b9f7b46;
    ram_cell[   15410] = 32'h0;  // 32'h026fb256;
    ram_cell[   15411] = 32'h0;  // 32'h1df9c2bc;
    ram_cell[   15412] = 32'h0;  // 32'hadc0bd78;
    ram_cell[   15413] = 32'h0;  // 32'h1e28c8b6;
    ram_cell[   15414] = 32'h0;  // 32'hecc68f75;
    ram_cell[   15415] = 32'h0;  // 32'h1b5c52a0;
    ram_cell[   15416] = 32'h0;  // 32'h550fa22a;
    ram_cell[   15417] = 32'h0;  // 32'ha12e6e72;
    ram_cell[   15418] = 32'h0;  // 32'h766126ce;
    ram_cell[   15419] = 32'h0;  // 32'h68e88c58;
    ram_cell[   15420] = 32'h0;  // 32'ha0e2e663;
    ram_cell[   15421] = 32'h0;  // 32'h14280e92;
    ram_cell[   15422] = 32'h0;  // 32'h47b5491f;
    ram_cell[   15423] = 32'h0;  // 32'h642560e0;
    ram_cell[   15424] = 32'h0;  // 32'ha81592d0;
    ram_cell[   15425] = 32'h0;  // 32'h76a3fc85;
    ram_cell[   15426] = 32'h0;  // 32'h70d985b7;
    ram_cell[   15427] = 32'h0;  // 32'h71a80cec;
    ram_cell[   15428] = 32'h0;  // 32'h5ddb5c03;
    ram_cell[   15429] = 32'h0;  // 32'hfdd0775c;
    ram_cell[   15430] = 32'h0;  // 32'hd45d474e;
    ram_cell[   15431] = 32'h0;  // 32'hb59148ef;
    ram_cell[   15432] = 32'h0;  // 32'h3f7189f7;
    ram_cell[   15433] = 32'h0;  // 32'h9502e95d;
    ram_cell[   15434] = 32'h0;  // 32'hdfc7efe3;
    ram_cell[   15435] = 32'h0;  // 32'h7f5b5160;
    ram_cell[   15436] = 32'h0;  // 32'hf37d2480;
    ram_cell[   15437] = 32'h0;  // 32'hc4e3bf63;
    ram_cell[   15438] = 32'h0;  // 32'h208b8a7c;
    ram_cell[   15439] = 32'h0;  // 32'h0246705e;
    ram_cell[   15440] = 32'h0;  // 32'h29bde62d;
    ram_cell[   15441] = 32'h0;  // 32'hf4bd93b1;
    ram_cell[   15442] = 32'h0;  // 32'heecbe050;
    ram_cell[   15443] = 32'h0;  // 32'h9cefde53;
    ram_cell[   15444] = 32'h0;  // 32'heb94dc97;
    ram_cell[   15445] = 32'h0;  // 32'h5de235b5;
    ram_cell[   15446] = 32'h0;  // 32'h52016842;
    ram_cell[   15447] = 32'h0;  // 32'hc935924d;
    ram_cell[   15448] = 32'h0;  // 32'hcdfa9c5a;
    ram_cell[   15449] = 32'h0;  // 32'h08acc5f6;
    ram_cell[   15450] = 32'h0;  // 32'h8782b9bb;
    ram_cell[   15451] = 32'h0;  // 32'h0b29de9f;
    ram_cell[   15452] = 32'h0;  // 32'h1b0dc158;
    ram_cell[   15453] = 32'h0;  // 32'h8f8d09ae;
    ram_cell[   15454] = 32'h0;  // 32'he4c499bc;
    ram_cell[   15455] = 32'h0;  // 32'h3a447828;
    ram_cell[   15456] = 32'h0;  // 32'h18860004;
    ram_cell[   15457] = 32'h0;  // 32'hc3ec4492;
    ram_cell[   15458] = 32'h0;  // 32'ha0b5315a;
    ram_cell[   15459] = 32'h0;  // 32'hf6605800;
    ram_cell[   15460] = 32'h0;  // 32'ha14b3f8a;
    ram_cell[   15461] = 32'h0;  // 32'h4ed542d6;
    ram_cell[   15462] = 32'h0;  // 32'h0942b27c;
    ram_cell[   15463] = 32'h0;  // 32'hc9cdce18;
    ram_cell[   15464] = 32'h0;  // 32'h5282d6b4;
    ram_cell[   15465] = 32'h0;  // 32'h2f11b4bd;
    ram_cell[   15466] = 32'h0;  // 32'h8e88a9c7;
    ram_cell[   15467] = 32'h0;  // 32'h6d8ccb27;
    ram_cell[   15468] = 32'h0;  // 32'hf68fd25a;
    ram_cell[   15469] = 32'h0;  // 32'h0d46bc3b;
    ram_cell[   15470] = 32'h0;  // 32'h15d0528f;
    ram_cell[   15471] = 32'h0;  // 32'h0e3b0f11;
    ram_cell[   15472] = 32'h0;  // 32'h1874c201;
    ram_cell[   15473] = 32'h0;  // 32'h8b232b38;
    ram_cell[   15474] = 32'h0;  // 32'h16f68e9d;
    ram_cell[   15475] = 32'h0;  // 32'h22a459fa;
    ram_cell[   15476] = 32'h0;  // 32'h489fd603;
    ram_cell[   15477] = 32'h0;  // 32'h10f61ecc;
    ram_cell[   15478] = 32'h0;  // 32'h7476a256;
    ram_cell[   15479] = 32'h0;  // 32'hb11e6e71;
    ram_cell[   15480] = 32'h0;  // 32'h26ba0659;
    ram_cell[   15481] = 32'h0;  // 32'h0ec91ddc;
    ram_cell[   15482] = 32'h0;  // 32'h8dd3bb34;
    ram_cell[   15483] = 32'h0;  // 32'h8117929b;
    ram_cell[   15484] = 32'h0;  // 32'h5ef38cda;
    ram_cell[   15485] = 32'h0;  // 32'h3c1ac772;
    ram_cell[   15486] = 32'h0;  // 32'hd8a2eab3;
    ram_cell[   15487] = 32'h0;  // 32'hcbb825bf;
    ram_cell[   15488] = 32'h0;  // 32'h5119c5a2;
    ram_cell[   15489] = 32'h0;  // 32'h0b3290b1;
    ram_cell[   15490] = 32'h0;  // 32'h369dd4e8;
    ram_cell[   15491] = 32'h0;  // 32'h27de01d4;
    ram_cell[   15492] = 32'h0;  // 32'h586d21ba;
    ram_cell[   15493] = 32'h0;  // 32'hbb75f112;
    ram_cell[   15494] = 32'h0;  // 32'h38b7f154;
    ram_cell[   15495] = 32'h0;  // 32'h0a2b1740;
    ram_cell[   15496] = 32'h0;  // 32'h16f58838;
    ram_cell[   15497] = 32'h0;  // 32'h83a54c55;
    ram_cell[   15498] = 32'h0;  // 32'h0b88b2d0;
    ram_cell[   15499] = 32'h0;  // 32'h379884b4;
    ram_cell[   15500] = 32'h0;  // 32'h286ba2ea;
    ram_cell[   15501] = 32'h0;  // 32'h9441ad15;
    ram_cell[   15502] = 32'h0;  // 32'h4ed3c7ca;
    ram_cell[   15503] = 32'h0;  // 32'h377525d9;
    ram_cell[   15504] = 32'h0;  // 32'h2df79ef2;
    ram_cell[   15505] = 32'h0;  // 32'hdcd04da8;
    ram_cell[   15506] = 32'h0;  // 32'h16e020a6;
    ram_cell[   15507] = 32'h0;  // 32'h874705fc;
    ram_cell[   15508] = 32'h0;  // 32'hdb4bbc7c;
    ram_cell[   15509] = 32'h0;  // 32'hf63e1308;
    ram_cell[   15510] = 32'h0;  // 32'hca309f49;
    ram_cell[   15511] = 32'h0;  // 32'h44107146;
    ram_cell[   15512] = 32'h0;  // 32'h59a6463e;
    ram_cell[   15513] = 32'h0;  // 32'h6bbb1049;
    ram_cell[   15514] = 32'h0;  // 32'h7eab833f;
    ram_cell[   15515] = 32'h0;  // 32'hb2e87edd;
    ram_cell[   15516] = 32'h0;  // 32'h2f253421;
    ram_cell[   15517] = 32'h0;  // 32'h89767089;
    ram_cell[   15518] = 32'h0;  // 32'he2457cf8;
    ram_cell[   15519] = 32'h0;  // 32'h67f79aee;
    ram_cell[   15520] = 32'h0;  // 32'h183181b5;
    ram_cell[   15521] = 32'h0;  // 32'h71bb6a23;
    ram_cell[   15522] = 32'h0;  // 32'h8c09fa0b;
    ram_cell[   15523] = 32'h0;  // 32'h156510bd;
    ram_cell[   15524] = 32'h0;  // 32'hea064dae;
    ram_cell[   15525] = 32'h0;  // 32'h62ee11bf;
    ram_cell[   15526] = 32'h0;  // 32'h03e187e6;
    ram_cell[   15527] = 32'h0;  // 32'h9c4c5d52;
    ram_cell[   15528] = 32'h0;  // 32'haa46ed2f;
    ram_cell[   15529] = 32'h0;  // 32'h3c05ba44;
    ram_cell[   15530] = 32'h0;  // 32'h461cc5e2;
    ram_cell[   15531] = 32'h0;  // 32'h89ecd4e1;
    ram_cell[   15532] = 32'h0;  // 32'hdf179548;
    ram_cell[   15533] = 32'h0;  // 32'h1e3d923b;
    ram_cell[   15534] = 32'h0;  // 32'h0c6e2c7e;
    ram_cell[   15535] = 32'h0;  // 32'hd77c360b;
    ram_cell[   15536] = 32'h0;  // 32'he1e22705;
    ram_cell[   15537] = 32'h0;  // 32'hb4cbd2cc;
    ram_cell[   15538] = 32'h0;  // 32'he03fe81c;
    ram_cell[   15539] = 32'h0;  // 32'h6a797c95;
    ram_cell[   15540] = 32'h0;  // 32'hec8b9ef0;
    ram_cell[   15541] = 32'h0;  // 32'h1c528dec;
    ram_cell[   15542] = 32'h0;  // 32'h95d222d9;
    ram_cell[   15543] = 32'h0;  // 32'h1fc5c6bd;
    ram_cell[   15544] = 32'h0;  // 32'h18c300fa;
    ram_cell[   15545] = 32'h0;  // 32'hc222eb6e;
    ram_cell[   15546] = 32'h0;  // 32'hcf9f8a58;
    ram_cell[   15547] = 32'h0;  // 32'hf64cd69d;
    ram_cell[   15548] = 32'h0;  // 32'h8c4853e3;
    ram_cell[   15549] = 32'h0;  // 32'h7e0d978a;
    ram_cell[   15550] = 32'h0;  // 32'h2a3b0127;
    ram_cell[   15551] = 32'h0;  // 32'h1b5f9a9c;
    ram_cell[   15552] = 32'h0;  // 32'hbcd573db;
    ram_cell[   15553] = 32'h0;  // 32'h2a75092f;
    ram_cell[   15554] = 32'h0;  // 32'h45075603;
    ram_cell[   15555] = 32'h0;  // 32'h1f2f47a2;
    ram_cell[   15556] = 32'h0;  // 32'h064a8432;
    ram_cell[   15557] = 32'h0;  // 32'h9aed9c52;
    ram_cell[   15558] = 32'h0;  // 32'hccb3c828;
    ram_cell[   15559] = 32'h0;  // 32'he0f41a3a;
    ram_cell[   15560] = 32'h0;  // 32'h7d59c3f4;
    ram_cell[   15561] = 32'h0;  // 32'h4035a8e7;
    ram_cell[   15562] = 32'h0;  // 32'he41607a2;
    ram_cell[   15563] = 32'h0;  // 32'hef54d5e0;
    ram_cell[   15564] = 32'h0;  // 32'he600b137;
    ram_cell[   15565] = 32'h0;  // 32'hc8e7b2c1;
    ram_cell[   15566] = 32'h0;  // 32'h8fe0320f;
    ram_cell[   15567] = 32'h0;  // 32'h7a0b6c94;
    ram_cell[   15568] = 32'h0;  // 32'ha4da6b0d;
    ram_cell[   15569] = 32'h0;  // 32'h24f8c8e8;
    ram_cell[   15570] = 32'h0;  // 32'h0eb7309c;
    ram_cell[   15571] = 32'h0;  // 32'hfcbe3912;
    ram_cell[   15572] = 32'h0;  // 32'ha31241da;
    ram_cell[   15573] = 32'h0;  // 32'h1dc4ff20;
    ram_cell[   15574] = 32'h0;  // 32'h8db29b2c;
    ram_cell[   15575] = 32'h0;  // 32'h95807dcc;
    ram_cell[   15576] = 32'h0;  // 32'h530f493e;
    ram_cell[   15577] = 32'h0;  // 32'hc7e49ab1;
    ram_cell[   15578] = 32'h0;  // 32'h1a7274ed;
    ram_cell[   15579] = 32'h0;  // 32'hb22d9f72;
    ram_cell[   15580] = 32'h0;  // 32'he7c3e0af;
    ram_cell[   15581] = 32'h0;  // 32'h21c6e0ca;
    ram_cell[   15582] = 32'h0;  // 32'he319bed6;
    ram_cell[   15583] = 32'h0;  // 32'h62a7af79;
    ram_cell[   15584] = 32'h0;  // 32'ha86f1403;
    ram_cell[   15585] = 32'h0;  // 32'ha008d445;
    ram_cell[   15586] = 32'h0;  // 32'h61f2f204;
    ram_cell[   15587] = 32'h0;  // 32'h1048a2a5;
    ram_cell[   15588] = 32'h0;  // 32'h77c91345;
    ram_cell[   15589] = 32'h0;  // 32'h691f3e1b;
    ram_cell[   15590] = 32'h0;  // 32'hc9ef47b5;
    ram_cell[   15591] = 32'h0;  // 32'h3ae09244;
    ram_cell[   15592] = 32'h0;  // 32'hf3a0232e;
    ram_cell[   15593] = 32'h0;  // 32'h22751548;
    ram_cell[   15594] = 32'h0;  // 32'hf61c6c9c;
    ram_cell[   15595] = 32'h0;  // 32'hbd53329f;
    ram_cell[   15596] = 32'h0;  // 32'h93804aaf;
    ram_cell[   15597] = 32'h0;  // 32'h59cf7d93;
    ram_cell[   15598] = 32'h0;  // 32'h564ac6b5;
    ram_cell[   15599] = 32'h0;  // 32'h967e7943;
    ram_cell[   15600] = 32'h0;  // 32'ha8ace5d9;
    ram_cell[   15601] = 32'h0;  // 32'h05f26091;
    ram_cell[   15602] = 32'h0;  // 32'hba366c1a;
    ram_cell[   15603] = 32'h0;  // 32'hc20e7785;
    ram_cell[   15604] = 32'h0;  // 32'hab6d99ea;
    ram_cell[   15605] = 32'h0;  // 32'hbc112de7;
    ram_cell[   15606] = 32'h0;  // 32'h7253bcb6;
    ram_cell[   15607] = 32'h0;  // 32'h76a5b712;
    ram_cell[   15608] = 32'h0;  // 32'h4beb055c;
    ram_cell[   15609] = 32'h0;  // 32'hd689d7bf;
    ram_cell[   15610] = 32'h0;  // 32'hf770a1c8;
    ram_cell[   15611] = 32'h0;  // 32'hfe6076df;
    ram_cell[   15612] = 32'h0;  // 32'ha8f4f812;
    ram_cell[   15613] = 32'h0;  // 32'h35fa2388;
    ram_cell[   15614] = 32'h0;  // 32'h78ff0241;
    ram_cell[   15615] = 32'h0;  // 32'hda49dd84;
    ram_cell[   15616] = 32'h0;  // 32'h94109423;
    ram_cell[   15617] = 32'h0;  // 32'h48d2c6e4;
    ram_cell[   15618] = 32'h0;  // 32'ha201b6df;
    ram_cell[   15619] = 32'h0;  // 32'hb9812b43;
    ram_cell[   15620] = 32'h0;  // 32'h6205c6ee;
    ram_cell[   15621] = 32'h0;  // 32'h9aa01d41;
    ram_cell[   15622] = 32'h0;  // 32'h440cc7df;
    ram_cell[   15623] = 32'h0;  // 32'hb5d3c028;
    ram_cell[   15624] = 32'h0;  // 32'hbc88dab9;
    ram_cell[   15625] = 32'h0;  // 32'h8db6418d;
    ram_cell[   15626] = 32'h0;  // 32'h0375a47a;
    ram_cell[   15627] = 32'h0;  // 32'h0c4037d4;
    ram_cell[   15628] = 32'h0;  // 32'h6d182241;
    ram_cell[   15629] = 32'h0;  // 32'he6b91908;
    ram_cell[   15630] = 32'h0;  // 32'hea1cc3cf;
    ram_cell[   15631] = 32'h0;  // 32'hd55fce40;
    ram_cell[   15632] = 32'h0;  // 32'h87531e9e;
    ram_cell[   15633] = 32'h0;  // 32'hfeb02699;
    ram_cell[   15634] = 32'h0;  // 32'h85897b4b;
    ram_cell[   15635] = 32'h0;  // 32'h874f7f7a;
    ram_cell[   15636] = 32'h0;  // 32'hd369e8de;
    ram_cell[   15637] = 32'h0;  // 32'h7bfbcc28;
    ram_cell[   15638] = 32'h0;  // 32'h85a5143c;
    ram_cell[   15639] = 32'h0;  // 32'hba9df449;
    ram_cell[   15640] = 32'h0;  // 32'h8f870878;
    ram_cell[   15641] = 32'h0;  // 32'h49874d61;
    ram_cell[   15642] = 32'h0;  // 32'h55d89137;
    ram_cell[   15643] = 32'h0;  // 32'hc03ea36a;
    ram_cell[   15644] = 32'h0;  // 32'hbda2f0c8;
    ram_cell[   15645] = 32'h0;  // 32'h6d2e1103;
    ram_cell[   15646] = 32'h0;  // 32'ha237dbac;
    ram_cell[   15647] = 32'h0;  // 32'hc8105faf;
    ram_cell[   15648] = 32'h0;  // 32'h8af4893a;
    ram_cell[   15649] = 32'h0;  // 32'ha45d76fe;
    ram_cell[   15650] = 32'h0;  // 32'h33b2a994;
    ram_cell[   15651] = 32'h0;  // 32'hf5c036fb;
    ram_cell[   15652] = 32'h0;  // 32'h163cb29a;
    ram_cell[   15653] = 32'h0;  // 32'h3bf2825e;
    ram_cell[   15654] = 32'h0;  // 32'hacc5e007;
    ram_cell[   15655] = 32'h0;  // 32'heffe2992;
    ram_cell[   15656] = 32'h0;  // 32'ha5c611fe;
    ram_cell[   15657] = 32'h0;  // 32'hdde0c1c5;
    ram_cell[   15658] = 32'h0;  // 32'h4196ac36;
    ram_cell[   15659] = 32'h0;  // 32'h4ff0fac6;
    ram_cell[   15660] = 32'h0;  // 32'h0c916fe2;
    ram_cell[   15661] = 32'h0;  // 32'h9af29e02;
    ram_cell[   15662] = 32'h0;  // 32'hb17953a6;
    ram_cell[   15663] = 32'h0;  // 32'hf47040e4;
    ram_cell[   15664] = 32'h0;  // 32'h469437a7;
    ram_cell[   15665] = 32'h0;  // 32'h51da7559;
    ram_cell[   15666] = 32'h0;  // 32'hc53922e4;
    ram_cell[   15667] = 32'h0;  // 32'he8793bb1;
    ram_cell[   15668] = 32'h0;  // 32'h11ee937d;
    ram_cell[   15669] = 32'h0;  // 32'heac74583;
    ram_cell[   15670] = 32'h0;  // 32'h1e5e935e;
    ram_cell[   15671] = 32'h0;  // 32'h44278f3d;
    ram_cell[   15672] = 32'h0;  // 32'h798737ae;
    ram_cell[   15673] = 32'h0;  // 32'h8aaaec9f;
    ram_cell[   15674] = 32'h0;  // 32'hc68e73df;
    ram_cell[   15675] = 32'h0;  // 32'hc5b6cdee;
    ram_cell[   15676] = 32'h0;  // 32'h55cd710c;
    ram_cell[   15677] = 32'h0;  // 32'h2ce29fb4;
    ram_cell[   15678] = 32'h0;  // 32'hbb04e523;
    ram_cell[   15679] = 32'h0;  // 32'h0ba8f4c1;
    ram_cell[   15680] = 32'h0;  // 32'hd2b4a3ba;
    ram_cell[   15681] = 32'h0;  // 32'h9837963e;
    ram_cell[   15682] = 32'h0;  // 32'h0512d2e0;
    ram_cell[   15683] = 32'h0;  // 32'hc80fbbcf;
    ram_cell[   15684] = 32'h0;  // 32'h9807242b;
    ram_cell[   15685] = 32'h0;  // 32'hfcfacd47;
    ram_cell[   15686] = 32'h0;  // 32'h95435572;
    ram_cell[   15687] = 32'h0;  // 32'ha98dbc68;
    ram_cell[   15688] = 32'h0;  // 32'h5ad7131f;
    ram_cell[   15689] = 32'h0;  // 32'h106f2e5a;
    ram_cell[   15690] = 32'h0;  // 32'h11a724c3;
    ram_cell[   15691] = 32'h0;  // 32'hce02765f;
    ram_cell[   15692] = 32'h0;  // 32'h8ec951d0;
    ram_cell[   15693] = 32'h0;  // 32'hf8411736;
    ram_cell[   15694] = 32'h0;  // 32'h568f65ee;
    ram_cell[   15695] = 32'h0;  // 32'h8366e0e2;
    ram_cell[   15696] = 32'h0;  // 32'h1febaaba;
    ram_cell[   15697] = 32'h0;  // 32'h55758b54;
    ram_cell[   15698] = 32'h0;  // 32'h25adfe0f;
    ram_cell[   15699] = 32'h0;  // 32'ha0be34c9;
    ram_cell[   15700] = 32'h0;  // 32'hf8e7743b;
    ram_cell[   15701] = 32'h0;  // 32'h3531b310;
    ram_cell[   15702] = 32'h0;  // 32'h7afa7a91;
    ram_cell[   15703] = 32'h0;  // 32'ha17c389a;
    ram_cell[   15704] = 32'h0;  // 32'hb8c6514a;
    ram_cell[   15705] = 32'h0;  // 32'h0e326902;
    ram_cell[   15706] = 32'h0;  // 32'hee45d5d6;
    ram_cell[   15707] = 32'h0;  // 32'h9513df0c;
    ram_cell[   15708] = 32'h0;  // 32'h3d2e3828;
    ram_cell[   15709] = 32'h0;  // 32'h89dce2b6;
    ram_cell[   15710] = 32'h0;  // 32'h51432285;
    ram_cell[   15711] = 32'h0;  // 32'h129280de;
    ram_cell[   15712] = 32'h0;  // 32'h0b3a9eb4;
    ram_cell[   15713] = 32'h0;  // 32'h9036df48;
    ram_cell[   15714] = 32'h0;  // 32'he78239ef;
    ram_cell[   15715] = 32'h0;  // 32'h5da7f211;
    ram_cell[   15716] = 32'h0;  // 32'hb49396f4;
    ram_cell[   15717] = 32'h0;  // 32'ha01e8504;
    ram_cell[   15718] = 32'h0;  // 32'h379aad0f;
    ram_cell[   15719] = 32'h0;  // 32'he9533496;
    ram_cell[   15720] = 32'h0;  // 32'h59b4f332;
    ram_cell[   15721] = 32'h0;  // 32'h549f984d;
    ram_cell[   15722] = 32'h0;  // 32'h5ab314bd;
    ram_cell[   15723] = 32'h0;  // 32'h2c4d5d2b;
    ram_cell[   15724] = 32'h0;  // 32'hbd377467;
    ram_cell[   15725] = 32'h0;  // 32'hc31d6995;
    ram_cell[   15726] = 32'h0;  // 32'hfd871c13;
    ram_cell[   15727] = 32'h0;  // 32'hee3fc8e5;
    ram_cell[   15728] = 32'h0;  // 32'h4a41b657;
    ram_cell[   15729] = 32'h0;  // 32'hffa57a56;
    ram_cell[   15730] = 32'h0;  // 32'hd193c1c0;
    ram_cell[   15731] = 32'h0;  // 32'ha944b5fa;
    ram_cell[   15732] = 32'h0;  // 32'h6beebdc7;
    ram_cell[   15733] = 32'h0;  // 32'h4a326988;
    ram_cell[   15734] = 32'h0;  // 32'h842485fe;
    ram_cell[   15735] = 32'h0;  // 32'he52c5aa8;
    ram_cell[   15736] = 32'h0;  // 32'h81106b43;
    ram_cell[   15737] = 32'h0;  // 32'h4447f202;
    ram_cell[   15738] = 32'h0;  // 32'h3b787028;
    ram_cell[   15739] = 32'h0;  // 32'hf7adba23;
    ram_cell[   15740] = 32'h0;  // 32'h31075864;
    ram_cell[   15741] = 32'h0;  // 32'h73a6fd94;
    ram_cell[   15742] = 32'h0;  // 32'h6eadd128;
    ram_cell[   15743] = 32'h0;  // 32'h2abe1132;
    ram_cell[   15744] = 32'h0;  // 32'h87ecded3;
    ram_cell[   15745] = 32'h0;  // 32'hff3dad6d;
    ram_cell[   15746] = 32'h0;  // 32'hf9c61ae3;
    ram_cell[   15747] = 32'h0;  // 32'hb8f47ed5;
    ram_cell[   15748] = 32'h0;  // 32'h5a12e6dd;
    ram_cell[   15749] = 32'h0;  // 32'h365e9c0a;
    ram_cell[   15750] = 32'h0;  // 32'hfc7e1051;
    ram_cell[   15751] = 32'h0;  // 32'h7898d97f;
    ram_cell[   15752] = 32'h0;  // 32'h91169582;
    ram_cell[   15753] = 32'h0;  // 32'hd3829002;
    ram_cell[   15754] = 32'h0;  // 32'h3f373742;
    ram_cell[   15755] = 32'h0;  // 32'haf7f5970;
    ram_cell[   15756] = 32'h0;  // 32'hed1ef504;
    ram_cell[   15757] = 32'h0;  // 32'h8c91eaba;
    ram_cell[   15758] = 32'h0;  // 32'h31477539;
    ram_cell[   15759] = 32'h0;  // 32'ha33dfc55;
    ram_cell[   15760] = 32'h0;  // 32'h87deff5a;
    ram_cell[   15761] = 32'h0;  // 32'hd505297d;
    ram_cell[   15762] = 32'h0;  // 32'h7f4c3311;
    ram_cell[   15763] = 32'h0;  // 32'h09bf2e15;
    ram_cell[   15764] = 32'h0;  // 32'h48d347cf;
    ram_cell[   15765] = 32'h0;  // 32'haa848de3;
    ram_cell[   15766] = 32'h0;  // 32'hc60fd421;
    ram_cell[   15767] = 32'h0;  // 32'h73c6b1ca;
    ram_cell[   15768] = 32'h0;  // 32'hd836efc5;
    ram_cell[   15769] = 32'h0;  // 32'hafa0a904;
    ram_cell[   15770] = 32'h0;  // 32'hdae07720;
    ram_cell[   15771] = 32'h0;  // 32'hb27cfca5;
    ram_cell[   15772] = 32'h0;  // 32'h3adfd1c2;
    ram_cell[   15773] = 32'h0;  // 32'h6d97cfe5;
    ram_cell[   15774] = 32'h0;  // 32'h13077f81;
    ram_cell[   15775] = 32'h0;  // 32'h06f047d9;
    ram_cell[   15776] = 32'h0;  // 32'h480fae5f;
    ram_cell[   15777] = 32'h0;  // 32'h88310b85;
    ram_cell[   15778] = 32'h0;  // 32'h997336b6;
    ram_cell[   15779] = 32'h0;  // 32'h2fafeb17;
    ram_cell[   15780] = 32'h0;  // 32'hba74340c;
    ram_cell[   15781] = 32'h0;  // 32'ha52744cc;
    ram_cell[   15782] = 32'h0;  // 32'h308648b3;
    ram_cell[   15783] = 32'h0;  // 32'h00bf2af3;
    ram_cell[   15784] = 32'h0;  // 32'h8d12436d;
    ram_cell[   15785] = 32'h0;  // 32'hd7f5a85d;
    ram_cell[   15786] = 32'h0;  // 32'hc0a1b546;
    ram_cell[   15787] = 32'h0;  // 32'hd7f99bca;
    ram_cell[   15788] = 32'h0;  // 32'h7299f883;
    ram_cell[   15789] = 32'h0;  // 32'h86ce31b7;
    ram_cell[   15790] = 32'h0;  // 32'h9327cccf;
    ram_cell[   15791] = 32'h0;  // 32'h32bb4e6d;
    ram_cell[   15792] = 32'h0;  // 32'h81892e34;
    ram_cell[   15793] = 32'h0;  // 32'h1f929eb0;
    ram_cell[   15794] = 32'h0;  // 32'h7b6a94ed;
    ram_cell[   15795] = 32'h0;  // 32'hd7276eff;
    ram_cell[   15796] = 32'h0;  // 32'h78865d67;
    ram_cell[   15797] = 32'h0;  // 32'h391bea83;
    ram_cell[   15798] = 32'h0;  // 32'hd8800b44;
    ram_cell[   15799] = 32'h0;  // 32'h21fa5e41;
    ram_cell[   15800] = 32'h0;  // 32'h3c788f1e;
    ram_cell[   15801] = 32'h0;  // 32'h8be088a1;
    ram_cell[   15802] = 32'h0;  // 32'had4132a7;
    ram_cell[   15803] = 32'h0;  // 32'h45aea03f;
    ram_cell[   15804] = 32'h0;  // 32'h2acca737;
    ram_cell[   15805] = 32'h0;  // 32'h4326b007;
    ram_cell[   15806] = 32'h0;  // 32'h57f5fc66;
    ram_cell[   15807] = 32'h0;  // 32'h3fd4c8c9;
    ram_cell[   15808] = 32'h0;  // 32'h3b5848ec;
    ram_cell[   15809] = 32'h0;  // 32'hf8c77fd7;
    ram_cell[   15810] = 32'h0;  // 32'hcd40d141;
    ram_cell[   15811] = 32'h0;  // 32'h79754254;
    ram_cell[   15812] = 32'h0;  // 32'h57280f4e;
    ram_cell[   15813] = 32'h0;  // 32'h88bac2fc;
    ram_cell[   15814] = 32'h0;  // 32'h1f10c0e9;
    ram_cell[   15815] = 32'h0;  // 32'heca3fb75;
    ram_cell[   15816] = 32'h0;  // 32'h6ebb2ab9;
    ram_cell[   15817] = 32'h0;  // 32'h02a8117a;
    ram_cell[   15818] = 32'h0;  // 32'h9c60e482;
    ram_cell[   15819] = 32'h0;  // 32'h9a8fab72;
    ram_cell[   15820] = 32'h0;  // 32'h6a0656e2;
    ram_cell[   15821] = 32'h0;  // 32'h46b02ad0;
    ram_cell[   15822] = 32'h0;  // 32'h14a76ff3;
    ram_cell[   15823] = 32'h0;  // 32'h1f1a7556;
    ram_cell[   15824] = 32'h0;  // 32'h03fd6024;
    ram_cell[   15825] = 32'h0;  // 32'h46ef4022;
    ram_cell[   15826] = 32'h0;  // 32'h7cf51aec;
    ram_cell[   15827] = 32'h0;  // 32'h84a79386;
    ram_cell[   15828] = 32'h0;  // 32'h49b824bc;
    ram_cell[   15829] = 32'h0;  // 32'ha23cd458;
    ram_cell[   15830] = 32'h0;  // 32'hf4d659d8;
    ram_cell[   15831] = 32'h0;  // 32'h1d84f327;
    ram_cell[   15832] = 32'h0;  // 32'h1d39f797;
    ram_cell[   15833] = 32'h0;  // 32'h6405c09c;
    ram_cell[   15834] = 32'h0;  // 32'h3a3de915;
    ram_cell[   15835] = 32'h0;  // 32'h11d37721;
    ram_cell[   15836] = 32'h0;  // 32'hb3891246;
    ram_cell[   15837] = 32'h0;  // 32'h0f66f890;
    ram_cell[   15838] = 32'h0;  // 32'h5ae1c4f0;
    ram_cell[   15839] = 32'h0;  // 32'h4e588cfc;
    ram_cell[   15840] = 32'h0;  // 32'hf64a3884;
    ram_cell[   15841] = 32'h0;  // 32'h17db6aff;
    ram_cell[   15842] = 32'h0;  // 32'he38085f8;
    ram_cell[   15843] = 32'h0;  // 32'h99ed36ab;
    ram_cell[   15844] = 32'h0;  // 32'h4eec0087;
    ram_cell[   15845] = 32'h0;  // 32'he673f5d2;
    ram_cell[   15846] = 32'h0;  // 32'hd2280916;
    ram_cell[   15847] = 32'h0;  // 32'h680c0c4a;
    ram_cell[   15848] = 32'h0;  // 32'h4c957c5f;
    ram_cell[   15849] = 32'h0;  // 32'hfe31cfdc;
    ram_cell[   15850] = 32'h0;  // 32'h1c4d1810;
    ram_cell[   15851] = 32'h0;  // 32'hdf912403;
    ram_cell[   15852] = 32'h0;  // 32'hf7fd2a42;
    ram_cell[   15853] = 32'h0;  // 32'h2dab6a37;
    ram_cell[   15854] = 32'h0;  // 32'hcbbaf489;
    ram_cell[   15855] = 32'h0;  // 32'h2ea3b2c0;
    ram_cell[   15856] = 32'h0;  // 32'h62a9cd5e;
    ram_cell[   15857] = 32'h0;  // 32'h237d9ffa;
    ram_cell[   15858] = 32'h0;  // 32'hac9e1623;
    ram_cell[   15859] = 32'h0;  // 32'h3551c9ee;
    ram_cell[   15860] = 32'h0;  // 32'he5aca931;
    ram_cell[   15861] = 32'h0;  // 32'hb9e4c2c9;
    ram_cell[   15862] = 32'h0;  // 32'h45b30c6b;
    ram_cell[   15863] = 32'h0;  // 32'ha1c09b78;
    ram_cell[   15864] = 32'h0;  // 32'h3bc2a222;
    ram_cell[   15865] = 32'h0;  // 32'h0a450b68;
    ram_cell[   15866] = 32'h0;  // 32'h4e813833;
    ram_cell[   15867] = 32'h0;  // 32'h72716995;
    ram_cell[   15868] = 32'h0;  // 32'h45a4e8af;
    ram_cell[   15869] = 32'h0;  // 32'hbd56c0f5;
    ram_cell[   15870] = 32'h0;  // 32'h0307b7b8;
    ram_cell[   15871] = 32'h0;  // 32'h431f3c4f;
    ram_cell[   15872] = 32'h0;  // 32'h3c9459d4;
    ram_cell[   15873] = 32'h0;  // 32'heca596fe;
    ram_cell[   15874] = 32'h0;  // 32'h75230603;
    ram_cell[   15875] = 32'h0;  // 32'h4ede9be5;
    ram_cell[   15876] = 32'h0;  // 32'h0acec417;
    ram_cell[   15877] = 32'h0;  // 32'he291c046;
    ram_cell[   15878] = 32'h0;  // 32'h286fad85;
    ram_cell[   15879] = 32'h0;  // 32'h17bfc794;
    ram_cell[   15880] = 32'h0;  // 32'h06bea336;
    ram_cell[   15881] = 32'h0;  // 32'h242092c7;
    ram_cell[   15882] = 32'h0;  // 32'h1be842b6;
    ram_cell[   15883] = 32'h0;  // 32'h6cc0d7fa;
    ram_cell[   15884] = 32'h0;  // 32'heed4e648;
    ram_cell[   15885] = 32'h0;  // 32'hc36d02e8;
    ram_cell[   15886] = 32'h0;  // 32'hf69cd617;
    ram_cell[   15887] = 32'h0;  // 32'h5f90bf76;
    ram_cell[   15888] = 32'h0;  // 32'hdc225d30;
    ram_cell[   15889] = 32'h0;  // 32'h1d766898;
    ram_cell[   15890] = 32'h0;  // 32'h91ded69e;
    ram_cell[   15891] = 32'h0;  // 32'h9df8c59e;
    ram_cell[   15892] = 32'h0;  // 32'hca7ec868;
    ram_cell[   15893] = 32'h0;  // 32'he4b11732;
    ram_cell[   15894] = 32'h0;  // 32'h1dee9590;
    ram_cell[   15895] = 32'h0;  // 32'h1d9c1360;
    ram_cell[   15896] = 32'h0;  // 32'h60966cc8;
    ram_cell[   15897] = 32'h0;  // 32'h2dd7cdb0;
    ram_cell[   15898] = 32'h0;  // 32'hd5483161;
    ram_cell[   15899] = 32'h0;  // 32'h0fad949d;
    ram_cell[   15900] = 32'h0;  // 32'h20c2ebb3;
    ram_cell[   15901] = 32'h0;  // 32'h7dcf397d;
    ram_cell[   15902] = 32'h0;  // 32'h781b5798;
    ram_cell[   15903] = 32'h0;  // 32'h8952b2db;
    ram_cell[   15904] = 32'h0;  // 32'h78ae7411;
    ram_cell[   15905] = 32'h0;  // 32'hf23e4099;
    ram_cell[   15906] = 32'h0;  // 32'ha417903f;
    ram_cell[   15907] = 32'h0;  // 32'h78a5d486;
    ram_cell[   15908] = 32'h0;  // 32'h16fc4813;
    ram_cell[   15909] = 32'h0;  // 32'hb7e05b3a;
    ram_cell[   15910] = 32'h0;  // 32'hdbd43cbc;
    ram_cell[   15911] = 32'h0;  // 32'h5f23b327;
    ram_cell[   15912] = 32'h0;  // 32'h5bc973d8;
    ram_cell[   15913] = 32'h0;  // 32'h7c03d508;
    ram_cell[   15914] = 32'h0;  // 32'h92a802e1;
    ram_cell[   15915] = 32'h0;  // 32'h37743d0b;
    ram_cell[   15916] = 32'h0;  // 32'hcbee4444;
    ram_cell[   15917] = 32'h0;  // 32'he5fc50d2;
    ram_cell[   15918] = 32'h0;  // 32'h32606248;
    ram_cell[   15919] = 32'h0;  // 32'h2baf3fd7;
    ram_cell[   15920] = 32'h0;  // 32'ha40c41d6;
    ram_cell[   15921] = 32'h0;  // 32'h75c0b2ee;
    ram_cell[   15922] = 32'h0;  // 32'heb726f44;
    ram_cell[   15923] = 32'h0;  // 32'h6019ff18;
    ram_cell[   15924] = 32'h0;  // 32'h8a2e7225;
    ram_cell[   15925] = 32'h0;  // 32'h42eac89b;
    ram_cell[   15926] = 32'h0;  // 32'h8298954e;
    ram_cell[   15927] = 32'h0;  // 32'h756eb100;
    ram_cell[   15928] = 32'h0;  // 32'hf1b6a64c;
    ram_cell[   15929] = 32'h0;  // 32'h0726b1bf;
    ram_cell[   15930] = 32'h0;  // 32'h6503c34d;
    ram_cell[   15931] = 32'h0;  // 32'h62717124;
    ram_cell[   15932] = 32'h0;  // 32'h22472688;
    ram_cell[   15933] = 32'h0;  // 32'hfd1d697a;
    ram_cell[   15934] = 32'h0;  // 32'h3e9b1863;
    ram_cell[   15935] = 32'h0;  // 32'h501899b4;
    ram_cell[   15936] = 32'h0;  // 32'h027c66d8;
    ram_cell[   15937] = 32'h0;  // 32'h7cf03830;
    ram_cell[   15938] = 32'h0;  // 32'h73f5a66f;
    ram_cell[   15939] = 32'h0;  // 32'h3479fe01;
    ram_cell[   15940] = 32'h0;  // 32'h17be5c48;
    ram_cell[   15941] = 32'h0;  // 32'h46431b8d;
    ram_cell[   15942] = 32'h0;  // 32'h56dfa150;
    ram_cell[   15943] = 32'h0;  // 32'h0859f1ac;
    ram_cell[   15944] = 32'h0;  // 32'h94c4c10a;
    ram_cell[   15945] = 32'h0;  // 32'hf0291bd1;
    ram_cell[   15946] = 32'h0;  // 32'h8c2b91b0;
    ram_cell[   15947] = 32'h0;  // 32'hac8c3a1e;
    ram_cell[   15948] = 32'h0;  // 32'h3b87c185;
    ram_cell[   15949] = 32'h0;  // 32'h7264ed1a;
    ram_cell[   15950] = 32'h0;  // 32'h7a0578cd;
    ram_cell[   15951] = 32'h0;  // 32'h6c27bf1f;
    ram_cell[   15952] = 32'h0;  // 32'hb1464c0a;
    ram_cell[   15953] = 32'h0;  // 32'h14002422;
    ram_cell[   15954] = 32'h0;  // 32'h6ad656f9;
    ram_cell[   15955] = 32'h0;  // 32'h8f84d261;
    ram_cell[   15956] = 32'h0;  // 32'h8e36414a;
    ram_cell[   15957] = 32'h0;  // 32'he36dbc7b;
    ram_cell[   15958] = 32'h0;  // 32'h3827624a;
    ram_cell[   15959] = 32'h0;  // 32'h3f80530e;
    ram_cell[   15960] = 32'h0;  // 32'h791c9de5;
    ram_cell[   15961] = 32'h0;  // 32'h2b992715;
    ram_cell[   15962] = 32'h0;  // 32'h202a4ad1;
    ram_cell[   15963] = 32'h0;  // 32'h1d39b615;
    ram_cell[   15964] = 32'h0;  // 32'h77ab4d3d;
    ram_cell[   15965] = 32'h0;  // 32'he12e6698;
    ram_cell[   15966] = 32'h0;  // 32'h87c3aab4;
    ram_cell[   15967] = 32'h0;  // 32'h19a5d661;
    ram_cell[   15968] = 32'h0;  // 32'h2dcaaeec;
    ram_cell[   15969] = 32'h0;  // 32'ha06e7d98;
    ram_cell[   15970] = 32'h0;  // 32'h2e8e9e7d;
    ram_cell[   15971] = 32'h0;  // 32'he2c21b5e;
    ram_cell[   15972] = 32'h0;  // 32'h8ecc81d5;
    ram_cell[   15973] = 32'h0;  // 32'h6cb021dd;
    ram_cell[   15974] = 32'h0;  // 32'h27e065a1;
    ram_cell[   15975] = 32'h0;  // 32'h16491b43;
    ram_cell[   15976] = 32'h0;  // 32'hc98c876f;
    ram_cell[   15977] = 32'h0;  // 32'h8bf76c69;
    ram_cell[   15978] = 32'h0;  // 32'had0b8ba7;
    ram_cell[   15979] = 32'h0;  // 32'hf40c0c24;
    ram_cell[   15980] = 32'h0;  // 32'h4a7642e9;
    ram_cell[   15981] = 32'h0;  // 32'h1a976a3e;
    ram_cell[   15982] = 32'h0;  // 32'h0b8643cc;
    ram_cell[   15983] = 32'h0;  // 32'he8354341;
    ram_cell[   15984] = 32'h0;  // 32'h4e31b83d;
    ram_cell[   15985] = 32'h0;  // 32'h16f264a0;
    ram_cell[   15986] = 32'h0;  // 32'h24b5f089;
    ram_cell[   15987] = 32'h0;  // 32'h1906a511;
    ram_cell[   15988] = 32'h0;  // 32'haee0e13e;
    ram_cell[   15989] = 32'h0;  // 32'h9eca5a40;
    ram_cell[   15990] = 32'h0;  // 32'hae5bed3a;
    ram_cell[   15991] = 32'h0;  // 32'he86b78e7;
    ram_cell[   15992] = 32'h0;  // 32'he6d4f888;
    ram_cell[   15993] = 32'h0;  // 32'h24aa1d3e;
    ram_cell[   15994] = 32'h0;  // 32'h53506bf0;
    ram_cell[   15995] = 32'h0;  // 32'hae3dc9d7;
    ram_cell[   15996] = 32'h0;  // 32'h936d3ec0;
    ram_cell[   15997] = 32'h0;  // 32'h666028aa;
    ram_cell[   15998] = 32'h0;  // 32'hdd51b3ee;
    ram_cell[   15999] = 32'h0;  // 32'h612b60e6;
    ram_cell[   16000] = 32'h0;  // 32'h63622aef;
    ram_cell[   16001] = 32'h0;  // 32'hb1d671cd;
    ram_cell[   16002] = 32'h0;  // 32'hb7607c9e;
    ram_cell[   16003] = 32'h0;  // 32'h0c274757;
    ram_cell[   16004] = 32'h0;  // 32'h45541eca;
    ram_cell[   16005] = 32'h0;  // 32'he330f026;
    ram_cell[   16006] = 32'h0;  // 32'hc37dacd4;
    ram_cell[   16007] = 32'h0;  // 32'h376d1c9c;
    ram_cell[   16008] = 32'h0;  // 32'h02720cf7;
    ram_cell[   16009] = 32'h0;  // 32'h7c4d98f8;
    ram_cell[   16010] = 32'h0;  // 32'h48d5337f;
    ram_cell[   16011] = 32'h0;  // 32'h006b1af5;
    ram_cell[   16012] = 32'h0;  // 32'hbdb5eb8e;
    ram_cell[   16013] = 32'h0;  // 32'h094d54e9;
    ram_cell[   16014] = 32'h0;  // 32'hd3cbd46e;
    ram_cell[   16015] = 32'h0;  // 32'he5c7425e;
    ram_cell[   16016] = 32'h0;  // 32'h40251123;
    ram_cell[   16017] = 32'h0;  // 32'h60c3e947;
    ram_cell[   16018] = 32'h0;  // 32'h14831f27;
    ram_cell[   16019] = 32'h0;  // 32'h5ac38b09;
    ram_cell[   16020] = 32'h0;  // 32'h4943eae4;
    ram_cell[   16021] = 32'h0;  // 32'h9057927d;
    ram_cell[   16022] = 32'h0;  // 32'h689293e2;
    ram_cell[   16023] = 32'h0;  // 32'hd20c6dd7;
    ram_cell[   16024] = 32'h0;  // 32'hc337212d;
    ram_cell[   16025] = 32'h0;  // 32'hd72bcd02;
    ram_cell[   16026] = 32'h0;  // 32'hdc621527;
    ram_cell[   16027] = 32'h0;  // 32'hbe0c3603;
    ram_cell[   16028] = 32'h0;  // 32'h78637f07;
    ram_cell[   16029] = 32'h0;  // 32'h9e414305;
    ram_cell[   16030] = 32'h0;  // 32'h46a803e0;
    ram_cell[   16031] = 32'h0;  // 32'h1e55eba2;
    ram_cell[   16032] = 32'h0;  // 32'hd0d9c1d9;
    ram_cell[   16033] = 32'h0;  // 32'h5e87d40e;
    ram_cell[   16034] = 32'h0;  // 32'h7cbb22ad;
    ram_cell[   16035] = 32'h0;  // 32'h3ec3244f;
    ram_cell[   16036] = 32'h0;  // 32'h00416285;
    ram_cell[   16037] = 32'h0;  // 32'h222d5ab8;
    ram_cell[   16038] = 32'h0;  // 32'h678bcded;
    ram_cell[   16039] = 32'h0;  // 32'hd0733b57;
    ram_cell[   16040] = 32'h0;  // 32'h3332e18d;
    ram_cell[   16041] = 32'h0;  // 32'h9f304055;
    ram_cell[   16042] = 32'h0;  // 32'h62c99244;
    ram_cell[   16043] = 32'h0;  // 32'h7d48148a;
    ram_cell[   16044] = 32'h0;  // 32'h66513b2d;
    ram_cell[   16045] = 32'h0;  // 32'h47c671b5;
    ram_cell[   16046] = 32'h0;  // 32'hea66682b;
    ram_cell[   16047] = 32'h0;  // 32'h6695a346;
    ram_cell[   16048] = 32'h0;  // 32'h13ff30cb;
    ram_cell[   16049] = 32'h0;  // 32'h01514079;
    ram_cell[   16050] = 32'h0;  // 32'h54983c14;
    ram_cell[   16051] = 32'h0;  // 32'h8b58b3cc;
    ram_cell[   16052] = 32'h0;  // 32'h37aca51e;
    ram_cell[   16053] = 32'h0;  // 32'h25e70713;
    ram_cell[   16054] = 32'h0;  // 32'h37578da6;
    ram_cell[   16055] = 32'h0;  // 32'h94c0d6e1;
    ram_cell[   16056] = 32'h0;  // 32'h1786a3ec;
    ram_cell[   16057] = 32'h0;  // 32'h27d86dd6;
    ram_cell[   16058] = 32'h0;  // 32'hb2138ad9;
    ram_cell[   16059] = 32'h0;  // 32'hcfb943e7;
    ram_cell[   16060] = 32'h0;  // 32'h10c6dc37;
    ram_cell[   16061] = 32'h0;  // 32'hb854ce5f;
    ram_cell[   16062] = 32'h0;  // 32'hd7e711a2;
    ram_cell[   16063] = 32'h0;  // 32'h333d3276;
    ram_cell[   16064] = 32'h0;  // 32'h114631e5;
    ram_cell[   16065] = 32'h0;  // 32'hca6ce004;
    ram_cell[   16066] = 32'h0;  // 32'h7f7620a7;
    ram_cell[   16067] = 32'h0;  // 32'h0c7a0f24;
    ram_cell[   16068] = 32'h0;  // 32'h6f2feb27;
    ram_cell[   16069] = 32'h0;  // 32'hf0a51346;
    ram_cell[   16070] = 32'h0;  // 32'hdd5be7cd;
    ram_cell[   16071] = 32'h0;  // 32'h76544fb6;
    ram_cell[   16072] = 32'h0;  // 32'h4e30939e;
    ram_cell[   16073] = 32'h0;  // 32'hd2d002a5;
    ram_cell[   16074] = 32'h0;  // 32'he6e56509;
    ram_cell[   16075] = 32'h0;  // 32'h0c002242;
    ram_cell[   16076] = 32'h0;  // 32'hda72a276;
    ram_cell[   16077] = 32'h0;  // 32'h18c1c48a;
    ram_cell[   16078] = 32'h0;  // 32'h4ccadcc9;
    ram_cell[   16079] = 32'h0;  // 32'h1f5258e4;
    ram_cell[   16080] = 32'h0;  // 32'h34ddf68b;
    ram_cell[   16081] = 32'h0;  // 32'hf61adc53;
    ram_cell[   16082] = 32'h0;  // 32'hfcb4b4c4;
    ram_cell[   16083] = 32'h0;  // 32'hb298b4c9;
    ram_cell[   16084] = 32'h0;  // 32'h94ff08dc;
    ram_cell[   16085] = 32'h0;  // 32'h2d1a92ce;
    ram_cell[   16086] = 32'h0;  // 32'hfb65938c;
    ram_cell[   16087] = 32'h0;  // 32'hd8510829;
    ram_cell[   16088] = 32'h0;  // 32'he23014a3;
    ram_cell[   16089] = 32'h0;  // 32'hf2aa3d4b;
    ram_cell[   16090] = 32'h0;  // 32'h6073b9d5;
    ram_cell[   16091] = 32'h0;  // 32'hf4e4bbcf;
    ram_cell[   16092] = 32'h0;  // 32'hcd9b0dc5;
    ram_cell[   16093] = 32'h0;  // 32'h062d6fda;
    ram_cell[   16094] = 32'h0;  // 32'he145dc58;
    ram_cell[   16095] = 32'h0;  // 32'hed905793;
    ram_cell[   16096] = 32'h0;  // 32'h56184855;
    ram_cell[   16097] = 32'h0;  // 32'habc9210f;
    ram_cell[   16098] = 32'h0;  // 32'h1d72aeb4;
    ram_cell[   16099] = 32'h0;  // 32'hafc91b9f;
    ram_cell[   16100] = 32'h0;  // 32'h3b85be8b;
    ram_cell[   16101] = 32'h0;  // 32'he84509e4;
    ram_cell[   16102] = 32'h0;  // 32'hcecaeef5;
    ram_cell[   16103] = 32'h0;  // 32'h7e1780ef;
    ram_cell[   16104] = 32'h0;  // 32'h09d8728e;
    ram_cell[   16105] = 32'h0;  // 32'ha3cb7d08;
    ram_cell[   16106] = 32'h0;  // 32'h947cbed2;
    ram_cell[   16107] = 32'h0;  // 32'hb8c39e04;
    ram_cell[   16108] = 32'h0;  // 32'hb23fc552;
    ram_cell[   16109] = 32'h0;  // 32'haa2f739a;
    ram_cell[   16110] = 32'h0;  // 32'h1daae815;
    ram_cell[   16111] = 32'h0;  // 32'h2b3ac748;
    ram_cell[   16112] = 32'h0;  // 32'h9515e715;
    ram_cell[   16113] = 32'h0;  // 32'haed20f67;
    ram_cell[   16114] = 32'h0;  // 32'hbda96124;
    ram_cell[   16115] = 32'h0;  // 32'h11e4204f;
    ram_cell[   16116] = 32'h0;  // 32'hda01865f;
    ram_cell[   16117] = 32'h0;  // 32'hd4a639e4;
    ram_cell[   16118] = 32'h0;  // 32'ha1ad86b7;
    ram_cell[   16119] = 32'h0;  // 32'hb8ca48bc;
    ram_cell[   16120] = 32'h0;  // 32'hdb0d3acf;
    ram_cell[   16121] = 32'h0;  // 32'hccda31ab;
    ram_cell[   16122] = 32'h0;  // 32'h9662bee1;
    ram_cell[   16123] = 32'h0;  // 32'h852896b9;
    ram_cell[   16124] = 32'h0;  // 32'h84aa5813;
    ram_cell[   16125] = 32'h0;  // 32'h6e630f47;
    ram_cell[   16126] = 32'h0;  // 32'he124fcfd;
    ram_cell[   16127] = 32'h0;  // 32'h304ed3ef;
    ram_cell[   16128] = 32'h0;  // 32'hcbe5e26d;
    ram_cell[   16129] = 32'h0;  // 32'h7ee549cd;
    ram_cell[   16130] = 32'h0;  // 32'hf4f29f73;
    ram_cell[   16131] = 32'h0;  // 32'hbba60f90;
    ram_cell[   16132] = 32'h0;  // 32'hf5b53ee1;
    ram_cell[   16133] = 32'h0;  // 32'h2dd0f7bb;
    ram_cell[   16134] = 32'h0;  // 32'hadfa1865;
    ram_cell[   16135] = 32'h0;  // 32'he637fb3e;
    ram_cell[   16136] = 32'h0;  // 32'h94ae6709;
    ram_cell[   16137] = 32'h0;  // 32'h230d6d32;
    ram_cell[   16138] = 32'h0;  // 32'h5199ce64;
    ram_cell[   16139] = 32'h0;  // 32'hd5db85f5;
    ram_cell[   16140] = 32'h0;  // 32'h1e1a524d;
    ram_cell[   16141] = 32'h0;  // 32'hf4905925;
    ram_cell[   16142] = 32'h0;  // 32'h56cb2091;
    ram_cell[   16143] = 32'h0;  // 32'h156f5b85;
    ram_cell[   16144] = 32'h0;  // 32'h465daf28;
    ram_cell[   16145] = 32'h0;  // 32'h0871ace5;
    ram_cell[   16146] = 32'h0;  // 32'h03352396;
    ram_cell[   16147] = 32'h0;  // 32'h56cb35f0;
    ram_cell[   16148] = 32'h0;  // 32'h894f50b4;
    ram_cell[   16149] = 32'h0;  // 32'h9719e3d4;
    ram_cell[   16150] = 32'h0;  // 32'h8e7ccb22;
    ram_cell[   16151] = 32'h0;  // 32'h94d86230;
    ram_cell[   16152] = 32'h0;  // 32'hb1b635e5;
    ram_cell[   16153] = 32'h0;  // 32'hce39c0ac;
    ram_cell[   16154] = 32'h0;  // 32'h9fb70113;
    ram_cell[   16155] = 32'h0;  // 32'hbc7062f0;
    ram_cell[   16156] = 32'h0;  // 32'ha46efa57;
    ram_cell[   16157] = 32'h0;  // 32'h049f9279;
    ram_cell[   16158] = 32'h0;  // 32'hb6a869b1;
    ram_cell[   16159] = 32'h0;  // 32'h1289dbe5;
    ram_cell[   16160] = 32'h0;  // 32'h31476493;
    ram_cell[   16161] = 32'h0;  // 32'hac658f7f;
    ram_cell[   16162] = 32'h0;  // 32'h11711289;
    ram_cell[   16163] = 32'h0;  // 32'hfa2d4c65;
    ram_cell[   16164] = 32'h0;  // 32'h270987da;
    ram_cell[   16165] = 32'h0;  // 32'ha0594526;
    ram_cell[   16166] = 32'h0;  // 32'hbe7cae22;
    ram_cell[   16167] = 32'h0;  // 32'hae571925;
    ram_cell[   16168] = 32'h0;  // 32'h92cba53d;
    ram_cell[   16169] = 32'h0;  // 32'hdf0c5ec0;
    ram_cell[   16170] = 32'h0;  // 32'h76e86f4b;
    ram_cell[   16171] = 32'h0;  // 32'h844e35ff;
    ram_cell[   16172] = 32'h0;  // 32'haea04e18;
    ram_cell[   16173] = 32'h0;  // 32'h8663a8d8;
    ram_cell[   16174] = 32'h0;  // 32'hc3c45aba;
    ram_cell[   16175] = 32'h0;  // 32'h486973b8;
    ram_cell[   16176] = 32'h0;  // 32'h9ec34428;
    ram_cell[   16177] = 32'h0;  // 32'h83bb016a;
    ram_cell[   16178] = 32'h0;  // 32'h99bd2e80;
    ram_cell[   16179] = 32'h0;  // 32'hb025dae0;
    ram_cell[   16180] = 32'h0;  // 32'h2c18240c;
    ram_cell[   16181] = 32'h0;  // 32'hc0e61afe;
    ram_cell[   16182] = 32'h0;  // 32'h687e252e;
    ram_cell[   16183] = 32'h0;  // 32'h6de49449;
    ram_cell[   16184] = 32'h0;  // 32'hb6173a6b;
    ram_cell[   16185] = 32'h0;  // 32'hdb851eb0;
    ram_cell[   16186] = 32'h0;  // 32'hacbf8b28;
    ram_cell[   16187] = 32'h0;  // 32'h8be19784;
    ram_cell[   16188] = 32'h0;  // 32'hb12d2154;
    ram_cell[   16189] = 32'h0;  // 32'h28e4071c;
    ram_cell[   16190] = 32'h0;  // 32'h19cb4af4;
    ram_cell[   16191] = 32'h0;  // 32'h61edf81c;
    ram_cell[   16192] = 32'h0;  // 32'h070e2372;
    ram_cell[   16193] = 32'h0;  // 32'h4e902243;
    ram_cell[   16194] = 32'h0;  // 32'h55d5c2b8;
    ram_cell[   16195] = 32'h0;  // 32'h06b8b1fb;
    ram_cell[   16196] = 32'h0;  // 32'h678994b0;
    ram_cell[   16197] = 32'h0;  // 32'h2d4b4813;
    ram_cell[   16198] = 32'h0;  // 32'h28f58a86;
    ram_cell[   16199] = 32'h0;  // 32'h5196a8ea;
    ram_cell[   16200] = 32'h0;  // 32'h2af0ae4f;
    ram_cell[   16201] = 32'h0;  // 32'h0d4ada45;
    ram_cell[   16202] = 32'h0;  // 32'h6ba069fa;
    ram_cell[   16203] = 32'h0;  // 32'h136039f2;
    ram_cell[   16204] = 32'h0;  // 32'h095a46cf;
    ram_cell[   16205] = 32'h0;  // 32'h949d9c2d;
    ram_cell[   16206] = 32'h0;  // 32'h1b030421;
    ram_cell[   16207] = 32'h0;  // 32'h4946de60;
    ram_cell[   16208] = 32'h0;  // 32'hc28151ce;
    ram_cell[   16209] = 32'h0;  // 32'h0dcc7446;
    ram_cell[   16210] = 32'h0;  // 32'ha349d13e;
    ram_cell[   16211] = 32'h0;  // 32'hd99ef094;
    ram_cell[   16212] = 32'h0;  // 32'h962222f4;
    ram_cell[   16213] = 32'h0;  // 32'hd902e001;
    ram_cell[   16214] = 32'h0;  // 32'h5160b194;
    ram_cell[   16215] = 32'h0;  // 32'hddf16305;
    ram_cell[   16216] = 32'h0;  // 32'hd31a601d;
    ram_cell[   16217] = 32'h0;  // 32'h4b9013a1;
    ram_cell[   16218] = 32'h0;  // 32'h3f1ec258;
    ram_cell[   16219] = 32'h0;  // 32'hc413b081;
    ram_cell[   16220] = 32'h0;  // 32'hd8279c36;
    ram_cell[   16221] = 32'h0;  // 32'h0ac7ca28;
    ram_cell[   16222] = 32'h0;  // 32'h5d2aa824;
    ram_cell[   16223] = 32'h0;  // 32'h0b23c588;
    ram_cell[   16224] = 32'h0;  // 32'h2d2aafec;
    ram_cell[   16225] = 32'h0;  // 32'hc8209eef;
    ram_cell[   16226] = 32'h0;  // 32'hfa6729cc;
    ram_cell[   16227] = 32'h0;  // 32'h1bfbe114;
    ram_cell[   16228] = 32'h0;  // 32'h9432ee9f;
    ram_cell[   16229] = 32'h0;  // 32'h99dfb573;
    ram_cell[   16230] = 32'h0;  // 32'h3ecdae55;
    ram_cell[   16231] = 32'h0;  // 32'hba502f80;
    ram_cell[   16232] = 32'h0;  // 32'hfa9c38a7;
    ram_cell[   16233] = 32'h0;  // 32'hb46994c4;
    ram_cell[   16234] = 32'h0;  // 32'h9d1876d7;
    ram_cell[   16235] = 32'h0;  // 32'h7ef0cf17;
    ram_cell[   16236] = 32'h0;  // 32'h4648d1b8;
    ram_cell[   16237] = 32'h0;  // 32'h479ac556;
    ram_cell[   16238] = 32'h0;  // 32'h9716e914;
    ram_cell[   16239] = 32'h0;  // 32'h5d62da23;
    ram_cell[   16240] = 32'h0;  // 32'h2ce1f304;
    ram_cell[   16241] = 32'h0;  // 32'hf68fcd17;
    ram_cell[   16242] = 32'h0;  // 32'he7d4e64e;
    ram_cell[   16243] = 32'h0;  // 32'hda3d33bb;
    ram_cell[   16244] = 32'h0;  // 32'hfe90378b;
    ram_cell[   16245] = 32'h0;  // 32'h25370c44;
    ram_cell[   16246] = 32'h0;  // 32'h3556f135;
    ram_cell[   16247] = 32'h0;  // 32'hcb69f750;
    ram_cell[   16248] = 32'h0;  // 32'h5c1136e1;
    ram_cell[   16249] = 32'h0;  // 32'h958776b5;
    ram_cell[   16250] = 32'h0;  // 32'hcbe12ef1;
    ram_cell[   16251] = 32'h0;  // 32'habee8970;
    ram_cell[   16252] = 32'h0;  // 32'h53a788d5;
    ram_cell[   16253] = 32'h0;  // 32'h71fab03a;
    ram_cell[   16254] = 32'h0;  // 32'h78d4efd8;
    ram_cell[   16255] = 32'h0;  // 32'h2c2f9f54;
    ram_cell[   16256] = 32'h0;  // 32'h46135100;
    ram_cell[   16257] = 32'h0;  // 32'hd9460248;
    ram_cell[   16258] = 32'h0;  // 32'h2e9b1713;
    ram_cell[   16259] = 32'h0;  // 32'h6a3ae969;
    ram_cell[   16260] = 32'h0;  // 32'h9bb6acc6;
    ram_cell[   16261] = 32'h0;  // 32'hf6a052fc;
    ram_cell[   16262] = 32'h0;  // 32'hea44b25f;
    ram_cell[   16263] = 32'h0;  // 32'h160b36d0;
    ram_cell[   16264] = 32'h0;  // 32'h6486b757;
    ram_cell[   16265] = 32'h0;  // 32'h91d71d8a;
    ram_cell[   16266] = 32'h0;  // 32'h29a1fdb1;
    ram_cell[   16267] = 32'h0;  // 32'hb2b43345;
    ram_cell[   16268] = 32'h0;  // 32'hc388ea22;
    ram_cell[   16269] = 32'h0;  // 32'hc7dd097a;
    ram_cell[   16270] = 32'h0;  // 32'h4ea594f8;
    ram_cell[   16271] = 32'h0;  // 32'h31b0e881;
    ram_cell[   16272] = 32'h0;  // 32'hef0fed2c;
    ram_cell[   16273] = 32'h0;  // 32'hbb0ca420;
    ram_cell[   16274] = 32'h0;  // 32'hbc03e5a2;
    ram_cell[   16275] = 32'h0;  // 32'hfeac2a38;
    ram_cell[   16276] = 32'h0;  // 32'ha8d25f54;
    ram_cell[   16277] = 32'h0;  // 32'h79180e1d;
    ram_cell[   16278] = 32'h0;  // 32'heff39aa2;
    ram_cell[   16279] = 32'h0;  // 32'h2032ec71;
    ram_cell[   16280] = 32'h0;  // 32'h5b1b8493;
    ram_cell[   16281] = 32'h0;  // 32'h4f77a3fb;
    ram_cell[   16282] = 32'h0;  // 32'h6c6553c0;
    ram_cell[   16283] = 32'h0;  // 32'h90768b29;
    ram_cell[   16284] = 32'h0;  // 32'h1f292b10;
    ram_cell[   16285] = 32'h0;  // 32'hc40c2a2e;
    ram_cell[   16286] = 32'h0;  // 32'h40b88f66;
    ram_cell[   16287] = 32'h0;  // 32'he1a97b2b;
    ram_cell[   16288] = 32'h0;  // 32'hb0615a6f;
    ram_cell[   16289] = 32'h0;  // 32'h8328e247;
    ram_cell[   16290] = 32'h0;  // 32'h5b40650d;
    ram_cell[   16291] = 32'h0;  // 32'h5b851abd;
    ram_cell[   16292] = 32'h0;  // 32'h30d50c34;
    ram_cell[   16293] = 32'h0;  // 32'h4dcafcbd;
    ram_cell[   16294] = 32'h0;  // 32'h4dc864ee;
    ram_cell[   16295] = 32'h0;  // 32'h8e79bb43;
    ram_cell[   16296] = 32'h0;  // 32'he6502cc3;
    ram_cell[   16297] = 32'h0;  // 32'h218bb1ab;
    ram_cell[   16298] = 32'h0;  // 32'hbbde4771;
    ram_cell[   16299] = 32'h0;  // 32'h09e3f65f;
    ram_cell[   16300] = 32'h0;  // 32'h7c322354;
    ram_cell[   16301] = 32'h0;  // 32'h0ce28907;
    ram_cell[   16302] = 32'h0;  // 32'h1285c331;
    ram_cell[   16303] = 32'h0;  // 32'hb4c26e5d;
    ram_cell[   16304] = 32'h0;  // 32'h059ac7f0;
    ram_cell[   16305] = 32'h0;  // 32'hd76883a1;
    ram_cell[   16306] = 32'h0;  // 32'h83876541;
    ram_cell[   16307] = 32'h0;  // 32'h2f85bbf1;
    ram_cell[   16308] = 32'h0;  // 32'hfb2c1b65;
    ram_cell[   16309] = 32'h0;  // 32'h2d709829;
    ram_cell[   16310] = 32'h0;  // 32'h92ebe697;
    ram_cell[   16311] = 32'h0;  // 32'h984639f1;
    ram_cell[   16312] = 32'h0;  // 32'hcbafad99;
    ram_cell[   16313] = 32'h0;  // 32'h155b56e3;
    ram_cell[   16314] = 32'h0;  // 32'h6982c061;
    ram_cell[   16315] = 32'h0;  // 32'hce2adb4c;
    ram_cell[   16316] = 32'h0;  // 32'h4a5e97a0;
    ram_cell[   16317] = 32'h0;  // 32'h14b47c48;
    ram_cell[   16318] = 32'h0;  // 32'hdd579db4;
    ram_cell[   16319] = 32'h0;  // 32'hf74393ac;
    ram_cell[   16320] = 32'h0;  // 32'h2a58e3b1;
    ram_cell[   16321] = 32'h0;  // 32'h31fd8f3b;
    ram_cell[   16322] = 32'h0;  // 32'hc4cd012e;
    ram_cell[   16323] = 32'h0;  // 32'hbc808052;
    ram_cell[   16324] = 32'h0;  // 32'hbf304677;
    ram_cell[   16325] = 32'h0;  // 32'h85dcebb2;
    ram_cell[   16326] = 32'h0;  // 32'hc843d83b;
    ram_cell[   16327] = 32'h0;  // 32'h8a604535;
    ram_cell[   16328] = 32'h0;  // 32'hf046d6b4;
    ram_cell[   16329] = 32'h0;  // 32'hf5432db4;
    ram_cell[   16330] = 32'h0;  // 32'h53ba9614;
    ram_cell[   16331] = 32'h0;  // 32'h120a719c;
    ram_cell[   16332] = 32'h0;  // 32'hee4ef6c4;
    ram_cell[   16333] = 32'h0;  // 32'h64a9945f;
    ram_cell[   16334] = 32'h0;  // 32'h486b0ba8;
    ram_cell[   16335] = 32'h0;  // 32'hfe23d90c;
    ram_cell[   16336] = 32'h0;  // 32'hba83e9e0;
    ram_cell[   16337] = 32'h0;  // 32'hcebc9058;
    ram_cell[   16338] = 32'h0;  // 32'h5e7c6b63;
    ram_cell[   16339] = 32'h0;  // 32'hca130085;
    ram_cell[   16340] = 32'h0;  // 32'hfd6f1b1e;
    ram_cell[   16341] = 32'h0;  // 32'hf7c1d6d6;
    ram_cell[   16342] = 32'h0;  // 32'h844fbfd0;
    ram_cell[   16343] = 32'h0;  // 32'h4d7dfa08;
    ram_cell[   16344] = 32'h0;  // 32'h70c8d52f;
    ram_cell[   16345] = 32'h0;  // 32'hd83463ab;
    ram_cell[   16346] = 32'h0;  // 32'h1bd8ae83;
    ram_cell[   16347] = 32'h0;  // 32'he6c4d890;
    ram_cell[   16348] = 32'h0;  // 32'h56e072b4;
    ram_cell[   16349] = 32'h0;  // 32'hc2b1e560;
    ram_cell[   16350] = 32'h0;  // 32'h7e856238;
    ram_cell[   16351] = 32'h0;  // 32'he13bdaa9;
    ram_cell[   16352] = 32'h0;  // 32'h0a9546b8;
    ram_cell[   16353] = 32'h0;  // 32'h414be9b8;
    ram_cell[   16354] = 32'h0;  // 32'h8e94fba6;
    ram_cell[   16355] = 32'h0;  // 32'h390b1d40;
    ram_cell[   16356] = 32'h0;  // 32'ha06d197c;
    ram_cell[   16357] = 32'h0;  // 32'h9f26d03c;
    ram_cell[   16358] = 32'h0;  // 32'hb7897d76;
    ram_cell[   16359] = 32'h0;  // 32'h272b7757;
    ram_cell[   16360] = 32'h0;  // 32'h76f3064b;
    ram_cell[   16361] = 32'h0;  // 32'h69918af0;
    ram_cell[   16362] = 32'h0;  // 32'haea54374;
    ram_cell[   16363] = 32'h0;  // 32'h07b1158e;
    ram_cell[   16364] = 32'h0;  // 32'h8dce3c6f;
    ram_cell[   16365] = 32'h0;  // 32'h70a642be;
    ram_cell[   16366] = 32'h0;  // 32'h3cb8788d;
    ram_cell[   16367] = 32'h0;  // 32'h06271d11;
    ram_cell[   16368] = 32'h0;  // 32'h79b78680;
    ram_cell[   16369] = 32'h0;  // 32'hc55b4f9f;
    ram_cell[   16370] = 32'h0;  // 32'h1aa4d9ae;
    ram_cell[   16371] = 32'h0;  // 32'h6a400868;
    ram_cell[   16372] = 32'h0;  // 32'h048e88b0;
    ram_cell[   16373] = 32'h0;  // 32'hff53112d;
    ram_cell[   16374] = 32'h0;  // 32'hf72a10f9;
    ram_cell[   16375] = 32'h0;  // 32'h715f462b;
    ram_cell[   16376] = 32'h0;  // 32'h35640203;
    ram_cell[   16377] = 32'h0;  // 32'h0a48f7cd;
    ram_cell[   16378] = 32'h0;  // 32'h0588448c;
    ram_cell[   16379] = 32'h0;  // 32'h9b8545e0;
    ram_cell[   16380] = 32'h0;  // 32'h1d23aa5c;
    ram_cell[   16381] = 32'h0;  // 32'ha116cf31;
    ram_cell[   16382] = 32'h0;  // 32'ha740c532;
    ram_cell[   16383] = 32'h0;  // 32'h29506d4a;
    // src matrix A
    ram_cell[   16384] = 32'h135fa3a6;
    ram_cell[   16385] = 32'he69a6e57;
    ram_cell[   16386] = 32'h3363e113;
    ram_cell[   16387] = 32'hefad56f2;
    ram_cell[   16388] = 32'h7cc2210a;
    ram_cell[   16389] = 32'he7f1e80a;
    ram_cell[   16390] = 32'h0e389271;
    ram_cell[   16391] = 32'h4a8cf755;
    ram_cell[   16392] = 32'h6f048ae0;
    ram_cell[   16393] = 32'hfc51570b;
    ram_cell[   16394] = 32'h813b0217;
    ram_cell[   16395] = 32'h9bf685be;
    ram_cell[   16396] = 32'h105f097d;
    ram_cell[   16397] = 32'h50fc8cce;
    ram_cell[   16398] = 32'hb48ed25f;
    ram_cell[   16399] = 32'h971f8ee0;
    ram_cell[   16400] = 32'h0dcee96f;
    ram_cell[   16401] = 32'h109a3384;
    ram_cell[   16402] = 32'hdb2a375a;
    ram_cell[   16403] = 32'h42a4967f;
    ram_cell[   16404] = 32'hc6e73407;
    ram_cell[   16405] = 32'h0db42bd2;
    ram_cell[   16406] = 32'h5bc09a59;
    ram_cell[   16407] = 32'h9bf8d743;
    ram_cell[   16408] = 32'h340c8f3a;
    ram_cell[   16409] = 32'h4714f297;
    ram_cell[   16410] = 32'h4b48bf51;
    ram_cell[   16411] = 32'h956571c3;
    ram_cell[   16412] = 32'h1685df39;
    ram_cell[   16413] = 32'h6ec1fd16;
    ram_cell[   16414] = 32'hd3e76eba;
    ram_cell[   16415] = 32'h9a7e779c;
    ram_cell[   16416] = 32'hd7d7adce;
    ram_cell[   16417] = 32'h5b8bb97e;
    ram_cell[   16418] = 32'hc71615ff;
    ram_cell[   16419] = 32'h33727223;
    ram_cell[   16420] = 32'h19b5b46c;
    ram_cell[   16421] = 32'h61fe07bf;
    ram_cell[   16422] = 32'hb7933fef;
    ram_cell[   16423] = 32'h01111855;
    ram_cell[   16424] = 32'ha13cf90c;
    ram_cell[   16425] = 32'hc84fad7d;
    ram_cell[   16426] = 32'h3e0d3940;
    ram_cell[   16427] = 32'h2d87f4e6;
    ram_cell[   16428] = 32'had893f35;
    ram_cell[   16429] = 32'hb39361d3;
    ram_cell[   16430] = 32'h011b46fb;
    ram_cell[   16431] = 32'h5027ea8c;
    ram_cell[   16432] = 32'h33f1de67;
    ram_cell[   16433] = 32'h0dece294;
    ram_cell[   16434] = 32'h8ae6cc42;
    ram_cell[   16435] = 32'h769f1545;
    ram_cell[   16436] = 32'h94d85c81;
    ram_cell[   16437] = 32'h02dcc656;
    ram_cell[   16438] = 32'h77dcfc93;
    ram_cell[   16439] = 32'h829cea53;
    ram_cell[   16440] = 32'hc6796d7c;
    ram_cell[   16441] = 32'hd8d0d34c;
    ram_cell[   16442] = 32'h2f69bfd0;
    ram_cell[   16443] = 32'h1b0ecc02;
    ram_cell[   16444] = 32'hcd833e1a;
    ram_cell[   16445] = 32'heb27b25a;
    ram_cell[   16446] = 32'hc606280d;
    ram_cell[   16447] = 32'hfdc45d57;
    ram_cell[   16448] = 32'h6d073fc1;
    ram_cell[   16449] = 32'h7fb761bb;
    ram_cell[   16450] = 32'h87167d59;
    ram_cell[   16451] = 32'h6bb69172;
    ram_cell[   16452] = 32'hfb0aa1a3;
    ram_cell[   16453] = 32'h7d44f56d;
    ram_cell[   16454] = 32'hb86087b4;
    ram_cell[   16455] = 32'h205f18b5;
    ram_cell[   16456] = 32'h73f1f908;
    ram_cell[   16457] = 32'hc2757136;
    ram_cell[   16458] = 32'hebb3f7ff;
    ram_cell[   16459] = 32'hee4a222b;
    ram_cell[   16460] = 32'hb8fa3563;
    ram_cell[   16461] = 32'h142d1963;
    ram_cell[   16462] = 32'h35df3b18;
    ram_cell[   16463] = 32'h1d2f0b66;
    ram_cell[   16464] = 32'habb3be54;
    ram_cell[   16465] = 32'h3975d9b9;
    ram_cell[   16466] = 32'h15f6b0e3;
    ram_cell[   16467] = 32'ha23444e6;
    ram_cell[   16468] = 32'haa208af7;
    ram_cell[   16469] = 32'h1426e663;
    ram_cell[   16470] = 32'hbdfd17ee;
    ram_cell[   16471] = 32'h5368c285;
    ram_cell[   16472] = 32'hd15be047;
    ram_cell[   16473] = 32'hd7c31f29;
    ram_cell[   16474] = 32'hbe06c1ce;
    ram_cell[   16475] = 32'ha10e705b;
    ram_cell[   16476] = 32'h1a76f9b8;
    ram_cell[   16477] = 32'h4aac875b;
    ram_cell[   16478] = 32'hd8d8a623;
    ram_cell[   16479] = 32'h9cadcbea;
    ram_cell[   16480] = 32'h03c71774;
    ram_cell[   16481] = 32'hf1a0de56;
    ram_cell[   16482] = 32'hcb3e4345;
    ram_cell[   16483] = 32'hf9ba2ce5;
    ram_cell[   16484] = 32'hce9eced5;
    ram_cell[   16485] = 32'hb05ed850;
    ram_cell[   16486] = 32'hd869a2ac;
    ram_cell[   16487] = 32'h3766bccd;
    ram_cell[   16488] = 32'h41269659;
    ram_cell[   16489] = 32'h4c4faed4;
    ram_cell[   16490] = 32'h98e4af51;
    ram_cell[   16491] = 32'h73eb25e4;
    ram_cell[   16492] = 32'h0e2db478;
    ram_cell[   16493] = 32'h633e9fa6;
    ram_cell[   16494] = 32'h782e3c0b;
    ram_cell[   16495] = 32'hd8fcc178;
    ram_cell[   16496] = 32'h6421e1e8;
    ram_cell[   16497] = 32'heb245532;
    ram_cell[   16498] = 32'hf2f9fbb5;
    ram_cell[   16499] = 32'h4a458616;
    ram_cell[   16500] = 32'h6c59d084;
    ram_cell[   16501] = 32'hc250a3ef;
    ram_cell[   16502] = 32'h2cf530fe;
    ram_cell[   16503] = 32'h3601c063;
    ram_cell[   16504] = 32'h3a5e4651;
    ram_cell[   16505] = 32'h83a3385c;
    ram_cell[   16506] = 32'h4ce955e1;
    ram_cell[   16507] = 32'h66b52f31;
    ram_cell[   16508] = 32'h3af0b672;
    ram_cell[   16509] = 32'hc8264f6c;
    ram_cell[   16510] = 32'hba310936;
    ram_cell[   16511] = 32'hc9b3d6d9;
    ram_cell[   16512] = 32'hf0fa42b6;
    ram_cell[   16513] = 32'h45bf9d0c;
    ram_cell[   16514] = 32'h26838fc2;
    ram_cell[   16515] = 32'hed7ea381;
    ram_cell[   16516] = 32'hfa54025d;
    ram_cell[   16517] = 32'h6914e927;
    ram_cell[   16518] = 32'hed93ac00;
    ram_cell[   16519] = 32'h1ef1d322;
    ram_cell[   16520] = 32'h79ebb57e;
    ram_cell[   16521] = 32'h23b6725d;
    ram_cell[   16522] = 32'h7f0295ac;
    ram_cell[   16523] = 32'h9b15936b;
    ram_cell[   16524] = 32'hcb9a7a0f;
    ram_cell[   16525] = 32'h540e816e;
    ram_cell[   16526] = 32'hd8c25be0;
    ram_cell[   16527] = 32'hc84e8597;
    ram_cell[   16528] = 32'hd3378fe1;
    ram_cell[   16529] = 32'he0c28e7f;
    ram_cell[   16530] = 32'h789a34a2;
    ram_cell[   16531] = 32'h4316373f;
    ram_cell[   16532] = 32'h6d13b236;
    ram_cell[   16533] = 32'hf8c6ff23;
    ram_cell[   16534] = 32'h57a9204f;
    ram_cell[   16535] = 32'ha6955e43;
    ram_cell[   16536] = 32'hdabd2f85;
    ram_cell[   16537] = 32'hbdd57b75;
    ram_cell[   16538] = 32'h260d16da;
    ram_cell[   16539] = 32'hf07de7a6;
    ram_cell[   16540] = 32'hde25d204;
    ram_cell[   16541] = 32'h6e9bda4c;
    ram_cell[   16542] = 32'h90f50fa4;
    ram_cell[   16543] = 32'ha1b2ded2;
    ram_cell[   16544] = 32'h2e905440;
    ram_cell[   16545] = 32'hd17c1356;
    ram_cell[   16546] = 32'h1d2ec368;
    ram_cell[   16547] = 32'h8e7872fd;
    ram_cell[   16548] = 32'h10058121;
    ram_cell[   16549] = 32'h2d0273b6;
    ram_cell[   16550] = 32'hf3759b8c;
    ram_cell[   16551] = 32'h0c48a5a4;
    ram_cell[   16552] = 32'hbb92f0a5;
    ram_cell[   16553] = 32'h790b257d;
    ram_cell[   16554] = 32'he2986b25;
    ram_cell[   16555] = 32'h54c16202;
    ram_cell[   16556] = 32'he68b02a4;
    ram_cell[   16557] = 32'hc92d23d8;
    ram_cell[   16558] = 32'h0feb5b94;
    ram_cell[   16559] = 32'h26f84b2b;
    ram_cell[   16560] = 32'h715c9f0d;
    ram_cell[   16561] = 32'h12b87cb8;
    ram_cell[   16562] = 32'hdba9ef78;
    ram_cell[   16563] = 32'h590756b8;
    ram_cell[   16564] = 32'h949ec4d5;
    ram_cell[   16565] = 32'hcdfb9c28;
    ram_cell[   16566] = 32'hd82999d3;
    ram_cell[   16567] = 32'h888c005e;
    ram_cell[   16568] = 32'h6a694826;
    ram_cell[   16569] = 32'h230a9625;
    ram_cell[   16570] = 32'h66d21014;
    ram_cell[   16571] = 32'h00a35e5c;
    ram_cell[   16572] = 32'h0fd26e72;
    ram_cell[   16573] = 32'h40b33e30;
    ram_cell[   16574] = 32'h2329b47d;
    ram_cell[   16575] = 32'hf9ee7a6d;
    ram_cell[   16576] = 32'hb91ad112;
    ram_cell[   16577] = 32'h605b3964;
    ram_cell[   16578] = 32'h976ca99d;
    ram_cell[   16579] = 32'hb76cbb6d;
    ram_cell[   16580] = 32'ha2a5b706;
    ram_cell[   16581] = 32'hcb8dd25d;
    ram_cell[   16582] = 32'h083d47e6;
    ram_cell[   16583] = 32'h738b18ee;
    ram_cell[   16584] = 32'hdbe587b1;
    ram_cell[   16585] = 32'hbc504b81;
    ram_cell[   16586] = 32'h98cf39c8;
    ram_cell[   16587] = 32'haf3f641d;
    ram_cell[   16588] = 32'had3e037f;
    ram_cell[   16589] = 32'hef9667ef;
    ram_cell[   16590] = 32'h81fc4967;
    ram_cell[   16591] = 32'h1a138d88;
    ram_cell[   16592] = 32'hc9e068ec;
    ram_cell[   16593] = 32'h117bce2d;
    ram_cell[   16594] = 32'h9c5b2b96;
    ram_cell[   16595] = 32'h6cf3102d;
    ram_cell[   16596] = 32'h3783362e;
    ram_cell[   16597] = 32'h04964254;
    ram_cell[   16598] = 32'hb77d3d9d;
    ram_cell[   16599] = 32'h45a46890;
    ram_cell[   16600] = 32'h5d4a33f9;
    ram_cell[   16601] = 32'h3b79cd1d;
    ram_cell[   16602] = 32'h86214214;
    ram_cell[   16603] = 32'h19dc558d;
    ram_cell[   16604] = 32'hf5da635c;
    ram_cell[   16605] = 32'h6a19c6d0;
    ram_cell[   16606] = 32'h2d44fa0b;
    ram_cell[   16607] = 32'hfaf3bb7c;
    ram_cell[   16608] = 32'h2ba2504f;
    ram_cell[   16609] = 32'heee86083;
    ram_cell[   16610] = 32'hb464bfad;
    ram_cell[   16611] = 32'hcd3454b8;
    ram_cell[   16612] = 32'hfd106fb4;
    ram_cell[   16613] = 32'h182a4539;
    ram_cell[   16614] = 32'hdd1143ad;
    ram_cell[   16615] = 32'h6b536706;
    ram_cell[   16616] = 32'h206fe575;
    ram_cell[   16617] = 32'he34a6f4b;
    ram_cell[   16618] = 32'hec8cdc2c;
    ram_cell[   16619] = 32'h2b785f0a;
    ram_cell[   16620] = 32'he2f29ed2;
    ram_cell[   16621] = 32'h3822b452;
    ram_cell[   16622] = 32'hf9efbd35;
    ram_cell[   16623] = 32'habd69847;
    ram_cell[   16624] = 32'h7df45ee2;
    ram_cell[   16625] = 32'h331fc427;
    ram_cell[   16626] = 32'h205bb9db;
    ram_cell[   16627] = 32'he1a50a1c;
    ram_cell[   16628] = 32'hf0542aba;
    ram_cell[   16629] = 32'h10cc10c3;
    ram_cell[   16630] = 32'h0ad24b99;
    ram_cell[   16631] = 32'he1a4307b;
    ram_cell[   16632] = 32'hfaa2525f;
    ram_cell[   16633] = 32'hdb882e90;
    ram_cell[   16634] = 32'h5fa0558a;
    ram_cell[   16635] = 32'h4aaf0dca;
    ram_cell[   16636] = 32'h6ec98bff;
    ram_cell[   16637] = 32'h55122481;
    ram_cell[   16638] = 32'h05cca9c7;
    ram_cell[   16639] = 32'h0a471c8c;
    ram_cell[   16640] = 32'h893011c6;
    ram_cell[   16641] = 32'hb0d40d72;
    ram_cell[   16642] = 32'hd3a3faae;
    ram_cell[   16643] = 32'h3b0c57af;
    ram_cell[   16644] = 32'h0fa4bff3;
    ram_cell[   16645] = 32'hde5a3987;
    ram_cell[   16646] = 32'h2d1050e6;
    ram_cell[   16647] = 32'h41e5ba68;
    ram_cell[   16648] = 32'hfe71b5f1;
    ram_cell[   16649] = 32'h2f97c4b0;
    ram_cell[   16650] = 32'h610c11e8;
    ram_cell[   16651] = 32'hc894b00a;
    ram_cell[   16652] = 32'h7b3980df;
    ram_cell[   16653] = 32'hfc320a15;
    ram_cell[   16654] = 32'h8fc5981b;
    ram_cell[   16655] = 32'h6a1291be;
    ram_cell[   16656] = 32'hb1a60743;
    ram_cell[   16657] = 32'hfa514e20;
    ram_cell[   16658] = 32'h9e469710;
    ram_cell[   16659] = 32'hd9f76ed5;
    ram_cell[   16660] = 32'h0c4afcfe;
    ram_cell[   16661] = 32'h591e1225;
    ram_cell[   16662] = 32'h955b2b66;
    ram_cell[   16663] = 32'h6be73176;
    ram_cell[   16664] = 32'hbf3b1d07;
    ram_cell[   16665] = 32'hf7df4703;
    ram_cell[   16666] = 32'h98263120;
    ram_cell[   16667] = 32'h94480274;
    ram_cell[   16668] = 32'h4be648e0;
    ram_cell[   16669] = 32'habf71ac3;
    ram_cell[   16670] = 32'h4bf0b7fa;
    ram_cell[   16671] = 32'hb302e0f0;
    ram_cell[   16672] = 32'h890faaf4;
    ram_cell[   16673] = 32'hd1c22c78;
    ram_cell[   16674] = 32'h20f89996;
    ram_cell[   16675] = 32'ha00fa541;
    ram_cell[   16676] = 32'h58939ada;
    ram_cell[   16677] = 32'h73536d2d;
    ram_cell[   16678] = 32'hab6e4c36;
    ram_cell[   16679] = 32'h6a1d5932;
    ram_cell[   16680] = 32'h471b5d7e;
    ram_cell[   16681] = 32'hc3ba3b71;
    ram_cell[   16682] = 32'h3866d64f;
    ram_cell[   16683] = 32'hc78f0692;
    ram_cell[   16684] = 32'he56e5512;
    ram_cell[   16685] = 32'hbf943ade;
    ram_cell[   16686] = 32'h8839a3a3;
    ram_cell[   16687] = 32'h1befcf61;
    ram_cell[   16688] = 32'h6b303edf;
    ram_cell[   16689] = 32'h363facbf;
    ram_cell[   16690] = 32'h040986aa;
    ram_cell[   16691] = 32'hff01da9c;
    ram_cell[   16692] = 32'h76cfa5b5;
    ram_cell[   16693] = 32'h3da60260;
    ram_cell[   16694] = 32'h40c0c254;
    ram_cell[   16695] = 32'h654758c3;
    ram_cell[   16696] = 32'heebf1356;
    ram_cell[   16697] = 32'h53455cde;
    ram_cell[   16698] = 32'hee71107f;
    ram_cell[   16699] = 32'h9c02a7a7;
    ram_cell[   16700] = 32'h8127df09;
    ram_cell[   16701] = 32'h1c53b97d;
    ram_cell[   16702] = 32'h470caee6;
    ram_cell[   16703] = 32'h54a1d770;
    ram_cell[   16704] = 32'h7b2973ba;
    ram_cell[   16705] = 32'h8684fe18;
    ram_cell[   16706] = 32'h3fe488c2;
    ram_cell[   16707] = 32'hfb484bab;
    ram_cell[   16708] = 32'hca44f156;
    ram_cell[   16709] = 32'hf2bb995b;
    ram_cell[   16710] = 32'h53779624;
    ram_cell[   16711] = 32'h464089e9;
    ram_cell[   16712] = 32'h33900b2c;
    ram_cell[   16713] = 32'he171265d;
    ram_cell[   16714] = 32'h970d405d;
    ram_cell[   16715] = 32'h250e34b2;
    ram_cell[   16716] = 32'h92568c85;
    ram_cell[   16717] = 32'hd26e7e33;
    ram_cell[   16718] = 32'hb16b906c;
    ram_cell[   16719] = 32'hd67dcead;
    ram_cell[   16720] = 32'h7477b708;
    ram_cell[   16721] = 32'h8524ba8e;
    ram_cell[   16722] = 32'h286290e4;
    ram_cell[   16723] = 32'h5fae8504;
    ram_cell[   16724] = 32'hbe60bbd6;
    ram_cell[   16725] = 32'h0598fdc2;
    ram_cell[   16726] = 32'hb2f74ab7;
    ram_cell[   16727] = 32'h222b3e54;
    ram_cell[   16728] = 32'hbe626ca3;
    ram_cell[   16729] = 32'h0ce75537;
    ram_cell[   16730] = 32'hde94cff8;
    ram_cell[   16731] = 32'h8757f43c;
    ram_cell[   16732] = 32'hdf61b46f;
    ram_cell[   16733] = 32'hba2ee8c5;
    ram_cell[   16734] = 32'h40d60722;
    ram_cell[   16735] = 32'hb6394df1;
    ram_cell[   16736] = 32'h23253e10;
    ram_cell[   16737] = 32'heb8747bb;
    ram_cell[   16738] = 32'h841a88f9;
    ram_cell[   16739] = 32'h553eca9a;
    ram_cell[   16740] = 32'h61a98105;
    ram_cell[   16741] = 32'ha7b49826;
    ram_cell[   16742] = 32'hc7e8f825;
    ram_cell[   16743] = 32'h1c92c144;
    ram_cell[   16744] = 32'h6e28aa2a;
    ram_cell[   16745] = 32'h4c73822d;
    ram_cell[   16746] = 32'h29b68c58;
    ram_cell[   16747] = 32'h4c929389;
    ram_cell[   16748] = 32'h83a958d1;
    ram_cell[   16749] = 32'h722b8b95;
    ram_cell[   16750] = 32'hcf53b692;
    ram_cell[   16751] = 32'h0a76314e;
    ram_cell[   16752] = 32'h9ec19d7f;
    ram_cell[   16753] = 32'hffc67daa;
    ram_cell[   16754] = 32'hce6482d0;
    ram_cell[   16755] = 32'hf587a8ca;
    ram_cell[   16756] = 32'h88dda85f;
    ram_cell[   16757] = 32'hb8a73402;
    ram_cell[   16758] = 32'h7661c387;
    ram_cell[   16759] = 32'h52242306;
    ram_cell[   16760] = 32'hd779252a;
    ram_cell[   16761] = 32'h7882c9dc;
    ram_cell[   16762] = 32'h35e35a10;
    ram_cell[   16763] = 32'hfd6637f6;
    ram_cell[   16764] = 32'h4acfcb1b;
    ram_cell[   16765] = 32'h037acb30;
    ram_cell[   16766] = 32'hc7425a32;
    ram_cell[   16767] = 32'hf7f4223e;
    ram_cell[   16768] = 32'h503f5746;
    ram_cell[   16769] = 32'hc3ccafa4;
    ram_cell[   16770] = 32'h8517befc;
    ram_cell[   16771] = 32'hd6aeeff0;
    ram_cell[   16772] = 32'ha1e0138d;
    ram_cell[   16773] = 32'h3e88782c;
    ram_cell[   16774] = 32'h45466905;
    ram_cell[   16775] = 32'h87196021;
    ram_cell[   16776] = 32'h9bea4c48;
    ram_cell[   16777] = 32'h20e3e6ee;
    ram_cell[   16778] = 32'h72bde09d;
    ram_cell[   16779] = 32'h58da40af;
    ram_cell[   16780] = 32'h11c51e5d;
    ram_cell[   16781] = 32'hc864d149;
    ram_cell[   16782] = 32'h9e840580;
    ram_cell[   16783] = 32'h12238010;
    ram_cell[   16784] = 32'h4c84a625;
    ram_cell[   16785] = 32'he87eb0c3;
    ram_cell[   16786] = 32'h668fc742;
    ram_cell[   16787] = 32'hc5aa5d33;
    ram_cell[   16788] = 32'hc242f236;
    ram_cell[   16789] = 32'h04ca0902;
    ram_cell[   16790] = 32'hb6a42630;
    ram_cell[   16791] = 32'h5af19a09;
    ram_cell[   16792] = 32'hd2b57d13;
    ram_cell[   16793] = 32'h564eb1b5;
    ram_cell[   16794] = 32'h7f292555;
    ram_cell[   16795] = 32'h1698c363;
    ram_cell[   16796] = 32'h0d525e0d;
    ram_cell[   16797] = 32'h6a8a1bb4;
    ram_cell[   16798] = 32'haf731384;
    ram_cell[   16799] = 32'h499fef48;
    ram_cell[   16800] = 32'hf3a21c47;
    ram_cell[   16801] = 32'h475d14b3;
    ram_cell[   16802] = 32'h7227e088;
    ram_cell[   16803] = 32'h0242e1d8;
    ram_cell[   16804] = 32'haf361539;
    ram_cell[   16805] = 32'hf7a450d1;
    ram_cell[   16806] = 32'he20ac62c;
    ram_cell[   16807] = 32'h7cdbe7c1;
    ram_cell[   16808] = 32'h98752dcd;
    ram_cell[   16809] = 32'h95c2245c;
    ram_cell[   16810] = 32'h6a160c81;
    ram_cell[   16811] = 32'h1edf28d8;
    ram_cell[   16812] = 32'h9b365806;
    ram_cell[   16813] = 32'hd18c4149;
    ram_cell[   16814] = 32'h8523107c;
    ram_cell[   16815] = 32'hd36de134;
    ram_cell[   16816] = 32'h674f8bc9;
    ram_cell[   16817] = 32'h693817e1;
    ram_cell[   16818] = 32'h0f9e8776;
    ram_cell[   16819] = 32'ha26237e1;
    ram_cell[   16820] = 32'h245b434c;
    ram_cell[   16821] = 32'h8b0872a9;
    ram_cell[   16822] = 32'h1509273d;
    ram_cell[   16823] = 32'h1468372e;
    ram_cell[   16824] = 32'h9cf88581;
    ram_cell[   16825] = 32'hc108b247;
    ram_cell[   16826] = 32'hf1d370ee;
    ram_cell[   16827] = 32'h208d2b19;
    ram_cell[   16828] = 32'hc5560b3b;
    ram_cell[   16829] = 32'hc3e4c17f;
    ram_cell[   16830] = 32'h2ab67060;
    ram_cell[   16831] = 32'h6d4e4fbd;
    ram_cell[   16832] = 32'h8907c83a;
    ram_cell[   16833] = 32'h6441c9ae;
    ram_cell[   16834] = 32'hdce1ff0b;
    ram_cell[   16835] = 32'hb0e2edb6;
    ram_cell[   16836] = 32'h987ab527;
    ram_cell[   16837] = 32'hcd91ceff;
    ram_cell[   16838] = 32'h334af240;
    ram_cell[   16839] = 32'hc2988701;
    ram_cell[   16840] = 32'h688056cc;
    ram_cell[   16841] = 32'hcbace6e2;
    ram_cell[   16842] = 32'h7253ad28;
    ram_cell[   16843] = 32'h0d345716;
    ram_cell[   16844] = 32'h837d324f;
    ram_cell[   16845] = 32'h6f039742;
    ram_cell[   16846] = 32'hf1d373ac;
    ram_cell[   16847] = 32'h82e40007;
    ram_cell[   16848] = 32'h26d8d5aa;
    ram_cell[   16849] = 32'hf1d6f4f0;
    ram_cell[   16850] = 32'ha7b8169a;
    ram_cell[   16851] = 32'hfa8c93e2;
    ram_cell[   16852] = 32'h41c36e4b;
    ram_cell[   16853] = 32'h703c7c5f;
    ram_cell[   16854] = 32'h27564a13;
    ram_cell[   16855] = 32'h9f176719;
    ram_cell[   16856] = 32'h085d274d;
    ram_cell[   16857] = 32'hdc02a955;
    ram_cell[   16858] = 32'h84656c6c;
    ram_cell[   16859] = 32'hf9387ea4;
    ram_cell[   16860] = 32'h090c8be4;
    ram_cell[   16861] = 32'hf5cc8373;
    ram_cell[   16862] = 32'h562d2c22;
    ram_cell[   16863] = 32'h9e62aaf6;
    ram_cell[   16864] = 32'h8ae439ad;
    ram_cell[   16865] = 32'hc8e62c61;
    ram_cell[   16866] = 32'h03118949;
    ram_cell[   16867] = 32'h41bde2c0;
    ram_cell[   16868] = 32'h62a4bf75;
    ram_cell[   16869] = 32'hf3eaca26;
    ram_cell[   16870] = 32'h5d8c24af;
    ram_cell[   16871] = 32'h49194636;
    ram_cell[   16872] = 32'h434814f5;
    ram_cell[   16873] = 32'h309b9c80;
    ram_cell[   16874] = 32'h8a883b7c;
    ram_cell[   16875] = 32'h3edc1d29;
    ram_cell[   16876] = 32'hcde46700;
    ram_cell[   16877] = 32'h2ad191ef;
    ram_cell[   16878] = 32'hd5796adb;
    ram_cell[   16879] = 32'hce682e37;
    ram_cell[   16880] = 32'hcfc55bf4;
    ram_cell[   16881] = 32'h23b16a91;
    ram_cell[   16882] = 32'h7d62cf90;
    ram_cell[   16883] = 32'h4377173e;
    ram_cell[   16884] = 32'h93743acd;
    ram_cell[   16885] = 32'h2247bd6c;
    ram_cell[   16886] = 32'hc6b95b4d;
    ram_cell[   16887] = 32'h913a1a46;
    ram_cell[   16888] = 32'h94bf7e01;
    ram_cell[   16889] = 32'hf33ac9c2;
    ram_cell[   16890] = 32'hefbc4edc;
    ram_cell[   16891] = 32'he28d573f;
    ram_cell[   16892] = 32'hd3913089;
    ram_cell[   16893] = 32'h3bf6e8d4;
    ram_cell[   16894] = 32'hda0aeb16;
    ram_cell[   16895] = 32'h48926487;
    ram_cell[   16896] = 32'h1ef71d24;
    ram_cell[   16897] = 32'h718cc729;
    ram_cell[   16898] = 32'hcef0c3fa;
    ram_cell[   16899] = 32'h03fbb3b4;
    ram_cell[   16900] = 32'h56b320b6;
    ram_cell[   16901] = 32'h0986f202;
    ram_cell[   16902] = 32'hda520faf;
    ram_cell[   16903] = 32'hb2742565;
    ram_cell[   16904] = 32'hf802f2cc;
    ram_cell[   16905] = 32'h74823636;
    ram_cell[   16906] = 32'hf48914a8;
    ram_cell[   16907] = 32'h3bf3673f;
    ram_cell[   16908] = 32'h82414ffb;
    ram_cell[   16909] = 32'h8bd500eb;
    ram_cell[   16910] = 32'hb0292c05;
    ram_cell[   16911] = 32'hc38211af;
    ram_cell[   16912] = 32'ha3e2bfdf;
    ram_cell[   16913] = 32'hf1821082;
    ram_cell[   16914] = 32'h7bf28ffb;
    ram_cell[   16915] = 32'h1c4ed95a;
    ram_cell[   16916] = 32'h2ed6b0f9;
    ram_cell[   16917] = 32'h955d32f3;
    ram_cell[   16918] = 32'h1cfca2fe;
    ram_cell[   16919] = 32'hed1ea10e;
    ram_cell[   16920] = 32'h0124b9f2;
    ram_cell[   16921] = 32'h7fa4f08d;
    ram_cell[   16922] = 32'heb391f0e;
    ram_cell[   16923] = 32'h47a903c6;
    ram_cell[   16924] = 32'h4ab33fd5;
    ram_cell[   16925] = 32'h924f8cf6;
    ram_cell[   16926] = 32'h5daad54f;
    ram_cell[   16927] = 32'h97ac07c4;
    ram_cell[   16928] = 32'h58f4edfa;
    ram_cell[   16929] = 32'h7e420e6d;
    ram_cell[   16930] = 32'h341509ea;
    ram_cell[   16931] = 32'hdf8e16ed;
    ram_cell[   16932] = 32'hd2ac1acd;
    ram_cell[   16933] = 32'h7746b85e;
    ram_cell[   16934] = 32'h91e7dedc;
    ram_cell[   16935] = 32'h16b8916d;
    ram_cell[   16936] = 32'h4bdf1d74;
    ram_cell[   16937] = 32'h3da66b94;
    ram_cell[   16938] = 32'h5fe4e5d0;
    ram_cell[   16939] = 32'h7a3671f9;
    ram_cell[   16940] = 32'h9d591047;
    ram_cell[   16941] = 32'h1262258d;
    ram_cell[   16942] = 32'h6d2290d9;
    ram_cell[   16943] = 32'hfcf6027c;
    ram_cell[   16944] = 32'h34e3ab65;
    ram_cell[   16945] = 32'h01e47494;
    ram_cell[   16946] = 32'h78d916bf;
    ram_cell[   16947] = 32'h06cdf43f;
    ram_cell[   16948] = 32'hbb854436;
    ram_cell[   16949] = 32'hfe6bf3d7;
    ram_cell[   16950] = 32'hd626578d;
    ram_cell[   16951] = 32'hc8bd8877;
    ram_cell[   16952] = 32'hf8d58c10;
    ram_cell[   16953] = 32'h4f5a928a;
    ram_cell[   16954] = 32'h8f1bc1ca;
    ram_cell[   16955] = 32'h9039edd9;
    ram_cell[   16956] = 32'hcc8603d1;
    ram_cell[   16957] = 32'hd496bf38;
    ram_cell[   16958] = 32'hb03f3e7d;
    ram_cell[   16959] = 32'h2f91d80c;
    ram_cell[   16960] = 32'hfd85e1d8;
    ram_cell[   16961] = 32'h0a72a34c;
    ram_cell[   16962] = 32'h34a7ff27;
    ram_cell[   16963] = 32'h2e71c99d;
    ram_cell[   16964] = 32'h0ad8500e;
    ram_cell[   16965] = 32'hac909f4b;
    ram_cell[   16966] = 32'he12a00c9;
    ram_cell[   16967] = 32'h0952e002;
    ram_cell[   16968] = 32'h1243fe06;
    ram_cell[   16969] = 32'h830d9239;
    ram_cell[   16970] = 32'h6e31a58b;
    ram_cell[   16971] = 32'ha0bc52de;
    ram_cell[   16972] = 32'hb3f4e668;
    ram_cell[   16973] = 32'h15be75f8;
    ram_cell[   16974] = 32'h29b16567;
    ram_cell[   16975] = 32'hbc8a6f32;
    ram_cell[   16976] = 32'h8dd2bc0e;
    ram_cell[   16977] = 32'hfaa0f4f4;
    ram_cell[   16978] = 32'h0bf56a26;
    ram_cell[   16979] = 32'h51ada65a;
    ram_cell[   16980] = 32'h7cadbb91;
    ram_cell[   16981] = 32'hc90edeea;
    ram_cell[   16982] = 32'hcd29c8b0;
    ram_cell[   16983] = 32'h6dd89590;
    ram_cell[   16984] = 32'h1ab4496d;
    ram_cell[   16985] = 32'h68d0c93c;
    ram_cell[   16986] = 32'h469c5e8d;
    ram_cell[   16987] = 32'h0e5bfbeb;
    ram_cell[   16988] = 32'h753e09fa;
    ram_cell[   16989] = 32'h47a0ac88;
    ram_cell[   16990] = 32'h57809e5c;
    ram_cell[   16991] = 32'he1ae36d2;
    ram_cell[   16992] = 32'h6094cc7b;
    ram_cell[   16993] = 32'h058cb41a;
    ram_cell[   16994] = 32'hc14a106b;
    ram_cell[   16995] = 32'hd8e58d93;
    ram_cell[   16996] = 32'h431c1d9c;
    ram_cell[   16997] = 32'hc314f4a1;
    ram_cell[   16998] = 32'hf918b496;
    ram_cell[   16999] = 32'h67dc1e39;
    ram_cell[   17000] = 32'h04294776;
    ram_cell[   17001] = 32'h2dbb0778;
    ram_cell[   17002] = 32'h58cea04f;
    ram_cell[   17003] = 32'h42b67141;
    ram_cell[   17004] = 32'h1827988d;
    ram_cell[   17005] = 32'h90c05830;
    ram_cell[   17006] = 32'ha57c1277;
    ram_cell[   17007] = 32'h64c1ed7a;
    ram_cell[   17008] = 32'h75893e29;
    ram_cell[   17009] = 32'h74bae5c1;
    ram_cell[   17010] = 32'hea3f1ff2;
    ram_cell[   17011] = 32'hfe66d146;
    ram_cell[   17012] = 32'h83267f13;
    ram_cell[   17013] = 32'haad6961e;
    ram_cell[   17014] = 32'h2ff74564;
    ram_cell[   17015] = 32'h112087ca;
    ram_cell[   17016] = 32'h550d85eb;
    ram_cell[   17017] = 32'h1766d9a5;
    ram_cell[   17018] = 32'hbd209aed;
    ram_cell[   17019] = 32'h4b8238c3;
    ram_cell[   17020] = 32'h7ba8bc45;
    ram_cell[   17021] = 32'h10e879a6;
    ram_cell[   17022] = 32'heb22a88b;
    ram_cell[   17023] = 32'h63072c75;
    ram_cell[   17024] = 32'hb482dabb;
    ram_cell[   17025] = 32'hc65feaeb;
    ram_cell[   17026] = 32'h30b8caef;
    ram_cell[   17027] = 32'h0a9e8e6e;
    ram_cell[   17028] = 32'haf5303f8;
    ram_cell[   17029] = 32'h898f9c60;
    ram_cell[   17030] = 32'h5879ca26;
    ram_cell[   17031] = 32'hfba75668;
    ram_cell[   17032] = 32'he54fdd2c;
    ram_cell[   17033] = 32'hd9834940;
    ram_cell[   17034] = 32'h1db522e8;
    ram_cell[   17035] = 32'h6c2afd8a;
    ram_cell[   17036] = 32'he4ed50e3;
    ram_cell[   17037] = 32'h990da0c8;
    ram_cell[   17038] = 32'h2ef949cd;
    ram_cell[   17039] = 32'hc2b5ae69;
    ram_cell[   17040] = 32'h339dd17e;
    ram_cell[   17041] = 32'h88a7eb9d;
    ram_cell[   17042] = 32'h6954a25e;
    ram_cell[   17043] = 32'hfca11882;
    ram_cell[   17044] = 32'h7f727e26;
    ram_cell[   17045] = 32'h38f374d3;
    ram_cell[   17046] = 32'hb081dff8;
    ram_cell[   17047] = 32'hef0f202f;
    ram_cell[   17048] = 32'h7f94198e;
    ram_cell[   17049] = 32'hc5a206bf;
    ram_cell[   17050] = 32'hafeb2b56;
    ram_cell[   17051] = 32'hbf7e5add;
    ram_cell[   17052] = 32'hfa4df228;
    ram_cell[   17053] = 32'hee43047b;
    ram_cell[   17054] = 32'hb356b744;
    ram_cell[   17055] = 32'h3295a8c0;
    ram_cell[   17056] = 32'h167e2880;
    ram_cell[   17057] = 32'h79e2ab3e;
    ram_cell[   17058] = 32'h676893b7;
    ram_cell[   17059] = 32'h3bfa7d1a;
    ram_cell[   17060] = 32'h45ae3e36;
    ram_cell[   17061] = 32'h09dafe33;
    ram_cell[   17062] = 32'h019f29e1;
    ram_cell[   17063] = 32'h3d3c87b9;
    ram_cell[   17064] = 32'hb2766f7e;
    ram_cell[   17065] = 32'hc33dc93e;
    ram_cell[   17066] = 32'h24add37d;
    ram_cell[   17067] = 32'hdea0e45b;
    ram_cell[   17068] = 32'h6a702014;
    ram_cell[   17069] = 32'h04c25ab8;
    ram_cell[   17070] = 32'h2e998bcc;
    ram_cell[   17071] = 32'h4d280dba;
    ram_cell[   17072] = 32'hfead9ce1;
    ram_cell[   17073] = 32'h673be5a7;
    ram_cell[   17074] = 32'haf340fbd;
    ram_cell[   17075] = 32'h522e9a8c;
    ram_cell[   17076] = 32'hc7b21953;
    ram_cell[   17077] = 32'hbc4b7e0f;
    ram_cell[   17078] = 32'h7bac270a;
    ram_cell[   17079] = 32'hab0e020b;
    ram_cell[   17080] = 32'ha2ccf5ef;
    ram_cell[   17081] = 32'h1f8c2be9;
    ram_cell[   17082] = 32'h9becaf3b;
    ram_cell[   17083] = 32'h35f032f1;
    ram_cell[   17084] = 32'he72ce56b;
    ram_cell[   17085] = 32'h7aa6fea5;
    ram_cell[   17086] = 32'hf910035a;
    ram_cell[   17087] = 32'hd652b8cc;
    ram_cell[   17088] = 32'h5c3a498f;
    ram_cell[   17089] = 32'h27eba048;
    ram_cell[   17090] = 32'haf04ba83;
    ram_cell[   17091] = 32'h9cdcad63;
    ram_cell[   17092] = 32'h29fe816e;
    ram_cell[   17093] = 32'h60819924;
    ram_cell[   17094] = 32'h36147af0;
    ram_cell[   17095] = 32'hd6e3d717;
    ram_cell[   17096] = 32'h800a8b81;
    ram_cell[   17097] = 32'h86144504;
    ram_cell[   17098] = 32'h0c859d58;
    ram_cell[   17099] = 32'hc99ef15e;
    ram_cell[   17100] = 32'hd141c0db;
    ram_cell[   17101] = 32'hd62a7ef8;
    ram_cell[   17102] = 32'h0a34d387;
    ram_cell[   17103] = 32'h49a10c91;
    ram_cell[   17104] = 32'hb9679ce8;
    ram_cell[   17105] = 32'he6469c86;
    ram_cell[   17106] = 32'h8e0b2a9c;
    ram_cell[   17107] = 32'he14159a6;
    ram_cell[   17108] = 32'h96541234;
    ram_cell[   17109] = 32'h95287083;
    ram_cell[   17110] = 32'h0055a550;
    ram_cell[   17111] = 32'hd40c4ede;
    ram_cell[   17112] = 32'h838aa16d;
    ram_cell[   17113] = 32'h57581904;
    ram_cell[   17114] = 32'h3d2464be;
    ram_cell[   17115] = 32'ha5bc3510;
    ram_cell[   17116] = 32'hb50cfb58;
    ram_cell[   17117] = 32'hcd9e5dbe;
    ram_cell[   17118] = 32'h8fabeddc;
    ram_cell[   17119] = 32'h29923e3c;
    ram_cell[   17120] = 32'h19487baa;
    ram_cell[   17121] = 32'h51803d2b;
    ram_cell[   17122] = 32'he4c37754;
    ram_cell[   17123] = 32'ha7f30685;
    ram_cell[   17124] = 32'h3c6b7c67;
    ram_cell[   17125] = 32'h3ef9f3c4;
    ram_cell[   17126] = 32'hee60f7dd;
    ram_cell[   17127] = 32'h52f3585e;
    ram_cell[   17128] = 32'ha27a8c6a;
    ram_cell[   17129] = 32'h800bfd32;
    ram_cell[   17130] = 32'h2331400f;
    ram_cell[   17131] = 32'he5332af8;
    ram_cell[   17132] = 32'h20445836;
    ram_cell[   17133] = 32'h82c2a718;
    ram_cell[   17134] = 32'h99111d8c;
    ram_cell[   17135] = 32'h5d959ad3;
    ram_cell[   17136] = 32'h5649f0c7;
    ram_cell[   17137] = 32'h27c1459d;
    ram_cell[   17138] = 32'h3daab101;
    ram_cell[   17139] = 32'h22dac171;
    ram_cell[   17140] = 32'h2d0f9f16;
    ram_cell[   17141] = 32'hbb577022;
    ram_cell[   17142] = 32'h37b7e86f;
    ram_cell[   17143] = 32'hb5e95065;
    ram_cell[   17144] = 32'ha3a49b35;
    ram_cell[   17145] = 32'hc99fb5db;
    ram_cell[   17146] = 32'h953b65a5;
    ram_cell[   17147] = 32'h4c9c6fa3;
    ram_cell[   17148] = 32'hf12f1280;
    ram_cell[   17149] = 32'h6adc0102;
    ram_cell[   17150] = 32'h3da7c9be;
    ram_cell[   17151] = 32'hca5110ea;
    ram_cell[   17152] = 32'h31d355cb;
    ram_cell[   17153] = 32'h979ab7d1;
    ram_cell[   17154] = 32'hd4e617a2;
    ram_cell[   17155] = 32'he5b5e3fe;
    ram_cell[   17156] = 32'hab1ab15e;
    ram_cell[   17157] = 32'h55bdb69e;
    ram_cell[   17158] = 32'h9457e844;
    ram_cell[   17159] = 32'h9ecc1591;
    ram_cell[   17160] = 32'h19585b72;
    ram_cell[   17161] = 32'h8307108b;
    ram_cell[   17162] = 32'he2e7a4f6;
    ram_cell[   17163] = 32'hae6edc8d;
    ram_cell[   17164] = 32'hac5a11c7;
    ram_cell[   17165] = 32'h448d06b5;
    ram_cell[   17166] = 32'hb021067d;
    ram_cell[   17167] = 32'h9553041b;
    ram_cell[   17168] = 32'hf469c6e2;
    ram_cell[   17169] = 32'h5c2b208d;
    ram_cell[   17170] = 32'h133c870d;
    ram_cell[   17171] = 32'he2bb0b39;
    ram_cell[   17172] = 32'h9353ff06;
    ram_cell[   17173] = 32'h8db1b9e5;
    ram_cell[   17174] = 32'hef457d52;
    ram_cell[   17175] = 32'hf83a7f8d;
    ram_cell[   17176] = 32'hdc4feb8e;
    ram_cell[   17177] = 32'hc8526dd1;
    ram_cell[   17178] = 32'h017251cb;
    ram_cell[   17179] = 32'he5421396;
    ram_cell[   17180] = 32'h93c4a2aa;
    ram_cell[   17181] = 32'h7420960c;
    ram_cell[   17182] = 32'hbebc83ae;
    ram_cell[   17183] = 32'h03aedc1d;
    ram_cell[   17184] = 32'hf1e78fac;
    ram_cell[   17185] = 32'h2e1abfa4;
    ram_cell[   17186] = 32'hbc08444c;
    ram_cell[   17187] = 32'h508a3484;
    ram_cell[   17188] = 32'he7c9d48d;
    ram_cell[   17189] = 32'h38383e8a;
    ram_cell[   17190] = 32'h7eb18d5a;
    ram_cell[   17191] = 32'h5ff73ae3;
    ram_cell[   17192] = 32'hbf742311;
    ram_cell[   17193] = 32'haeb7da2f;
    ram_cell[   17194] = 32'h02fce7e4;
    ram_cell[   17195] = 32'h85d87869;
    ram_cell[   17196] = 32'h33115880;
    ram_cell[   17197] = 32'h9538d19e;
    ram_cell[   17198] = 32'hfef7a284;
    ram_cell[   17199] = 32'hf4ecd78a;
    ram_cell[   17200] = 32'h2f43bcab;
    ram_cell[   17201] = 32'h6f1d37fe;
    ram_cell[   17202] = 32'hba216c2e;
    ram_cell[   17203] = 32'h38f912ee;
    ram_cell[   17204] = 32'h101d8a2e;
    ram_cell[   17205] = 32'hdfee766d;
    ram_cell[   17206] = 32'h76202a6f;
    ram_cell[   17207] = 32'h392f945b;
    ram_cell[   17208] = 32'h407562fa;
    ram_cell[   17209] = 32'h6ea7ae44;
    ram_cell[   17210] = 32'h537711ed;
    ram_cell[   17211] = 32'hda18778a;
    ram_cell[   17212] = 32'h148c4ddf;
    ram_cell[   17213] = 32'hc85aaf50;
    ram_cell[   17214] = 32'h7d34bd0b;
    ram_cell[   17215] = 32'h715c19ec;
    ram_cell[   17216] = 32'h9c76431f;
    ram_cell[   17217] = 32'hf76e9aa6;
    ram_cell[   17218] = 32'h08fcb4ad;
    ram_cell[   17219] = 32'h3934d8bf;
    ram_cell[   17220] = 32'h5cb20123;
    ram_cell[   17221] = 32'h599db21c;
    ram_cell[   17222] = 32'hfd14113d;
    ram_cell[   17223] = 32'h7b70f30a;
    ram_cell[   17224] = 32'hb0044b72;
    ram_cell[   17225] = 32'he4b50f14;
    ram_cell[   17226] = 32'h8de8622c;
    ram_cell[   17227] = 32'hcdd598e9;
    ram_cell[   17228] = 32'h307e2056;
    ram_cell[   17229] = 32'h7abb51ad;
    ram_cell[   17230] = 32'hb516268a;
    ram_cell[   17231] = 32'h4ac44e9c;
    ram_cell[   17232] = 32'h4fb57a26;
    ram_cell[   17233] = 32'hd68c81ee;
    ram_cell[   17234] = 32'h7537f66d;
    ram_cell[   17235] = 32'h2e108d9c;
    ram_cell[   17236] = 32'h52bbbf37;
    ram_cell[   17237] = 32'hf68217c7;
    ram_cell[   17238] = 32'he9acdb90;
    ram_cell[   17239] = 32'h3217e42b;
    ram_cell[   17240] = 32'h6a500229;
    ram_cell[   17241] = 32'hbac38507;
    ram_cell[   17242] = 32'h54437ad7;
    ram_cell[   17243] = 32'h330c8ef9;
    ram_cell[   17244] = 32'h61f6c9c2;
    ram_cell[   17245] = 32'h2dca0f36;
    ram_cell[   17246] = 32'hd111032b;
    ram_cell[   17247] = 32'hc923cc22;
    ram_cell[   17248] = 32'h702193c4;
    ram_cell[   17249] = 32'h939b0564;
    ram_cell[   17250] = 32'ha9075997;
    ram_cell[   17251] = 32'h26f92d3e;
    ram_cell[   17252] = 32'h543aa94f;
    ram_cell[   17253] = 32'he12a7ab9;
    ram_cell[   17254] = 32'he64cd70a;
    ram_cell[   17255] = 32'h21442f8b;
    ram_cell[   17256] = 32'h64deb74c;
    ram_cell[   17257] = 32'h0b7bc9d9;
    ram_cell[   17258] = 32'hb3684e35;
    ram_cell[   17259] = 32'h7c9608d5;
    ram_cell[   17260] = 32'he20fa5e8;
    ram_cell[   17261] = 32'hec3fbd4e;
    ram_cell[   17262] = 32'h63634ba9;
    ram_cell[   17263] = 32'h2f462106;
    ram_cell[   17264] = 32'hfba4e7a0;
    ram_cell[   17265] = 32'h7c5d28ed;
    ram_cell[   17266] = 32'hd89333b7;
    ram_cell[   17267] = 32'h2fba6cc6;
    ram_cell[   17268] = 32'h7dc3d7e8;
    ram_cell[   17269] = 32'heb3724f2;
    ram_cell[   17270] = 32'h62491d83;
    ram_cell[   17271] = 32'h9b6996b8;
    ram_cell[   17272] = 32'h779dcf91;
    ram_cell[   17273] = 32'hd94b60de;
    ram_cell[   17274] = 32'hbddc04ef;
    ram_cell[   17275] = 32'h4d32c700;
    ram_cell[   17276] = 32'hf9667eb7;
    ram_cell[   17277] = 32'haa529dd8;
    ram_cell[   17278] = 32'h773ca898;
    ram_cell[   17279] = 32'hff786fe5;
    ram_cell[   17280] = 32'h3c26dd61;
    ram_cell[   17281] = 32'h9eac7193;
    ram_cell[   17282] = 32'h68526e43;
    ram_cell[   17283] = 32'hc058ecff;
    ram_cell[   17284] = 32'hab7b7b55;
    ram_cell[   17285] = 32'h0ce825bb;
    ram_cell[   17286] = 32'he5ce3f8d;
    ram_cell[   17287] = 32'h304bee2b;
    ram_cell[   17288] = 32'h8ea4fdc8;
    ram_cell[   17289] = 32'h41c4224e;
    ram_cell[   17290] = 32'hced2c3c7;
    ram_cell[   17291] = 32'hd06b639e;
    ram_cell[   17292] = 32'h3a3008c6;
    ram_cell[   17293] = 32'hd3abc334;
    ram_cell[   17294] = 32'h7affad91;
    ram_cell[   17295] = 32'hf126abff;
    ram_cell[   17296] = 32'h23c4e3b8;
    ram_cell[   17297] = 32'h3ddd0865;
    ram_cell[   17298] = 32'h82fe2199;
    ram_cell[   17299] = 32'hbc037c12;
    ram_cell[   17300] = 32'h552d5305;
    ram_cell[   17301] = 32'h49123a57;
    ram_cell[   17302] = 32'h89b302ff;
    ram_cell[   17303] = 32'h07c2d8d4;
    ram_cell[   17304] = 32'h6a8a5827;
    ram_cell[   17305] = 32'h544a5022;
    ram_cell[   17306] = 32'h5f7d9d75;
    ram_cell[   17307] = 32'haf46d45e;
    ram_cell[   17308] = 32'he18b27b9;
    ram_cell[   17309] = 32'h9eacc1de;
    ram_cell[   17310] = 32'ha89c5487;
    ram_cell[   17311] = 32'h65ec8e48;
    ram_cell[   17312] = 32'h1c71331b;
    ram_cell[   17313] = 32'hb6d25ce6;
    ram_cell[   17314] = 32'hc20f5623;
    ram_cell[   17315] = 32'h9d534021;
    ram_cell[   17316] = 32'h84324318;
    ram_cell[   17317] = 32'hf6f1c71d;
    ram_cell[   17318] = 32'h3d575ebe;
    ram_cell[   17319] = 32'h30949c56;
    ram_cell[   17320] = 32'h6996e789;
    ram_cell[   17321] = 32'h187925f1;
    ram_cell[   17322] = 32'hd75363ce;
    ram_cell[   17323] = 32'h33dcd97d;
    ram_cell[   17324] = 32'h2fe6c60b;
    ram_cell[   17325] = 32'h129ca445;
    ram_cell[   17326] = 32'h598c12d9;
    ram_cell[   17327] = 32'h6ba717e0;
    ram_cell[   17328] = 32'h08840c53;
    ram_cell[   17329] = 32'h33e8ad31;
    ram_cell[   17330] = 32'h522fe41e;
    ram_cell[   17331] = 32'hb7f4b7ac;
    ram_cell[   17332] = 32'he2d0fe0e;
    ram_cell[   17333] = 32'h3f7d0034;
    ram_cell[   17334] = 32'hcc8d7b02;
    ram_cell[   17335] = 32'h6c6f7cb3;
    ram_cell[   17336] = 32'h2b68805e;
    ram_cell[   17337] = 32'h7b132d84;
    ram_cell[   17338] = 32'haa6a25d2;
    ram_cell[   17339] = 32'he310be58;
    ram_cell[   17340] = 32'hf3bd9ca0;
    ram_cell[   17341] = 32'hd8c52039;
    ram_cell[   17342] = 32'haae2d80c;
    ram_cell[   17343] = 32'h989e7062;
    ram_cell[   17344] = 32'h88de0170;
    ram_cell[   17345] = 32'h5e9bd6f2;
    ram_cell[   17346] = 32'h09ca9085;
    ram_cell[   17347] = 32'h287ba6b9;
    ram_cell[   17348] = 32'h88861c91;
    ram_cell[   17349] = 32'h3f08e37c;
    ram_cell[   17350] = 32'heca952f9;
    ram_cell[   17351] = 32'h0cfa7778;
    ram_cell[   17352] = 32'h6af7e245;
    ram_cell[   17353] = 32'h8ec58f7a;
    ram_cell[   17354] = 32'hb35d1dd3;
    ram_cell[   17355] = 32'hcd7508bb;
    ram_cell[   17356] = 32'hd16d6537;
    ram_cell[   17357] = 32'ha93f653e;
    ram_cell[   17358] = 32'h9e70bce3;
    ram_cell[   17359] = 32'he520b512;
    ram_cell[   17360] = 32'hd8026834;
    ram_cell[   17361] = 32'h7b7c38f8;
    ram_cell[   17362] = 32'he764610c;
    ram_cell[   17363] = 32'h35157bab;
    ram_cell[   17364] = 32'hc0b29d28;
    ram_cell[   17365] = 32'h2aa3f4ba;
    ram_cell[   17366] = 32'h35a7e40c;
    ram_cell[   17367] = 32'hc54b4351;
    ram_cell[   17368] = 32'hd5ab821c;
    ram_cell[   17369] = 32'h4ab39576;
    ram_cell[   17370] = 32'ha3a2a3fa;
    ram_cell[   17371] = 32'hcdb5333e;
    ram_cell[   17372] = 32'hc83f072a;
    ram_cell[   17373] = 32'he8cc2e7d;
    ram_cell[   17374] = 32'h3ed3f72d;
    ram_cell[   17375] = 32'hd273a0ba;
    ram_cell[   17376] = 32'hcd3a1790;
    ram_cell[   17377] = 32'hb8c4bd04;
    ram_cell[   17378] = 32'h317a0d6b;
    ram_cell[   17379] = 32'hf419c03c;
    ram_cell[   17380] = 32'h9c91124b;
    ram_cell[   17381] = 32'hcdaa27c6;
    ram_cell[   17382] = 32'hbd2282e0;
    ram_cell[   17383] = 32'hf23b48b8;
    ram_cell[   17384] = 32'h4f5ea29b;
    ram_cell[   17385] = 32'hbeb563e3;
    ram_cell[   17386] = 32'h9fe6ed03;
    ram_cell[   17387] = 32'hc1a7f793;
    ram_cell[   17388] = 32'ha6b464a3;
    ram_cell[   17389] = 32'h07658465;
    ram_cell[   17390] = 32'he08c9700;
    ram_cell[   17391] = 32'h4ef8b0f1;
    ram_cell[   17392] = 32'h4fb630fd;
    ram_cell[   17393] = 32'hd65742cd;
    ram_cell[   17394] = 32'h1724cf8e;
    ram_cell[   17395] = 32'hed4f850b;
    ram_cell[   17396] = 32'h267fe947;
    ram_cell[   17397] = 32'hd8c3b53a;
    ram_cell[   17398] = 32'hb14b727b;
    ram_cell[   17399] = 32'hd4a9185f;
    ram_cell[   17400] = 32'h57d56d63;
    ram_cell[   17401] = 32'hb7c831b3;
    ram_cell[   17402] = 32'hd0c5094e;
    ram_cell[   17403] = 32'h5e22fc73;
    ram_cell[   17404] = 32'h61dfd15d;
    ram_cell[   17405] = 32'he6e267d1;
    ram_cell[   17406] = 32'ha0091fbd;
    ram_cell[   17407] = 32'h60c595c8;
    ram_cell[   17408] = 32'h2d0bbc9b;
    ram_cell[   17409] = 32'hfcd5c76f;
    ram_cell[   17410] = 32'h6fb2af06;
    ram_cell[   17411] = 32'h633d2d59;
    ram_cell[   17412] = 32'h58998880;
    ram_cell[   17413] = 32'ha290bc38;
    ram_cell[   17414] = 32'hcae53dca;
    ram_cell[   17415] = 32'h52527de5;
    ram_cell[   17416] = 32'hcf42435d;
    ram_cell[   17417] = 32'hf4a904f6;
    ram_cell[   17418] = 32'h71c12d1f;
    ram_cell[   17419] = 32'ha8c5c5d6;
    ram_cell[   17420] = 32'ha7d56b21;
    ram_cell[   17421] = 32'hab3b4bf0;
    ram_cell[   17422] = 32'hb93ce7f6;
    ram_cell[   17423] = 32'h6c146e32;
    ram_cell[   17424] = 32'heab37714;
    ram_cell[   17425] = 32'hf88bb8c2;
    ram_cell[   17426] = 32'h718cc470;
    ram_cell[   17427] = 32'hc1105ad4;
    ram_cell[   17428] = 32'h387323d2;
    ram_cell[   17429] = 32'hbfc7ffb1;
    ram_cell[   17430] = 32'ha20872e5;
    ram_cell[   17431] = 32'hd5714d14;
    ram_cell[   17432] = 32'h115c1a9b;
    ram_cell[   17433] = 32'h7362100e;
    ram_cell[   17434] = 32'h507b04ec;
    ram_cell[   17435] = 32'hf9c0be9f;
    ram_cell[   17436] = 32'h57f022d3;
    ram_cell[   17437] = 32'h9b62cb54;
    ram_cell[   17438] = 32'h72bf0a1d;
    ram_cell[   17439] = 32'he4c55bb6;
    ram_cell[   17440] = 32'h3aa4975b;
    ram_cell[   17441] = 32'ha13c2507;
    ram_cell[   17442] = 32'he166d031;
    ram_cell[   17443] = 32'h1294a33e;
    ram_cell[   17444] = 32'hb3022d20;
    ram_cell[   17445] = 32'h0a0fdd03;
    ram_cell[   17446] = 32'h2de35ace;
    ram_cell[   17447] = 32'hdb7fe537;
    ram_cell[   17448] = 32'hecb93074;
    ram_cell[   17449] = 32'h41026b08;
    ram_cell[   17450] = 32'hf48fb3d6;
    ram_cell[   17451] = 32'h1d7042b7;
    ram_cell[   17452] = 32'ha4e26ffa;
    ram_cell[   17453] = 32'h8c085900;
    ram_cell[   17454] = 32'h16498644;
    ram_cell[   17455] = 32'hb6ad1e40;
    ram_cell[   17456] = 32'h097b1dc7;
    ram_cell[   17457] = 32'h40a86cff;
    ram_cell[   17458] = 32'h2f3365e8;
    ram_cell[   17459] = 32'hcc0e998d;
    ram_cell[   17460] = 32'h089ea5e6;
    ram_cell[   17461] = 32'ha63fa023;
    ram_cell[   17462] = 32'h65c020c8;
    ram_cell[   17463] = 32'h2ca1bc8e;
    ram_cell[   17464] = 32'h8d1030db;
    ram_cell[   17465] = 32'hc12e5218;
    ram_cell[   17466] = 32'h60b82ee0;
    ram_cell[   17467] = 32'h93db0945;
    ram_cell[   17468] = 32'he84d89fd;
    ram_cell[   17469] = 32'h287fac23;
    ram_cell[   17470] = 32'h0b284962;
    ram_cell[   17471] = 32'hdbaf5da3;
    ram_cell[   17472] = 32'h4d375bb5;
    ram_cell[   17473] = 32'h24c3927b;
    ram_cell[   17474] = 32'hd26b143d;
    ram_cell[   17475] = 32'h0dc8d96c;
    ram_cell[   17476] = 32'h554f474e;
    ram_cell[   17477] = 32'h2ec74ee8;
    ram_cell[   17478] = 32'hcb65ea10;
    ram_cell[   17479] = 32'hb239cd5d;
    ram_cell[   17480] = 32'h79997a62;
    ram_cell[   17481] = 32'h909d7838;
    ram_cell[   17482] = 32'h18fe2b11;
    ram_cell[   17483] = 32'h589c57ae;
    ram_cell[   17484] = 32'hd2eae7e5;
    ram_cell[   17485] = 32'hdca925b4;
    ram_cell[   17486] = 32'h92c85284;
    ram_cell[   17487] = 32'h5fcff5cf;
    ram_cell[   17488] = 32'hed9346ab;
    ram_cell[   17489] = 32'h376037a2;
    ram_cell[   17490] = 32'hd2f41c8d;
    ram_cell[   17491] = 32'h59a9dcb2;
    ram_cell[   17492] = 32'hb8b778c1;
    ram_cell[   17493] = 32'h9cf1f3d7;
    ram_cell[   17494] = 32'hd72af199;
    ram_cell[   17495] = 32'hc248e2e4;
    ram_cell[   17496] = 32'h91ff17f6;
    ram_cell[   17497] = 32'h87a0600b;
    ram_cell[   17498] = 32'h397a8f06;
    ram_cell[   17499] = 32'h500c1ba4;
    ram_cell[   17500] = 32'hc6889366;
    ram_cell[   17501] = 32'h45b984fc;
    ram_cell[   17502] = 32'h74a914cd;
    ram_cell[   17503] = 32'hc71da6b3;
    ram_cell[   17504] = 32'h7bf92689;
    ram_cell[   17505] = 32'heac30c92;
    ram_cell[   17506] = 32'h4ca0480d;
    ram_cell[   17507] = 32'h6ed18a2f;
    ram_cell[   17508] = 32'h9ecc5442;
    ram_cell[   17509] = 32'hbb0abe92;
    ram_cell[   17510] = 32'h69b3e37c;
    ram_cell[   17511] = 32'h851f10f8;
    ram_cell[   17512] = 32'h1dedd3e8;
    ram_cell[   17513] = 32'hb67719bd;
    ram_cell[   17514] = 32'h830154d5;
    ram_cell[   17515] = 32'h350ce85e;
    ram_cell[   17516] = 32'h8f14c3b1;
    ram_cell[   17517] = 32'h22461efe;
    ram_cell[   17518] = 32'hba97b2bd;
    ram_cell[   17519] = 32'h4f0d3fe4;
    ram_cell[   17520] = 32'h176b898e;
    ram_cell[   17521] = 32'hd9368b71;
    ram_cell[   17522] = 32'h067c97f6;
    ram_cell[   17523] = 32'ha5f1f529;
    ram_cell[   17524] = 32'h08809c14;
    ram_cell[   17525] = 32'h769f5855;
    ram_cell[   17526] = 32'h8a7ccf38;
    ram_cell[   17527] = 32'h09473df2;
    ram_cell[   17528] = 32'hc3ce3c74;
    ram_cell[   17529] = 32'h8bdc1050;
    ram_cell[   17530] = 32'h7b8f399a;
    ram_cell[   17531] = 32'hd9dd2c5e;
    ram_cell[   17532] = 32'hbfbf4516;
    ram_cell[   17533] = 32'h782b504b;
    ram_cell[   17534] = 32'hf0e2f4c1;
    ram_cell[   17535] = 32'ha5495426;
    ram_cell[   17536] = 32'heaea5e0b;
    ram_cell[   17537] = 32'h45e9d2c4;
    ram_cell[   17538] = 32'h7ebce45f;
    ram_cell[   17539] = 32'h1ae90338;
    ram_cell[   17540] = 32'h27e3f946;
    ram_cell[   17541] = 32'ha38d27e6;
    ram_cell[   17542] = 32'hcea64a04;
    ram_cell[   17543] = 32'ha786e270;
    ram_cell[   17544] = 32'h4b6b2803;
    ram_cell[   17545] = 32'he548b943;
    ram_cell[   17546] = 32'h1a39bb50;
    ram_cell[   17547] = 32'hef2a0d28;
    ram_cell[   17548] = 32'h14061655;
    ram_cell[   17549] = 32'h0e713dcb;
    ram_cell[   17550] = 32'h97120fde;
    ram_cell[   17551] = 32'h32b1bed8;
    ram_cell[   17552] = 32'h4fd03700;
    ram_cell[   17553] = 32'h9566f745;
    ram_cell[   17554] = 32'hb02f0e68;
    ram_cell[   17555] = 32'h644fcf04;
    ram_cell[   17556] = 32'h225265f4;
    ram_cell[   17557] = 32'h1b422c7b;
    ram_cell[   17558] = 32'h33f91c2a;
    ram_cell[   17559] = 32'h12af99b5;
    ram_cell[   17560] = 32'hc535db36;
    ram_cell[   17561] = 32'hfaa8ebde;
    ram_cell[   17562] = 32'h035317bf;
    ram_cell[   17563] = 32'h0e95add8;
    ram_cell[   17564] = 32'h6753968d;
    ram_cell[   17565] = 32'h88f1c896;
    ram_cell[   17566] = 32'h9500d060;
    ram_cell[   17567] = 32'h1bc92595;
    ram_cell[   17568] = 32'h28e29b3e;
    ram_cell[   17569] = 32'h8d0e3378;
    ram_cell[   17570] = 32'h34447090;
    ram_cell[   17571] = 32'h62d4158a;
    ram_cell[   17572] = 32'h38741725;
    ram_cell[   17573] = 32'h7c84c2b5;
    ram_cell[   17574] = 32'hcc591cf9;
    ram_cell[   17575] = 32'h49c92cf4;
    ram_cell[   17576] = 32'h658d6e67;
    ram_cell[   17577] = 32'h13e36654;
    ram_cell[   17578] = 32'hedd88c8e;
    ram_cell[   17579] = 32'hda7b4ca5;
    ram_cell[   17580] = 32'h13677fbf;
    ram_cell[   17581] = 32'hc3728f6e;
    ram_cell[   17582] = 32'ha76dfe31;
    ram_cell[   17583] = 32'h37fa87b9;
    ram_cell[   17584] = 32'hda6b1849;
    ram_cell[   17585] = 32'hb170b25d;
    ram_cell[   17586] = 32'h343c1306;
    ram_cell[   17587] = 32'h990ed7b8;
    ram_cell[   17588] = 32'h2a63e808;
    ram_cell[   17589] = 32'hb8cf3fb3;
    ram_cell[   17590] = 32'hea7fcec6;
    ram_cell[   17591] = 32'h3940c0e1;
    ram_cell[   17592] = 32'h6607affb;
    ram_cell[   17593] = 32'haec32dcc;
    ram_cell[   17594] = 32'h81371246;
    ram_cell[   17595] = 32'hdda07182;
    ram_cell[   17596] = 32'h368e152f;
    ram_cell[   17597] = 32'he1d98343;
    ram_cell[   17598] = 32'h52c5e7ae;
    ram_cell[   17599] = 32'h666e8fed;
    ram_cell[   17600] = 32'h36f6d0c5;
    ram_cell[   17601] = 32'hc06f8d81;
    ram_cell[   17602] = 32'hcb9f0285;
    ram_cell[   17603] = 32'hf02ac89b;
    ram_cell[   17604] = 32'h8d5c507d;
    ram_cell[   17605] = 32'h0cc60808;
    ram_cell[   17606] = 32'h05bdb45f;
    ram_cell[   17607] = 32'h91a90ea9;
    ram_cell[   17608] = 32'ha78f5402;
    ram_cell[   17609] = 32'ha9941b93;
    ram_cell[   17610] = 32'hb94bda72;
    ram_cell[   17611] = 32'hf77312dc;
    ram_cell[   17612] = 32'h79f1d602;
    ram_cell[   17613] = 32'h553f756d;
    ram_cell[   17614] = 32'h309049b4;
    ram_cell[   17615] = 32'hccd8fd5f;
    ram_cell[   17616] = 32'hc04a110a;
    ram_cell[   17617] = 32'h2fd3844b;
    ram_cell[   17618] = 32'h0953f074;
    ram_cell[   17619] = 32'h30056cdd;
    ram_cell[   17620] = 32'h9e9bfbd9;
    ram_cell[   17621] = 32'ha13701a8;
    ram_cell[   17622] = 32'h837f8160;
    ram_cell[   17623] = 32'h302c9792;
    ram_cell[   17624] = 32'h388c7407;
    ram_cell[   17625] = 32'he979814d;
    ram_cell[   17626] = 32'hb4ea4158;
    ram_cell[   17627] = 32'hbb944cab;
    ram_cell[   17628] = 32'hc7e0c521;
    ram_cell[   17629] = 32'h9277d4b4;
    ram_cell[   17630] = 32'ha55426a1;
    ram_cell[   17631] = 32'hd6ded3b0;
    ram_cell[   17632] = 32'h32e2bea7;
    ram_cell[   17633] = 32'hae2a1106;
    ram_cell[   17634] = 32'hee3ef2eb;
    ram_cell[   17635] = 32'hecd1e4ca;
    ram_cell[   17636] = 32'h442e9135;
    ram_cell[   17637] = 32'h596d5183;
    ram_cell[   17638] = 32'hcbec40a5;
    ram_cell[   17639] = 32'h0e405f3a;
    ram_cell[   17640] = 32'h8b63cb6c;
    ram_cell[   17641] = 32'he418a7ef;
    ram_cell[   17642] = 32'h54740827;
    ram_cell[   17643] = 32'h108c32e8;
    ram_cell[   17644] = 32'h1dc342c0;
    ram_cell[   17645] = 32'hd54865d1;
    ram_cell[   17646] = 32'h57d2af38;
    ram_cell[   17647] = 32'h1ab29837;
    ram_cell[   17648] = 32'h344b0d76;
    ram_cell[   17649] = 32'h95fa44ba;
    ram_cell[   17650] = 32'hb99506b7;
    ram_cell[   17651] = 32'h8ce2a231;
    ram_cell[   17652] = 32'h871d4760;
    ram_cell[   17653] = 32'hc7c874a8;
    ram_cell[   17654] = 32'h5b454111;
    ram_cell[   17655] = 32'h7b0eff70;
    ram_cell[   17656] = 32'h6df743d5;
    ram_cell[   17657] = 32'he5f09aec;
    ram_cell[   17658] = 32'h566a55ed;
    ram_cell[   17659] = 32'h135d015f;
    ram_cell[   17660] = 32'h786c68a4;
    ram_cell[   17661] = 32'hd701a750;
    ram_cell[   17662] = 32'h2b2082e2;
    ram_cell[   17663] = 32'ha0d5ca77;
    ram_cell[   17664] = 32'h121cdb05;
    ram_cell[   17665] = 32'h9ef0d68e;
    ram_cell[   17666] = 32'h8c2ffcbb;
    ram_cell[   17667] = 32'hc1bf9ba8;
    ram_cell[   17668] = 32'h13bf3f28;
    ram_cell[   17669] = 32'h29c7b71d;
    ram_cell[   17670] = 32'h1aff7fb6;
    ram_cell[   17671] = 32'hbd8084ac;
    ram_cell[   17672] = 32'h4c7ca8c6;
    ram_cell[   17673] = 32'hb03675f1;
    ram_cell[   17674] = 32'hde0472cc;
    ram_cell[   17675] = 32'haf412997;
    ram_cell[   17676] = 32'h42a51b63;
    ram_cell[   17677] = 32'hfb08d036;
    ram_cell[   17678] = 32'h67006935;
    ram_cell[   17679] = 32'h3488f42d;
    ram_cell[   17680] = 32'h4f6a6205;
    ram_cell[   17681] = 32'hf677d05b;
    ram_cell[   17682] = 32'hd0bdc791;
    ram_cell[   17683] = 32'h37f427c0;
    ram_cell[   17684] = 32'h88d1ff98;
    ram_cell[   17685] = 32'h479e708f;
    ram_cell[   17686] = 32'h1e25bdcd;
    ram_cell[   17687] = 32'h1db5d1ae;
    ram_cell[   17688] = 32'hc125eecf;
    ram_cell[   17689] = 32'h761e4625;
    ram_cell[   17690] = 32'h32013625;
    ram_cell[   17691] = 32'h56a68183;
    ram_cell[   17692] = 32'h43bae53f;
    ram_cell[   17693] = 32'h81e1817c;
    ram_cell[   17694] = 32'hbbf366c1;
    ram_cell[   17695] = 32'hb45f4441;
    ram_cell[   17696] = 32'h7de3db10;
    ram_cell[   17697] = 32'hca7849a3;
    ram_cell[   17698] = 32'h3a7b55fe;
    ram_cell[   17699] = 32'h76231c89;
    ram_cell[   17700] = 32'h4f3def1a;
    ram_cell[   17701] = 32'hc8a72e8c;
    ram_cell[   17702] = 32'hc98e13ce;
    ram_cell[   17703] = 32'hd1139d81;
    ram_cell[   17704] = 32'hf3c8c8e1;
    ram_cell[   17705] = 32'h165c4c31;
    ram_cell[   17706] = 32'hfe2b5620;
    ram_cell[   17707] = 32'hda768b2b;
    ram_cell[   17708] = 32'h3f3199da;
    ram_cell[   17709] = 32'h1b0a8ade;
    ram_cell[   17710] = 32'h87f649e7;
    ram_cell[   17711] = 32'h31523726;
    ram_cell[   17712] = 32'hf377c083;
    ram_cell[   17713] = 32'hb2732b67;
    ram_cell[   17714] = 32'hdfdfba40;
    ram_cell[   17715] = 32'hded1334d;
    ram_cell[   17716] = 32'h3844a18d;
    ram_cell[   17717] = 32'h4d1aeb99;
    ram_cell[   17718] = 32'hd93bd701;
    ram_cell[   17719] = 32'h8cbbad3f;
    ram_cell[   17720] = 32'h1a645880;
    ram_cell[   17721] = 32'h3f552b2c;
    ram_cell[   17722] = 32'h6b40d8aa;
    ram_cell[   17723] = 32'hb534aa3d;
    ram_cell[   17724] = 32'hb9d3341d;
    ram_cell[   17725] = 32'h5ef18525;
    ram_cell[   17726] = 32'h9d6f467b;
    ram_cell[   17727] = 32'hc868ef0c;
    ram_cell[   17728] = 32'hc363848b;
    ram_cell[   17729] = 32'h942a9cde;
    ram_cell[   17730] = 32'h8a512018;
    ram_cell[   17731] = 32'he80c6cc4;
    ram_cell[   17732] = 32'h2b6a6b3e;
    ram_cell[   17733] = 32'hcbd19317;
    ram_cell[   17734] = 32'h5482748e;
    ram_cell[   17735] = 32'h8bfc51c2;
    ram_cell[   17736] = 32'h06daec36;
    ram_cell[   17737] = 32'hba561e55;
    ram_cell[   17738] = 32'h16b3b2ed;
    ram_cell[   17739] = 32'h5d83509b;
    ram_cell[   17740] = 32'hc6de8fb1;
    ram_cell[   17741] = 32'ha1558f41;
    ram_cell[   17742] = 32'he0b0cd0e;
    ram_cell[   17743] = 32'h944ef188;
    ram_cell[   17744] = 32'h5f27b23c;
    ram_cell[   17745] = 32'hb2709dee;
    ram_cell[   17746] = 32'hd4f07a16;
    ram_cell[   17747] = 32'h7e32679b;
    ram_cell[   17748] = 32'h84fbbee6;
    ram_cell[   17749] = 32'h46ee332d;
    ram_cell[   17750] = 32'hb7101a21;
    ram_cell[   17751] = 32'h86ff2bf7;
    ram_cell[   17752] = 32'hdcc413dc;
    ram_cell[   17753] = 32'ha782b49b;
    ram_cell[   17754] = 32'haf1ed67d;
    ram_cell[   17755] = 32'h420a5782;
    ram_cell[   17756] = 32'h631f494c;
    ram_cell[   17757] = 32'hda74d819;
    ram_cell[   17758] = 32'h34bc058c;
    ram_cell[   17759] = 32'h606673f5;
    ram_cell[   17760] = 32'hddfc1cea;
    ram_cell[   17761] = 32'h192a8c91;
    ram_cell[   17762] = 32'h9d56ea01;
    ram_cell[   17763] = 32'h67df2dca;
    ram_cell[   17764] = 32'h98567c43;
    ram_cell[   17765] = 32'h3c94519e;
    ram_cell[   17766] = 32'h83913113;
    ram_cell[   17767] = 32'he3b40d53;
    ram_cell[   17768] = 32'h974fca86;
    ram_cell[   17769] = 32'h5c95c5e6;
    ram_cell[   17770] = 32'h501e27cd;
    ram_cell[   17771] = 32'h0b812021;
    ram_cell[   17772] = 32'hff466e5d;
    ram_cell[   17773] = 32'hf6fd99e0;
    ram_cell[   17774] = 32'h976a4b52;
    ram_cell[   17775] = 32'hd12d01e7;
    ram_cell[   17776] = 32'had499ede;
    ram_cell[   17777] = 32'he0771cbd;
    ram_cell[   17778] = 32'hf37c915d;
    ram_cell[   17779] = 32'h11383b1e;
    ram_cell[   17780] = 32'h5ba70b99;
    ram_cell[   17781] = 32'h1f6b4088;
    ram_cell[   17782] = 32'hb549d6e2;
    ram_cell[   17783] = 32'h27d998f2;
    ram_cell[   17784] = 32'hcf36bd17;
    ram_cell[   17785] = 32'hdb1468a6;
    ram_cell[   17786] = 32'hf94b1e97;
    ram_cell[   17787] = 32'hec404ba3;
    ram_cell[   17788] = 32'hbd8c19f0;
    ram_cell[   17789] = 32'he10c7001;
    ram_cell[   17790] = 32'h0ad495f2;
    ram_cell[   17791] = 32'h9dce2816;
    ram_cell[   17792] = 32'hf87c0181;
    ram_cell[   17793] = 32'hdbe68089;
    ram_cell[   17794] = 32'h222db902;
    ram_cell[   17795] = 32'h83b75f9f;
    ram_cell[   17796] = 32'h5b42a090;
    ram_cell[   17797] = 32'h55fc1112;
    ram_cell[   17798] = 32'hf1559fdf;
    ram_cell[   17799] = 32'hbfdc70ba;
    ram_cell[   17800] = 32'hc751a666;
    ram_cell[   17801] = 32'habfe72b8;
    ram_cell[   17802] = 32'hc3ab5541;
    ram_cell[   17803] = 32'h1776cbc4;
    ram_cell[   17804] = 32'hfb02a6a3;
    ram_cell[   17805] = 32'h05356937;
    ram_cell[   17806] = 32'h2193899c;
    ram_cell[   17807] = 32'hbf3b7b36;
    ram_cell[   17808] = 32'h22779456;
    ram_cell[   17809] = 32'hfbb213de;
    ram_cell[   17810] = 32'had45b0f3;
    ram_cell[   17811] = 32'h318881a9;
    ram_cell[   17812] = 32'h9289abd0;
    ram_cell[   17813] = 32'h2ff894ae;
    ram_cell[   17814] = 32'hc763435f;
    ram_cell[   17815] = 32'hb0f0b092;
    ram_cell[   17816] = 32'h538df1ff;
    ram_cell[   17817] = 32'h8e096524;
    ram_cell[   17818] = 32'h2b613da0;
    ram_cell[   17819] = 32'h3584116c;
    ram_cell[   17820] = 32'h9e8be044;
    ram_cell[   17821] = 32'h5022410e;
    ram_cell[   17822] = 32'h287301a0;
    ram_cell[   17823] = 32'hfe338435;
    ram_cell[   17824] = 32'h294857f2;
    ram_cell[   17825] = 32'h2579d6f5;
    ram_cell[   17826] = 32'h678681d8;
    ram_cell[   17827] = 32'h7bcd5f36;
    ram_cell[   17828] = 32'h35825a9b;
    ram_cell[   17829] = 32'h4252d91d;
    ram_cell[   17830] = 32'h5775e2cd;
    ram_cell[   17831] = 32'h8400f7a3;
    ram_cell[   17832] = 32'hd28ce628;
    ram_cell[   17833] = 32'hcaef5f51;
    ram_cell[   17834] = 32'h97fce1d1;
    ram_cell[   17835] = 32'h4466c54c;
    ram_cell[   17836] = 32'h2a4cfbba;
    ram_cell[   17837] = 32'hf3aaafa5;
    ram_cell[   17838] = 32'haa778636;
    ram_cell[   17839] = 32'ha6076527;
    ram_cell[   17840] = 32'he0f8c74b;
    ram_cell[   17841] = 32'h5fe549a0;
    ram_cell[   17842] = 32'h480ced2e;
    ram_cell[   17843] = 32'hac5a835a;
    ram_cell[   17844] = 32'hf348b043;
    ram_cell[   17845] = 32'hd856c48e;
    ram_cell[   17846] = 32'h448fba8b;
    ram_cell[   17847] = 32'h98a7070c;
    ram_cell[   17848] = 32'hfd184e00;
    ram_cell[   17849] = 32'hcc2b07cf;
    ram_cell[   17850] = 32'h1bebe731;
    ram_cell[   17851] = 32'hd7378a2b;
    ram_cell[   17852] = 32'hf480d000;
    ram_cell[   17853] = 32'h28de1818;
    ram_cell[   17854] = 32'h206ec7bc;
    ram_cell[   17855] = 32'hab50cd1a;
    ram_cell[   17856] = 32'h536b2b94;
    ram_cell[   17857] = 32'h5b0ae31c;
    ram_cell[   17858] = 32'h76cb1e08;
    ram_cell[   17859] = 32'h34d3b148;
    ram_cell[   17860] = 32'h004ef353;
    ram_cell[   17861] = 32'h09111238;
    ram_cell[   17862] = 32'h645451f8;
    ram_cell[   17863] = 32'ha295c294;
    ram_cell[   17864] = 32'ha4ceb1df;
    ram_cell[   17865] = 32'h7c100a29;
    ram_cell[   17866] = 32'h61c4fd21;
    ram_cell[   17867] = 32'h8868d4d3;
    ram_cell[   17868] = 32'h6eec0683;
    ram_cell[   17869] = 32'h46a8ca1e;
    ram_cell[   17870] = 32'h5d63c2be;
    ram_cell[   17871] = 32'h6194847f;
    ram_cell[   17872] = 32'hd98ce70a;
    ram_cell[   17873] = 32'h724592a3;
    ram_cell[   17874] = 32'h52f8d730;
    ram_cell[   17875] = 32'h337885a5;
    ram_cell[   17876] = 32'h0c4d5bf1;
    ram_cell[   17877] = 32'ha3986674;
    ram_cell[   17878] = 32'h3f93a946;
    ram_cell[   17879] = 32'h8e33b375;
    ram_cell[   17880] = 32'h7273ddca;
    ram_cell[   17881] = 32'h91cb2402;
    ram_cell[   17882] = 32'h50305c4e;
    ram_cell[   17883] = 32'h9d08c2b1;
    ram_cell[   17884] = 32'hb8fbbbf7;
    ram_cell[   17885] = 32'h0ab97c5f;
    ram_cell[   17886] = 32'hb2af608e;
    ram_cell[   17887] = 32'h704e5eb5;
    ram_cell[   17888] = 32'hc558fdd1;
    ram_cell[   17889] = 32'h8d2cf664;
    ram_cell[   17890] = 32'hb84c9c1c;
    ram_cell[   17891] = 32'h25b3478b;
    ram_cell[   17892] = 32'h08d82526;
    ram_cell[   17893] = 32'h15a2e5de;
    ram_cell[   17894] = 32'hd67f0f06;
    ram_cell[   17895] = 32'h2500fe7a;
    ram_cell[   17896] = 32'h51fc1dd9;
    ram_cell[   17897] = 32'hd42c4b1c;
    ram_cell[   17898] = 32'hdaa425a8;
    ram_cell[   17899] = 32'hb5d600d4;
    ram_cell[   17900] = 32'h9500f976;
    ram_cell[   17901] = 32'h0a64f868;
    ram_cell[   17902] = 32'h281a3240;
    ram_cell[   17903] = 32'h5b5abb2e;
    ram_cell[   17904] = 32'h1185ceaa;
    ram_cell[   17905] = 32'hd48775c1;
    ram_cell[   17906] = 32'hbc2efe6f;
    ram_cell[   17907] = 32'h5bb6b320;
    ram_cell[   17908] = 32'hbe4e7ff4;
    ram_cell[   17909] = 32'hbbc68a9a;
    ram_cell[   17910] = 32'h8a0d3cbe;
    ram_cell[   17911] = 32'h5a60f312;
    ram_cell[   17912] = 32'hf6ffdf5b;
    ram_cell[   17913] = 32'h683eee4d;
    ram_cell[   17914] = 32'h41d554d8;
    ram_cell[   17915] = 32'h131835d5;
    ram_cell[   17916] = 32'he0554153;
    ram_cell[   17917] = 32'hc22145c6;
    ram_cell[   17918] = 32'hb6f6dfe7;
    ram_cell[   17919] = 32'h328779d5;
    ram_cell[   17920] = 32'h1a336497;
    ram_cell[   17921] = 32'h8f576ffd;
    ram_cell[   17922] = 32'ha093e62c;
    ram_cell[   17923] = 32'h0c1aef40;
    ram_cell[   17924] = 32'hdae9fade;
    ram_cell[   17925] = 32'h29963233;
    ram_cell[   17926] = 32'hfc2631a0;
    ram_cell[   17927] = 32'h837ba046;
    ram_cell[   17928] = 32'hf8851ce7;
    ram_cell[   17929] = 32'h7b33a381;
    ram_cell[   17930] = 32'hd125688f;
    ram_cell[   17931] = 32'hb8565612;
    ram_cell[   17932] = 32'hb0f73956;
    ram_cell[   17933] = 32'h002b8249;
    ram_cell[   17934] = 32'h3668c24a;
    ram_cell[   17935] = 32'hf1d85b67;
    ram_cell[   17936] = 32'h77a02cdb;
    ram_cell[   17937] = 32'h2cc96470;
    ram_cell[   17938] = 32'h2853b8ed;
    ram_cell[   17939] = 32'h331195d6;
    ram_cell[   17940] = 32'hcc9bd0a9;
    ram_cell[   17941] = 32'h2ab0bb86;
    ram_cell[   17942] = 32'heeef71d8;
    ram_cell[   17943] = 32'he3a0d1b7;
    ram_cell[   17944] = 32'ha52f5800;
    ram_cell[   17945] = 32'h5e58c6a9;
    ram_cell[   17946] = 32'h528120be;
    ram_cell[   17947] = 32'h1172aa09;
    ram_cell[   17948] = 32'haa5bc8f5;
    ram_cell[   17949] = 32'hcaf2b109;
    ram_cell[   17950] = 32'ha2661d9e;
    ram_cell[   17951] = 32'h5bdaa739;
    ram_cell[   17952] = 32'h6118614f;
    ram_cell[   17953] = 32'h0b014aef;
    ram_cell[   17954] = 32'h489104ae;
    ram_cell[   17955] = 32'h8c05c39c;
    ram_cell[   17956] = 32'h3a28ee1c;
    ram_cell[   17957] = 32'h4e49f7ee;
    ram_cell[   17958] = 32'hbedab32f;
    ram_cell[   17959] = 32'hedd43c96;
    ram_cell[   17960] = 32'hff59e143;
    ram_cell[   17961] = 32'h17247f2a;
    ram_cell[   17962] = 32'h847a469b;
    ram_cell[   17963] = 32'hc947c8ca;
    ram_cell[   17964] = 32'hb1053f4c;
    ram_cell[   17965] = 32'he5f5b030;
    ram_cell[   17966] = 32'hcd67f919;
    ram_cell[   17967] = 32'hdd094624;
    ram_cell[   17968] = 32'h9e627c69;
    ram_cell[   17969] = 32'hb01ee1af;
    ram_cell[   17970] = 32'h29611f80;
    ram_cell[   17971] = 32'hccfa2c9f;
    ram_cell[   17972] = 32'hf0e704d2;
    ram_cell[   17973] = 32'hb21a829f;
    ram_cell[   17974] = 32'h3c7536fb;
    ram_cell[   17975] = 32'h4c767e1e;
    ram_cell[   17976] = 32'hee0594e8;
    ram_cell[   17977] = 32'hbf73bf4a;
    ram_cell[   17978] = 32'hdfaeeb5e;
    ram_cell[   17979] = 32'h74d79f22;
    ram_cell[   17980] = 32'h162ee949;
    ram_cell[   17981] = 32'hc53e7461;
    ram_cell[   17982] = 32'hc973b9de;
    ram_cell[   17983] = 32'h87cca0c1;
    ram_cell[   17984] = 32'he74866c3;
    ram_cell[   17985] = 32'hdd61d22f;
    ram_cell[   17986] = 32'h9cb217b4;
    ram_cell[   17987] = 32'ha5c3b477;
    ram_cell[   17988] = 32'h3a796b3e;
    ram_cell[   17989] = 32'ha3187caa;
    ram_cell[   17990] = 32'h9b136e34;
    ram_cell[   17991] = 32'h8f7ff267;
    ram_cell[   17992] = 32'h62141c22;
    ram_cell[   17993] = 32'hbe1f911f;
    ram_cell[   17994] = 32'h6cd58b35;
    ram_cell[   17995] = 32'h3248e2c4;
    ram_cell[   17996] = 32'hc0b7d22e;
    ram_cell[   17997] = 32'hf3625018;
    ram_cell[   17998] = 32'h55cc3d97;
    ram_cell[   17999] = 32'h813fa129;
    ram_cell[   18000] = 32'h387724ad;
    ram_cell[   18001] = 32'h6b7c9454;
    ram_cell[   18002] = 32'h192cb23d;
    ram_cell[   18003] = 32'h6585ac38;
    ram_cell[   18004] = 32'h4a4f6860;
    ram_cell[   18005] = 32'h0f0fe7f2;
    ram_cell[   18006] = 32'hfc1472bc;
    ram_cell[   18007] = 32'h6fddddd1;
    ram_cell[   18008] = 32'h436f5dbe;
    ram_cell[   18009] = 32'h71bf4c50;
    ram_cell[   18010] = 32'h0e8d1b18;
    ram_cell[   18011] = 32'h399a7f13;
    ram_cell[   18012] = 32'hfac55290;
    ram_cell[   18013] = 32'h92b62d72;
    ram_cell[   18014] = 32'hf70940b3;
    ram_cell[   18015] = 32'h3c6a9253;
    ram_cell[   18016] = 32'h785ce641;
    ram_cell[   18017] = 32'h74216d30;
    ram_cell[   18018] = 32'h4c72b56e;
    ram_cell[   18019] = 32'hb9608cfc;
    ram_cell[   18020] = 32'h244dc912;
    ram_cell[   18021] = 32'h2dcc6f33;
    ram_cell[   18022] = 32'h9b8b8d4f;
    ram_cell[   18023] = 32'he5898eda;
    ram_cell[   18024] = 32'hfda8a993;
    ram_cell[   18025] = 32'hc441becb;
    ram_cell[   18026] = 32'h26ee2a3e;
    ram_cell[   18027] = 32'h30c6aa44;
    ram_cell[   18028] = 32'h1abad0a5;
    ram_cell[   18029] = 32'h3f097ee1;
    ram_cell[   18030] = 32'h9126a7d6;
    ram_cell[   18031] = 32'h500f3689;
    ram_cell[   18032] = 32'h1533b9d4;
    ram_cell[   18033] = 32'h679a34e5;
    ram_cell[   18034] = 32'h72d01e20;
    ram_cell[   18035] = 32'hcc4797e1;
    ram_cell[   18036] = 32'h0e9529f0;
    ram_cell[   18037] = 32'h8e840970;
    ram_cell[   18038] = 32'h8d52040e;
    ram_cell[   18039] = 32'h5691794e;
    ram_cell[   18040] = 32'h2a4a7444;
    ram_cell[   18041] = 32'hb79800de;
    ram_cell[   18042] = 32'hc7191cd0;
    ram_cell[   18043] = 32'hf2e184c4;
    ram_cell[   18044] = 32'h41a9b862;
    ram_cell[   18045] = 32'h0eff1cb3;
    ram_cell[   18046] = 32'h78034a27;
    ram_cell[   18047] = 32'hc1d54ebd;
    ram_cell[   18048] = 32'hd414828c;
    ram_cell[   18049] = 32'h4cfbd3b1;
    ram_cell[   18050] = 32'hcdc526ea;
    ram_cell[   18051] = 32'h8fe9d7cb;
    ram_cell[   18052] = 32'h9851a8b7;
    ram_cell[   18053] = 32'h2a4e653b;
    ram_cell[   18054] = 32'hb95b3f48;
    ram_cell[   18055] = 32'hfdb7b2d2;
    ram_cell[   18056] = 32'hb9f71155;
    ram_cell[   18057] = 32'h607e25b0;
    ram_cell[   18058] = 32'hc23e371b;
    ram_cell[   18059] = 32'h7c724476;
    ram_cell[   18060] = 32'h086167e4;
    ram_cell[   18061] = 32'hb8969326;
    ram_cell[   18062] = 32'hc64a4237;
    ram_cell[   18063] = 32'h58e223e4;
    ram_cell[   18064] = 32'h485f3c5a;
    ram_cell[   18065] = 32'h29f87c87;
    ram_cell[   18066] = 32'hb2a7f903;
    ram_cell[   18067] = 32'h4d51d2b2;
    ram_cell[   18068] = 32'hd3cb4094;
    ram_cell[   18069] = 32'h48ef43ec;
    ram_cell[   18070] = 32'h4a372c84;
    ram_cell[   18071] = 32'h8b37f6f4;
    ram_cell[   18072] = 32'h2988b05d;
    ram_cell[   18073] = 32'h1ac40cf5;
    ram_cell[   18074] = 32'hb1e6fb6c;
    ram_cell[   18075] = 32'h9a359a77;
    ram_cell[   18076] = 32'habfaa827;
    ram_cell[   18077] = 32'hfa33f126;
    ram_cell[   18078] = 32'hdeeae648;
    ram_cell[   18079] = 32'hd5b367a5;
    ram_cell[   18080] = 32'h3983e219;
    ram_cell[   18081] = 32'h9a394a9a;
    ram_cell[   18082] = 32'h1b24ea46;
    ram_cell[   18083] = 32'h4f6ed57f;
    ram_cell[   18084] = 32'h44d5fb09;
    ram_cell[   18085] = 32'h1a451c53;
    ram_cell[   18086] = 32'h750ad880;
    ram_cell[   18087] = 32'hb1b7c157;
    ram_cell[   18088] = 32'ha1984537;
    ram_cell[   18089] = 32'hc7afa171;
    ram_cell[   18090] = 32'h8da2c1c3;
    ram_cell[   18091] = 32'h4453fa44;
    ram_cell[   18092] = 32'hfa476600;
    ram_cell[   18093] = 32'h3e21b557;
    ram_cell[   18094] = 32'h83940b15;
    ram_cell[   18095] = 32'h5bbbc780;
    ram_cell[   18096] = 32'h9f7a4d5e;
    ram_cell[   18097] = 32'hc50fab44;
    ram_cell[   18098] = 32'h1eac1653;
    ram_cell[   18099] = 32'h70f0881a;
    ram_cell[   18100] = 32'h769badbc;
    ram_cell[   18101] = 32'h9213cefb;
    ram_cell[   18102] = 32'h99834c25;
    ram_cell[   18103] = 32'h3eac8b1c;
    ram_cell[   18104] = 32'h42b58f19;
    ram_cell[   18105] = 32'hf2853bcd;
    ram_cell[   18106] = 32'h8bf0e153;
    ram_cell[   18107] = 32'hce38fcc6;
    ram_cell[   18108] = 32'heb4c84f3;
    ram_cell[   18109] = 32'hd4406fc0;
    ram_cell[   18110] = 32'h8880fdf1;
    ram_cell[   18111] = 32'h4a9333d5;
    ram_cell[   18112] = 32'ha003699b;
    ram_cell[   18113] = 32'h1cb169f0;
    ram_cell[   18114] = 32'h52a1d7cb;
    ram_cell[   18115] = 32'hbc7250fd;
    ram_cell[   18116] = 32'h5d171ece;
    ram_cell[   18117] = 32'h2c31ba98;
    ram_cell[   18118] = 32'hcee1f533;
    ram_cell[   18119] = 32'he1bcdbcb;
    ram_cell[   18120] = 32'h10702a62;
    ram_cell[   18121] = 32'h34398796;
    ram_cell[   18122] = 32'ha6a894c3;
    ram_cell[   18123] = 32'h2c63f18d;
    ram_cell[   18124] = 32'h30f5ef68;
    ram_cell[   18125] = 32'h8dbf41f1;
    ram_cell[   18126] = 32'h84adb49c;
    ram_cell[   18127] = 32'h2b517ac3;
    ram_cell[   18128] = 32'hc19f7124;
    ram_cell[   18129] = 32'h2d4af6e1;
    ram_cell[   18130] = 32'hd4f44d11;
    ram_cell[   18131] = 32'h49ba6722;
    ram_cell[   18132] = 32'hf6326a32;
    ram_cell[   18133] = 32'ha3369871;
    ram_cell[   18134] = 32'h13c64974;
    ram_cell[   18135] = 32'hab69a731;
    ram_cell[   18136] = 32'h4ba3a59b;
    ram_cell[   18137] = 32'h9b884475;
    ram_cell[   18138] = 32'hec96505d;
    ram_cell[   18139] = 32'ha03bdae9;
    ram_cell[   18140] = 32'h57e28a34;
    ram_cell[   18141] = 32'hd210a703;
    ram_cell[   18142] = 32'h69352bb0;
    ram_cell[   18143] = 32'h17284bbb;
    ram_cell[   18144] = 32'he36414ea;
    ram_cell[   18145] = 32'h0bb5b684;
    ram_cell[   18146] = 32'h43c2824b;
    ram_cell[   18147] = 32'h4ed16298;
    ram_cell[   18148] = 32'h15adb87b;
    ram_cell[   18149] = 32'haa392525;
    ram_cell[   18150] = 32'h7dca80b3;
    ram_cell[   18151] = 32'hc3741057;
    ram_cell[   18152] = 32'h300290bb;
    ram_cell[   18153] = 32'h8c9874d3;
    ram_cell[   18154] = 32'h66164752;
    ram_cell[   18155] = 32'h5ff20ded;
    ram_cell[   18156] = 32'h3d1c1755;
    ram_cell[   18157] = 32'h12eeed3a;
    ram_cell[   18158] = 32'h22b1e463;
    ram_cell[   18159] = 32'h32544b28;
    ram_cell[   18160] = 32'hdb54667c;
    ram_cell[   18161] = 32'h908794ce;
    ram_cell[   18162] = 32'hc94fd868;
    ram_cell[   18163] = 32'h993e41af;
    ram_cell[   18164] = 32'h38dadadd;
    ram_cell[   18165] = 32'ha5f89e30;
    ram_cell[   18166] = 32'h9ae42b5f;
    ram_cell[   18167] = 32'hd5d318dc;
    ram_cell[   18168] = 32'h0b91c809;
    ram_cell[   18169] = 32'h88220504;
    ram_cell[   18170] = 32'h4942d3da;
    ram_cell[   18171] = 32'hd2e8de50;
    ram_cell[   18172] = 32'h5bcb371d;
    ram_cell[   18173] = 32'ha158188b;
    ram_cell[   18174] = 32'hb3eec912;
    ram_cell[   18175] = 32'hddbeb86e;
    ram_cell[   18176] = 32'h575b9e21;
    ram_cell[   18177] = 32'h59c97c04;
    ram_cell[   18178] = 32'h0496cb90;
    ram_cell[   18179] = 32'h705be613;
    ram_cell[   18180] = 32'he5df3bb5;
    ram_cell[   18181] = 32'h357f804c;
    ram_cell[   18182] = 32'h8f1c4011;
    ram_cell[   18183] = 32'h73d9ffa6;
    ram_cell[   18184] = 32'h8ceb36e8;
    ram_cell[   18185] = 32'h8525ffcd;
    ram_cell[   18186] = 32'h543f044c;
    ram_cell[   18187] = 32'hed3aa072;
    ram_cell[   18188] = 32'hc019ed78;
    ram_cell[   18189] = 32'h6fa9b1b6;
    ram_cell[   18190] = 32'hecea86a4;
    ram_cell[   18191] = 32'h1d7e50f5;
    ram_cell[   18192] = 32'h2fca9476;
    ram_cell[   18193] = 32'h00cd47c5;
    ram_cell[   18194] = 32'h9a35f6ab;
    ram_cell[   18195] = 32'h35d4339b;
    ram_cell[   18196] = 32'h93076f9d;
    ram_cell[   18197] = 32'hcd679735;
    ram_cell[   18198] = 32'h0d6d0420;
    ram_cell[   18199] = 32'h35bc9a8c;
    ram_cell[   18200] = 32'hde1f148b;
    ram_cell[   18201] = 32'h03a71a20;
    ram_cell[   18202] = 32'h48e471bf;
    ram_cell[   18203] = 32'h2e05df03;
    ram_cell[   18204] = 32'h4e5288c4;
    ram_cell[   18205] = 32'h7606c2eb;
    ram_cell[   18206] = 32'h40068f88;
    ram_cell[   18207] = 32'h4aec4cd1;
    ram_cell[   18208] = 32'hbfed4606;
    ram_cell[   18209] = 32'h50bf065e;
    ram_cell[   18210] = 32'h0e0989be;
    ram_cell[   18211] = 32'hd03b1f16;
    ram_cell[   18212] = 32'h3a19d50c;
    ram_cell[   18213] = 32'he3af29f4;
    ram_cell[   18214] = 32'h380ac810;
    ram_cell[   18215] = 32'hdfbcc550;
    ram_cell[   18216] = 32'h7637d6a4;
    ram_cell[   18217] = 32'h1f2a8671;
    ram_cell[   18218] = 32'h1acd7582;
    ram_cell[   18219] = 32'h74da275b;
    ram_cell[   18220] = 32'h97bf930c;
    ram_cell[   18221] = 32'h6efe96b8;
    ram_cell[   18222] = 32'h7af2cab0;
    ram_cell[   18223] = 32'h77d0436d;
    ram_cell[   18224] = 32'hb2ccdfab;
    ram_cell[   18225] = 32'h80ac6eb8;
    ram_cell[   18226] = 32'h6481080a;
    ram_cell[   18227] = 32'h38b5671f;
    ram_cell[   18228] = 32'h47f51cea;
    ram_cell[   18229] = 32'ha1d7cba6;
    ram_cell[   18230] = 32'h5574e32e;
    ram_cell[   18231] = 32'h602cfa5a;
    ram_cell[   18232] = 32'ha36f2da1;
    ram_cell[   18233] = 32'hb86c37eb;
    ram_cell[   18234] = 32'he22b1780;
    ram_cell[   18235] = 32'h3a3c9a0a;
    ram_cell[   18236] = 32'h3cac6bd1;
    ram_cell[   18237] = 32'hfd9edd87;
    ram_cell[   18238] = 32'hb07be073;
    ram_cell[   18239] = 32'ha9f8edda;
    ram_cell[   18240] = 32'hcd1253df;
    ram_cell[   18241] = 32'h8ebe2ba6;
    ram_cell[   18242] = 32'hc1d7131f;
    ram_cell[   18243] = 32'h2b54cedf;
    ram_cell[   18244] = 32'hc555d63d;
    ram_cell[   18245] = 32'h7047bae2;
    ram_cell[   18246] = 32'hfa0ab101;
    ram_cell[   18247] = 32'h947ad08e;
    ram_cell[   18248] = 32'ha129881b;
    ram_cell[   18249] = 32'hef414b00;
    ram_cell[   18250] = 32'h260f6604;
    ram_cell[   18251] = 32'h81695026;
    ram_cell[   18252] = 32'h8d941ba7;
    ram_cell[   18253] = 32'hd19ad197;
    ram_cell[   18254] = 32'hfdb105ec;
    ram_cell[   18255] = 32'h0a0dab6c;
    ram_cell[   18256] = 32'hd03398c0;
    ram_cell[   18257] = 32'h1734a16c;
    ram_cell[   18258] = 32'hfd818fff;
    ram_cell[   18259] = 32'h44d15582;
    ram_cell[   18260] = 32'h83106450;
    ram_cell[   18261] = 32'h6ec8c563;
    ram_cell[   18262] = 32'h075489ac;
    ram_cell[   18263] = 32'h7e354b01;
    ram_cell[   18264] = 32'h10862299;
    ram_cell[   18265] = 32'h7aefaebe;
    ram_cell[   18266] = 32'h19471c09;
    ram_cell[   18267] = 32'h3e79ebd9;
    ram_cell[   18268] = 32'ha84f03f8;
    ram_cell[   18269] = 32'h4e55a92f;
    ram_cell[   18270] = 32'h262381cc;
    ram_cell[   18271] = 32'h9c600b9f;
    ram_cell[   18272] = 32'h7d565fd2;
    ram_cell[   18273] = 32'hf51b2f5d;
    ram_cell[   18274] = 32'h1bfedc26;
    ram_cell[   18275] = 32'h0e1869d5;
    ram_cell[   18276] = 32'h647f865d;
    ram_cell[   18277] = 32'h20cb29e4;
    ram_cell[   18278] = 32'h98ace247;
    ram_cell[   18279] = 32'h79a3657a;
    ram_cell[   18280] = 32'h0eb5324f;
    ram_cell[   18281] = 32'h201d4207;
    ram_cell[   18282] = 32'h5137035a;
    ram_cell[   18283] = 32'h31b0dca0;
    ram_cell[   18284] = 32'h37f4c05d;
    ram_cell[   18285] = 32'hcebe3888;
    ram_cell[   18286] = 32'hf68e1fa9;
    ram_cell[   18287] = 32'h72c3f71d;
    ram_cell[   18288] = 32'ha00ae75e;
    ram_cell[   18289] = 32'h2fbd849c;
    ram_cell[   18290] = 32'h8c6c2e9a;
    ram_cell[   18291] = 32'h60cbec27;
    ram_cell[   18292] = 32'h5fbfc707;
    ram_cell[   18293] = 32'h9042aa76;
    ram_cell[   18294] = 32'h1ecc1a85;
    ram_cell[   18295] = 32'hcede846e;
    ram_cell[   18296] = 32'hccb79dce;
    ram_cell[   18297] = 32'ha1cf61cb;
    ram_cell[   18298] = 32'hbc758e80;
    ram_cell[   18299] = 32'h2d237bb4;
    ram_cell[   18300] = 32'h17b832af;
    ram_cell[   18301] = 32'ha97ecdcb;
    ram_cell[   18302] = 32'h4b047d02;
    ram_cell[   18303] = 32'hccf25b92;
    ram_cell[   18304] = 32'he5ce1c3f;
    ram_cell[   18305] = 32'h0f8bcf0b;
    ram_cell[   18306] = 32'h20296361;
    ram_cell[   18307] = 32'h30970496;
    ram_cell[   18308] = 32'h356589f5;
    ram_cell[   18309] = 32'heb1927e0;
    ram_cell[   18310] = 32'h8e39cc8e;
    ram_cell[   18311] = 32'hea620e95;
    ram_cell[   18312] = 32'h4a1c3481;
    ram_cell[   18313] = 32'ha7b0fa41;
    ram_cell[   18314] = 32'he7f8581c;
    ram_cell[   18315] = 32'h8b54abd3;
    ram_cell[   18316] = 32'h19c3bc90;
    ram_cell[   18317] = 32'hf5dae3d8;
    ram_cell[   18318] = 32'h77a15dee;
    ram_cell[   18319] = 32'hc2f1a676;
    ram_cell[   18320] = 32'h505574ad;
    ram_cell[   18321] = 32'he8132dc8;
    ram_cell[   18322] = 32'h53f9f0ed;
    ram_cell[   18323] = 32'h4ccb885b;
    ram_cell[   18324] = 32'h9e21ae66;
    ram_cell[   18325] = 32'ha3b29835;
    ram_cell[   18326] = 32'h2eb06d35;
    ram_cell[   18327] = 32'h36dfa99f;
    ram_cell[   18328] = 32'h7a7a89dd;
    ram_cell[   18329] = 32'hee842470;
    ram_cell[   18330] = 32'h8c8c5c36;
    ram_cell[   18331] = 32'h8b057500;
    ram_cell[   18332] = 32'hd55128f3;
    ram_cell[   18333] = 32'h51648954;
    ram_cell[   18334] = 32'he2fae186;
    ram_cell[   18335] = 32'h6c4881de;
    ram_cell[   18336] = 32'h30a13372;
    ram_cell[   18337] = 32'h241c464d;
    ram_cell[   18338] = 32'hfaf10c3f;
    ram_cell[   18339] = 32'hc5c9ef7c;
    ram_cell[   18340] = 32'h8343505e;
    ram_cell[   18341] = 32'hd9972595;
    ram_cell[   18342] = 32'h724d3725;
    ram_cell[   18343] = 32'h0514e562;
    ram_cell[   18344] = 32'h349b9017;
    ram_cell[   18345] = 32'h807ff131;
    ram_cell[   18346] = 32'he8cda6e9;
    ram_cell[   18347] = 32'h7344e988;
    ram_cell[   18348] = 32'h77ba2ca4;
    ram_cell[   18349] = 32'h12be34f7;
    ram_cell[   18350] = 32'he841ffbb;
    ram_cell[   18351] = 32'h12d40d4b;
    ram_cell[   18352] = 32'h32e37423;
    ram_cell[   18353] = 32'hdca37ffc;
    ram_cell[   18354] = 32'h663c8102;
    ram_cell[   18355] = 32'hdbe3104d;
    ram_cell[   18356] = 32'hafea2a28;
    ram_cell[   18357] = 32'hb65d9594;
    ram_cell[   18358] = 32'h3f60fe72;
    ram_cell[   18359] = 32'hde46efab;
    ram_cell[   18360] = 32'hdd49ea24;
    ram_cell[   18361] = 32'h5394790e;
    ram_cell[   18362] = 32'h46476de9;
    ram_cell[   18363] = 32'h37437670;
    ram_cell[   18364] = 32'h902cf107;
    ram_cell[   18365] = 32'h620f0db1;
    ram_cell[   18366] = 32'he4a6af12;
    ram_cell[   18367] = 32'haebc98fb;
    ram_cell[   18368] = 32'h6b6cead7;
    ram_cell[   18369] = 32'h4cae1cc9;
    ram_cell[   18370] = 32'h193f00f1;
    ram_cell[   18371] = 32'hc0eca39e;
    ram_cell[   18372] = 32'h54ce860b;
    ram_cell[   18373] = 32'h9a9b6b79;
    ram_cell[   18374] = 32'h9ea688c7;
    ram_cell[   18375] = 32'h9e26cde7;
    ram_cell[   18376] = 32'h8816796c;
    ram_cell[   18377] = 32'h2dfc9fc9;
    ram_cell[   18378] = 32'h9541a2c6;
    ram_cell[   18379] = 32'h2aa22dc1;
    ram_cell[   18380] = 32'hec86e982;
    ram_cell[   18381] = 32'h0390b945;
    ram_cell[   18382] = 32'h7d07b5e3;
    ram_cell[   18383] = 32'h93f0c5c3;
    ram_cell[   18384] = 32'h5b58fcdc;
    ram_cell[   18385] = 32'h3c076ce4;
    ram_cell[   18386] = 32'ha01896ec;
    ram_cell[   18387] = 32'hf540ec85;
    ram_cell[   18388] = 32'hb21b2fcc;
    ram_cell[   18389] = 32'h3e0d02ba;
    ram_cell[   18390] = 32'hf408c20e;
    ram_cell[   18391] = 32'hdd5149ba;
    ram_cell[   18392] = 32'h8dee997b;
    ram_cell[   18393] = 32'h10241c10;
    ram_cell[   18394] = 32'h33be24db;
    ram_cell[   18395] = 32'he0b419d2;
    ram_cell[   18396] = 32'h5ddddb29;
    ram_cell[   18397] = 32'hac09f37e;
    ram_cell[   18398] = 32'hd1168c9b;
    ram_cell[   18399] = 32'h035e6063;
    ram_cell[   18400] = 32'h33033eb5;
    ram_cell[   18401] = 32'hdcbc941d;
    ram_cell[   18402] = 32'hb896b5ac;
    ram_cell[   18403] = 32'h298ad604;
    ram_cell[   18404] = 32'ha8b61c6a;
    ram_cell[   18405] = 32'he4df0c0c;
    ram_cell[   18406] = 32'h7649c30a;
    ram_cell[   18407] = 32'ha162b7b1;
    ram_cell[   18408] = 32'h90fb793c;
    ram_cell[   18409] = 32'hba123944;
    ram_cell[   18410] = 32'h360ac7fa;
    ram_cell[   18411] = 32'h1b743b50;
    ram_cell[   18412] = 32'hd948d73e;
    ram_cell[   18413] = 32'h2ea95a2b;
    ram_cell[   18414] = 32'hc78f0dca;
    ram_cell[   18415] = 32'h84d2dfe5;
    ram_cell[   18416] = 32'h6b15d230;
    ram_cell[   18417] = 32'hd146372a;
    ram_cell[   18418] = 32'hc2dd00ac;
    ram_cell[   18419] = 32'hc8c1f153;
    ram_cell[   18420] = 32'h9515dc84;
    ram_cell[   18421] = 32'hbbdd4e8b;
    ram_cell[   18422] = 32'hc6b21927;
    ram_cell[   18423] = 32'h1a78d355;
    ram_cell[   18424] = 32'h46c0d49a;
    ram_cell[   18425] = 32'h2d8eab27;
    ram_cell[   18426] = 32'h563baf94;
    ram_cell[   18427] = 32'h34c35014;
    ram_cell[   18428] = 32'h056fefe7;
    ram_cell[   18429] = 32'h5fe7bb49;
    ram_cell[   18430] = 32'hadb98c9b;
    ram_cell[   18431] = 32'h2d540036;
    ram_cell[   18432] = 32'hb9185131;
    ram_cell[   18433] = 32'hbb064209;
    ram_cell[   18434] = 32'h9ac82241;
    ram_cell[   18435] = 32'h0c0206bd;
    ram_cell[   18436] = 32'hd90eb0ee;
    ram_cell[   18437] = 32'he23c614a;
    ram_cell[   18438] = 32'h59a42875;
    ram_cell[   18439] = 32'h848f0543;
    ram_cell[   18440] = 32'h73db2535;
    ram_cell[   18441] = 32'hb6d0233b;
    ram_cell[   18442] = 32'ha70d6837;
    ram_cell[   18443] = 32'ha5e5463e;
    ram_cell[   18444] = 32'hc63a11a2;
    ram_cell[   18445] = 32'h546a65ae;
    ram_cell[   18446] = 32'h93447503;
    ram_cell[   18447] = 32'h14daae26;
    ram_cell[   18448] = 32'hbc9dde71;
    ram_cell[   18449] = 32'hd9305763;
    ram_cell[   18450] = 32'hd35d9422;
    ram_cell[   18451] = 32'h8636db9c;
    ram_cell[   18452] = 32'h0df2b588;
    ram_cell[   18453] = 32'h097b483a;
    ram_cell[   18454] = 32'haf7cdb9e;
    ram_cell[   18455] = 32'ha219947b;
    ram_cell[   18456] = 32'h35a8b6ee;
    ram_cell[   18457] = 32'h791d3e40;
    ram_cell[   18458] = 32'hfb6214de;
    ram_cell[   18459] = 32'h85c33313;
    ram_cell[   18460] = 32'hae13bf42;
    ram_cell[   18461] = 32'h8b9c9676;
    ram_cell[   18462] = 32'ha37dbec9;
    ram_cell[   18463] = 32'h4f1ad947;
    ram_cell[   18464] = 32'hae9bbdd6;
    ram_cell[   18465] = 32'hcb92f6c5;
    ram_cell[   18466] = 32'h073c317b;
    ram_cell[   18467] = 32'h81b620f5;
    ram_cell[   18468] = 32'h7aaecb9b;
    ram_cell[   18469] = 32'ha57d16a9;
    ram_cell[   18470] = 32'h1b1994a2;
    ram_cell[   18471] = 32'h2416274c;
    ram_cell[   18472] = 32'h8457a66f;
    ram_cell[   18473] = 32'h2cbad613;
    ram_cell[   18474] = 32'h9e6f6be7;
    ram_cell[   18475] = 32'h17b65e95;
    ram_cell[   18476] = 32'hb65112ed;
    ram_cell[   18477] = 32'heefe0623;
    ram_cell[   18478] = 32'hece9b4c7;
    ram_cell[   18479] = 32'h367a14c1;
    ram_cell[   18480] = 32'hf8f1fc4e;
    ram_cell[   18481] = 32'h068aab8b;
    ram_cell[   18482] = 32'hfe108fd6;
    ram_cell[   18483] = 32'h2a5b9d5d;
    ram_cell[   18484] = 32'h6058d69d;
    ram_cell[   18485] = 32'h79ad4ae1;
    ram_cell[   18486] = 32'h1924674c;
    ram_cell[   18487] = 32'h74399282;
    ram_cell[   18488] = 32'h9a7aa53a;
    ram_cell[   18489] = 32'hb6ac2f93;
    ram_cell[   18490] = 32'h77689762;
    ram_cell[   18491] = 32'h36be1711;
    ram_cell[   18492] = 32'h009ef02f;
    ram_cell[   18493] = 32'hcb8cf19f;
    ram_cell[   18494] = 32'h75a9b512;
    ram_cell[   18495] = 32'h051bbf09;
    ram_cell[   18496] = 32'h3f9fea0b;
    ram_cell[   18497] = 32'h56508ad9;
    ram_cell[   18498] = 32'h23e728da;
    ram_cell[   18499] = 32'h5cf1b2ac;
    ram_cell[   18500] = 32'h49261c89;
    ram_cell[   18501] = 32'h06ea9d01;
    ram_cell[   18502] = 32'hbbd0fbee;
    ram_cell[   18503] = 32'h8bd59bb2;
    ram_cell[   18504] = 32'h6fd73db7;
    ram_cell[   18505] = 32'hd7aea74c;
    ram_cell[   18506] = 32'h6bf12f1f;
    ram_cell[   18507] = 32'h91b291f7;
    ram_cell[   18508] = 32'heaac7880;
    ram_cell[   18509] = 32'h968860db;
    ram_cell[   18510] = 32'heecb8e5d;
    ram_cell[   18511] = 32'h9b22ad4b;
    ram_cell[   18512] = 32'hac75a5fa;
    ram_cell[   18513] = 32'h7f87fc0c;
    ram_cell[   18514] = 32'h176814ab;
    ram_cell[   18515] = 32'ha9775ea2;
    ram_cell[   18516] = 32'h0fc65e71;
    ram_cell[   18517] = 32'h4ca056eb;
    ram_cell[   18518] = 32'h52605c40;
    ram_cell[   18519] = 32'haeef859d;
    ram_cell[   18520] = 32'hfe767950;
    ram_cell[   18521] = 32'h878fffff;
    ram_cell[   18522] = 32'h159db583;
    ram_cell[   18523] = 32'h3413f41f;
    ram_cell[   18524] = 32'h3102b33c;
    ram_cell[   18525] = 32'h9c554450;
    ram_cell[   18526] = 32'h12e9dd0c;
    ram_cell[   18527] = 32'h4184e678;
    ram_cell[   18528] = 32'h9b219861;
    ram_cell[   18529] = 32'hfce8193e;
    ram_cell[   18530] = 32'h28035796;
    ram_cell[   18531] = 32'ha8345a8a;
    ram_cell[   18532] = 32'haf1e399b;
    ram_cell[   18533] = 32'hc7873f11;
    ram_cell[   18534] = 32'h5c2f2ac1;
    ram_cell[   18535] = 32'h15ad0340;
    ram_cell[   18536] = 32'ha621bb81;
    ram_cell[   18537] = 32'h0ba03983;
    ram_cell[   18538] = 32'h869cc43c;
    ram_cell[   18539] = 32'h1c2f28dc;
    ram_cell[   18540] = 32'h949c884e;
    ram_cell[   18541] = 32'h2d506c4f;
    ram_cell[   18542] = 32'h3e78d763;
    ram_cell[   18543] = 32'h67a9f9a2;
    ram_cell[   18544] = 32'hd666562e;
    ram_cell[   18545] = 32'h6a9fe013;
    ram_cell[   18546] = 32'h76ff9afa;
    ram_cell[   18547] = 32'h36d3beb6;
    ram_cell[   18548] = 32'h18a0bc9b;
    ram_cell[   18549] = 32'h044e57f4;
    ram_cell[   18550] = 32'hf8a83351;
    ram_cell[   18551] = 32'h1a95405d;
    ram_cell[   18552] = 32'h8128f347;
    ram_cell[   18553] = 32'h3b8c43ce;
    ram_cell[   18554] = 32'hfd9c3fa1;
    ram_cell[   18555] = 32'h18c65e55;
    ram_cell[   18556] = 32'h5c4fb48a;
    ram_cell[   18557] = 32'he9a60d9c;
    ram_cell[   18558] = 32'hb0d8fe8d;
    ram_cell[   18559] = 32'hce842c03;
    ram_cell[   18560] = 32'h6c7562b0;
    ram_cell[   18561] = 32'h455dd2a1;
    ram_cell[   18562] = 32'h2a229015;
    ram_cell[   18563] = 32'h38d60359;
    ram_cell[   18564] = 32'h7c7704c4;
    ram_cell[   18565] = 32'hf9e90061;
    ram_cell[   18566] = 32'hbcacf9f4;
    ram_cell[   18567] = 32'h0c40978d;
    ram_cell[   18568] = 32'h150ac40a;
    ram_cell[   18569] = 32'h63ae1501;
    ram_cell[   18570] = 32'h2669a528;
    ram_cell[   18571] = 32'h92d6f941;
    ram_cell[   18572] = 32'h2c6b914c;
    ram_cell[   18573] = 32'h5f834494;
    ram_cell[   18574] = 32'h1fec82db;
    ram_cell[   18575] = 32'hf579b9c0;
    ram_cell[   18576] = 32'h9a28565a;
    ram_cell[   18577] = 32'hd9fccf65;
    ram_cell[   18578] = 32'h8f749d41;
    ram_cell[   18579] = 32'h3bf72309;
    ram_cell[   18580] = 32'h1ad47596;
    ram_cell[   18581] = 32'he399fa90;
    ram_cell[   18582] = 32'h024258f7;
    ram_cell[   18583] = 32'h2e8ef90a;
    ram_cell[   18584] = 32'h3653a83f;
    ram_cell[   18585] = 32'h60e459d1;
    ram_cell[   18586] = 32'hed0fb32d;
    ram_cell[   18587] = 32'h32ee2a31;
    ram_cell[   18588] = 32'hfc515771;
    ram_cell[   18589] = 32'hdb4e3b85;
    ram_cell[   18590] = 32'he38e2e43;
    ram_cell[   18591] = 32'h56667252;
    ram_cell[   18592] = 32'h0b5843d0;
    ram_cell[   18593] = 32'h4cba972e;
    ram_cell[   18594] = 32'h1ed82c2f;
    ram_cell[   18595] = 32'h14f011e3;
    ram_cell[   18596] = 32'h485df854;
    ram_cell[   18597] = 32'ha9a6d2e0;
    ram_cell[   18598] = 32'h20a27a65;
    ram_cell[   18599] = 32'h87c5c113;
    ram_cell[   18600] = 32'he8f552c3;
    ram_cell[   18601] = 32'hee2f9734;
    ram_cell[   18602] = 32'he5da8023;
    ram_cell[   18603] = 32'h25083d6a;
    ram_cell[   18604] = 32'h4a01a63d;
    ram_cell[   18605] = 32'h5b13adb2;
    ram_cell[   18606] = 32'h43b5f5eb;
    ram_cell[   18607] = 32'h3e1da7cf;
    ram_cell[   18608] = 32'hb9cee18b;
    ram_cell[   18609] = 32'he0c41d56;
    ram_cell[   18610] = 32'h876fd650;
    ram_cell[   18611] = 32'h4a01fbd0;
    ram_cell[   18612] = 32'h4989b563;
    ram_cell[   18613] = 32'h6c3b4a0e;
    ram_cell[   18614] = 32'h83b2cbb3;
    ram_cell[   18615] = 32'he40131a2;
    ram_cell[   18616] = 32'h53be40e5;
    ram_cell[   18617] = 32'hcca6808f;
    ram_cell[   18618] = 32'h40492ec2;
    ram_cell[   18619] = 32'hcbe60490;
    ram_cell[   18620] = 32'hc493fe8f;
    ram_cell[   18621] = 32'h5a3c3587;
    ram_cell[   18622] = 32'h196d48b7;
    ram_cell[   18623] = 32'h54bf0ae2;
    ram_cell[   18624] = 32'hdd7f0b51;
    ram_cell[   18625] = 32'h3d8fbe7c;
    ram_cell[   18626] = 32'h99c6d073;
    ram_cell[   18627] = 32'h35d54e07;
    ram_cell[   18628] = 32'h2b224471;
    ram_cell[   18629] = 32'h8ae62b2d;
    ram_cell[   18630] = 32'h7fd3b5a3;
    ram_cell[   18631] = 32'he3509ab8;
    ram_cell[   18632] = 32'h409cea98;
    ram_cell[   18633] = 32'h7d8ca6a7;
    ram_cell[   18634] = 32'h59e7c997;
    ram_cell[   18635] = 32'h8ba0079e;
    ram_cell[   18636] = 32'hecf465a6;
    ram_cell[   18637] = 32'hb2b70ae7;
    ram_cell[   18638] = 32'h824724f3;
    ram_cell[   18639] = 32'h0e862c98;
    ram_cell[   18640] = 32'h325451a2;
    ram_cell[   18641] = 32'hea79c8a0;
    ram_cell[   18642] = 32'haebf92f3;
    ram_cell[   18643] = 32'h0ef35b75;
    ram_cell[   18644] = 32'hf06a5273;
    ram_cell[   18645] = 32'h9f3eaa0e;
    ram_cell[   18646] = 32'h3a1344a9;
    ram_cell[   18647] = 32'h33a73986;
    ram_cell[   18648] = 32'h5d060352;
    ram_cell[   18649] = 32'h17d06d5a;
    ram_cell[   18650] = 32'hdce95e59;
    ram_cell[   18651] = 32'hdf57ecb8;
    ram_cell[   18652] = 32'h941b2f7d;
    ram_cell[   18653] = 32'hffbf3bdb;
    ram_cell[   18654] = 32'h2b864160;
    ram_cell[   18655] = 32'ha38a8308;
    ram_cell[   18656] = 32'h6ad81dc5;
    ram_cell[   18657] = 32'hc01ecffb;
    ram_cell[   18658] = 32'h8a7d438a;
    ram_cell[   18659] = 32'habd5c67c;
    ram_cell[   18660] = 32'hf5bbfcfe;
    ram_cell[   18661] = 32'h8be4f6c4;
    ram_cell[   18662] = 32'h480cc925;
    ram_cell[   18663] = 32'h181b1134;
    ram_cell[   18664] = 32'hd1068e76;
    ram_cell[   18665] = 32'h2fac9e98;
    ram_cell[   18666] = 32'h1491badf;
    ram_cell[   18667] = 32'h1c2d15ab;
    ram_cell[   18668] = 32'hcfa5a786;
    ram_cell[   18669] = 32'h33afba2c;
    ram_cell[   18670] = 32'h59ab1ce0;
    ram_cell[   18671] = 32'ha1b0d614;
    ram_cell[   18672] = 32'hffe10be1;
    ram_cell[   18673] = 32'h2fb49b87;
    ram_cell[   18674] = 32'h1c197b69;
    ram_cell[   18675] = 32'hab4cb9fa;
    ram_cell[   18676] = 32'h4ae0e99c;
    ram_cell[   18677] = 32'h83f8dcfa;
    ram_cell[   18678] = 32'hb2873d33;
    ram_cell[   18679] = 32'ha23bdcf2;
    ram_cell[   18680] = 32'h828eedce;
    ram_cell[   18681] = 32'h52ccea43;
    ram_cell[   18682] = 32'h10228c5d;
    ram_cell[   18683] = 32'hd4bf79c8;
    ram_cell[   18684] = 32'h4b166773;
    ram_cell[   18685] = 32'h15bdf30b;
    ram_cell[   18686] = 32'hcf7c7332;
    ram_cell[   18687] = 32'h9cf3eeab;
    ram_cell[   18688] = 32'h41cda17a;
    ram_cell[   18689] = 32'h691620d6;
    ram_cell[   18690] = 32'hf4b44b88;
    ram_cell[   18691] = 32'hba79eeb3;
    ram_cell[   18692] = 32'h46f1e485;
    ram_cell[   18693] = 32'ha909acd0;
    ram_cell[   18694] = 32'h4e94b91e;
    ram_cell[   18695] = 32'h09d8e6cf;
    ram_cell[   18696] = 32'he9ff638d;
    ram_cell[   18697] = 32'h8ce90e43;
    ram_cell[   18698] = 32'hcb24798b;
    ram_cell[   18699] = 32'h86397390;
    ram_cell[   18700] = 32'heaf300bc;
    ram_cell[   18701] = 32'h2b3d5c46;
    ram_cell[   18702] = 32'hc0b6c428;
    ram_cell[   18703] = 32'h31a9f0f7;
    ram_cell[   18704] = 32'h7f0bdd64;
    ram_cell[   18705] = 32'hc21f0526;
    ram_cell[   18706] = 32'h63ccfa28;
    ram_cell[   18707] = 32'h916cee73;
    ram_cell[   18708] = 32'h5287c099;
    ram_cell[   18709] = 32'hc80689f0;
    ram_cell[   18710] = 32'h928af452;
    ram_cell[   18711] = 32'h578f549f;
    ram_cell[   18712] = 32'hbe8b53e4;
    ram_cell[   18713] = 32'hc8557180;
    ram_cell[   18714] = 32'h311a299d;
    ram_cell[   18715] = 32'h084ac60c;
    ram_cell[   18716] = 32'h3ec9cbda;
    ram_cell[   18717] = 32'h4f7ee06b;
    ram_cell[   18718] = 32'he5b356f7;
    ram_cell[   18719] = 32'h1e3c6c3c;
    ram_cell[   18720] = 32'h3375cbdb;
    ram_cell[   18721] = 32'hb5b6658b;
    ram_cell[   18722] = 32'h096f258e;
    ram_cell[   18723] = 32'hcd04a3e1;
    ram_cell[   18724] = 32'h517fffee;
    ram_cell[   18725] = 32'h01afe580;
    ram_cell[   18726] = 32'hc5ded930;
    ram_cell[   18727] = 32'h2afa016a;
    ram_cell[   18728] = 32'hfb6f2007;
    ram_cell[   18729] = 32'he810f8e2;
    ram_cell[   18730] = 32'hf4b1c001;
    ram_cell[   18731] = 32'hfb87880a;
    ram_cell[   18732] = 32'hb574ebdb;
    ram_cell[   18733] = 32'h193f18c7;
    ram_cell[   18734] = 32'h5b6ab21c;
    ram_cell[   18735] = 32'hf72dc827;
    ram_cell[   18736] = 32'h445c38fd;
    ram_cell[   18737] = 32'hcbe2981b;
    ram_cell[   18738] = 32'hff45961b;
    ram_cell[   18739] = 32'h97323ffe;
    ram_cell[   18740] = 32'hde7eea7b;
    ram_cell[   18741] = 32'h1d0b9e07;
    ram_cell[   18742] = 32'h678d87b7;
    ram_cell[   18743] = 32'hc5fab262;
    ram_cell[   18744] = 32'h82d46232;
    ram_cell[   18745] = 32'h07d074ce;
    ram_cell[   18746] = 32'h6ddeed02;
    ram_cell[   18747] = 32'h51b90241;
    ram_cell[   18748] = 32'hcefca8da;
    ram_cell[   18749] = 32'hfbc6ed56;
    ram_cell[   18750] = 32'hc4612e7a;
    ram_cell[   18751] = 32'h646ab37e;
    ram_cell[   18752] = 32'hcc778a8a;
    ram_cell[   18753] = 32'ha17009a5;
    ram_cell[   18754] = 32'h0e83f873;
    ram_cell[   18755] = 32'h88940175;
    ram_cell[   18756] = 32'hffd5106d;
    ram_cell[   18757] = 32'h6819e834;
    ram_cell[   18758] = 32'hfa4dda17;
    ram_cell[   18759] = 32'h85146f8e;
    ram_cell[   18760] = 32'h41728b47;
    ram_cell[   18761] = 32'h2686130d;
    ram_cell[   18762] = 32'hc713a6fc;
    ram_cell[   18763] = 32'hb6c4e31d;
    ram_cell[   18764] = 32'h04a67974;
    ram_cell[   18765] = 32'h2d4113f1;
    ram_cell[   18766] = 32'hd64302a9;
    ram_cell[   18767] = 32'h252ad664;
    ram_cell[   18768] = 32'hcbfe3719;
    ram_cell[   18769] = 32'h1462cb54;
    ram_cell[   18770] = 32'hd9848548;
    ram_cell[   18771] = 32'h6383441c;
    ram_cell[   18772] = 32'h843621be;
    ram_cell[   18773] = 32'h28b64ce5;
    ram_cell[   18774] = 32'h01c507e5;
    ram_cell[   18775] = 32'hc86fc04d;
    ram_cell[   18776] = 32'h98bd43c3;
    ram_cell[   18777] = 32'h7ffd5e78;
    ram_cell[   18778] = 32'hd310830c;
    ram_cell[   18779] = 32'h706e8738;
    ram_cell[   18780] = 32'h62933211;
    ram_cell[   18781] = 32'hab1256ed;
    ram_cell[   18782] = 32'h34d856fc;
    ram_cell[   18783] = 32'habca0de8;
    ram_cell[   18784] = 32'hebee0675;
    ram_cell[   18785] = 32'hf6fd1afc;
    ram_cell[   18786] = 32'hb5651315;
    ram_cell[   18787] = 32'hbff971d0;
    ram_cell[   18788] = 32'h93b20e03;
    ram_cell[   18789] = 32'h3cacdc0e;
    ram_cell[   18790] = 32'h8e7e4318;
    ram_cell[   18791] = 32'h9ba51835;
    ram_cell[   18792] = 32'h3c59c8d5;
    ram_cell[   18793] = 32'hc6a467b7;
    ram_cell[   18794] = 32'hc90a8cb0;
    ram_cell[   18795] = 32'h8bcb9ac2;
    ram_cell[   18796] = 32'h53e9f412;
    ram_cell[   18797] = 32'h2bfb41cd;
    ram_cell[   18798] = 32'h4d50bd96;
    ram_cell[   18799] = 32'h9be8a167;
    ram_cell[   18800] = 32'h493e4b77;
    ram_cell[   18801] = 32'h9c65034f;
    ram_cell[   18802] = 32'h68470dac;
    ram_cell[   18803] = 32'hee622e50;
    ram_cell[   18804] = 32'hbfc8ee8f;
    ram_cell[   18805] = 32'hf454cc0b;
    ram_cell[   18806] = 32'ha1cb49e6;
    ram_cell[   18807] = 32'hfe71f514;
    ram_cell[   18808] = 32'hb95ab291;
    ram_cell[   18809] = 32'h4064bf86;
    ram_cell[   18810] = 32'h722b124b;
    ram_cell[   18811] = 32'h6f74b8bc;
    ram_cell[   18812] = 32'h8cc10709;
    ram_cell[   18813] = 32'h58410b97;
    ram_cell[   18814] = 32'haee4c4d4;
    ram_cell[   18815] = 32'h20b33df9;
    ram_cell[   18816] = 32'hc528a91d;
    ram_cell[   18817] = 32'hc4bfb430;
    ram_cell[   18818] = 32'hab49a5ec;
    ram_cell[   18819] = 32'h6b2975c2;
    ram_cell[   18820] = 32'had5e39e7;
    ram_cell[   18821] = 32'hf513fb36;
    ram_cell[   18822] = 32'hb04e616f;
    ram_cell[   18823] = 32'h6aaa8ccb;
    ram_cell[   18824] = 32'h91d40361;
    ram_cell[   18825] = 32'h3888d08f;
    ram_cell[   18826] = 32'hdffcd74d;
    ram_cell[   18827] = 32'hdce0fd4e;
    ram_cell[   18828] = 32'h59abd139;
    ram_cell[   18829] = 32'hcaa7a57c;
    ram_cell[   18830] = 32'hf78f9beb;
    ram_cell[   18831] = 32'hf06e64f9;
    ram_cell[   18832] = 32'ha36e3841;
    ram_cell[   18833] = 32'hd7efca67;
    ram_cell[   18834] = 32'ha2772eae;
    ram_cell[   18835] = 32'h763fc5c6;
    ram_cell[   18836] = 32'h918a68f3;
    ram_cell[   18837] = 32'h1c2f3909;
    ram_cell[   18838] = 32'h4452da28;
    ram_cell[   18839] = 32'hbeb0d5af;
    ram_cell[   18840] = 32'hb396ca02;
    ram_cell[   18841] = 32'h441bdfdd;
    ram_cell[   18842] = 32'hd567ade8;
    ram_cell[   18843] = 32'hee0d62b9;
    ram_cell[   18844] = 32'h9311a42b;
    ram_cell[   18845] = 32'hba62849c;
    ram_cell[   18846] = 32'h7ad52efe;
    ram_cell[   18847] = 32'h380be2b9;
    ram_cell[   18848] = 32'h2e6ba25e;
    ram_cell[   18849] = 32'h43bc5726;
    ram_cell[   18850] = 32'h93412fdd;
    ram_cell[   18851] = 32'hbc45cba5;
    ram_cell[   18852] = 32'h0ffd1cbb;
    ram_cell[   18853] = 32'h2e720ffd;
    ram_cell[   18854] = 32'h921f012e;
    ram_cell[   18855] = 32'h7c7ab5f2;
    ram_cell[   18856] = 32'h1c31386d;
    ram_cell[   18857] = 32'h34a62c12;
    ram_cell[   18858] = 32'hd54f5d28;
    ram_cell[   18859] = 32'h6e70a33f;
    ram_cell[   18860] = 32'hdec20a0a;
    ram_cell[   18861] = 32'h0f2e5b28;
    ram_cell[   18862] = 32'h541195ff;
    ram_cell[   18863] = 32'h4f0cd18b;
    ram_cell[   18864] = 32'h7a331b8f;
    ram_cell[   18865] = 32'h84121457;
    ram_cell[   18866] = 32'h37662e1e;
    ram_cell[   18867] = 32'h0e9b0229;
    ram_cell[   18868] = 32'h8b78e929;
    ram_cell[   18869] = 32'h5fdb32ea;
    ram_cell[   18870] = 32'h693b875d;
    ram_cell[   18871] = 32'hdae9c76e;
    ram_cell[   18872] = 32'h916e7360;
    ram_cell[   18873] = 32'he2616d3d;
    ram_cell[   18874] = 32'h1839a4ca;
    ram_cell[   18875] = 32'h160cec49;
    ram_cell[   18876] = 32'hac4af4bc;
    ram_cell[   18877] = 32'h1dd0d9f3;
    ram_cell[   18878] = 32'h9c86ac63;
    ram_cell[   18879] = 32'h5501d20e;
    ram_cell[   18880] = 32'h329f7dbd;
    ram_cell[   18881] = 32'h88716d52;
    ram_cell[   18882] = 32'h5782f641;
    ram_cell[   18883] = 32'h2218e95f;
    ram_cell[   18884] = 32'he8b75891;
    ram_cell[   18885] = 32'h3377d378;
    ram_cell[   18886] = 32'h39520c71;
    ram_cell[   18887] = 32'h5dd5e3a4;
    ram_cell[   18888] = 32'hbb75771e;
    ram_cell[   18889] = 32'h3fa71a20;
    ram_cell[   18890] = 32'hf48190b5;
    ram_cell[   18891] = 32'h85eeb823;
    ram_cell[   18892] = 32'hdbff6fff;
    ram_cell[   18893] = 32'h9cf83869;
    ram_cell[   18894] = 32'h6ea8a82f;
    ram_cell[   18895] = 32'hc7bc1891;
    ram_cell[   18896] = 32'h69153bcf;
    ram_cell[   18897] = 32'ha70669d9;
    ram_cell[   18898] = 32'hde61255e;
    ram_cell[   18899] = 32'haf446c1c;
    ram_cell[   18900] = 32'h720c70fc;
    ram_cell[   18901] = 32'hbbefd980;
    ram_cell[   18902] = 32'hf082b264;
    ram_cell[   18903] = 32'h92fed86c;
    ram_cell[   18904] = 32'hb82c1591;
    ram_cell[   18905] = 32'h599b977c;
    ram_cell[   18906] = 32'h4a103733;
    ram_cell[   18907] = 32'h5edd5b8c;
    ram_cell[   18908] = 32'hc84b49ec;
    ram_cell[   18909] = 32'h7aa4d97d;
    ram_cell[   18910] = 32'hb0bb8d1b;
    ram_cell[   18911] = 32'h26712261;
    ram_cell[   18912] = 32'h16af81b3;
    ram_cell[   18913] = 32'hc2a2af14;
    ram_cell[   18914] = 32'h5e944eb3;
    ram_cell[   18915] = 32'h56d7c020;
    ram_cell[   18916] = 32'hfa347c75;
    ram_cell[   18917] = 32'hb138b88f;
    ram_cell[   18918] = 32'hf3776935;
    ram_cell[   18919] = 32'h52c7cc92;
    ram_cell[   18920] = 32'h5f20a7a2;
    ram_cell[   18921] = 32'hca92f458;
    ram_cell[   18922] = 32'h013a2f57;
    ram_cell[   18923] = 32'he13b3b7c;
    ram_cell[   18924] = 32'h16d50488;
    ram_cell[   18925] = 32'h398d9485;
    ram_cell[   18926] = 32'hf448d7aa;
    ram_cell[   18927] = 32'h5471e2e2;
    ram_cell[   18928] = 32'h12ff7945;
    ram_cell[   18929] = 32'hc3b0e125;
    ram_cell[   18930] = 32'h75796c2b;
    ram_cell[   18931] = 32'h245133d6;
    ram_cell[   18932] = 32'h666515c3;
    ram_cell[   18933] = 32'h7361955b;
    ram_cell[   18934] = 32'h57f3e5cb;
    ram_cell[   18935] = 32'h5b0dedae;
    ram_cell[   18936] = 32'hc41abc1e;
    ram_cell[   18937] = 32'h68b23573;
    ram_cell[   18938] = 32'h4655f30c;
    ram_cell[   18939] = 32'h3f6823ed;
    ram_cell[   18940] = 32'hfb94a780;
    ram_cell[   18941] = 32'ha8933dc3;
    ram_cell[   18942] = 32'h40919b44;
    ram_cell[   18943] = 32'h9697e7dc;
    ram_cell[   18944] = 32'h261595dc;
    ram_cell[   18945] = 32'h4013cb1e;
    ram_cell[   18946] = 32'h9476cd02;
    ram_cell[   18947] = 32'hff1a1c58;
    ram_cell[   18948] = 32'h247ac95c;
    ram_cell[   18949] = 32'h63fa00c4;
    ram_cell[   18950] = 32'h00d41323;
    ram_cell[   18951] = 32'h7ff56ea1;
    ram_cell[   18952] = 32'had7721dc;
    ram_cell[   18953] = 32'h15d504ef;
    ram_cell[   18954] = 32'h64c768fa;
    ram_cell[   18955] = 32'hfd4cbe7f;
    ram_cell[   18956] = 32'ha5be9fdc;
    ram_cell[   18957] = 32'hffa4a3c1;
    ram_cell[   18958] = 32'hbce03bcf;
    ram_cell[   18959] = 32'h9ffc3214;
    ram_cell[   18960] = 32'h1f80923e;
    ram_cell[   18961] = 32'haf36eb6e;
    ram_cell[   18962] = 32'h77259989;
    ram_cell[   18963] = 32'h963f296e;
    ram_cell[   18964] = 32'hd5730f73;
    ram_cell[   18965] = 32'hbcbe0335;
    ram_cell[   18966] = 32'h714b2bbb;
    ram_cell[   18967] = 32'h20e54118;
    ram_cell[   18968] = 32'h3ae55c22;
    ram_cell[   18969] = 32'hf1baf427;
    ram_cell[   18970] = 32'hd2792566;
    ram_cell[   18971] = 32'h4d1a5fc3;
    ram_cell[   18972] = 32'h08088ec6;
    ram_cell[   18973] = 32'hddac4692;
    ram_cell[   18974] = 32'h73b4b1ed;
    ram_cell[   18975] = 32'hbafc3de4;
    ram_cell[   18976] = 32'h0968808b;
    ram_cell[   18977] = 32'ha0ce44b1;
    ram_cell[   18978] = 32'hbd16bf5e;
    ram_cell[   18979] = 32'h6c5a6fe3;
    ram_cell[   18980] = 32'h0e2ca298;
    ram_cell[   18981] = 32'h77986109;
    ram_cell[   18982] = 32'h18105840;
    ram_cell[   18983] = 32'hfdb92904;
    ram_cell[   18984] = 32'h036251ba;
    ram_cell[   18985] = 32'hb636b517;
    ram_cell[   18986] = 32'h9e990ca9;
    ram_cell[   18987] = 32'h2f860642;
    ram_cell[   18988] = 32'h09eddbc7;
    ram_cell[   18989] = 32'h0ac7ca8a;
    ram_cell[   18990] = 32'h56e1d09a;
    ram_cell[   18991] = 32'h6a9cdcdd;
    ram_cell[   18992] = 32'h8cb5ccfe;
    ram_cell[   18993] = 32'h5f4bf2ea;
    ram_cell[   18994] = 32'h2ffb553b;
    ram_cell[   18995] = 32'h595cf5f1;
    ram_cell[   18996] = 32'h37b321c8;
    ram_cell[   18997] = 32'h650b6298;
    ram_cell[   18998] = 32'he057719b;
    ram_cell[   18999] = 32'h0f4b29d8;
    ram_cell[   19000] = 32'h4287e0da;
    ram_cell[   19001] = 32'h2bb4bf9e;
    ram_cell[   19002] = 32'hc9c29099;
    ram_cell[   19003] = 32'h87d14aaa;
    ram_cell[   19004] = 32'h0ee4c02b;
    ram_cell[   19005] = 32'hbfab60ae;
    ram_cell[   19006] = 32'habe91dc1;
    ram_cell[   19007] = 32'h3d44bc3b;
    ram_cell[   19008] = 32'h47d56202;
    ram_cell[   19009] = 32'h3ec47683;
    ram_cell[   19010] = 32'hf73396b2;
    ram_cell[   19011] = 32'h7f85bc60;
    ram_cell[   19012] = 32'h8004036e;
    ram_cell[   19013] = 32'hbf5add9a;
    ram_cell[   19014] = 32'h5c41f1d4;
    ram_cell[   19015] = 32'h467ec9e7;
    ram_cell[   19016] = 32'h293abbe1;
    ram_cell[   19017] = 32'he9719d2a;
    ram_cell[   19018] = 32'ha7baebb8;
    ram_cell[   19019] = 32'h9ad7b477;
    ram_cell[   19020] = 32'h8bd789e2;
    ram_cell[   19021] = 32'h664dbef3;
    ram_cell[   19022] = 32'h51e8f25e;
    ram_cell[   19023] = 32'he98921ea;
    ram_cell[   19024] = 32'hafbff2a5;
    ram_cell[   19025] = 32'hf1af1111;
    ram_cell[   19026] = 32'hfc32a2c9;
    ram_cell[   19027] = 32'h6bc521f2;
    ram_cell[   19028] = 32'hb86c87fc;
    ram_cell[   19029] = 32'hd6a72306;
    ram_cell[   19030] = 32'h4740d465;
    ram_cell[   19031] = 32'h0a4acd11;
    ram_cell[   19032] = 32'h4889a461;
    ram_cell[   19033] = 32'hb3e51f97;
    ram_cell[   19034] = 32'h59ad4d5e;
    ram_cell[   19035] = 32'h952a3d21;
    ram_cell[   19036] = 32'h958ed2e6;
    ram_cell[   19037] = 32'hc697f5b9;
    ram_cell[   19038] = 32'h5cfe551e;
    ram_cell[   19039] = 32'h125fa1de;
    ram_cell[   19040] = 32'hc01b8f4b;
    ram_cell[   19041] = 32'h452d417d;
    ram_cell[   19042] = 32'h18229091;
    ram_cell[   19043] = 32'h8f0704b4;
    ram_cell[   19044] = 32'hf6df9c2a;
    ram_cell[   19045] = 32'h3bc265a6;
    ram_cell[   19046] = 32'h637a1792;
    ram_cell[   19047] = 32'h3c1991fc;
    ram_cell[   19048] = 32'h901efdf9;
    ram_cell[   19049] = 32'h2da6fb20;
    ram_cell[   19050] = 32'he4443ac1;
    ram_cell[   19051] = 32'h961350ea;
    ram_cell[   19052] = 32'hfde8b2b1;
    ram_cell[   19053] = 32'h297e7daa;
    ram_cell[   19054] = 32'h9d6b80b1;
    ram_cell[   19055] = 32'he25f0ef0;
    ram_cell[   19056] = 32'h67a362e7;
    ram_cell[   19057] = 32'h58348f95;
    ram_cell[   19058] = 32'ha8ab5aa6;
    ram_cell[   19059] = 32'h1d433c3f;
    ram_cell[   19060] = 32'ha353b23d;
    ram_cell[   19061] = 32'h993a14ce;
    ram_cell[   19062] = 32'hf4940f64;
    ram_cell[   19063] = 32'h648b862e;
    ram_cell[   19064] = 32'hfb7beb60;
    ram_cell[   19065] = 32'h598d9867;
    ram_cell[   19066] = 32'h8a302e4c;
    ram_cell[   19067] = 32'he6d41a70;
    ram_cell[   19068] = 32'hb90f9082;
    ram_cell[   19069] = 32'h0bcaa466;
    ram_cell[   19070] = 32'h77844513;
    ram_cell[   19071] = 32'hc0cf881c;
    ram_cell[   19072] = 32'hfc9e2087;
    ram_cell[   19073] = 32'h660a032d;
    ram_cell[   19074] = 32'h87ee9648;
    ram_cell[   19075] = 32'h1908e538;
    ram_cell[   19076] = 32'hf583d749;
    ram_cell[   19077] = 32'he87cf9dd;
    ram_cell[   19078] = 32'h27dba523;
    ram_cell[   19079] = 32'h21fce62b;
    ram_cell[   19080] = 32'h9dbb281d;
    ram_cell[   19081] = 32'h88ce567b;
    ram_cell[   19082] = 32'hc9e0c0d4;
    ram_cell[   19083] = 32'h4b8cf285;
    ram_cell[   19084] = 32'hadf15eca;
    ram_cell[   19085] = 32'h760c7fb6;
    ram_cell[   19086] = 32'h71584bb3;
    ram_cell[   19087] = 32'h6b2a6d8b;
    ram_cell[   19088] = 32'h93983a72;
    ram_cell[   19089] = 32'h06111344;
    ram_cell[   19090] = 32'h9ec2542e;
    ram_cell[   19091] = 32'h9671a9b8;
    ram_cell[   19092] = 32'hc1495638;
    ram_cell[   19093] = 32'h4a66b90c;
    ram_cell[   19094] = 32'h3fac68d5;
    ram_cell[   19095] = 32'hc072da9a;
    ram_cell[   19096] = 32'hbbe8f779;
    ram_cell[   19097] = 32'h62f7159a;
    ram_cell[   19098] = 32'hc37b977d;
    ram_cell[   19099] = 32'h9dbe7508;
    ram_cell[   19100] = 32'h9d69a669;
    ram_cell[   19101] = 32'h92ceb6e5;
    ram_cell[   19102] = 32'h2edd4512;
    ram_cell[   19103] = 32'h33c1218f;
    ram_cell[   19104] = 32'ha1d55f2f;
    ram_cell[   19105] = 32'h7142b1c9;
    ram_cell[   19106] = 32'hed905369;
    ram_cell[   19107] = 32'h6b21c9a5;
    ram_cell[   19108] = 32'h74df98bf;
    ram_cell[   19109] = 32'h0ab5bdb7;
    ram_cell[   19110] = 32'h55af1c66;
    ram_cell[   19111] = 32'h6649d869;
    ram_cell[   19112] = 32'h3e92b0e7;
    ram_cell[   19113] = 32'h2c0c4ad6;
    ram_cell[   19114] = 32'h08e8c977;
    ram_cell[   19115] = 32'hdd0d366e;
    ram_cell[   19116] = 32'hbaeb63d6;
    ram_cell[   19117] = 32'ha873ac84;
    ram_cell[   19118] = 32'h0a2cd91e;
    ram_cell[   19119] = 32'h161504f0;
    ram_cell[   19120] = 32'hd4701420;
    ram_cell[   19121] = 32'hc50b0642;
    ram_cell[   19122] = 32'h7eae0299;
    ram_cell[   19123] = 32'h72780120;
    ram_cell[   19124] = 32'hbf2e055a;
    ram_cell[   19125] = 32'h70ce4a8a;
    ram_cell[   19126] = 32'hb6581935;
    ram_cell[   19127] = 32'hd0608233;
    ram_cell[   19128] = 32'h33d4b883;
    ram_cell[   19129] = 32'h333a4264;
    ram_cell[   19130] = 32'he653def1;
    ram_cell[   19131] = 32'h83c327b9;
    ram_cell[   19132] = 32'hb145264b;
    ram_cell[   19133] = 32'hbb9527cb;
    ram_cell[   19134] = 32'h0b7f2116;
    ram_cell[   19135] = 32'ha9d012b4;
    ram_cell[   19136] = 32'h9812a0d5;
    ram_cell[   19137] = 32'h547bd538;
    ram_cell[   19138] = 32'h870796a7;
    ram_cell[   19139] = 32'ha4584a54;
    ram_cell[   19140] = 32'h2b1d1ad1;
    ram_cell[   19141] = 32'h5b0de44c;
    ram_cell[   19142] = 32'h6e844f3f;
    ram_cell[   19143] = 32'hc2d27469;
    ram_cell[   19144] = 32'h02b286a0;
    ram_cell[   19145] = 32'h5813c9c6;
    ram_cell[   19146] = 32'h1b5dd9bb;
    ram_cell[   19147] = 32'h2b6c1f81;
    ram_cell[   19148] = 32'hde45f58e;
    ram_cell[   19149] = 32'h20867cf5;
    ram_cell[   19150] = 32'h2b9ed106;
    ram_cell[   19151] = 32'h34f7c47a;
    ram_cell[   19152] = 32'h7070ca36;
    ram_cell[   19153] = 32'h3d73bec0;
    ram_cell[   19154] = 32'hec3e6fe0;
    ram_cell[   19155] = 32'hd4859d28;
    ram_cell[   19156] = 32'hd18d7940;
    ram_cell[   19157] = 32'h4ab40f62;
    ram_cell[   19158] = 32'h512f594d;
    ram_cell[   19159] = 32'ha70d6dc0;
    ram_cell[   19160] = 32'hf7b3e9ef;
    ram_cell[   19161] = 32'h87299dc6;
    ram_cell[   19162] = 32'hc78d4658;
    ram_cell[   19163] = 32'h2d82c1d6;
    ram_cell[   19164] = 32'h4dd9531c;
    ram_cell[   19165] = 32'h39daeb4f;
    ram_cell[   19166] = 32'hbc6b4c58;
    ram_cell[   19167] = 32'h820be664;
    ram_cell[   19168] = 32'h765a3c5b;
    ram_cell[   19169] = 32'h8094c7c2;
    ram_cell[   19170] = 32'h0414d0f6;
    ram_cell[   19171] = 32'h6d9c153a;
    ram_cell[   19172] = 32'h99fa608c;
    ram_cell[   19173] = 32'heaffceba;
    ram_cell[   19174] = 32'hd73c4a59;
    ram_cell[   19175] = 32'hcbfdcb19;
    ram_cell[   19176] = 32'ha4c0407b;
    ram_cell[   19177] = 32'h35fb6967;
    ram_cell[   19178] = 32'hd4d86fe4;
    ram_cell[   19179] = 32'hbed1853d;
    ram_cell[   19180] = 32'h3366bcd9;
    ram_cell[   19181] = 32'hb0936f96;
    ram_cell[   19182] = 32'hfc4f09fb;
    ram_cell[   19183] = 32'ha83a8d78;
    ram_cell[   19184] = 32'h7544ad3f;
    ram_cell[   19185] = 32'hc334c5f4;
    ram_cell[   19186] = 32'he49bb01d;
    ram_cell[   19187] = 32'hfbb962b7;
    ram_cell[   19188] = 32'hfa067a0d;
    ram_cell[   19189] = 32'h10be1462;
    ram_cell[   19190] = 32'h2bd01e4c;
    ram_cell[   19191] = 32'h1ccde8d9;
    ram_cell[   19192] = 32'h4ec94736;
    ram_cell[   19193] = 32'h9f4958e1;
    ram_cell[   19194] = 32'hb16efef5;
    ram_cell[   19195] = 32'hb32af24b;
    ram_cell[   19196] = 32'ha1b95533;
    ram_cell[   19197] = 32'h70988358;
    ram_cell[   19198] = 32'h988b77b9;
    ram_cell[   19199] = 32'hbfbf570d;
    ram_cell[   19200] = 32'h9fe576ca;
    ram_cell[   19201] = 32'hf04776fd;
    ram_cell[   19202] = 32'hde21b583;
    ram_cell[   19203] = 32'h78e53d55;
    ram_cell[   19204] = 32'h15e269bc;
    ram_cell[   19205] = 32'hd7427235;
    ram_cell[   19206] = 32'h5545f647;
    ram_cell[   19207] = 32'h74c10302;
    ram_cell[   19208] = 32'h8b8de661;
    ram_cell[   19209] = 32'hef23e9fa;
    ram_cell[   19210] = 32'hdd92eb21;
    ram_cell[   19211] = 32'h8b638254;
    ram_cell[   19212] = 32'hadc1cd62;
    ram_cell[   19213] = 32'h2dff816b;
    ram_cell[   19214] = 32'h2bf35b6e;
    ram_cell[   19215] = 32'h135b7eb6;
    ram_cell[   19216] = 32'h99d1efdf;
    ram_cell[   19217] = 32'h4410a901;
    ram_cell[   19218] = 32'h78efac3a;
    ram_cell[   19219] = 32'h48d64929;
    ram_cell[   19220] = 32'hb91594f3;
    ram_cell[   19221] = 32'h0cd8703e;
    ram_cell[   19222] = 32'h366f5729;
    ram_cell[   19223] = 32'h8fa5d059;
    ram_cell[   19224] = 32'h20286290;
    ram_cell[   19225] = 32'hed250dfd;
    ram_cell[   19226] = 32'h06979e1e;
    ram_cell[   19227] = 32'h40c9cfe0;
    ram_cell[   19228] = 32'hfede9b66;
    ram_cell[   19229] = 32'h40a7aa2e;
    ram_cell[   19230] = 32'hd58aae4b;
    ram_cell[   19231] = 32'hb35894f8;
    ram_cell[   19232] = 32'hed2786d7;
    ram_cell[   19233] = 32'hfeb92fda;
    ram_cell[   19234] = 32'h09735a06;
    ram_cell[   19235] = 32'h8809481d;
    ram_cell[   19236] = 32'h8133559a;
    ram_cell[   19237] = 32'h5acb61f2;
    ram_cell[   19238] = 32'h7cc05bf6;
    ram_cell[   19239] = 32'hdad41045;
    ram_cell[   19240] = 32'hecbb7f1d;
    ram_cell[   19241] = 32'ha972ee64;
    ram_cell[   19242] = 32'ha00be562;
    ram_cell[   19243] = 32'hc90b1f65;
    ram_cell[   19244] = 32'h1c7cc8e6;
    ram_cell[   19245] = 32'hd919cd32;
    ram_cell[   19246] = 32'h27405d9e;
    ram_cell[   19247] = 32'h04198972;
    ram_cell[   19248] = 32'h042d6dc8;
    ram_cell[   19249] = 32'h3d1f5632;
    ram_cell[   19250] = 32'h025fdd8f;
    ram_cell[   19251] = 32'h3cf7fa99;
    ram_cell[   19252] = 32'hb7b9c0ac;
    ram_cell[   19253] = 32'hefb88e2e;
    ram_cell[   19254] = 32'hdde69199;
    ram_cell[   19255] = 32'h1e39321e;
    ram_cell[   19256] = 32'h854d93ed;
    ram_cell[   19257] = 32'h94bbb460;
    ram_cell[   19258] = 32'h36310f53;
    ram_cell[   19259] = 32'h5eb3e01c;
    ram_cell[   19260] = 32'h72fd87a8;
    ram_cell[   19261] = 32'h28a6edd9;
    ram_cell[   19262] = 32'h6d9e7654;
    ram_cell[   19263] = 32'h397bf606;
    ram_cell[   19264] = 32'h912cc86b;
    ram_cell[   19265] = 32'h65eb72d9;
    ram_cell[   19266] = 32'h36045c6b;
    ram_cell[   19267] = 32'h186285fb;
    ram_cell[   19268] = 32'h9f1f4033;
    ram_cell[   19269] = 32'h9607da46;
    ram_cell[   19270] = 32'hdaea810a;
    ram_cell[   19271] = 32'ha7a0ced4;
    ram_cell[   19272] = 32'h3f2fecd7;
    ram_cell[   19273] = 32'hb14cf8e1;
    ram_cell[   19274] = 32'h657cf054;
    ram_cell[   19275] = 32'hcd531853;
    ram_cell[   19276] = 32'h6061fb49;
    ram_cell[   19277] = 32'h536647d9;
    ram_cell[   19278] = 32'h722d3364;
    ram_cell[   19279] = 32'h8ce725ba;
    ram_cell[   19280] = 32'h983b35f3;
    ram_cell[   19281] = 32'h7503f1fb;
    ram_cell[   19282] = 32'hd4f54617;
    ram_cell[   19283] = 32'h9dbfed25;
    ram_cell[   19284] = 32'h95e18a81;
    ram_cell[   19285] = 32'hac7f536c;
    ram_cell[   19286] = 32'h1834e2e4;
    ram_cell[   19287] = 32'h243c739c;
    ram_cell[   19288] = 32'h3fc8fb3c;
    ram_cell[   19289] = 32'h5cecb11c;
    ram_cell[   19290] = 32'h2843c19e;
    ram_cell[   19291] = 32'h3aa5b43f;
    ram_cell[   19292] = 32'h24033e88;
    ram_cell[   19293] = 32'ha0fd6105;
    ram_cell[   19294] = 32'h27172934;
    ram_cell[   19295] = 32'h8238d22f;
    ram_cell[   19296] = 32'hdafbc2ce;
    ram_cell[   19297] = 32'ha63291f2;
    ram_cell[   19298] = 32'hb0b66c1e;
    ram_cell[   19299] = 32'h39313fb1;
    ram_cell[   19300] = 32'hce0f0edf;
    ram_cell[   19301] = 32'hbab30516;
    ram_cell[   19302] = 32'hda1fdbb5;
    ram_cell[   19303] = 32'h4e2d1571;
    ram_cell[   19304] = 32'h69ac0963;
    ram_cell[   19305] = 32'h35151e17;
    ram_cell[   19306] = 32'h99778c98;
    ram_cell[   19307] = 32'hf8ff7f87;
    ram_cell[   19308] = 32'hfd6d1000;
    ram_cell[   19309] = 32'hb8bd1578;
    ram_cell[   19310] = 32'hff08032e;
    ram_cell[   19311] = 32'hda70ff40;
    ram_cell[   19312] = 32'hbe3568bf;
    ram_cell[   19313] = 32'h76913d69;
    ram_cell[   19314] = 32'h8a286843;
    ram_cell[   19315] = 32'hb89762df;
    ram_cell[   19316] = 32'h77c5c91b;
    ram_cell[   19317] = 32'h7a7aa937;
    ram_cell[   19318] = 32'h41fa32f4;
    ram_cell[   19319] = 32'haed5bf9a;
    ram_cell[   19320] = 32'h729161a3;
    ram_cell[   19321] = 32'hfc72af47;
    ram_cell[   19322] = 32'h134fa638;
    ram_cell[   19323] = 32'h4189385e;
    ram_cell[   19324] = 32'h0b65fd83;
    ram_cell[   19325] = 32'h4aff9580;
    ram_cell[   19326] = 32'h676f7de6;
    ram_cell[   19327] = 32'h2f54e4c1;
    ram_cell[   19328] = 32'heddc3b09;
    ram_cell[   19329] = 32'hfe6157a4;
    ram_cell[   19330] = 32'hc759278a;
    ram_cell[   19331] = 32'h4a310426;
    ram_cell[   19332] = 32'hd3a147ba;
    ram_cell[   19333] = 32'h4e8f119c;
    ram_cell[   19334] = 32'ha8efa9d9;
    ram_cell[   19335] = 32'h9bddc98b;
    ram_cell[   19336] = 32'h9313684f;
    ram_cell[   19337] = 32'he2688fbb;
    ram_cell[   19338] = 32'h35010a20;
    ram_cell[   19339] = 32'h3af47c6f;
    ram_cell[   19340] = 32'h76252751;
    ram_cell[   19341] = 32'hcdd21946;
    ram_cell[   19342] = 32'h966f5f1c;
    ram_cell[   19343] = 32'hf0e17162;
    ram_cell[   19344] = 32'hee4692ea;
    ram_cell[   19345] = 32'h800f36d1;
    ram_cell[   19346] = 32'h6883162e;
    ram_cell[   19347] = 32'hf2c8763c;
    ram_cell[   19348] = 32'h4571b8eb;
    ram_cell[   19349] = 32'h5383463f;
    ram_cell[   19350] = 32'h84aa0d21;
    ram_cell[   19351] = 32'h73c6b899;
    ram_cell[   19352] = 32'hfcc64ce2;
    ram_cell[   19353] = 32'hf96e131a;
    ram_cell[   19354] = 32'he7a72ae5;
    ram_cell[   19355] = 32'hbf0bcd16;
    ram_cell[   19356] = 32'h8b7370e8;
    ram_cell[   19357] = 32'h7a2bb3ef;
    ram_cell[   19358] = 32'h656d8b9c;
    ram_cell[   19359] = 32'h9d519ec5;
    ram_cell[   19360] = 32'hbbffd2fc;
    ram_cell[   19361] = 32'h86cf29d9;
    ram_cell[   19362] = 32'h55a05ba1;
    ram_cell[   19363] = 32'h9fd7ca4b;
    ram_cell[   19364] = 32'hd83a5ff5;
    ram_cell[   19365] = 32'h728347d6;
    ram_cell[   19366] = 32'h84203e0a;
    ram_cell[   19367] = 32'h14d732eb;
    ram_cell[   19368] = 32'h96f98f1a;
    ram_cell[   19369] = 32'h8890837f;
    ram_cell[   19370] = 32'hdcc813aa;
    ram_cell[   19371] = 32'h4f82af61;
    ram_cell[   19372] = 32'hc0547f3f;
    ram_cell[   19373] = 32'h630084f9;
    ram_cell[   19374] = 32'h0fe5f621;
    ram_cell[   19375] = 32'h084463e8;
    ram_cell[   19376] = 32'hb90ae083;
    ram_cell[   19377] = 32'h9fd07987;
    ram_cell[   19378] = 32'h8e17ddb1;
    ram_cell[   19379] = 32'h38b0efca;
    ram_cell[   19380] = 32'ha968a94e;
    ram_cell[   19381] = 32'h4ea78859;
    ram_cell[   19382] = 32'hf1b3f74b;
    ram_cell[   19383] = 32'h4aee349a;
    ram_cell[   19384] = 32'h7caf9fec;
    ram_cell[   19385] = 32'h54cc9afd;
    ram_cell[   19386] = 32'hf92f0373;
    ram_cell[   19387] = 32'h40b830ff;
    ram_cell[   19388] = 32'hf57bf62a;
    ram_cell[   19389] = 32'h146cb5f6;
    ram_cell[   19390] = 32'h3569181c;
    ram_cell[   19391] = 32'hc426c177;
    ram_cell[   19392] = 32'h3abe67ae;
    ram_cell[   19393] = 32'h2d127b17;
    ram_cell[   19394] = 32'hb8835883;
    ram_cell[   19395] = 32'hf7114811;
    ram_cell[   19396] = 32'h098dc63d;
    ram_cell[   19397] = 32'h0de85ca7;
    ram_cell[   19398] = 32'h99f1aeb0;
    ram_cell[   19399] = 32'ha26370c6;
    ram_cell[   19400] = 32'h8f64817f;
    ram_cell[   19401] = 32'h1781bf98;
    ram_cell[   19402] = 32'h8162c46d;
    ram_cell[   19403] = 32'hafe95c1d;
    ram_cell[   19404] = 32'h175bdc42;
    ram_cell[   19405] = 32'hab8b02ee;
    ram_cell[   19406] = 32'hce1fbcc6;
    ram_cell[   19407] = 32'hce74e6a0;
    ram_cell[   19408] = 32'h6f61929d;
    ram_cell[   19409] = 32'h4781fbb9;
    ram_cell[   19410] = 32'he035b3da;
    ram_cell[   19411] = 32'hc7b3b82a;
    ram_cell[   19412] = 32'habf2c806;
    ram_cell[   19413] = 32'h23a14ee2;
    ram_cell[   19414] = 32'he915d712;
    ram_cell[   19415] = 32'hd268c73f;
    ram_cell[   19416] = 32'hbf201579;
    ram_cell[   19417] = 32'h3fe8e6b4;
    ram_cell[   19418] = 32'hbad6c490;
    ram_cell[   19419] = 32'h926aa27f;
    ram_cell[   19420] = 32'hfbb8dd0e;
    ram_cell[   19421] = 32'h0aff1f8d;
    ram_cell[   19422] = 32'h1f025bda;
    ram_cell[   19423] = 32'h3f84c912;
    ram_cell[   19424] = 32'hd3a456bf;
    ram_cell[   19425] = 32'hef0fd48d;
    ram_cell[   19426] = 32'h310bfbd7;
    ram_cell[   19427] = 32'h80b5b296;
    ram_cell[   19428] = 32'hd4551c8e;
    ram_cell[   19429] = 32'h1d0543f2;
    ram_cell[   19430] = 32'h46489629;
    ram_cell[   19431] = 32'hc5704bcd;
    ram_cell[   19432] = 32'hba2f4322;
    ram_cell[   19433] = 32'h9529bc3f;
    ram_cell[   19434] = 32'h833609d0;
    ram_cell[   19435] = 32'hde1a3c88;
    ram_cell[   19436] = 32'h3e6e01d7;
    ram_cell[   19437] = 32'ha6221991;
    ram_cell[   19438] = 32'h3420b7e7;
    ram_cell[   19439] = 32'h7fde7610;
    ram_cell[   19440] = 32'h6c82eb6c;
    ram_cell[   19441] = 32'h26483809;
    ram_cell[   19442] = 32'h97497156;
    ram_cell[   19443] = 32'h4bcaa827;
    ram_cell[   19444] = 32'h60f41b87;
    ram_cell[   19445] = 32'hb1a4034a;
    ram_cell[   19446] = 32'hbf7f137d;
    ram_cell[   19447] = 32'h42ddbc22;
    ram_cell[   19448] = 32'ha7da7396;
    ram_cell[   19449] = 32'h3506b511;
    ram_cell[   19450] = 32'h987ad3a3;
    ram_cell[   19451] = 32'h6188c075;
    ram_cell[   19452] = 32'hd80da0a8;
    ram_cell[   19453] = 32'h5f67ab87;
    ram_cell[   19454] = 32'hd6fa3e2d;
    ram_cell[   19455] = 32'h159a51d4;
    ram_cell[   19456] = 32'h23668981;
    ram_cell[   19457] = 32'h5468ad47;
    ram_cell[   19458] = 32'hb86b2ba8;
    ram_cell[   19459] = 32'hffbd482e;
    ram_cell[   19460] = 32'h7ff7b48f;
    ram_cell[   19461] = 32'hf93be4c8;
    ram_cell[   19462] = 32'h472cf587;
    ram_cell[   19463] = 32'h765f2995;
    ram_cell[   19464] = 32'h9bb1532d;
    ram_cell[   19465] = 32'h62f2c8b0;
    ram_cell[   19466] = 32'h45d2aebb;
    ram_cell[   19467] = 32'h15b47429;
    ram_cell[   19468] = 32'hd84020ca;
    ram_cell[   19469] = 32'h52ff56f2;
    ram_cell[   19470] = 32'h8533df63;
    ram_cell[   19471] = 32'h328a1ef6;
    ram_cell[   19472] = 32'h299b874a;
    ram_cell[   19473] = 32'h69d7c23d;
    ram_cell[   19474] = 32'h5e245b59;
    ram_cell[   19475] = 32'h266c3605;
    ram_cell[   19476] = 32'h9e0844a3;
    ram_cell[   19477] = 32'h2139c58f;
    ram_cell[   19478] = 32'h6d4be665;
    ram_cell[   19479] = 32'h570393fc;
    ram_cell[   19480] = 32'hfbdb7ac1;
    ram_cell[   19481] = 32'hf4be2f42;
    ram_cell[   19482] = 32'haa8770d2;
    ram_cell[   19483] = 32'h0f388f4f;
    ram_cell[   19484] = 32'ha0bdd17f;
    ram_cell[   19485] = 32'ha23a1f9b;
    ram_cell[   19486] = 32'h7c8ad013;
    ram_cell[   19487] = 32'hdc954fe5;
    ram_cell[   19488] = 32'hb2ee2ba4;
    ram_cell[   19489] = 32'hd236921c;
    ram_cell[   19490] = 32'h553d701e;
    ram_cell[   19491] = 32'h24fc6df1;
    ram_cell[   19492] = 32'h0aaf9fdd;
    ram_cell[   19493] = 32'h2eba442d;
    ram_cell[   19494] = 32'hfc5674bb;
    ram_cell[   19495] = 32'h3b88a69a;
    ram_cell[   19496] = 32'h8ab85678;
    ram_cell[   19497] = 32'hd0c128d2;
    ram_cell[   19498] = 32'hd0f82ca9;
    ram_cell[   19499] = 32'h223bf61f;
    ram_cell[   19500] = 32'h57d91173;
    ram_cell[   19501] = 32'hdf56951f;
    ram_cell[   19502] = 32'hcf3a5b87;
    ram_cell[   19503] = 32'h69280bd3;
    ram_cell[   19504] = 32'h8966dae4;
    ram_cell[   19505] = 32'hbe65d86f;
    ram_cell[   19506] = 32'hfd11e1f2;
    ram_cell[   19507] = 32'h56452302;
    ram_cell[   19508] = 32'hd8245759;
    ram_cell[   19509] = 32'h5032d897;
    ram_cell[   19510] = 32'h5b0ef59f;
    ram_cell[   19511] = 32'h29095727;
    ram_cell[   19512] = 32'he5d7b54f;
    ram_cell[   19513] = 32'h9acecfca;
    ram_cell[   19514] = 32'hcb93b4e3;
    ram_cell[   19515] = 32'hc787077f;
    ram_cell[   19516] = 32'h82e20e73;
    ram_cell[   19517] = 32'h5621ceb7;
    ram_cell[   19518] = 32'h99cec752;
    ram_cell[   19519] = 32'h1a4a06aa;
    ram_cell[   19520] = 32'h2835dbad;
    ram_cell[   19521] = 32'h53c0210a;
    ram_cell[   19522] = 32'h03607109;
    ram_cell[   19523] = 32'hbc94c464;
    ram_cell[   19524] = 32'hdac5a1a1;
    ram_cell[   19525] = 32'h0d471509;
    ram_cell[   19526] = 32'h951e47ac;
    ram_cell[   19527] = 32'hb8cb0bff;
    ram_cell[   19528] = 32'ha441a7f3;
    ram_cell[   19529] = 32'h8880b1f5;
    ram_cell[   19530] = 32'h1641f769;
    ram_cell[   19531] = 32'hbd9be53d;
    ram_cell[   19532] = 32'hf23087ef;
    ram_cell[   19533] = 32'h907d789d;
    ram_cell[   19534] = 32'hf00b3fd6;
    ram_cell[   19535] = 32'h48f0c8c6;
    ram_cell[   19536] = 32'h17e4c802;
    ram_cell[   19537] = 32'h114d5fab;
    ram_cell[   19538] = 32'h50b38087;
    ram_cell[   19539] = 32'h41ccecfa;
    ram_cell[   19540] = 32'hcc803fc1;
    ram_cell[   19541] = 32'h3d33fe28;
    ram_cell[   19542] = 32'h4923794d;
    ram_cell[   19543] = 32'hda560467;
    ram_cell[   19544] = 32'hb47732c1;
    ram_cell[   19545] = 32'hf7a70326;
    ram_cell[   19546] = 32'ha1ac60f6;
    ram_cell[   19547] = 32'h431e4b35;
    ram_cell[   19548] = 32'hfefcaf7c;
    ram_cell[   19549] = 32'hdfa9addc;
    ram_cell[   19550] = 32'h41ee4824;
    ram_cell[   19551] = 32'hb5bc5255;
    ram_cell[   19552] = 32'h258d906e;
    ram_cell[   19553] = 32'h4a6da90f;
    ram_cell[   19554] = 32'h68dc01c2;
    ram_cell[   19555] = 32'hfc377ca0;
    ram_cell[   19556] = 32'h4029e833;
    ram_cell[   19557] = 32'h8f4780cf;
    ram_cell[   19558] = 32'h817d890f;
    ram_cell[   19559] = 32'h28a9fd7f;
    ram_cell[   19560] = 32'hb14b8833;
    ram_cell[   19561] = 32'hca53fd8a;
    ram_cell[   19562] = 32'hbd18d7f8;
    ram_cell[   19563] = 32'ha5383e1e;
    ram_cell[   19564] = 32'hadebade6;
    ram_cell[   19565] = 32'hc95f7d13;
    ram_cell[   19566] = 32'hccb8e2c2;
    ram_cell[   19567] = 32'h01426aa8;
    ram_cell[   19568] = 32'h43f1dd4a;
    ram_cell[   19569] = 32'h73e11add;
    ram_cell[   19570] = 32'hd9497e9a;
    ram_cell[   19571] = 32'h4665fbcb;
    ram_cell[   19572] = 32'hcb8aeafc;
    ram_cell[   19573] = 32'hc8a7864a;
    ram_cell[   19574] = 32'h350778ce;
    ram_cell[   19575] = 32'h0cc4bd99;
    ram_cell[   19576] = 32'h7c0651b1;
    ram_cell[   19577] = 32'hb26b83f5;
    ram_cell[   19578] = 32'h3bd88fb8;
    ram_cell[   19579] = 32'h4b25b84e;
    ram_cell[   19580] = 32'hbbff5775;
    ram_cell[   19581] = 32'h95281cf1;
    ram_cell[   19582] = 32'h4d49301c;
    ram_cell[   19583] = 32'hf152ecd8;
    ram_cell[   19584] = 32'h62fdd866;
    ram_cell[   19585] = 32'h9e66bbfc;
    ram_cell[   19586] = 32'hdfd6b080;
    ram_cell[   19587] = 32'h49a7d6e4;
    ram_cell[   19588] = 32'hd2e77391;
    ram_cell[   19589] = 32'h4fcf6613;
    ram_cell[   19590] = 32'hae7dc683;
    ram_cell[   19591] = 32'hcc2e6586;
    ram_cell[   19592] = 32'ha25670e2;
    ram_cell[   19593] = 32'h2423a5fa;
    ram_cell[   19594] = 32'ha5d889c4;
    ram_cell[   19595] = 32'h15193549;
    ram_cell[   19596] = 32'hff9b22d1;
    ram_cell[   19597] = 32'h4b5f74fa;
    ram_cell[   19598] = 32'h21391122;
    ram_cell[   19599] = 32'hecd81c88;
    ram_cell[   19600] = 32'h587ee2d1;
    ram_cell[   19601] = 32'h961742bb;
    ram_cell[   19602] = 32'hb4ff4db2;
    ram_cell[   19603] = 32'hc67fbae3;
    ram_cell[   19604] = 32'hb279d324;
    ram_cell[   19605] = 32'h4ae98ccd;
    ram_cell[   19606] = 32'h897fc95c;
    ram_cell[   19607] = 32'hc4a139cf;
    ram_cell[   19608] = 32'h5ce09702;
    ram_cell[   19609] = 32'hd0f218fd;
    ram_cell[   19610] = 32'hf4fc9a84;
    ram_cell[   19611] = 32'h76e519fe;
    ram_cell[   19612] = 32'h64d6dba3;
    ram_cell[   19613] = 32'hbe9075f6;
    ram_cell[   19614] = 32'h76c1aed1;
    ram_cell[   19615] = 32'h41379a9f;
    ram_cell[   19616] = 32'hb5f984a3;
    ram_cell[   19617] = 32'h3e11a88e;
    ram_cell[   19618] = 32'h9dfeb758;
    ram_cell[   19619] = 32'hd51fc9b5;
    ram_cell[   19620] = 32'h64b1f4b7;
    ram_cell[   19621] = 32'h574f7cef;
    ram_cell[   19622] = 32'h69b7dfc8;
    ram_cell[   19623] = 32'h7845ec75;
    ram_cell[   19624] = 32'hdf85d1d1;
    ram_cell[   19625] = 32'hecf6737b;
    ram_cell[   19626] = 32'h7529a37f;
    ram_cell[   19627] = 32'ha16d7e2a;
    ram_cell[   19628] = 32'h31ea795a;
    ram_cell[   19629] = 32'h2d4ad8e4;
    ram_cell[   19630] = 32'h4a55dd7a;
    ram_cell[   19631] = 32'h83cd8ed6;
    ram_cell[   19632] = 32'hd5f35b16;
    ram_cell[   19633] = 32'h7ae874c2;
    ram_cell[   19634] = 32'hcfdd30ed;
    ram_cell[   19635] = 32'hbd73ee7b;
    ram_cell[   19636] = 32'h94de7cc2;
    ram_cell[   19637] = 32'h42dcb8ec;
    ram_cell[   19638] = 32'he76c2e8a;
    ram_cell[   19639] = 32'hf0c90af9;
    ram_cell[   19640] = 32'h387b5b75;
    ram_cell[   19641] = 32'ha3024085;
    ram_cell[   19642] = 32'h28819673;
    ram_cell[   19643] = 32'he267ae2e;
    ram_cell[   19644] = 32'h86af961c;
    ram_cell[   19645] = 32'hd70983af;
    ram_cell[   19646] = 32'h54b7d805;
    ram_cell[   19647] = 32'h3091f0f3;
    ram_cell[   19648] = 32'h638922a4;
    ram_cell[   19649] = 32'h12869aa3;
    ram_cell[   19650] = 32'h28fc22dc;
    ram_cell[   19651] = 32'h6e425847;
    ram_cell[   19652] = 32'h10017185;
    ram_cell[   19653] = 32'h0db82199;
    ram_cell[   19654] = 32'h3715a535;
    ram_cell[   19655] = 32'hdea170f2;
    ram_cell[   19656] = 32'h95cd6210;
    ram_cell[   19657] = 32'h373a60f6;
    ram_cell[   19658] = 32'he7837017;
    ram_cell[   19659] = 32'h0333a8da;
    ram_cell[   19660] = 32'h43d4c77f;
    ram_cell[   19661] = 32'hc0021425;
    ram_cell[   19662] = 32'hb1d4c2de;
    ram_cell[   19663] = 32'hff7d44a0;
    ram_cell[   19664] = 32'h6d3a91f3;
    ram_cell[   19665] = 32'h4d1a5b46;
    ram_cell[   19666] = 32'h015f9c8b;
    ram_cell[   19667] = 32'h515d7177;
    ram_cell[   19668] = 32'hd790cdce;
    ram_cell[   19669] = 32'h797ce144;
    ram_cell[   19670] = 32'h65373d56;
    ram_cell[   19671] = 32'hb6ddd0bb;
    ram_cell[   19672] = 32'hbf60f103;
    ram_cell[   19673] = 32'h0d9b11b2;
    ram_cell[   19674] = 32'hdf9694b6;
    ram_cell[   19675] = 32'hce2d7c37;
    ram_cell[   19676] = 32'hea908df0;
    ram_cell[   19677] = 32'h06818be8;
    ram_cell[   19678] = 32'h18b6416d;
    ram_cell[   19679] = 32'h55699793;
    ram_cell[   19680] = 32'h082eec74;
    ram_cell[   19681] = 32'he311105d;
    ram_cell[   19682] = 32'h9bc50420;
    ram_cell[   19683] = 32'h07a2fae7;
    ram_cell[   19684] = 32'h7576c0be;
    ram_cell[   19685] = 32'hcb3cc8ed;
    ram_cell[   19686] = 32'h0a5a2cbd;
    ram_cell[   19687] = 32'h2d66e702;
    ram_cell[   19688] = 32'hdc5b3db1;
    ram_cell[   19689] = 32'hcc6a641b;
    ram_cell[   19690] = 32'hd79a87d1;
    ram_cell[   19691] = 32'h7d553702;
    ram_cell[   19692] = 32'h4a2f42cf;
    ram_cell[   19693] = 32'h6d53b3cc;
    ram_cell[   19694] = 32'hdd9e17f8;
    ram_cell[   19695] = 32'he849592f;
    ram_cell[   19696] = 32'hf98e3c9b;
    ram_cell[   19697] = 32'h5b77cc38;
    ram_cell[   19698] = 32'h52aa5c20;
    ram_cell[   19699] = 32'h04084bd9;
    ram_cell[   19700] = 32'h2cee39a6;
    ram_cell[   19701] = 32'h15c0403e;
    ram_cell[   19702] = 32'h990075c4;
    ram_cell[   19703] = 32'h0fe00d14;
    ram_cell[   19704] = 32'ha4023a94;
    ram_cell[   19705] = 32'h6ce07b05;
    ram_cell[   19706] = 32'h3cb3fb80;
    ram_cell[   19707] = 32'h33351d8c;
    ram_cell[   19708] = 32'h659e5e55;
    ram_cell[   19709] = 32'hdadf65f5;
    ram_cell[   19710] = 32'hca48b0e3;
    ram_cell[   19711] = 32'h0a9d092c;
    ram_cell[   19712] = 32'hab3d687d;
    ram_cell[   19713] = 32'h60b79c7c;
    ram_cell[   19714] = 32'h85e49fc6;
    ram_cell[   19715] = 32'h1eb02a86;
    ram_cell[   19716] = 32'h70cac46b;
    ram_cell[   19717] = 32'h31e28dd8;
    ram_cell[   19718] = 32'hb797b87d;
    ram_cell[   19719] = 32'h262e9a3a;
    ram_cell[   19720] = 32'ha7e86807;
    ram_cell[   19721] = 32'hcad92fc7;
    ram_cell[   19722] = 32'hbb8f00cd;
    ram_cell[   19723] = 32'h2d8ba74b;
    ram_cell[   19724] = 32'hc2a4a48a;
    ram_cell[   19725] = 32'hc9661346;
    ram_cell[   19726] = 32'hb55b0034;
    ram_cell[   19727] = 32'h58e9efa3;
    ram_cell[   19728] = 32'ha0159d8c;
    ram_cell[   19729] = 32'hb46d6d88;
    ram_cell[   19730] = 32'h08cd59e9;
    ram_cell[   19731] = 32'h9f159225;
    ram_cell[   19732] = 32'he5c792a5;
    ram_cell[   19733] = 32'hc92d8086;
    ram_cell[   19734] = 32'h78ad945f;
    ram_cell[   19735] = 32'h3c6536d1;
    ram_cell[   19736] = 32'hcaf6ee41;
    ram_cell[   19737] = 32'ha0af4178;
    ram_cell[   19738] = 32'h79b9570a;
    ram_cell[   19739] = 32'haf7beb9d;
    ram_cell[   19740] = 32'h9930b010;
    ram_cell[   19741] = 32'h4f9fd5d8;
    ram_cell[   19742] = 32'h4fb15a4c;
    ram_cell[   19743] = 32'h4af81ac7;
    ram_cell[   19744] = 32'h0eb7488c;
    ram_cell[   19745] = 32'h77b2905e;
    ram_cell[   19746] = 32'h6df19a08;
    ram_cell[   19747] = 32'he586bbca;
    ram_cell[   19748] = 32'h123a9c69;
    ram_cell[   19749] = 32'hbb06cc29;
    ram_cell[   19750] = 32'h0e9f0789;
    ram_cell[   19751] = 32'h94b80295;
    ram_cell[   19752] = 32'h16f725f9;
    ram_cell[   19753] = 32'h6e9fe7e3;
    ram_cell[   19754] = 32'h04dde9c3;
    ram_cell[   19755] = 32'h8f27e353;
    ram_cell[   19756] = 32'he3d7a091;
    ram_cell[   19757] = 32'h32e36237;
    ram_cell[   19758] = 32'h16c654a7;
    ram_cell[   19759] = 32'h40746e5e;
    ram_cell[   19760] = 32'hedf6dab5;
    ram_cell[   19761] = 32'heb2bbea2;
    ram_cell[   19762] = 32'h5072a0a6;
    ram_cell[   19763] = 32'hf46b837b;
    ram_cell[   19764] = 32'h2273f67a;
    ram_cell[   19765] = 32'hba0b0f37;
    ram_cell[   19766] = 32'hc3db182c;
    ram_cell[   19767] = 32'h671b5899;
    ram_cell[   19768] = 32'h1dfda285;
    ram_cell[   19769] = 32'hee5e1845;
    ram_cell[   19770] = 32'h75f7309f;
    ram_cell[   19771] = 32'h41d36bcb;
    ram_cell[   19772] = 32'hbeb6a4e8;
    ram_cell[   19773] = 32'h3ea53ddf;
    ram_cell[   19774] = 32'h387c6c66;
    ram_cell[   19775] = 32'h60377336;
    ram_cell[   19776] = 32'h99f981d0;
    ram_cell[   19777] = 32'h1780d838;
    ram_cell[   19778] = 32'hdab21430;
    ram_cell[   19779] = 32'hb86290b2;
    ram_cell[   19780] = 32'he98b2bc6;
    ram_cell[   19781] = 32'h36d25fbe;
    ram_cell[   19782] = 32'h2464533a;
    ram_cell[   19783] = 32'h2bf1cea8;
    ram_cell[   19784] = 32'h7382d9ff;
    ram_cell[   19785] = 32'ha890e0da;
    ram_cell[   19786] = 32'h4331a8d6;
    ram_cell[   19787] = 32'hfd16f46c;
    ram_cell[   19788] = 32'h76e7decb;
    ram_cell[   19789] = 32'h93fd8ad2;
    ram_cell[   19790] = 32'hca60019e;
    ram_cell[   19791] = 32'h97f40d2e;
    ram_cell[   19792] = 32'h0fe34c76;
    ram_cell[   19793] = 32'hb88c9da5;
    ram_cell[   19794] = 32'hcf411da0;
    ram_cell[   19795] = 32'hbe48d4c3;
    ram_cell[   19796] = 32'h1b3f3219;
    ram_cell[   19797] = 32'h0caa40f0;
    ram_cell[   19798] = 32'hb29ba940;
    ram_cell[   19799] = 32'h47f6fc40;
    ram_cell[   19800] = 32'he90d4695;
    ram_cell[   19801] = 32'h09177aed;
    ram_cell[   19802] = 32'h62dfc761;
    ram_cell[   19803] = 32'h023152c4;
    ram_cell[   19804] = 32'h7097910b;
    ram_cell[   19805] = 32'hf71fc442;
    ram_cell[   19806] = 32'h79efccfe;
    ram_cell[   19807] = 32'h9560c17b;
    ram_cell[   19808] = 32'h4d33b49e;
    ram_cell[   19809] = 32'hbf900a37;
    ram_cell[   19810] = 32'h4da425a4;
    ram_cell[   19811] = 32'hb843d769;
    ram_cell[   19812] = 32'hfe33de32;
    ram_cell[   19813] = 32'ha403b1f1;
    ram_cell[   19814] = 32'h33529d83;
    ram_cell[   19815] = 32'h3f2540f1;
    ram_cell[   19816] = 32'hc968f711;
    ram_cell[   19817] = 32'h4c2fae40;
    ram_cell[   19818] = 32'h0edb35b8;
    ram_cell[   19819] = 32'h66cd3dce;
    ram_cell[   19820] = 32'h99185a36;
    ram_cell[   19821] = 32'hf7ebe502;
    ram_cell[   19822] = 32'heedadf3f;
    ram_cell[   19823] = 32'h705f1539;
    ram_cell[   19824] = 32'ha48c8a71;
    ram_cell[   19825] = 32'h2865bbe1;
    ram_cell[   19826] = 32'hcc0edbf0;
    ram_cell[   19827] = 32'h27994990;
    ram_cell[   19828] = 32'had6a2f25;
    ram_cell[   19829] = 32'h7e7163fb;
    ram_cell[   19830] = 32'h21c529d9;
    ram_cell[   19831] = 32'hb08afd03;
    ram_cell[   19832] = 32'h1fe9aabc;
    ram_cell[   19833] = 32'ha3977e8b;
    ram_cell[   19834] = 32'h7ae2844f;
    ram_cell[   19835] = 32'h554e3495;
    ram_cell[   19836] = 32'h642ee238;
    ram_cell[   19837] = 32'hdd258d7d;
    ram_cell[   19838] = 32'hcde65099;
    ram_cell[   19839] = 32'hdd633ece;
    ram_cell[   19840] = 32'h124ccec0;
    ram_cell[   19841] = 32'hfab7c51a;
    ram_cell[   19842] = 32'hf262bdc0;
    ram_cell[   19843] = 32'ha96a789a;
    ram_cell[   19844] = 32'h53dc93c9;
    ram_cell[   19845] = 32'h0b7df142;
    ram_cell[   19846] = 32'h6eba3911;
    ram_cell[   19847] = 32'h22bb619c;
    ram_cell[   19848] = 32'h5b558b4b;
    ram_cell[   19849] = 32'hce4ad965;
    ram_cell[   19850] = 32'h632ba526;
    ram_cell[   19851] = 32'h57dc58b6;
    ram_cell[   19852] = 32'he7fa5144;
    ram_cell[   19853] = 32'hec4e0e50;
    ram_cell[   19854] = 32'hfb8e1548;
    ram_cell[   19855] = 32'h86dbe026;
    ram_cell[   19856] = 32'h36cc0abc;
    ram_cell[   19857] = 32'h593e9f68;
    ram_cell[   19858] = 32'h2ebee031;
    ram_cell[   19859] = 32'hea97fdc4;
    ram_cell[   19860] = 32'h8bc612ce;
    ram_cell[   19861] = 32'h9c763753;
    ram_cell[   19862] = 32'h962784b9;
    ram_cell[   19863] = 32'h935dc451;
    ram_cell[   19864] = 32'h4ed1f2ee;
    ram_cell[   19865] = 32'h4f2c2690;
    ram_cell[   19866] = 32'h740ce1fc;
    ram_cell[   19867] = 32'h3588205d;
    ram_cell[   19868] = 32'h40827c08;
    ram_cell[   19869] = 32'h1c7004d9;
    ram_cell[   19870] = 32'h3a84bef7;
    ram_cell[   19871] = 32'hc2a17778;
    ram_cell[   19872] = 32'hadab138f;
    ram_cell[   19873] = 32'h5e0386c3;
    ram_cell[   19874] = 32'hf0faff9a;
    ram_cell[   19875] = 32'h8af95bb0;
    ram_cell[   19876] = 32'h292e818a;
    ram_cell[   19877] = 32'hb102b501;
    ram_cell[   19878] = 32'ha36a0f4a;
    ram_cell[   19879] = 32'h5bcefae2;
    ram_cell[   19880] = 32'h14697304;
    ram_cell[   19881] = 32'h2976b01c;
    ram_cell[   19882] = 32'hd9b1d1d7;
    ram_cell[   19883] = 32'hf0bf2b79;
    ram_cell[   19884] = 32'h803097b3;
    ram_cell[   19885] = 32'h7595d532;
    ram_cell[   19886] = 32'h62ef0240;
    ram_cell[   19887] = 32'ha3378a0f;
    ram_cell[   19888] = 32'h6e981f0d;
    ram_cell[   19889] = 32'hae3702ec;
    ram_cell[   19890] = 32'hf69f5e5d;
    ram_cell[   19891] = 32'h1e66df5d;
    ram_cell[   19892] = 32'h93592c2f;
    ram_cell[   19893] = 32'h59a1131c;
    ram_cell[   19894] = 32'hd6b29dbc;
    ram_cell[   19895] = 32'h48556992;
    ram_cell[   19896] = 32'hd3e4bbb3;
    ram_cell[   19897] = 32'h704fc3c9;
    ram_cell[   19898] = 32'h720cffb3;
    ram_cell[   19899] = 32'h6d8be7ee;
    ram_cell[   19900] = 32'h56ecbb0f;
    ram_cell[   19901] = 32'h22220f59;
    ram_cell[   19902] = 32'h0663d9b7;
    ram_cell[   19903] = 32'h2c454d12;
    ram_cell[   19904] = 32'he6ffea5c;
    ram_cell[   19905] = 32'hee6b088a;
    ram_cell[   19906] = 32'h8b2dfceb;
    ram_cell[   19907] = 32'hf77ef455;
    ram_cell[   19908] = 32'hbf8280ac;
    ram_cell[   19909] = 32'had4915a6;
    ram_cell[   19910] = 32'hd4136cf9;
    ram_cell[   19911] = 32'hb0b6d5f3;
    ram_cell[   19912] = 32'he1736ca3;
    ram_cell[   19913] = 32'h042f6275;
    ram_cell[   19914] = 32'h812b9e6c;
    ram_cell[   19915] = 32'h049de5ab;
    ram_cell[   19916] = 32'h0f79e4c2;
    ram_cell[   19917] = 32'h524b31da;
    ram_cell[   19918] = 32'h240f57e3;
    ram_cell[   19919] = 32'hf983cd2d;
    ram_cell[   19920] = 32'h466bda79;
    ram_cell[   19921] = 32'h44818888;
    ram_cell[   19922] = 32'h09f0a9d8;
    ram_cell[   19923] = 32'h06723345;
    ram_cell[   19924] = 32'hd068324c;
    ram_cell[   19925] = 32'h1f3a8909;
    ram_cell[   19926] = 32'hfb6c4966;
    ram_cell[   19927] = 32'h070c9364;
    ram_cell[   19928] = 32'h5fda8a8c;
    ram_cell[   19929] = 32'hcf7073f8;
    ram_cell[   19930] = 32'h4be87825;
    ram_cell[   19931] = 32'h852f2b65;
    ram_cell[   19932] = 32'h4837d60a;
    ram_cell[   19933] = 32'h830f209c;
    ram_cell[   19934] = 32'hd8251bc5;
    ram_cell[   19935] = 32'hf9a3e3ba;
    ram_cell[   19936] = 32'h3e753d97;
    ram_cell[   19937] = 32'hbfbbea0e;
    ram_cell[   19938] = 32'h596beeae;
    ram_cell[   19939] = 32'h8088603f;
    ram_cell[   19940] = 32'h35124ed6;
    ram_cell[   19941] = 32'hc7d766ea;
    ram_cell[   19942] = 32'hb1513eed;
    ram_cell[   19943] = 32'h2d62d4ff;
    ram_cell[   19944] = 32'h5d2772e1;
    ram_cell[   19945] = 32'he6b55a34;
    ram_cell[   19946] = 32'h52f5ee92;
    ram_cell[   19947] = 32'hbf004ebe;
    ram_cell[   19948] = 32'hfa1ca6cf;
    ram_cell[   19949] = 32'hc293aa40;
    ram_cell[   19950] = 32'h97c8e879;
    ram_cell[   19951] = 32'hb509940c;
    ram_cell[   19952] = 32'h26630145;
    ram_cell[   19953] = 32'h40e8b497;
    ram_cell[   19954] = 32'h1a13efed;
    ram_cell[   19955] = 32'h2b124891;
    ram_cell[   19956] = 32'hcc21127d;
    ram_cell[   19957] = 32'h17f4f644;
    ram_cell[   19958] = 32'hd30b8e40;
    ram_cell[   19959] = 32'h9a7e0a98;
    ram_cell[   19960] = 32'h605ea7a2;
    ram_cell[   19961] = 32'h635bbf1d;
    ram_cell[   19962] = 32'hf3270936;
    ram_cell[   19963] = 32'had1bd93d;
    ram_cell[   19964] = 32'h95d77bca;
    ram_cell[   19965] = 32'he319abff;
    ram_cell[   19966] = 32'hce1cb2c4;
    ram_cell[   19967] = 32'h1252c3ac;
    ram_cell[   19968] = 32'hf3796dc1;
    ram_cell[   19969] = 32'h61d88d92;
    ram_cell[   19970] = 32'h1d8185f8;
    ram_cell[   19971] = 32'h75582a43;
    ram_cell[   19972] = 32'hc8606a37;
    ram_cell[   19973] = 32'h33fdc905;
    ram_cell[   19974] = 32'h4946c768;
    ram_cell[   19975] = 32'h8d504165;
    ram_cell[   19976] = 32'h162fb1d8;
    ram_cell[   19977] = 32'ha9342527;
    ram_cell[   19978] = 32'h189da4a1;
    ram_cell[   19979] = 32'h97429150;
    ram_cell[   19980] = 32'hfae444e6;
    ram_cell[   19981] = 32'h91d875e7;
    ram_cell[   19982] = 32'hc6dc0b54;
    ram_cell[   19983] = 32'h35c6e591;
    ram_cell[   19984] = 32'h6c736591;
    ram_cell[   19985] = 32'h27f47847;
    ram_cell[   19986] = 32'h9d122124;
    ram_cell[   19987] = 32'h2f68d088;
    ram_cell[   19988] = 32'h66b962a0;
    ram_cell[   19989] = 32'h9d354c97;
    ram_cell[   19990] = 32'h39c35180;
    ram_cell[   19991] = 32'h708ef6fb;
    ram_cell[   19992] = 32'h3cf9e0fe;
    ram_cell[   19993] = 32'h942ebcc6;
    ram_cell[   19994] = 32'hc7c1bbbf;
    ram_cell[   19995] = 32'h4d1157ae;
    ram_cell[   19996] = 32'hf7b7258b;
    ram_cell[   19997] = 32'he64def66;
    ram_cell[   19998] = 32'hfa1cf5ca;
    ram_cell[   19999] = 32'h6a092647;
    ram_cell[   20000] = 32'hde92a14f;
    ram_cell[   20001] = 32'h894ebc94;
    ram_cell[   20002] = 32'h4bde626b;
    ram_cell[   20003] = 32'h09b4028d;
    ram_cell[   20004] = 32'h40bc6314;
    ram_cell[   20005] = 32'h946517b8;
    ram_cell[   20006] = 32'h4f68bde3;
    ram_cell[   20007] = 32'h89ec439f;
    ram_cell[   20008] = 32'h6054bd31;
    ram_cell[   20009] = 32'hafecf1bd;
    ram_cell[   20010] = 32'he38488d6;
    ram_cell[   20011] = 32'h0f3692de;
    ram_cell[   20012] = 32'hb9092d55;
    ram_cell[   20013] = 32'hfec24a02;
    ram_cell[   20014] = 32'h26838a1d;
    ram_cell[   20015] = 32'h472db4ce;
    ram_cell[   20016] = 32'h3faee942;
    ram_cell[   20017] = 32'h37555c28;
    ram_cell[   20018] = 32'h807f030e;
    ram_cell[   20019] = 32'h5b0a719a;
    ram_cell[   20020] = 32'hbda0122d;
    ram_cell[   20021] = 32'hb8a9a57a;
    ram_cell[   20022] = 32'hf5cd6612;
    ram_cell[   20023] = 32'h91c4465c;
    ram_cell[   20024] = 32'hdc8371be;
    ram_cell[   20025] = 32'h6f270cd4;
    ram_cell[   20026] = 32'h29bcb2c7;
    ram_cell[   20027] = 32'hcce5ff81;
    ram_cell[   20028] = 32'hf41bc19a;
    ram_cell[   20029] = 32'h42265bd5;
    ram_cell[   20030] = 32'hc081ead2;
    ram_cell[   20031] = 32'h17c46a97;
    ram_cell[   20032] = 32'h660e558a;
    ram_cell[   20033] = 32'haa597b3d;
    ram_cell[   20034] = 32'h74af04ee;
    ram_cell[   20035] = 32'h533d8c09;
    ram_cell[   20036] = 32'h7cce5cfd;
    ram_cell[   20037] = 32'h8f0c6e85;
    ram_cell[   20038] = 32'he9dbfdd1;
    ram_cell[   20039] = 32'hf86b2546;
    ram_cell[   20040] = 32'h1ff1c789;
    ram_cell[   20041] = 32'h5acd5fea;
    ram_cell[   20042] = 32'h63c33f6a;
    ram_cell[   20043] = 32'hc25f17b1;
    ram_cell[   20044] = 32'h53d01e3c;
    ram_cell[   20045] = 32'h0dcfb8a6;
    ram_cell[   20046] = 32'h3208bea6;
    ram_cell[   20047] = 32'h31dfcb6f;
    ram_cell[   20048] = 32'hce4407a5;
    ram_cell[   20049] = 32'ha9e194cc;
    ram_cell[   20050] = 32'h6e607097;
    ram_cell[   20051] = 32'h2a54b0b0;
    ram_cell[   20052] = 32'hf81ec3fd;
    ram_cell[   20053] = 32'h6a9419b0;
    ram_cell[   20054] = 32'hd5355017;
    ram_cell[   20055] = 32'ha947117e;
    ram_cell[   20056] = 32'h7aa260c0;
    ram_cell[   20057] = 32'hf7314a08;
    ram_cell[   20058] = 32'h12a418c4;
    ram_cell[   20059] = 32'h6c48e1fd;
    ram_cell[   20060] = 32'h920e7394;
    ram_cell[   20061] = 32'h2f73a9bc;
    ram_cell[   20062] = 32'hb9190cb8;
    ram_cell[   20063] = 32'h7079ac33;
    ram_cell[   20064] = 32'h55200173;
    ram_cell[   20065] = 32'h9ff7f35c;
    ram_cell[   20066] = 32'ha2c04d9f;
    ram_cell[   20067] = 32'h4235011c;
    ram_cell[   20068] = 32'h5b09dd39;
    ram_cell[   20069] = 32'h4bea9488;
    ram_cell[   20070] = 32'h4eab80ff;
    ram_cell[   20071] = 32'hfbae2a0f;
    ram_cell[   20072] = 32'hc8253286;
    ram_cell[   20073] = 32'h0464aae5;
    ram_cell[   20074] = 32'hd6c94396;
    ram_cell[   20075] = 32'h556e1401;
    ram_cell[   20076] = 32'h4efa6b36;
    ram_cell[   20077] = 32'he62bc093;
    ram_cell[   20078] = 32'h532fcd16;
    ram_cell[   20079] = 32'h817b4ce8;
    ram_cell[   20080] = 32'h70a1bfb5;
    ram_cell[   20081] = 32'h2b5ad045;
    ram_cell[   20082] = 32'h8857b24b;
    ram_cell[   20083] = 32'hd0d57ced;
    ram_cell[   20084] = 32'h42670e32;
    ram_cell[   20085] = 32'h93625cf0;
    ram_cell[   20086] = 32'h2015c72b;
    ram_cell[   20087] = 32'h38a06f1a;
    ram_cell[   20088] = 32'hd9df8c35;
    ram_cell[   20089] = 32'h895d4117;
    ram_cell[   20090] = 32'h410555a9;
    ram_cell[   20091] = 32'h3e32d9cc;
    ram_cell[   20092] = 32'hf0c58702;
    ram_cell[   20093] = 32'ha4cfe714;
    ram_cell[   20094] = 32'h0fc9ceb7;
    ram_cell[   20095] = 32'ha3001dfa;
    ram_cell[   20096] = 32'hb9f7af35;
    ram_cell[   20097] = 32'h40bd0f91;
    ram_cell[   20098] = 32'he70ed38f;
    ram_cell[   20099] = 32'h8c8c3b7a;
    ram_cell[   20100] = 32'hed327c5a;
    ram_cell[   20101] = 32'h8587ef28;
    ram_cell[   20102] = 32'h01395091;
    ram_cell[   20103] = 32'hc288969e;
    ram_cell[   20104] = 32'h13ab2d58;
    ram_cell[   20105] = 32'h2cf2c22f;
    ram_cell[   20106] = 32'h5b0f240f;
    ram_cell[   20107] = 32'h811fd874;
    ram_cell[   20108] = 32'h7d2c147b;
    ram_cell[   20109] = 32'hfd4a3453;
    ram_cell[   20110] = 32'hfd573d3d;
    ram_cell[   20111] = 32'h95f4fc43;
    ram_cell[   20112] = 32'hd1b3faa2;
    ram_cell[   20113] = 32'h3058616d;
    ram_cell[   20114] = 32'hfe3d8757;
    ram_cell[   20115] = 32'h6f970b23;
    ram_cell[   20116] = 32'h979b7279;
    ram_cell[   20117] = 32'hcde9204b;
    ram_cell[   20118] = 32'h99f70432;
    ram_cell[   20119] = 32'h679cbc01;
    ram_cell[   20120] = 32'hf70b00e5;
    ram_cell[   20121] = 32'h8a684c95;
    ram_cell[   20122] = 32'he49fdde6;
    ram_cell[   20123] = 32'h8772733e;
    ram_cell[   20124] = 32'hfdeb2f03;
    ram_cell[   20125] = 32'h5a636154;
    ram_cell[   20126] = 32'h0ce34af0;
    ram_cell[   20127] = 32'hd8f9eae4;
    ram_cell[   20128] = 32'hab72aa0c;
    ram_cell[   20129] = 32'h225dbf6e;
    ram_cell[   20130] = 32'h3e04be8c;
    ram_cell[   20131] = 32'h3bb03b66;
    ram_cell[   20132] = 32'h48435b7d;
    ram_cell[   20133] = 32'h4bab2121;
    ram_cell[   20134] = 32'h2c4f99cb;
    ram_cell[   20135] = 32'hc3ddb665;
    ram_cell[   20136] = 32'hb450d24e;
    ram_cell[   20137] = 32'h2bac8f6c;
    ram_cell[   20138] = 32'h5d04c26d;
    ram_cell[   20139] = 32'h96476a1a;
    ram_cell[   20140] = 32'ha2266b9e;
    ram_cell[   20141] = 32'h79a07861;
    ram_cell[   20142] = 32'h48156432;
    ram_cell[   20143] = 32'h1a75f247;
    ram_cell[   20144] = 32'hb98c291d;
    ram_cell[   20145] = 32'h159752b8;
    ram_cell[   20146] = 32'h0bd7d83a;
    ram_cell[   20147] = 32'hdbbb5928;
    ram_cell[   20148] = 32'h9a12c337;
    ram_cell[   20149] = 32'hc8885252;
    ram_cell[   20150] = 32'hb373ac96;
    ram_cell[   20151] = 32'h391025b9;
    ram_cell[   20152] = 32'h855f6030;
    ram_cell[   20153] = 32'h6f36b27b;
    ram_cell[   20154] = 32'h6ee56d60;
    ram_cell[   20155] = 32'hf9948a53;
    ram_cell[   20156] = 32'h8baa3d3b;
    ram_cell[   20157] = 32'hf9ab3a4d;
    ram_cell[   20158] = 32'h7f961249;
    ram_cell[   20159] = 32'hdac5cf6f;
    ram_cell[   20160] = 32'h29036302;
    ram_cell[   20161] = 32'h0228bea6;
    ram_cell[   20162] = 32'h799719c3;
    ram_cell[   20163] = 32'hdfb318d0;
    ram_cell[   20164] = 32'h427b83cb;
    ram_cell[   20165] = 32'hb40c98ec;
    ram_cell[   20166] = 32'hff2c6308;
    ram_cell[   20167] = 32'h6f4f3330;
    ram_cell[   20168] = 32'hf39e8f69;
    ram_cell[   20169] = 32'h0503e151;
    ram_cell[   20170] = 32'h05a027e4;
    ram_cell[   20171] = 32'he207bc0a;
    ram_cell[   20172] = 32'hd670d3bd;
    ram_cell[   20173] = 32'h61288e7f;
    ram_cell[   20174] = 32'hd8b09886;
    ram_cell[   20175] = 32'h345311ba;
    ram_cell[   20176] = 32'h414a27c2;
    ram_cell[   20177] = 32'h8c85670b;
    ram_cell[   20178] = 32'ha20b3b26;
    ram_cell[   20179] = 32'hd964643b;
    ram_cell[   20180] = 32'hdf8344e5;
    ram_cell[   20181] = 32'h03692216;
    ram_cell[   20182] = 32'h8787cbfb;
    ram_cell[   20183] = 32'ha941e9fb;
    ram_cell[   20184] = 32'h517531bb;
    ram_cell[   20185] = 32'h1f03850b;
    ram_cell[   20186] = 32'hb30a6007;
    ram_cell[   20187] = 32'h44b5b0b3;
    ram_cell[   20188] = 32'h0b3c8af0;
    ram_cell[   20189] = 32'hb552cd1b;
    ram_cell[   20190] = 32'hc53ed1f6;
    ram_cell[   20191] = 32'h896b99c7;
    ram_cell[   20192] = 32'hb0efc6ab;
    ram_cell[   20193] = 32'h1cf112e8;
    ram_cell[   20194] = 32'hcebec285;
    ram_cell[   20195] = 32'he46ae56f;
    ram_cell[   20196] = 32'h265fe935;
    ram_cell[   20197] = 32'hc5c34b86;
    ram_cell[   20198] = 32'h6ead49ac;
    ram_cell[   20199] = 32'hd51329e9;
    ram_cell[   20200] = 32'h6eeb91f8;
    ram_cell[   20201] = 32'hd37dacfa;
    ram_cell[   20202] = 32'h331f21ff;
    ram_cell[   20203] = 32'h58d3777a;
    ram_cell[   20204] = 32'h88cc9051;
    ram_cell[   20205] = 32'h18840b9a;
    ram_cell[   20206] = 32'ha9fea933;
    ram_cell[   20207] = 32'h72c5f09d;
    ram_cell[   20208] = 32'h6f4ca5ea;
    ram_cell[   20209] = 32'h2127415a;
    ram_cell[   20210] = 32'h4359912a;
    ram_cell[   20211] = 32'h4f6d732b;
    ram_cell[   20212] = 32'h0880d1f7;
    ram_cell[   20213] = 32'h77e64d1a;
    ram_cell[   20214] = 32'h5ac620b8;
    ram_cell[   20215] = 32'h45327f96;
    ram_cell[   20216] = 32'hb3149565;
    ram_cell[   20217] = 32'hcaa5dd28;
    ram_cell[   20218] = 32'h2e65355f;
    ram_cell[   20219] = 32'h3b905957;
    ram_cell[   20220] = 32'h1431e930;
    ram_cell[   20221] = 32'hb7ed26c8;
    ram_cell[   20222] = 32'h71b06f63;
    ram_cell[   20223] = 32'ha63c94f1;
    ram_cell[   20224] = 32'hca101f13;
    ram_cell[   20225] = 32'h9c1f061f;
    ram_cell[   20226] = 32'hcb8d9368;
    ram_cell[   20227] = 32'hfe71f4bb;
    ram_cell[   20228] = 32'h730daddc;
    ram_cell[   20229] = 32'h3348f65d;
    ram_cell[   20230] = 32'h4e04b9f2;
    ram_cell[   20231] = 32'h7367c12c;
    ram_cell[   20232] = 32'h68807ab6;
    ram_cell[   20233] = 32'h976d7dcd;
    ram_cell[   20234] = 32'h4a67f744;
    ram_cell[   20235] = 32'h0924b362;
    ram_cell[   20236] = 32'h9577aef2;
    ram_cell[   20237] = 32'h147cff3a;
    ram_cell[   20238] = 32'h8172273a;
    ram_cell[   20239] = 32'ha86182fe;
    ram_cell[   20240] = 32'h129b1e97;
    ram_cell[   20241] = 32'h0ee1e010;
    ram_cell[   20242] = 32'h36b2f3bb;
    ram_cell[   20243] = 32'h84f49986;
    ram_cell[   20244] = 32'ha1ead1b9;
    ram_cell[   20245] = 32'h9d9a43af;
    ram_cell[   20246] = 32'h524fa4d8;
    ram_cell[   20247] = 32'ha7dd7c97;
    ram_cell[   20248] = 32'h9f8422de;
    ram_cell[   20249] = 32'hfcf26783;
    ram_cell[   20250] = 32'haa3ab4e1;
    ram_cell[   20251] = 32'hc327feab;
    ram_cell[   20252] = 32'h65aa71ba;
    ram_cell[   20253] = 32'h51ad6d5f;
    ram_cell[   20254] = 32'h3c9da63b;
    ram_cell[   20255] = 32'h393dcc31;
    ram_cell[   20256] = 32'h0615db69;
    ram_cell[   20257] = 32'h319098dd;
    ram_cell[   20258] = 32'h33531ea6;
    ram_cell[   20259] = 32'hf178689d;
    ram_cell[   20260] = 32'h78d477f8;
    ram_cell[   20261] = 32'h0730f5a5;
    ram_cell[   20262] = 32'h4259b197;
    ram_cell[   20263] = 32'h3b74c13e;
    ram_cell[   20264] = 32'hcf37fcf2;
    ram_cell[   20265] = 32'h3e5db1de;
    ram_cell[   20266] = 32'hdb4a9958;
    ram_cell[   20267] = 32'h44585a47;
    ram_cell[   20268] = 32'hc9e0d956;
    ram_cell[   20269] = 32'h84cf12eb;
    ram_cell[   20270] = 32'h339e3066;
    ram_cell[   20271] = 32'he7480a3b;
    ram_cell[   20272] = 32'he5d407f4;
    ram_cell[   20273] = 32'hbe472068;
    ram_cell[   20274] = 32'h95e272b8;
    ram_cell[   20275] = 32'h654747f2;
    ram_cell[   20276] = 32'hcdccead3;
    ram_cell[   20277] = 32'hf22a233a;
    ram_cell[   20278] = 32'h6226b443;
    ram_cell[   20279] = 32'h512a18ef;
    ram_cell[   20280] = 32'h11d882cc;
    ram_cell[   20281] = 32'h10d7df2d;
    ram_cell[   20282] = 32'h4a375edd;
    ram_cell[   20283] = 32'hf476e5b1;
    ram_cell[   20284] = 32'h8dc2f98e;
    ram_cell[   20285] = 32'ha8a69286;
    ram_cell[   20286] = 32'ha5121e40;
    ram_cell[   20287] = 32'hfeceba03;
    ram_cell[   20288] = 32'h65441f26;
    ram_cell[   20289] = 32'h82d200bd;
    ram_cell[   20290] = 32'h20640fac;
    ram_cell[   20291] = 32'hf9777da1;
    ram_cell[   20292] = 32'hc70c6e66;
    ram_cell[   20293] = 32'h2811e150;
    ram_cell[   20294] = 32'h103a1fb2;
    ram_cell[   20295] = 32'h41324128;
    ram_cell[   20296] = 32'hb3720689;
    ram_cell[   20297] = 32'h09623bf3;
    ram_cell[   20298] = 32'h0d6a95b7;
    ram_cell[   20299] = 32'h05fdbbf3;
    ram_cell[   20300] = 32'hdcdef3a1;
    ram_cell[   20301] = 32'h0f0b1710;
    ram_cell[   20302] = 32'hc06f7396;
    ram_cell[   20303] = 32'h3dfaed57;
    ram_cell[   20304] = 32'h6be799de;
    ram_cell[   20305] = 32'hab74c476;
    ram_cell[   20306] = 32'h85c587c8;
    ram_cell[   20307] = 32'hce8cf603;
    ram_cell[   20308] = 32'hb4e0147a;
    ram_cell[   20309] = 32'hddc27b72;
    ram_cell[   20310] = 32'h8d184816;
    ram_cell[   20311] = 32'h82d1028d;
    ram_cell[   20312] = 32'hed5bad37;
    ram_cell[   20313] = 32'h77af0eb8;
    ram_cell[   20314] = 32'h94245583;
    ram_cell[   20315] = 32'h9815ede6;
    ram_cell[   20316] = 32'h76ba9d89;
    ram_cell[   20317] = 32'h8045afb5;
    ram_cell[   20318] = 32'h98d1106e;
    ram_cell[   20319] = 32'h6a805d5d;
    ram_cell[   20320] = 32'h3f5ec415;
    ram_cell[   20321] = 32'h77cd69ec;
    ram_cell[   20322] = 32'h615f0cfc;
    ram_cell[   20323] = 32'h01951081;
    ram_cell[   20324] = 32'h7124e722;
    ram_cell[   20325] = 32'hb1b6c1b8;
    ram_cell[   20326] = 32'hc1f6b244;
    ram_cell[   20327] = 32'hfe9e2106;
    ram_cell[   20328] = 32'hfe5de7b8;
    ram_cell[   20329] = 32'h0308d8ad;
    ram_cell[   20330] = 32'h12840052;
    ram_cell[   20331] = 32'h3ffefe81;
    ram_cell[   20332] = 32'hdf167d9a;
    ram_cell[   20333] = 32'h9dc8c7bc;
    ram_cell[   20334] = 32'hc00290c3;
    ram_cell[   20335] = 32'haa058da9;
    ram_cell[   20336] = 32'hfb79d09f;
    ram_cell[   20337] = 32'h6912bb88;
    ram_cell[   20338] = 32'had09bcc1;
    ram_cell[   20339] = 32'h97b2d500;
    ram_cell[   20340] = 32'h03950384;
    ram_cell[   20341] = 32'h07ffe60c;
    ram_cell[   20342] = 32'hda9465d2;
    ram_cell[   20343] = 32'hf13797df;
    ram_cell[   20344] = 32'hb65743c5;
    ram_cell[   20345] = 32'h58eb8e7a;
    ram_cell[   20346] = 32'h0977c972;
    ram_cell[   20347] = 32'h8af50723;
    ram_cell[   20348] = 32'h0a134339;
    ram_cell[   20349] = 32'hd020e0e6;
    ram_cell[   20350] = 32'hab7cadeb;
    ram_cell[   20351] = 32'h8a6da7b4;
    ram_cell[   20352] = 32'h8391ab7e;
    ram_cell[   20353] = 32'h0dfb0625;
    ram_cell[   20354] = 32'h964caaf5;
    ram_cell[   20355] = 32'h60ee5ee4;
    ram_cell[   20356] = 32'h5ed62ee4;
    ram_cell[   20357] = 32'h1e7f4549;
    ram_cell[   20358] = 32'h0343e833;
    ram_cell[   20359] = 32'hd0e45083;
    ram_cell[   20360] = 32'h8b97809b;
    ram_cell[   20361] = 32'h33a9ee44;
    ram_cell[   20362] = 32'h471aaa44;
    ram_cell[   20363] = 32'hb446f05c;
    ram_cell[   20364] = 32'h98e40661;
    ram_cell[   20365] = 32'hc015d8ad;
    ram_cell[   20366] = 32'h497bfcc7;
    ram_cell[   20367] = 32'h35d87e03;
    ram_cell[   20368] = 32'h1ae933db;
    ram_cell[   20369] = 32'h602282bf;
    ram_cell[   20370] = 32'h2d7d2a8c;
    ram_cell[   20371] = 32'h5227e5aa;
    ram_cell[   20372] = 32'h42c536d4;
    ram_cell[   20373] = 32'h4aa5a44e;
    ram_cell[   20374] = 32'hb537d896;
    ram_cell[   20375] = 32'h6ff30d7f;
    ram_cell[   20376] = 32'h4510c281;
    ram_cell[   20377] = 32'hf83de156;
    ram_cell[   20378] = 32'h05e7d1fd;
    ram_cell[   20379] = 32'h73623688;
    ram_cell[   20380] = 32'h058d0e22;
    ram_cell[   20381] = 32'h006d3311;
    ram_cell[   20382] = 32'h24e25b05;
    ram_cell[   20383] = 32'h6c014242;
    ram_cell[   20384] = 32'h1b858439;
    ram_cell[   20385] = 32'h38df9375;
    ram_cell[   20386] = 32'h16db7692;
    ram_cell[   20387] = 32'h2a324dab;
    ram_cell[   20388] = 32'hd74f898a;
    ram_cell[   20389] = 32'h03a593c0;
    ram_cell[   20390] = 32'h0dd6b873;
    ram_cell[   20391] = 32'h005cb00f;
    ram_cell[   20392] = 32'h2607924b;
    ram_cell[   20393] = 32'h36042686;
    ram_cell[   20394] = 32'h9ce6f8ab;
    ram_cell[   20395] = 32'hef24ffd3;
    ram_cell[   20396] = 32'h6e6ec981;
    ram_cell[   20397] = 32'h449c1c7d;
    ram_cell[   20398] = 32'h68a0953a;
    ram_cell[   20399] = 32'heeb8fbe7;
    ram_cell[   20400] = 32'h76cb9192;
    ram_cell[   20401] = 32'h18462ec9;
    ram_cell[   20402] = 32'h96793f49;
    ram_cell[   20403] = 32'h97717cde;
    ram_cell[   20404] = 32'h00f32bfd;
    ram_cell[   20405] = 32'h5cec4347;
    ram_cell[   20406] = 32'h4596add4;
    ram_cell[   20407] = 32'h92564208;
    ram_cell[   20408] = 32'h39e0d4aa;
    ram_cell[   20409] = 32'h70278d3f;
    ram_cell[   20410] = 32'h0c903f65;
    ram_cell[   20411] = 32'h6fb51c5e;
    ram_cell[   20412] = 32'ha3e56e6d;
    ram_cell[   20413] = 32'h230cc10e;
    ram_cell[   20414] = 32'hfb71cf75;
    ram_cell[   20415] = 32'h4d565c75;
    ram_cell[   20416] = 32'hf65af29a;
    ram_cell[   20417] = 32'hb2d1591d;
    ram_cell[   20418] = 32'hd7d6c624;
    ram_cell[   20419] = 32'hcc3638a0;
    ram_cell[   20420] = 32'h162c0794;
    ram_cell[   20421] = 32'h48d7b5d3;
    ram_cell[   20422] = 32'hf2032045;
    ram_cell[   20423] = 32'he300ba9c;
    ram_cell[   20424] = 32'hbfe31e76;
    ram_cell[   20425] = 32'h16b359c7;
    ram_cell[   20426] = 32'h73c7f281;
    ram_cell[   20427] = 32'h97c8c78a;
    ram_cell[   20428] = 32'h788cb898;
    ram_cell[   20429] = 32'h9d4eb37f;
    ram_cell[   20430] = 32'ha52dbb22;
    ram_cell[   20431] = 32'h9d0ab353;
    ram_cell[   20432] = 32'h8c53d243;
    ram_cell[   20433] = 32'hbc257b89;
    ram_cell[   20434] = 32'h0afe5abe;
    ram_cell[   20435] = 32'h74bc1e17;
    ram_cell[   20436] = 32'hafea4ffe;
    ram_cell[   20437] = 32'hd9f7d590;
    ram_cell[   20438] = 32'hb3b7e0b2;
    ram_cell[   20439] = 32'h17e50c77;
    ram_cell[   20440] = 32'h3a1c815f;
    ram_cell[   20441] = 32'h78e20cef;
    ram_cell[   20442] = 32'h26e29c85;
    ram_cell[   20443] = 32'h6550b201;
    ram_cell[   20444] = 32'h3969c1fc;
    ram_cell[   20445] = 32'h65ca616b;
    ram_cell[   20446] = 32'h9354a981;
    ram_cell[   20447] = 32'h1400e1b8;
    ram_cell[   20448] = 32'h164a7e70;
    ram_cell[   20449] = 32'h9940a579;
    ram_cell[   20450] = 32'h81fc89a5;
    ram_cell[   20451] = 32'he6ee31ef;
    ram_cell[   20452] = 32'hf169dbaf;
    ram_cell[   20453] = 32'hcbc3718b;
    ram_cell[   20454] = 32'hd9f056e8;
    ram_cell[   20455] = 32'hdeb94345;
    ram_cell[   20456] = 32'h505bdae5;
    ram_cell[   20457] = 32'hbd114494;
    ram_cell[   20458] = 32'h99e0ae27;
    ram_cell[   20459] = 32'hcd5fe894;
    ram_cell[   20460] = 32'h1bfdbc53;
    ram_cell[   20461] = 32'hd2263ce6;
    ram_cell[   20462] = 32'h09a54450;
    ram_cell[   20463] = 32'h3622b690;
    ram_cell[   20464] = 32'h91233c9f;
    ram_cell[   20465] = 32'hcbec25c6;
    ram_cell[   20466] = 32'h6462f627;
    ram_cell[   20467] = 32'hf8d5f0b3;
    ram_cell[   20468] = 32'h0695dafd;
    ram_cell[   20469] = 32'hd1ceefbd;
    ram_cell[   20470] = 32'h52655955;
    ram_cell[   20471] = 32'h39c678cb;
    ram_cell[   20472] = 32'ha0b903af;
    ram_cell[   20473] = 32'h12da35b5;
    ram_cell[   20474] = 32'hbd816b70;
    ram_cell[   20475] = 32'h5b67fd8a;
    ram_cell[   20476] = 32'ha785c620;
    ram_cell[   20477] = 32'h284d4390;
    ram_cell[   20478] = 32'h0dd11ced;
    ram_cell[   20479] = 32'h2052c3a3;
    ram_cell[   20480] = 32'h2f64015d;
    ram_cell[   20481] = 32'h763ad77c;
    ram_cell[   20482] = 32'hc3fdbef6;
    ram_cell[   20483] = 32'hc203c0c1;
    ram_cell[   20484] = 32'hb04d8171;
    ram_cell[   20485] = 32'h3fac3956;
    ram_cell[   20486] = 32'h047052a6;
    ram_cell[   20487] = 32'h9d67c2c3;
    ram_cell[   20488] = 32'h1105eb90;
    ram_cell[   20489] = 32'h156f98ef;
    ram_cell[   20490] = 32'h4ff3b62c;
    ram_cell[   20491] = 32'h5f8b56e0;
    ram_cell[   20492] = 32'hf2749c34;
    ram_cell[   20493] = 32'hd75a45c3;
    ram_cell[   20494] = 32'hc12c95e0;
    ram_cell[   20495] = 32'ha0db05cc;
    ram_cell[   20496] = 32'hc4bcf433;
    ram_cell[   20497] = 32'h368c8e14;
    ram_cell[   20498] = 32'he42ddbf2;
    ram_cell[   20499] = 32'h827a2127;
    ram_cell[   20500] = 32'h982f4702;
    ram_cell[   20501] = 32'hf5247cb4;
    ram_cell[   20502] = 32'hed9cb522;
    ram_cell[   20503] = 32'h19df783e;
    ram_cell[   20504] = 32'ha196bb48;
    ram_cell[   20505] = 32'h84700783;
    ram_cell[   20506] = 32'h327b4876;
    ram_cell[   20507] = 32'h723e5d9f;
    ram_cell[   20508] = 32'h4860848d;
    ram_cell[   20509] = 32'hd06bd035;
    ram_cell[   20510] = 32'hd62360c6;
    ram_cell[   20511] = 32'h5412180c;
    ram_cell[   20512] = 32'h11871806;
    ram_cell[   20513] = 32'h0a1bcee9;
    ram_cell[   20514] = 32'h6929f9fd;
    ram_cell[   20515] = 32'ha0daeaba;
    ram_cell[   20516] = 32'hc54dec54;
    ram_cell[   20517] = 32'hcca3d6c7;
    ram_cell[   20518] = 32'h2d5791d9;
    ram_cell[   20519] = 32'hd130dc35;
    ram_cell[   20520] = 32'h9828089b;
    ram_cell[   20521] = 32'hb8a5118f;
    ram_cell[   20522] = 32'h29a93db9;
    ram_cell[   20523] = 32'h0e87b3f2;
    ram_cell[   20524] = 32'h2c7c715f;
    ram_cell[   20525] = 32'h7405814f;
    ram_cell[   20526] = 32'h6312bfb8;
    ram_cell[   20527] = 32'h347df9f5;
    ram_cell[   20528] = 32'h8e200c71;
    ram_cell[   20529] = 32'hb54d8520;
    ram_cell[   20530] = 32'h0eac4fa1;
    ram_cell[   20531] = 32'h726f9f65;
    ram_cell[   20532] = 32'hef04d743;
    ram_cell[   20533] = 32'hc8d26954;
    ram_cell[   20534] = 32'h2105f134;
    ram_cell[   20535] = 32'h5c724493;
    ram_cell[   20536] = 32'h0b80ad0b;
    ram_cell[   20537] = 32'hca2bde52;
    ram_cell[   20538] = 32'h9446478d;
    ram_cell[   20539] = 32'hace8c523;
    ram_cell[   20540] = 32'h8e6a83cd;
    ram_cell[   20541] = 32'hda3b13ac;
    ram_cell[   20542] = 32'hcb1b3d77;
    ram_cell[   20543] = 32'h2b7b5c4d;
    ram_cell[   20544] = 32'hcbf3ac94;
    ram_cell[   20545] = 32'ha32a1c37;
    ram_cell[   20546] = 32'hc538cb44;
    ram_cell[   20547] = 32'h8d02ec85;
    ram_cell[   20548] = 32'hfd477f15;
    ram_cell[   20549] = 32'h9bb8706d;
    ram_cell[   20550] = 32'heb7ca705;
    ram_cell[   20551] = 32'h0fa444f9;
    ram_cell[   20552] = 32'h42cedabc;
    ram_cell[   20553] = 32'h96174b38;
    ram_cell[   20554] = 32'h385e3486;
    ram_cell[   20555] = 32'h9931ece0;
    ram_cell[   20556] = 32'h111c0177;
    ram_cell[   20557] = 32'ha67f3c93;
    ram_cell[   20558] = 32'h4623fed5;
    ram_cell[   20559] = 32'hb78ddf0e;
    ram_cell[   20560] = 32'hda74e2ee;
    ram_cell[   20561] = 32'h237659c8;
    ram_cell[   20562] = 32'h5a4e5bc7;
    ram_cell[   20563] = 32'h81379a58;
    ram_cell[   20564] = 32'h8d83f262;
    ram_cell[   20565] = 32'hea341d5d;
    ram_cell[   20566] = 32'h9dfbd1b5;
    ram_cell[   20567] = 32'hbb14e34b;
    ram_cell[   20568] = 32'hb2178cd8;
    ram_cell[   20569] = 32'h07a30c0f;
    ram_cell[   20570] = 32'he099cc29;
    ram_cell[   20571] = 32'h6f740919;
    ram_cell[   20572] = 32'haaba42fa;
    ram_cell[   20573] = 32'h09533fc2;
    ram_cell[   20574] = 32'h0a4eff9c;
    ram_cell[   20575] = 32'hb7e554dd;
    ram_cell[   20576] = 32'h0a17bf39;
    ram_cell[   20577] = 32'h01d59dbf;
    ram_cell[   20578] = 32'h1c4ded5b;
    ram_cell[   20579] = 32'h53dc7b2a;
    ram_cell[   20580] = 32'he78eddf6;
    ram_cell[   20581] = 32'h76fcbc2d;
    ram_cell[   20582] = 32'ha5f5dba4;
    ram_cell[   20583] = 32'hceda2f57;
    ram_cell[   20584] = 32'hd60ad181;
    ram_cell[   20585] = 32'h2b82e4cc;
    ram_cell[   20586] = 32'h82e66e4a;
    ram_cell[   20587] = 32'h790cf9cd;
    ram_cell[   20588] = 32'hccb5b5e2;
    ram_cell[   20589] = 32'h0e2d438e;
    ram_cell[   20590] = 32'h7e6b1abf;
    ram_cell[   20591] = 32'hdad63795;
    ram_cell[   20592] = 32'h15343a40;
    ram_cell[   20593] = 32'h72d34f72;
    ram_cell[   20594] = 32'h8313d65c;
    ram_cell[   20595] = 32'h0722fed9;
    ram_cell[   20596] = 32'h50a09516;
    ram_cell[   20597] = 32'h6a89df69;
    ram_cell[   20598] = 32'hdc675722;
    ram_cell[   20599] = 32'h95b88c9a;
    ram_cell[   20600] = 32'hde9cae79;
    ram_cell[   20601] = 32'h6ecde87a;
    ram_cell[   20602] = 32'hbed7db43;
    ram_cell[   20603] = 32'h586757db;
    ram_cell[   20604] = 32'hea702736;
    ram_cell[   20605] = 32'h6697e77b;
    ram_cell[   20606] = 32'h5173653a;
    ram_cell[   20607] = 32'ha4ca7c83;
    ram_cell[   20608] = 32'hee2847a6;
    ram_cell[   20609] = 32'hcc978e7e;
    ram_cell[   20610] = 32'h26470dcd;
    ram_cell[   20611] = 32'hca63636c;
    ram_cell[   20612] = 32'hd97e5eac;
    ram_cell[   20613] = 32'h63cf55f1;
    ram_cell[   20614] = 32'h5419500e;
    ram_cell[   20615] = 32'h9b824fc9;
    ram_cell[   20616] = 32'h587a004f;
    ram_cell[   20617] = 32'h289ac05c;
    ram_cell[   20618] = 32'h07daa0d8;
    ram_cell[   20619] = 32'h041f1728;
    ram_cell[   20620] = 32'ha04b1eed;
    ram_cell[   20621] = 32'h86674549;
    ram_cell[   20622] = 32'h13c04407;
    ram_cell[   20623] = 32'h6efab20c;
    ram_cell[   20624] = 32'h34d6c15f;
    ram_cell[   20625] = 32'h26891096;
    ram_cell[   20626] = 32'h1d8b001f;
    ram_cell[   20627] = 32'h48651634;
    ram_cell[   20628] = 32'h4377279f;
    ram_cell[   20629] = 32'hd0ddd031;
    ram_cell[   20630] = 32'hc43ca7a6;
    ram_cell[   20631] = 32'h9a3e06ba;
    ram_cell[   20632] = 32'h9810ba12;
    ram_cell[   20633] = 32'hfec130d7;
    ram_cell[   20634] = 32'hac409a5c;
    ram_cell[   20635] = 32'h96306134;
    ram_cell[   20636] = 32'hb2862ed8;
    ram_cell[   20637] = 32'hadef8680;
    ram_cell[   20638] = 32'h848584b4;
    ram_cell[   20639] = 32'hd4576a5b;
    ram_cell[   20640] = 32'h80993299;
    ram_cell[   20641] = 32'h3905f179;
    ram_cell[   20642] = 32'h0dc31230;
    ram_cell[   20643] = 32'h16e5f6f9;
    ram_cell[   20644] = 32'ha52a24a6;
    ram_cell[   20645] = 32'h9695d686;
    ram_cell[   20646] = 32'hc0448bcd;
    ram_cell[   20647] = 32'h85717774;
    ram_cell[   20648] = 32'h940b22a2;
    ram_cell[   20649] = 32'h6ae407c4;
    ram_cell[   20650] = 32'he765618d;
    ram_cell[   20651] = 32'hed5b73ed;
    ram_cell[   20652] = 32'h0b7b2ada;
    ram_cell[   20653] = 32'heff2d857;
    ram_cell[   20654] = 32'h2604f88a;
    ram_cell[   20655] = 32'h9f4eee5b;
    ram_cell[   20656] = 32'h4f0829b9;
    ram_cell[   20657] = 32'h01d0063b;
    ram_cell[   20658] = 32'hf5954a04;
    ram_cell[   20659] = 32'hbe323fab;
    ram_cell[   20660] = 32'h988df660;
    ram_cell[   20661] = 32'h5eaffada;
    ram_cell[   20662] = 32'h3fe1eaf7;
    ram_cell[   20663] = 32'h54eaeea4;
    ram_cell[   20664] = 32'h03257450;
    ram_cell[   20665] = 32'h7362f3f2;
    ram_cell[   20666] = 32'h245b1efb;
    ram_cell[   20667] = 32'hf1b15153;
    ram_cell[   20668] = 32'h385901c9;
    ram_cell[   20669] = 32'h72d3141e;
    ram_cell[   20670] = 32'hed948234;
    ram_cell[   20671] = 32'hc948e0dc;
    ram_cell[   20672] = 32'h744f5185;
    ram_cell[   20673] = 32'h5305e5b9;
    ram_cell[   20674] = 32'hc26e6f62;
    ram_cell[   20675] = 32'hc4ee4aa7;
    ram_cell[   20676] = 32'h79d712d3;
    ram_cell[   20677] = 32'h06d68fc9;
    ram_cell[   20678] = 32'ha5adac65;
    ram_cell[   20679] = 32'h94e261cb;
    ram_cell[   20680] = 32'hb4d3cfa9;
    ram_cell[   20681] = 32'hd07bc6c8;
    ram_cell[   20682] = 32'hab8557c1;
    ram_cell[   20683] = 32'h042c6004;
    ram_cell[   20684] = 32'h03e5ba3e;
    ram_cell[   20685] = 32'hebb823ce;
    ram_cell[   20686] = 32'h34dbc743;
    ram_cell[   20687] = 32'h53c6a2a0;
    ram_cell[   20688] = 32'he7d1de54;
    ram_cell[   20689] = 32'h51f6920d;
    ram_cell[   20690] = 32'he3a51936;
    ram_cell[   20691] = 32'h5bf07be5;
    ram_cell[   20692] = 32'h273bb1ab;
    ram_cell[   20693] = 32'hcd878f10;
    ram_cell[   20694] = 32'hc79adb5b;
    ram_cell[   20695] = 32'h08d0981c;
    ram_cell[   20696] = 32'h36076101;
    ram_cell[   20697] = 32'hdc58fc31;
    ram_cell[   20698] = 32'h68e63fbb;
    ram_cell[   20699] = 32'he1b88195;
    ram_cell[   20700] = 32'hf956e066;
    ram_cell[   20701] = 32'hb72423bf;
    ram_cell[   20702] = 32'hb8472af3;
    ram_cell[   20703] = 32'h7133934b;
    ram_cell[   20704] = 32'he02053da;
    ram_cell[   20705] = 32'hc4de5ead;
    ram_cell[   20706] = 32'he28fd0bb;
    ram_cell[   20707] = 32'h6a5bf74c;
    ram_cell[   20708] = 32'h2dc42db0;
    ram_cell[   20709] = 32'h0db65f65;
    ram_cell[   20710] = 32'h54cd11cb;
    ram_cell[   20711] = 32'hd17707bb;
    ram_cell[   20712] = 32'hc7d9e535;
    ram_cell[   20713] = 32'h5cd8c3d3;
    ram_cell[   20714] = 32'hba4150f4;
    ram_cell[   20715] = 32'h9673febe;
    ram_cell[   20716] = 32'h1514d964;
    ram_cell[   20717] = 32'hfa03a3f0;
    ram_cell[   20718] = 32'h562fd2ac;
    ram_cell[   20719] = 32'h3d38081e;
    ram_cell[   20720] = 32'h7070ce9e;
    ram_cell[   20721] = 32'h20601ab7;
    ram_cell[   20722] = 32'hca2456cf;
    ram_cell[   20723] = 32'hba5d0277;
    ram_cell[   20724] = 32'hfc199eda;
    ram_cell[   20725] = 32'hca01d27b;
    ram_cell[   20726] = 32'h9ebec75b;
    ram_cell[   20727] = 32'h2c5d82d2;
    ram_cell[   20728] = 32'hc37a75ee;
    ram_cell[   20729] = 32'h06e3af0e;
    ram_cell[   20730] = 32'hea61717b;
    ram_cell[   20731] = 32'h77e4bbf7;
    ram_cell[   20732] = 32'hfa6a5746;
    ram_cell[   20733] = 32'h418d5910;
    ram_cell[   20734] = 32'h04812d80;
    ram_cell[   20735] = 32'h33016cbd;
    ram_cell[   20736] = 32'hbce468d8;
    ram_cell[   20737] = 32'hca6d2907;
    ram_cell[   20738] = 32'hab2a88a1;
    ram_cell[   20739] = 32'h3f98a5d8;
    ram_cell[   20740] = 32'hfc534d85;
    ram_cell[   20741] = 32'ha2fa8a9e;
    ram_cell[   20742] = 32'h4ca74089;
    ram_cell[   20743] = 32'h3cf8e038;
    ram_cell[   20744] = 32'hd68b930d;
    ram_cell[   20745] = 32'h0697def6;
    ram_cell[   20746] = 32'h89d4b73a;
    ram_cell[   20747] = 32'hba958017;
    ram_cell[   20748] = 32'h87518b71;
    ram_cell[   20749] = 32'h3696d261;
    ram_cell[   20750] = 32'hec8d0ed1;
    ram_cell[   20751] = 32'h6141244e;
    ram_cell[   20752] = 32'hdc449628;
    ram_cell[   20753] = 32'h627e1d32;
    ram_cell[   20754] = 32'h378b8504;
    ram_cell[   20755] = 32'he18ddbb7;
    ram_cell[   20756] = 32'h6909a987;
    ram_cell[   20757] = 32'he3d24572;
    ram_cell[   20758] = 32'h6964a82d;
    ram_cell[   20759] = 32'hd9091185;
    ram_cell[   20760] = 32'h82c908ce;
    ram_cell[   20761] = 32'hf6f7a160;
    ram_cell[   20762] = 32'hb30f2ff3;
    ram_cell[   20763] = 32'h15182757;
    ram_cell[   20764] = 32'he4895a49;
    ram_cell[   20765] = 32'h142bd334;
    ram_cell[   20766] = 32'ha658aa0b;
    ram_cell[   20767] = 32'h1d4df8bd;
    ram_cell[   20768] = 32'hcbbd046c;
    ram_cell[   20769] = 32'h27981914;
    ram_cell[   20770] = 32'h1e0501b3;
    ram_cell[   20771] = 32'hb78c20ea;
    ram_cell[   20772] = 32'hcc2932c3;
    ram_cell[   20773] = 32'h58649d34;
    ram_cell[   20774] = 32'haa52617c;
    ram_cell[   20775] = 32'h8bf4a29a;
    ram_cell[   20776] = 32'h8b9f26ff;
    ram_cell[   20777] = 32'h58bbeeff;
    ram_cell[   20778] = 32'h6df6f5bc;
    ram_cell[   20779] = 32'h085c1995;
    ram_cell[   20780] = 32'h16bfe888;
    ram_cell[   20781] = 32'h0b2c403d;
    ram_cell[   20782] = 32'he90238c1;
    ram_cell[   20783] = 32'h5d55ff1b;
    ram_cell[   20784] = 32'he7508c17;
    ram_cell[   20785] = 32'hab0882a4;
    ram_cell[   20786] = 32'h83ea1157;
    ram_cell[   20787] = 32'h56b33f2f;
    ram_cell[   20788] = 32'h1c19d76f;
    ram_cell[   20789] = 32'hfdbafe78;
    ram_cell[   20790] = 32'h76cae9ec;
    ram_cell[   20791] = 32'h4d420a18;
    ram_cell[   20792] = 32'hc9e91c7b;
    ram_cell[   20793] = 32'hef3a9020;
    ram_cell[   20794] = 32'h6b2149a1;
    ram_cell[   20795] = 32'h134a229b;
    ram_cell[   20796] = 32'h16ce98c4;
    ram_cell[   20797] = 32'h6297b45e;
    ram_cell[   20798] = 32'h1c36863d;
    ram_cell[   20799] = 32'h7587d93e;
    ram_cell[   20800] = 32'h1220c32f;
    ram_cell[   20801] = 32'h2d5d8059;
    ram_cell[   20802] = 32'h716329d4;
    ram_cell[   20803] = 32'h64438b8c;
    ram_cell[   20804] = 32'hbf9e39e8;
    ram_cell[   20805] = 32'hd3948139;
    ram_cell[   20806] = 32'h21681372;
    ram_cell[   20807] = 32'hf126e61c;
    ram_cell[   20808] = 32'hd55511ff;
    ram_cell[   20809] = 32'hc30dd982;
    ram_cell[   20810] = 32'h1d4bc874;
    ram_cell[   20811] = 32'h0195fddf;
    ram_cell[   20812] = 32'h34b3a614;
    ram_cell[   20813] = 32'h42845cdb;
    ram_cell[   20814] = 32'h4644ddad;
    ram_cell[   20815] = 32'he71aa5de;
    ram_cell[   20816] = 32'ha5d9f43c;
    ram_cell[   20817] = 32'h3f7b06ec;
    ram_cell[   20818] = 32'h5dcc2f11;
    ram_cell[   20819] = 32'hcea2c519;
    ram_cell[   20820] = 32'hb1115e4d;
    ram_cell[   20821] = 32'h3e8f10c2;
    ram_cell[   20822] = 32'h5e39ffbc;
    ram_cell[   20823] = 32'h4a2d1129;
    ram_cell[   20824] = 32'h8f039422;
    ram_cell[   20825] = 32'h5c4aa7aa;
    ram_cell[   20826] = 32'hf660879f;
    ram_cell[   20827] = 32'h5ce4090d;
    ram_cell[   20828] = 32'hcdc74279;
    ram_cell[   20829] = 32'hd8c588b5;
    ram_cell[   20830] = 32'ha8789d7b;
    ram_cell[   20831] = 32'h6e94b710;
    ram_cell[   20832] = 32'h1c55a00b;
    ram_cell[   20833] = 32'h6a108b3f;
    ram_cell[   20834] = 32'h62d40647;
    ram_cell[   20835] = 32'he42a7448;
    ram_cell[   20836] = 32'h01c028f6;
    ram_cell[   20837] = 32'he9c93f33;
    ram_cell[   20838] = 32'hd2801296;
    ram_cell[   20839] = 32'hcb59b543;
    ram_cell[   20840] = 32'hf825c2dd;
    ram_cell[   20841] = 32'he97f6362;
    ram_cell[   20842] = 32'h4c118ce0;
    ram_cell[   20843] = 32'hb8cb0578;
    ram_cell[   20844] = 32'h423aeb11;
    ram_cell[   20845] = 32'h6fd9e30b;
    ram_cell[   20846] = 32'hdbc83fb3;
    ram_cell[   20847] = 32'hcbb2f1a4;
    ram_cell[   20848] = 32'h3f17bba6;
    ram_cell[   20849] = 32'h1e26081b;
    ram_cell[   20850] = 32'h165ddb8a;
    ram_cell[   20851] = 32'h9e654c5b;
    ram_cell[   20852] = 32'h4a418704;
    ram_cell[   20853] = 32'he3331cd7;
    ram_cell[   20854] = 32'h346cefab;
    ram_cell[   20855] = 32'hdfa70953;
    ram_cell[   20856] = 32'ha538eea8;
    ram_cell[   20857] = 32'h2c21a485;
    ram_cell[   20858] = 32'hcd6ac45d;
    ram_cell[   20859] = 32'h090985b2;
    ram_cell[   20860] = 32'h50b98a51;
    ram_cell[   20861] = 32'h9451b703;
    ram_cell[   20862] = 32'ha7e3430b;
    ram_cell[   20863] = 32'h92bfbb49;
    ram_cell[   20864] = 32'h099b4422;
    ram_cell[   20865] = 32'h6eba6bbe;
    ram_cell[   20866] = 32'hdac06ba8;
    ram_cell[   20867] = 32'h4cb04721;
    ram_cell[   20868] = 32'h5d37616d;
    ram_cell[   20869] = 32'h6f1f1175;
    ram_cell[   20870] = 32'haefb694f;
    ram_cell[   20871] = 32'hfd460fab;
    ram_cell[   20872] = 32'hddbeed1f;
    ram_cell[   20873] = 32'h736b9347;
    ram_cell[   20874] = 32'h8d17af58;
    ram_cell[   20875] = 32'hbc7d23ad;
    ram_cell[   20876] = 32'hc70d1165;
    ram_cell[   20877] = 32'h8d7c9791;
    ram_cell[   20878] = 32'h0addf16d;
    ram_cell[   20879] = 32'h680fd560;
    ram_cell[   20880] = 32'h3256451a;
    ram_cell[   20881] = 32'hf5871b9e;
    ram_cell[   20882] = 32'heb83650d;
    ram_cell[   20883] = 32'ha8e9aa7e;
    ram_cell[   20884] = 32'h4f04fa4b;
    ram_cell[   20885] = 32'h7560b28f;
    ram_cell[   20886] = 32'h514fb411;
    ram_cell[   20887] = 32'he77304b7;
    ram_cell[   20888] = 32'ha6c73420;
    ram_cell[   20889] = 32'h30c46676;
    ram_cell[   20890] = 32'h3ad6f36b;
    ram_cell[   20891] = 32'hf91cb68d;
    ram_cell[   20892] = 32'h629db9f0;
    ram_cell[   20893] = 32'h5c06d5f9;
    ram_cell[   20894] = 32'h6ec0b944;
    ram_cell[   20895] = 32'h3e621052;
    ram_cell[   20896] = 32'hd6c7fbe9;
    ram_cell[   20897] = 32'h3cd76c9b;
    ram_cell[   20898] = 32'h289768ff;
    ram_cell[   20899] = 32'h325cae48;
    ram_cell[   20900] = 32'h6874d982;
    ram_cell[   20901] = 32'he7cace8a;
    ram_cell[   20902] = 32'ha14c2472;
    ram_cell[   20903] = 32'ha24086f4;
    ram_cell[   20904] = 32'h40b151d3;
    ram_cell[   20905] = 32'hf75e21b2;
    ram_cell[   20906] = 32'h4638e2e9;
    ram_cell[   20907] = 32'h9710e0f7;
    ram_cell[   20908] = 32'h39bed5c3;
    ram_cell[   20909] = 32'hd730bed7;
    ram_cell[   20910] = 32'h9461d9e8;
    ram_cell[   20911] = 32'hdbf98ab3;
    ram_cell[   20912] = 32'h7a3999b0;
    ram_cell[   20913] = 32'ha1bdd7df;
    ram_cell[   20914] = 32'h3ec74cbc;
    ram_cell[   20915] = 32'hef135ea3;
    ram_cell[   20916] = 32'h1035a73b;
    ram_cell[   20917] = 32'h52f3b5ad;
    ram_cell[   20918] = 32'hbed1e3ae;
    ram_cell[   20919] = 32'hf03dc933;
    ram_cell[   20920] = 32'h766c1ddf;
    ram_cell[   20921] = 32'h84276549;
    ram_cell[   20922] = 32'h57c0e660;
    ram_cell[   20923] = 32'hea8932a6;
    ram_cell[   20924] = 32'h4b1cde49;
    ram_cell[   20925] = 32'h0c7beff8;
    ram_cell[   20926] = 32'hf638dedd;
    ram_cell[   20927] = 32'h46c2982e;
    ram_cell[   20928] = 32'hcccadf87;
    ram_cell[   20929] = 32'h6dd40932;
    ram_cell[   20930] = 32'h8281f62a;
    ram_cell[   20931] = 32'h4aa3e69f;
    ram_cell[   20932] = 32'he25dce46;
    ram_cell[   20933] = 32'he4b176c6;
    ram_cell[   20934] = 32'h68787b82;
    ram_cell[   20935] = 32'h64082eb4;
    ram_cell[   20936] = 32'hc2a7ad34;
    ram_cell[   20937] = 32'h8bf35c20;
    ram_cell[   20938] = 32'h7a2da07f;
    ram_cell[   20939] = 32'h31e3a4de;
    ram_cell[   20940] = 32'h827330a9;
    ram_cell[   20941] = 32'h8f2855ed;
    ram_cell[   20942] = 32'h5c21fb2f;
    ram_cell[   20943] = 32'haaaa5fbf;
    ram_cell[   20944] = 32'hd8c21bc3;
    ram_cell[   20945] = 32'h7c80c5e9;
    ram_cell[   20946] = 32'he8722c90;
    ram_cell[   20947] = 32'hc9cc1da2;
    ram_cell[   20948] = 32'h5999f15d;
    ram_cell[   20949] = 32'h426d8d59;
    ram_cell[   20950] = 32'h73e883f8;
    ram_cell[   20951] = 32'ha6b88c93;
    ram_cell[   20952] = 32'hcbbd3f6d;
    ram_cell[   20953] = 32'ha7ea4559;
    ram_cell[   20954] = 32'hca377851;
    ram_cell[   20955] = 32'hff414cab;
    ram_cell[   20956] = 32'h02596587;
    ram_cell[   20957] = 32'h11ed326c;
    ram_cell[   20958] = 32'h2e101489;
    ram_cell[   20959] = 32'hd1f27da8;
    ram_cell[   20960] = 32'h68057f96;
    ram_cell[   20961] = 32'heb9470ac;
    ram_cell[   20962] = 32'ha1872763;
    ram_cell[   20963] = 32'h9e42e2e7;
    ram_cell[   20964] = 32'h0424cd5c;
    ram_cell[   20965] = 32'h9113eac1;
    ram_cell[   20966] = 32'h6b99f5ef;
    ram_cell[   20967] = 32'h7bed0b0a;
    ram_cell[   20968] = 32'h64762908;
    ram_cell[   20969] = 32'h61c46856;
    ram_cell[   20970] = 32'h97782000;
    ram_cell[   20971] = 32'hf42fff28;
    ram_cell[   20972] = 32'h623c4526;
    ram_cell[   20973] = 32'h893a272f;
    ram_cell[   20974] = 32'h0a1d0892;
    ram_cell[   20975] = 32'ha61276a4;
    ram_cell[   20976] = 32'h0d2736bb;
    ram_cell[   20977] = 32'h110ef2a2;
    ram_cell[   20978] = 32'h64c3dd28;
    ram_cell[   20979] = 32'ha1f7ba75;
    ram_cell[   20980] = 32'h314560eb;
    ram_cell[   20981] = 32'h5facb6b0;
    ram_cell[   20982] = 32'h35cb302e;
    ram_cell[   20983] = 32'h9c4f5ec7;
    ram_cell[   20984] = 32'h9bacc164;
    ram_cell[   20985] = 32'h72882c09;
    ram_cell[   20986] = 32'h32b38caa;
    ram_cell[   20987] = 32'hdd0b63f1;
    ram_cell[   20988] = 32'hbc803790;
    ram_cell[   20989] = 32'h0d0cb91c;
    ram_cell[   20990] = 32'h4e7a3880;
    ram_cell[   20991] = 32'h3c7a3528;
    ram_cell[   20992] = 32'h2f59b9ec;
    ram_cell[   20993] = 32'hce495a2d;
    ram_cell[   20994] = 32'hb178419c;
    ram_cell[   20995] = 32'h53faa6a0;
    ram_cell[   20996] = 32'h2bd9416a;
    ram_cell[   20997] = 32'h6c3a3407;
    ram_cell[   20998] = 32'he09eac1c;
    ram_cell[   20999] = 32'hf2b615da;
    ram_cell[   21000] = 32'hd7b6c740;
    ram_cell[   21001] = 32'h09e1c525;
    ram_cell[   21002] = 32'ha922c6df;
    ram_cell[   21003] = 32'h918c3a32;
    ram_cell[   21004] = 32'h627d44cc;
    ram_cell[   21005] = 32'h97424ebf;
    ram_cell[   21006] = 32'hae99de43;
    ram_cell[   21007] = 32'he5dd470a;
    ram_cell[   21008] = 32'h489584be;
    ram_cell[   21009] = 32'hbc8d5060;
    ram_cell[   21010] = 32'hd244d27f;
    ram_cell[   21011] = 32'h727715dd;
    ram_cell[   21012] = 32'h4625c321;
    ram_cell[   21013] = 32'h2da8867b;
    ram_cell[   21014] = 32'hbecb0905;
    ram_cell[   21015] = 32'h390177fc;
    ram_cell[   21016] = 32'h777342ee;
    ram_cell[   21017] = 32'hd8b07227;
    ram_cell[   21018] = 32'hb69fc3f3;
    ram_cell[   21019] = 32'h2141e2ff;
    ram_cell[   21020] = 32'h2b299ee2;
    ram_cell[   21021] = 32'h3f488a51;
    ram_cell[   21022] = 32'hda15ca61;
    ram_cell[   21023] = 32'h56a9061e;
    ram_cell[   21024] = 32'hd888f4ce;
    ram_cell[   21025] = 32'hbc67b900;
    ram_cell[   21026] = 32'h7d901997;
    ram_cell[   21027] = 32'heae43add;
    ram_cell[   21028] = 32'h2f8095ff;
    ram_cell[   21029] = 32'h00bfee4b;
    ram_cell[   21030] = 32'hf2e6391e;
    ram_cell[   21031] = 32'hc4e79e55;
    ram_cell[   21032] = 32'h64c356bf;
    ram_cell[   21033] = 32'h7a16d3e2;
    ram_cell[   21034] = 32'hc27248c0;
    ram_cell[   21035] = 32'h43b1a771;
    ram_cell[   21036] = 32'h8dcffe1d;
    ram_cell[   21037] = 32'h7336c9e2;
    ram_cell[   21038] = 32'h49f44862;
    ram_cell[   21039] = 32'h38f2da18;
    ram_cell[   21040] = 32'hee9eb7d9;
    ram_cell[   21041] = 32'h50798344;
    ram_cell[   21042] = 32'hfe93490c;
    ram_cell[   21043] = 32'hd1e0dc70;
    ram_cell[   21044] = 32'h49fea5a3;
    ram_cell[   21045] = 32'h179f2670;
    ram_cell[   21046] = 32'h22c54b4f;
    ram_cell[   21047] = 32'hf7872a8f;
    ram_cell[   21048] = 32'h662162b5;
    ram_cell[   21049] = 32'h61196174;
    ram_cell[   21050] = 32'h35f64266;
    ram_cell[   21051] = 32'h4c44855b;
    ram_cell[   21052] = 32'h42b59058;
    ram_cell[   21053] = 32'he69d7ad7;
    ram_cell[   21054] = 32'h409c584d;
    ram_cell[   21055] = 32'h1a3f745f;
    ram_cell[   21056] = 32'h0992c039;
    ram_cell[   21057] = 32'h1cf2d001;
    ram_cell[   21058] = 32'hec0efbaf;
    ram_cell[   21059] = 32'he37933a2;
    ram_cell[   21060] = 32'h9bfda23a;
    ram_cell[   21061] = 32'hf1ad86d7;
    ram_cell[   21062] = 32'h4278c72e;
    ram_cell[   21063] = 32'h0bd38697;
    ram_cell[   21064] = 32'hb1ad3461;
    ram_cell[   21065] = 32'h697dd97e;
    ram_cell[   21066] = 32'he52c5479;
    ram_cell[   21067] = 32'h172cfb3e;
    ram_cell[   21068] = 32'h8e8652ac;
    ram_cell[   21069] = 32'hf4d4316f;
    ram_cell[   21070] = 32'habf3dbd3;
    ram_cell[   21071] = 32'h4d2a7ec0;
    ram_cell[   21072] = 32'haf92d346;
    ram_cell[   21073] = 32'h34fbc556;
    ram_cell[   21074] = 32'ha8dcea8d;
    ram_cell[   21075] = 32'h3bb9fabb;
    ram_cell[   21076] = 32'hd8b9c5af;
    ram_cell[   21077] = 32'h52d1a2cc;
    ram_cell[   21078] = 32'h0c0adcff;
    ram_cell[   21079] = 32'hdb9ee00d;
    ram_cell[   21080] = 32'h35403e55;
    ram_cell[   21081] = 32'h3fe4c260;
    ram_cell[   21082] = 32'hde5972b0;
    ram_cell[   21083] = 32'hbb8564d0;
    ram_cell[   21084] = 32'h60f97505;
    ram_cell[   21085] = 32'hd4e1eca8;
    ram_cell[   21086] = 32'h2ae81023;
    ram_cell[   21087] = 32'h1ef527cc;
    ram_cell[   21088] = 32'h2b1dcdf9;
    ram_cell[   21089] = 32'h17521e5e;
    ram_cell[   21090] = 32'hb49cd734;
    ram_cell[   21091] = 32'h8ea2f7c1;
    ram_cell[   21092] = 32'hf6352a50;
    ram_cell[   21093] = 32'hfb7d4116;
    ram_cell[   21094] = 32'h608f6a85;
    ram_cell[   21095] = 32'h82a5a942;
    ram_cell[   21096] = 32'h65a29cd5;
    ram_cell[   21097] = 32'h451c65b5;
    ram_cell[   21098] = 32'h669a6886;
    ram_cell[   21099] = 32'hbf03a725;
    ram_cell[   21100] = 32'h69b5e98b;
    ram_cell[   21101] = 32'he7693615;
    ram_cell[   21102] = 32'h57b2a1cc;
    ram_cell[   21103] = 32'h75ab2ae5;
    ram_cell[   21104] = 32'h497ed232;
    ram_cell[   21105] = 32'h7a0f2ba3;
    ram_cell[   21106] = 32'h97839ddb;
    ram_cell[   21107] = 32'h01a76d18;
    ram_cell[   21108] = 32'hf27f7772;
    ram_cell[   21109] = 32'hd68777d3;
    ram_cell[   21110] = 32'hc7b72bff;
    ram_cell[   21111] = 32'h0d80f3c7;
    ram_cell[   21112] = 32'h76a6664b;
    ram_cell[   21113] = 32'haefc8181;
    ram_cell[   21114] = 32'hcf75bd17;
    ram_cell[   21115] = 32'h26fa4974;
    ram_cell[   21116] = 32'h7cce76b0;
    ram_cell[   21117] = 32'hca4249b9;
    ram_cell[   21118] = 32'h573f39b8;
    ram_cell[   21119] = 32'habe980e4;
    ram_cell[   21120] = 32'h449260ca;
    ram_cell[   21121] = 32'hf1ee94e1;
    ram_cell[   21122] = 32'h1eb12db2;
    ram_cell[   21123] = 32'h2e3ebf2a;
    ram_cell[   21124] = 32'h947767a3;
    ram_cell[   21125] = 32'he3741485;
    ram_cell[   21126] = 32'hdbf3246b;
    ram_cell[   21127] = 32'hf02ff574;
    ram_cell[   21128] = 32'h0ee0a430;
    ram_cell[   21129] = 32'h102e9538;
    ram_cell[   21130] = 32'h3802cad9;
    ram_cell[   21131] = 32'h9de22952;
    ram_cell[   21132] = 32'hff88a683;
    ram_cell[   21133] = 32'hb572b177;
    ram_cell[   21134] = 32'hb60503a3;
    ram_cell[   21135] = 32'hf81b873c;
    ram_cell[   21136] = 32'h7295c753;
    ram_cell[   21137] = 32'h7201ef17;
    ram_cell[   21138] = 32'h4c1ce94b;
    ram_cell[   21139] = 32'h7b9afe61;
    ram_cell[   21140] = 32'h39497959;
    ram_cell[   21141] = 32'hd5ae7dd9;
    ram_cell[   21142] = 32'hc434be5f;
    ram_cell[   21143] = 32'hd5f29689;
    ram_cell[   21144] = 32'h854ed623;
    ram_cell[   21145] = 32'h2a7947a4;
    ram_cell[   21146] = 32'h9c11b596;
    ram_cell[   21147] = 32'h67094fac;
    ram_cell[   21148] = 32'h2dd5ed40;
    ram_cell[   21149] = 32'h79373d0c;
    ram_cell[   21150] = 32'h8acca7c7;
    ram_cell[   21151] = 32'h9aa656b5;
    ram_cell[   21152] = 32'h26e095e7;
    ram_cell[   21153] = 32'hdd9483bc;
    ram_cell[   21154] = 32'h7caff90e;
    ram_cell[   21155] = 32'h7e1fd852;
    ram_cell[   21156] = 32'hda95820c;
    ram_cell[   21157] = 32'heb291739;
    ram_cell[   21158] = 32'h6da13cd3;
    ram_cell[   21159] = 32'h43371d12;
    ram_cell[   21160] = 32'h35f4201c;
    ram_cell[   21161] = 32'h67583733;
    ram_cell[   21162] = 32'h88155037;
    ram_cell[   21163] = 32'h5bdba99b;
    ram_cell[   21164] = 32'h926800c4;
    ram_cell[   21165] = 32'h493f47d6;
    ram_cell[   21166] = 32'hf5b1fc09;
    ram_cell[   21167] = 32'h30f1f25c;
    ram_cell[   21168] = 32'ha327b60c;
    ram_cell[   21169] = 32'h8d9937d3;
    ram_cell[   21170] = 32'hfb5da0db;
    ram_cell[   21171] = 32'h8a7ba74a;
    ram_cell[   21172] = 32'h454c50cd;
    ram_cell[   21173] = 32'h08e758bf;
    ram_cell[   21174] = 32'h972ed581;
    ram_cell[   21175] = 32'hc1a7bd7f;
    ram_cell[   21176] = 32'he7052021;
    ram_cell[   21177] = 32'h93b0e131;
    ram_cell[   21178] = 32'h28b2000a;
    ram_cell[   21179] = 32'h18348c68;
    ram_cell[   21180] = 32'h6dc30d49;
    ram_cell[   21181] = 32'h20152a7f;
    ram_cell[   21182] = 32'hbf35e5b4;
    ram_cell[   21183] = 32'h0d0cb8e9;
    ram_cell[   21184] = 32'hbe9b8816;
    ram_cell[   21185] = 32'hf633f555;
    ram_cell[   21186] = 32'h6665c2d0;
    ram_cell[   21187] = 32'hedaf7448;
    ram_cell[   21188] = 32'h4e0247c8;
    ram_cell[   21189] = 32'h46d3b104;
    ram_cell[   21190] = 32'h5cc7137c;
    ram_cell[   21191] = 32'hb997510b;
    ram_cell[   21192] = 32'hfd520d86;
    ram_cell[   21193] = 32'hb65a49c3;
    ram_cell[   21194] = 32'h6a00792a;
    ram_cell[   21195] = 32'hb978cf4e;
    ram_cell[   21196] = 32'hbbd90fed;
    ram_cell[   21197] = 32'hfa719a71;
    ram_cell[   21198] = 32'h49ce9ff5;
    ram_cell[   21199] = 32'ha94ec447;
    ram_cell[   21200] = 32'he7eff42b;
    ram_cell[   21201] = 32'h83bfea83;
    ram_cell[   21202] = 32'h02e055b7;
    ram_cell[   21203] = 32'h94739aa2;
    ram_cell[   21204] = 32'h7dae387e;
    ram_cell[   21205] = 32'h036940d5;
    ram_cell[   21206] = 32'hb92b4df2;
    ram_cell[   21207] = 32'habb4b6a6;
    ram_cell[   21208] = 32'h649db6eb;
    ram_cell[   21209] = 32'h8838e7fb;
    ram_cell[   21210] = 32'h19ce4d12;
    ram_cell[   21211] = 32'h739743bf;
    ram_cell[   21212] = 32'h10099717;
    ram_cell[   21213] = 32'habfd2a62;
    ram_cell[   21214] = 32'h91e376f9;
    ram_cell[   21215] = 32'h3681cad4;
    ram_cell[   21216] = 32'h6840257b;
    ram_cell[   21217] = 32'h497ecb51;
    ram_cell[   21218] = 32'hf55611cf;
    ram_cell[   21219] = 32'h3cd3aff6;
    ram_cell[   21220] = 32'h6b1d79fb;
    ram_cell[   21221] = 32'hab0d866a;
    ram_cell[   21222] = 32'h542bf8ec;
    ram_cell[   21223] = 32'h6800b93f;
    ram_cell[   21224] = 32'h3cd9b994;
    ram_cell[   21225] = 32'h85c37ebe;
    ram_cell[   21226] = 32'hb664b6fe;
    ram_cell[   21227] = 32'h11bc7698;
    ram_cell[   21228] = 32'hbd9716b5;
    ram_cell[   21229] = 32'hda066250;
    ram_cell[   21230] = 32'hfc276bb6;
    ram_cell[   21231] = 32'ha703c727;
    ram_cell[   21232] = 32'h61a9b125;
    ram_cell[   21233] = 32'hcda88e32;
    ram_cell[   21234] = 32'h12e64052;
    ram_cell[   21235] = 32'h9275bee1;
    ram_cell[   21236] = 32'hd535080d;
    ram_cell[   21237] = 32'h0ac2784d;
    ram_cell[   21238] = 32'h90b99ad9;
    ram_cell[   21239] = 32'h31964cf6;
    ram_cell[   21240] = 32'h15bae44e;
    ram_cell[   21241] = 32'h4c7cc0fb;
    ram_cell[   21242] = 32'h3962ea68;
    ram_cell[   21243] = 32'h8410aa8a;
    ram_cell[   21244] = 32'h08b72be1;
    ram_cell[   21245] = 32'h592243ac;
    ram_cell[   21246] = 32'hdac17616;
    ram_cell[   21247] = 32'haccd7dca;
    ram_cell[   21248] = 32'h08e4705a;
    ram_cell[   21249] = 32'h1e73c0b3;
    ram_cell[   21250] = 32'hcacb7861;
    ram_cell[   21251] = 32'he7b6b26b;
    ram_cell[   21252] = 32'h49177959;
    ram_cell[   21253] = 32'h5ec7908c;
    ram_cell[   21254] = 32'h166e3a44;
    ram_cell[   21255] = 32'h5587452c;
    ram_cell[   21256] = 32'h74c5deb6;
    ram_cell[   21257] = 32'he5ed9205;
    ram_cell[   21258] = 32'h9ad92d8e;
    ram_cell[   21259] = 32'h5345bd8b;
    ram_cell[   21260] = 32'h92242d8c;
    ram_cell[   21261] = 32'h72c5ecaf;
    ram_cell[   21262] = 32'hfdf54217;
    ram_cell[   21263] = 32'h7f7a3ea5;
    ram_cell[   21264] = 32'h28024a88;
    ram_cell[   21265] = 32'h81d0d6b5;
    ram_cell[   21266] = 32'h8e6ad9cc;
    ram_cell[   21267] = 32'h51776050;
    ram_cell[   21268] = 32'hc2568204;
    ram_cell[   21269] = 32'ha1455794;
    ram_cell[   21270] = 32'h41ef0663;
    ram_cell[   21271] = 32'h9ba9765d;
    ram_cell[   21272] = 32'haa203fee;
    ram_cell[   21273] = 32'h38c8680d;
    ram_cell[   21274] = 32'hb8b0f4ad;
    ram_cell[   21275] = 32'h051fa4ff;
    ram_cell[   21276] = 32'h0331d548;
    ram_cell[   21277] = 32'h70d295ba;
    ram_cell[   21278] = 32'h6f3261c8;
    ram_cell[   21279] = 32'hfdf54c2a;
    ram_cell[   21280] = 32'h56a77246;
    ram_cell[   21281] = 32'h004b0fd0;
    ram_cell[   21282] = 32'hdfdda0c2;
    ram_cell[   21283] = 32'h683d0257;
    ram_cell[   21284] = 32'hff4fe355;
    ram_cell[   21285] = 32'h813bb33f;
    ram_cell[   21286] = 32'hd3afc5a1;
    ram_cell[   21287] = 32'h0ccba6ea;
    ram_cell[   21288] = 32'h0953fbce;
    ram_cell[   21289] = 32'h7127afad;
    ram_cell[   21290] = 32'h3121f690;
    ram_cell[   21291] = 32'hcb18eba4;
    ram_cell[   21292] = 32'hf101300a;
    ram_cell[   21293] = 32'h98cbb33e;
    ram_cell[   21294] = 32'hfa09c6d4;
    ram_cell[   21295] = 32'hfe72834e;
    ram_cell[   21296] = 32'hac02f5a8;
    ram_cell[   21297] = 32'hc6697983;
    ram_cell[   21298] = 32'he864aa66;
    ram_cell[   21299] = 32'h32e7d482;
    ram_cell[   21300] = 32'h84da642f;
    ram_cell[   21301] = 32'he6681e46;
    ram_cell[   21302] = 32'h364e548a;
    ram_cell[   21303] = 32'ha7afaecd;
    ram_cell[   21304] = 32'hd51fad1b;
    ram_cell[   21305] = 32'h889d4fb1;
    ram_cell[   21306] = 32'he988e0fc;
    ram_cell[   21307] = 32'hd2e73624;
    ram_cell[   21308] = 32'h37a980cb;
    ram_cell[   21309] = 32'h0aecdf5c;
    ram_cell[   21310] = 32'h66bcbbb5;
    ram_cell[   21311] = 32'h1f91e68f;
    ram_cell[   21312] = 32'ha2b3c468;
    ram_cell[   21313] = 32'h53590d58;
    ram_cell[   21314] = 32'hfaab8d30;
    ram_cell[   21315] = 32'h7c695d43;
    ram_cell[   21316] = 32'h155edf1e;
    ram_cell[   21317] = 32'h768bafb8;
    ram_cell[   21318] = 32'h1a290bcb;
    ram_cell[   21319] = 32'h57388a90;
    ram_cell[   21320] = 32'h73df4cdd;
    ram_cell[   21321] = 32'hdaf8b343;
    ram_cell[   21322] = 32'he9b3b513;
    ram_cell[   21323] = 32'he4dcae3c;
    ram_cell[   21324] = 32'h5334846f;
    ram_cell[   21325] = 32'h3b5183f5;
    ram_cell[   21326] = 32'h232faef8;
    ram_cell[   21327] = 32'h92fe55d4;
    ram_cell[   21328] = 32'h4ce3b018;
    ram_cell[   21329] = 32'h6b2bc0e8;
    ram_cell[   21330] = 32'h48c75eab;
    ram_cell[   21331] = 32'h9332b986;
    ram_cell[   21332] = 32'h32c69b0a;
    ram_cell[   21333] = 32'h95e3ce5a;
    ram_cell[   21334] = 32'haf31f463;
    ram_cell[   21335] = 32'hdce69a32;
    ram_cell[   21336] = 32'h7b78c1d9;
    ram_cell[   21337] = 32'h59efce24;
    ram_cell[   21338] = 32'h0386b8e7;
    ram_cell[   21339] = 32'hb48d6472;
    ram_cell[   21340] = 32'h698da2ee;
    ram_cell[   21341] = 32'h351f8fc8;
    ram_cell[   21342] = 32'hda01b970;
    ram_cell[   21343] = 32'hc185af90;
    ram_cell[   21344] = 32'hd1e1d49e;
    ram_cell[   21345] = 32'h04fc09b3;
    ram_cell[   21346] = 32'h3afd434e;
    ram_cell[   21347] = 32'h11d3a29f;
    ram_cell[   21348] = 32'h6d1cd8f5;
    ram_cell[   21349] = 32'hccf15b01;
    ram_cell[   21350] = 32'haa44ffe7;
    ram_cell[   21351] = 32'h586fe76c;
    ram_cell[   21352] = 32'hdf6eadbb;
    ram_cell[   21353] = 32'hd315cf52;
    ram_cell[   21354] = 32'hb7dc0559;
    ram_cell[   21355] = 32'h28131c88;
    ram_cell[   21356] = 32'h7cc2c237;
    ram_cell[   21357] = 32'h430938c7;
    ram_cell[   21358] = 32'hb1d1f64f;
    ram_cell[   21359] = 32'h34f58743;
    ram_cell[   21360] = 32'h843da3f4;
    ram_cell[   21361] = 32'h7e21c39d;
    ram_cell[   21362] = 32'h0d3e206e;
    ram_cell[   21363] = 32'h7f2d1fdd;
    ram_cell[   21364] = 32'he5af9337;
    ram_cell[   21365] = 32'h1c411e19;
    ram_cell[   21366] = 32'hff9abbf7;
    ram_cell[   21367] = 32'h9a9f6c0f;
    ram_cell[   21368] = 32'h441f990c;
    ram_cell[   21369] = 32'h9d08e1cf;
    ram_cell[   21370] = 32'ha0b384bf;
    ram_cell[   21371] = 32'h6e5fb5f4;
    ram_cell[   21372] = 32'h5283965c;
    ram_cell[   21373] = 32'h01a95761;
    ram_cell[   21374] = 32'h6bdf98f6;
    ram_cell[   21375] = 32'h0b6b5f73;
    ram_cell[   21376] = 32'h8e6b20ad;
    ram_cell[   21377] = 32'h511ba542;
    ram_cell[   21378] = 32'he7e1a4f9;
    ram_cell[   21379] = 32'h7d59f1d9;
    ram_cell[   21380] = 32'h80cea8cb;
    ram_cell[   21381] = 32'h0843dfd0;
    ram_cell[   21382] = 32'h19a2e970;
    ram_cell[   21383] = 32'h40ee88e6;
    ram_cell[   21384] = 32'h44e8447d;
    ram_cell[   21385] = 32'he883a4d0;
    ram_cell[   21386] = 32'h6d51c897;
    ram_cell[   21387] = 32'h723574b0;
    ram_cell[   21388] = 32'h56ad8275;
    ram_cell[   21389] = 32'h456c90de;
    ram_cell[   21390] = 32'hb9ae874e;
    ram_cell[   21391] = 32'h49098f77;
    ram_cell[   21392] = 32'hc5747f17;
    ram_cell[   21393] = 32'hfd60a2b5;
    ram_cell[   21394] = 32'hcf37822b;
    ram_cell[   21395] = 32'h488c6d31;
    ram_cell[   21396] = 32'h0046600c;
    ram_cell[   21397] = 32'h08bcd5ae;
    ram_cell[   21398] = 32'he1bedea0;
    ram_cell[   21399] = 32'h05d10faa;
    ram_cell[   21400] = 32'h760721c1;
    ram_cell[   21401] = 32'hce2ca6f6;
    ram_cell[   21402] = 32'h70aeac3b;
    ram_cell[   21403] = 32'h02f9d24e;
    ram_cell[   21404] = 32'h9932047c;
    ram_cell[   21405] = 32'hbf3de21f;
    ram_cell[   21406] = 32'h2af1b1d4;
    ram_cell[   21407] = 32'hd58dbbd7;
    ram_cell[   21408] = 32'hef987d5c;
    ram_cell[   21409] = 32'hcb6e5e34;
    ram_cell[   21410] = 32'h0065ec90;
    ram_cell[   21411] = 32'h627b53cd;
    ram_cell[   21412] = 32'hb2149204;
    ram_cell[   21413] = 32'h53c5d9bd;
    ram_cell[   21414] = 32'h86f7a002;
    ram_cell[   21415] = 32'h98f71803;
    ram_cell[   21416] = 32'h7210562b;
    ram_cell[   21417] = 32'h6f7aefac;
    ram_cell[   21418] = 32'hf43f056b;
    ram_cell[   21419] = 32'he5b07068;
    ram_cell[   21420] = 32'hdfb4dae9;
    ram_cell[   21421] = 32'hd7069c22;
    ram_cell[   21422] = 32'hd61306ba;
    ram_cell[   21423] = 32'hd0c613be;
    ram_cell[   21424] = 32'hfe30e691;
    ram_cell[   21425] = 32'h2b99a2ae;
    ram_cell[   21426] = 32'hdc088dea;
    ram_cell[   21427] = 32'he144aded;
    ram_cell[   21428] = 32'h90d0085b;
    ram_cell[   21429] = 32'h86ba6277;
    ram_cell[   21430] = 32'hf84d9e6c;
    ram_cell[   21431] = 32'h8aa8078e;
    ram_cell[   21432] = 32'h00ece0b1;
    ram_cell[   21433] = 32'h2dd302b6;
    ram_cell[   21434] = 32'hfb5dcfc2;
    ram_cell[   21435] = 32'h88dffa28;
    ram_cell[   21436] = 32'h547cdece;
    ram_cell[   21437] = 32'he0093297;
    ram_cell[   21438] = 32'heac77cc3;
    ram_cell[   21439] = 32'hca11dedc;
    ram_cell[   21440] = 32'h162fac8d;
    ram_cell[   21441] = 32'hdd04f740;
    ram_cell[   21442] = 32'h465e419e;
    ram_cell[   21443] = 32'h773c7bc6;
    ram_cell[   21444] = 32'h6e3b8c12;
    ram_cell[   21445] = 32'h6260cb98;
    ram_cell[   21446] = 32'ha29f1cf7;
    ram_cell[   21447] = 32'h6d8f0779;
    ram_cell[   21448] = 32'h491c1b40;
    ram_cell[   21449] = 32'h5d3e9e40;
    ram_cell[   21450] = 32'h8fd53a1d;
    ram_cell[   21451] = 32'he70a66c3;
    ram_cell[   21452] = 32'h4e11c1c3;
    ram_cell[   21453] = 32'hd9e64ea2;
    ram_cell[   21454] = 32'h48f93f8a;
    ram_cell[   21455] = 32'hcf776ffb;
    ram_cell[   21456] = 32'h7d229f7d;
    ram_cell[   21457] = 32'h1c4fa3f8;
    ram_cell[   21458] = 32'hfd2a5c28;
    ram_cell[   21459] = 32'h45d6ad90;
    ram_cell[   21460] = 32'ha57c2ac6;
    ram_cell[   21461] = 32'h04a4e41a;
    ram_cell[   21462] = 32'hd06d58d4;
    ram_cell[   21463] = 32'h42b5e96c;
    ram_cell[   21464] = 32'hdcfc5d20;
    ram_cell[   21465] = 32'h8b7a88fa;
    ram_cell[   21466] = 32'hf276c122;
    ram_cell[   21467] = 32'h9cd1a64a;
    ram_cell[   21468] = 32'hdeb01fef;
    ram_cell[   21469] = 32'h626c368f;
    ram_cell[   21470] = 32'h779ce677;
    ram_cell[   21471] = 32'h32ed9a38;
    ram_cell[   21472] = 32'h82c27c59;
    ram_cell[   21473] = 32'hc1c2b022;
    ram_cell[   21474] = 32'h3d5a6e66;
    ram_cell[   21475] = 32'h8d67a038;
    ram_cell[   21476] = 32'h5ce4eaa7;
    ram_cell[   21477] = 32'hb6721684;
    ram_cell[   21478] = 32'hd2787e32;
    ram_cell[   21479] = 32'h4cd199d0;
    ram_cell[   21480] = 32'he6d81a77;
    ram_cell[   21481] = 32'ha32fd29b;
    ram_cell[   21482] = 32'he9206dbe;
    ram_cell[   21483] = 32'h57773b70;
    ram_cell[   21484] = 32'h4b88e266;
    ram_cell[   21485] = 32'he228708d;
    ram_cell[   21486] = 32'haad95938;
    ram_cell[   21487] = 32'h55a429b8;
    ram_cell[   21488] = 32'hf437b536;
    ram_cell[   21489] = 32'h6aedf1eb;
    ram_cell[   21490] = 32'h9707a975;
    ram_cell[   21491] = 32'hc590d25f;
    ram_cell[   21492] = 32'h3dbd5722;
    ram_cell[   21493] = 32'hbed15891;
    ram_cell[   21494] = 32'h79056b4e;
    ram_cell[   21495] = 32'h65089b02;
    ram_cell[   21496] = 32'hfd0a53bc;
    ram_cell[   21497] = 32'ha0bb2145;
    ram_cell[   21498] = 32'h824cfa39;
    ram_cell[   21499] = 32'h98d65aef;
    ram_cell[   21500] = 32'he7cfa3da;
    ram_cell[   21501] = 32'h6932f84c;
    ram_cell[   21502] = 32'h363f9692;
    ram_cell[   21503] = 32'h46068d10;
    ram_cell[   21504] = 32'h69d943ad;
    ram_cell[   21505] = 32'h7ab5a0c0;
    ram_cell[   21506] = 32'h0944e888;
    ram_cell[   21507] = 32'h9daeac97;
    ram_cell[   21508] = 32'h6f8f36bc;
    ram_cell[   21509] = 32'h77c0bc1b;
    ram_cell[   21510] = 32'hc1951dd2;
    ram_cell[   21511] = 32'ha8d1b37b;
    ram_cell[   21512] = 32'h5950fae2;
    ram_cell[   21513] = 32'h10c844b2;
    ram_cell[   21514] = 32'h20bcc689;
    ram_cell[   21515] = 32'h26013ef8;
    ram_cell[   21516] = 32'ha832da42;
    ram_cell[   21517] = 32'hafb98163;
    ram_cell[   21518] = 32'h0b8edae5;
    ram_cell[   21519] = 32'h98fc69a9;
    ram_cell[   21520] = 32'h22fa8d47;
    ram_cell[   21521] = 32'hc834cd68;
    ram_cell[   21522] = 32'hbcb26a13;
    ram_cell[   21523] = 32'h07f4bc23;
    ram_cell[   21524] = 32'h86ae81b0;
    ram_cell[   21525] = 32'h5421b92f;
    ram_cell[   21526] = 32'h9cdb8580;
    ram_cell[   21527] = 32'h75e5d03d;
    ram_cell[   21528] = 32'h28354586;
    ram_cell[   21529] = 32'h8d0c3bbe;
    ram_cell[   21530] = 32'h0e5d6d01;
    ram_cell[   21531] = 32'h16d6abb0;
    ram_cell[   21532] = 32'h01eab3dc;
    ram_cell[   21533] = 32'h69986e83;
    ram_cell[   21534] = 32'h8ef2e669;
    ram_cell[   21535] = 32'h1bdfcc41;
    ram_cell[   21536] = 32'h7e080a76;
    ram_cell[   21537] = 32'h167721ee;
    ram_cell[   21538] = 32'hbcff1b7a;
    ram_cell[   21539] = 32'h5011d52e;
    ram_cell[   21540] = 32'h47bc7674;
    ram_cell[   21541] = 32'h42b5cbc2;
    ram_cell[   21542] = 32'hf48318de;
    ram_cell[   21543] = 32'h326cfb97;
    ram_cell[   21544] = 32'hcc6f50b6;
    ram_cell[   21545] = 32'h073bc251;
    ram_cell[   21546] = 32'hefacb0c2;
    ram_cell[   21547] = 32'ha74d1138;
    ram_cell[   21548] = 32'h1266c453;
    ram_cell[   21549] = 32'h0bcd37fe;
    ram_cell[   21550] = 32'he439982d;
    ram_cell[   21551] = 32'ha0df4205;
    ram_cell[   21552] = 32'heb331400;
    ram_cell[   21553] = 32'h7b07aed5;
    ram_cell[   21554] = 32'he87a4f98;
    ram_cell[   21555] = 32'he1f4e66f;
    ram_cell[   21556] = 32'hbd34e151;
    ram_cell[   21557] = 32'hbc5caafb;
    ram_cell[   21558] = 32'h0347ba00;
    ram_cell[   21559] = 32'hdf6bf02e;
    ram_cell[   21560] = 32'hccf03926;
    ram_cell[   21561] = 32'h43f63e78;
    ram_cell[   21562] = 32'hdcc96c7c;
    ram_cell[   21563] = 32'hd08ba3f4;
    ram_cell[   21564] = 32'h1949af62;
    ram_cell[   21565] = 32'h6b29eec8;
    ram_cell[   21566] = 32'h5c054698;
    ram_cell[   21567] = 32'h940a6a06;
    ram_cell[   21568] = 32'h8e71aed9;
    ram_cell[   21569] = 32'h727e4427;
    ram_cell[   21570] = 32'h994d5fca;
    ram_cell[   21571] = 32'h4b2d4e94;
    ram_cell[   21572] = 32'hc676581d;
    ram_cell[   21573] = 32'h5461e06d;
    ram_cell[   21574] = 32'h1d0f4710;
    ram_cell[   21575] = 32'haf80d413;
    ram_cell[   21576] = 32'h3751c92b;
    ram_cell[   21577] = 32'h2bcc518c;
    ram_cell[   21578] = 32'hd1c70783;
    ram_cell[   21579] = 32'ha1c51170;
    ram_cell[   21580] = 32'hb8a4e0bd;
    ram_cell[   21581] = 32'h9d4503eb;
    ram_cell[   21582] = 32'hce59093f;
    ram_cell[   21583] = 32'h75a85cd1;
    ram_cell[   21584] = 32'hebc3dc60;
    ram_cell[   21585] = 32'hc5abe67a;
    ram_cell[   21586] = 32'h1a2e9b48;
    ram_cell[   21587] = 32'hda357426;
    ram_cell[   21588] = 32'hdc5a2236;
    ram_cell[   21589] = 32'h818126f9;
    ram_cell[   21590] = 32'h2dc07b26;
    ram_cell[   21591] = 32'h430add37;
    ram_cell[   21592] = 32'h3bb65f34;
    ram_cell[   21593] = 32'haae0b942;
    ram_cell[   21594] = 32'h0f19923b;
    ram_cell[   21595] = 32'h954c40c6;
    ram_cell[   21596] = 32'h3ba95151;
    ram_cell[   21597] = 32'h37c23d41;
    ram_cell[   21598] = 32'hf9155a34;
    ram_cell[   21599] = 32'h5798b580;
    ram_cell[   21600] = 32'h0d473d34;
    ram_cell[   21601] = 32'h0789a24b;
    ram_cell[   21602] = 32'hc4bf7b7d;
    ram_cell[   21603] = 32'hc7c7195b;
    ram_cell[   21604] = 32'haed47648;
    ram_cell[   21605] = 32'h5266b8d6;
    ram_cell[   21606] = 32'h9ce864ff;
    ram_cell[   21607] = 32'h09a5e456;
    ram_cell[   21608] = 32'h4263a7e0;
    ram_cell[   21609] = 32'hb37efb31;
    ram_cell[   21610] = 32'h7c2576a2;
    ram_cell[   21611] = 32'h1901b02a;
    ram_cell[   21612] = 32'hcab0322d;
    ram_cell[   21613] = 32'h69303718;
    ram_cell[   21614] = 32'h8c05a367;
    ram_cell[   21615] = 32'hc0dc3b10;
    ram_cell[   21616] = 32'h789b1863;
    ram_cell[   21617] = 32'h5b91fa25;
    ram_cell[   21618] = 32'hbfbc0bc3;
    ram_cell[   21619] = 32'he69fe5c1;
    ram_cell[   21620] = 32'h12b36608;
    ram_cell[   21621] = 32'he07b7aab;
    ram_cell[   21622] = 32'h5459dcf1;
    ram_cell[   21623] = 32'h21d61779;
    ram_cell[   21624] = 32'hdf70a02d;
    ram_cell[   21625] = 32'hc95bf840;
    ram_cell[   21626] = 32'hbcec37fa;
    ram_cell[   21627] = 32'he4d962bc;
    ram_cell[   21628] = 32'he477f309;
    ram_cell[   21629] = 32'hf709453c;
    ram_cell[   21630] = 32'hd0121e96;
    ram_cell[   21631] = 32'ha9fe0c1b;
    ram_cell[   21632] = 32'h9db304ab;
    ram_cell[   21633] = 32'ha55ec3bd;
    ram_cell[   21634] = 32'h0bcce837;
    ram_cell[   21635] = 32'hd61fd77e;
    ram_cell[   21636] = 32'h1f84fe95;
    ram_cell[   21637] = 32'h37fc4b2c;
    ram_cell[   21638] = 32'hdb09bbea;
    ram_cell[   21639] = 32'h0ba21a5e;
    ram_cell[   21640] = 32'h20815c45;
    ram_cell[   21641] = 32'ha47d0eae;
    ram_cell[   21642] = 32'h2dd15f4c;
    ram_cell[   21643] = 32'hb3a377f0;
    ram_cell[   21644] = 32'h0ffcffd3;
    ram_cell[   21645] = 32'h6e468bcf;
    ram_cell[   21646] = 32'hf9f50416;
    ram_cell[   21647] = 32'h20c98b28;
    ram_cell[   21648] = 32'h28bba78f;
    ram_cell[   21649] = 32'h80ca56fd;
    ram_cell[   21650] = 32'h92bd2967;
    ram_cell[   21651] = 32'hb5c9483b;
    ram_cell[   21652] = 32'hcc80598b;
    ram_cell[   21653] = 32'h1191f47a;
    ram_cell[   21654] = 32'h79ac6787;
    ram_cell[   21655] = 32'h20f247a9;
    ram_cell[   21656] = 32'hd689040d;
    ram_cell[   21657] = 32'h1752859b;
    ram_cell[   21658] = 32'h554abae3;
    ram_cell[   21659] = 32'hb198e4fc;
    ram_cell[   21660] = 32'h2982ad31;
    ram_cell[   21661] = 32'hbd31120e;
    ram_cell[   21662] = 32'h05231500;
    ram_cell[   21663] = 32'h072a4b36;
    ram_cell[   21664] = 32'ha46d0664;
    ram_cell[   21665] = 32'h6e1f1007;
    ram_cell[   21666] = 32'h75c4ba7d;
    ram_cell[   21667] = 32'hc7801a07;
    ram_cell[   21668] = 32'hc90e2c95;
    ram_cell[   21669] = 32'h3852882d;
    ram_cell[   21670] = 32'hc868c319;
    ram_cell[   21671] = 32'hc4a4f18e;
    ram_cell[   21672] = 32'he3fc4fb0;
    ram_cell[   21673] = 32'h15279dbe;
    ram_cell[   21674] = 32'h797d204e;
    ram_cell[   21675] = 32'hafa60976;
    ram_cell[   21676] = 32'h331dfc30;
    ram_cell[   21677] = 32'hc8011298;
    ram_cell[   21678] = 32'h45df2fbc;
    ram_cell[   21679] = 32'h8176337b;
    ram_cell[   21680] = 32'he7887f55;
    ram_cell[   21681] = 32'h80d9633a;
    ram_cell[   21682] = 32'hbbad22aa;
    ram_cell[   21683] = 32'h21c8cdd1;
    ram_cell[   21684] = 32'hff9168e9;
    ram_cell[   21685] = 32'h7db90c8e;
    ram_cell[   21686] = 32'he6e6b064;
    ram_cell[   21687] = 32'h3220909a;
    ram_cell[   21688] = 32'ha16dcafc;
    ram_cell[   21689] = 32'h8c103aa5;
    ram_cell[   21690] = 32'h70407d17;
    ram_cell[   21691] = 32'hbf215775;
    ram_cell[   21692] = 32'heeec15bb;
    ram_cell[   21693] = 32'haf08a619;
    ram_cell[   21694] = 32'hd8598ea0;
    ram_cell[   21695] = 32'h95afb479;
    ram_cell[   21696] = 32'h2871b98c;
    ram_cell[   21697] = 32'h2aefa96e;
    ram_cell[   21698] = 32'hb7b6164e;
    ram_cell[   21699] = 32'h9aa3fd84;
    ram_cell[   21700] = 32'hb419ae29;
    ram_cell[   21701] = 32'h3bc43b01;
    ram_cell[   21702] = 32'he3f3c17c;
    ram_cell[   21703] = 32'hfb36f2a1;
    ram_cell[   21704] = 32'hcfb2824a;
    ram_cell[   21705] = 32'h467c7ad8;
    ram_cell[   21706] = 32'h4ad2ff30;
    ram_cell[   21707] = 32'h1efa1b2a;
    ram_cell[   21708] = 32'hc8cf26b8;
    ram_cell[   21709] = 32'h5550d5ea;
    ram_cell[   21710] = 32'h12f4e162;
    ram_cell[   21711] = 32'h07ab3aec;
    ram_cell[   21712] = 32'h2f45e122;
    ram_cell[   21713] = 32'h2e1a3913;
    ram_cell[   21714] = 32'h02b20fae;
    ram_cell[   21715] = 32'h9540abca;
    ram_cell[   21716] = 32'hdf97e7e7;
    ram_cell[   21717] = 32'h035a8640;
    ram_cell[   21718] = 32'hdd608a4b;
    ram_cell[   21719] = 32'h3e7455d5;
    ram_cell[   21720] = 32'h497666eb;
    ram_cell[   21721] = 32'h580decaf;
    ram_cell[   21722] = 32'hc965d398;
    ram_cell[   21723] = 32'h6970cfb0;
    ram_cell[   21724] = 32'h68d67b81;
    ram_cell[   21725] = 32'h353761a9;
    ram_cell[   21726] = 32'he52a4f88;
    ram_cell[   21727] = 32'hf2735296;
    ram_cell[   21728] = 32'h327db441;
    ram_cell[   21729] = 32'h94c3977b;
    ram_cell[   21730] = 32'h562e7cf9;
    ram_cell[   21731] = 32'h797c95d7;
    ram_cell[   21732] = 32'hc40da67e;
    ram_cell[   21733] = 32'h9a40a685;
    ram_cell[   21734] = 32'h715a249d;
    ram_cell[   21735] = 32'h6dd5c440;
    ram_cell[   21736] = 32'h61296a39;
    ram_cell[   21737] = 32'h2111be7f;
    ram_cell[   21738] = 32'h5b13e569;
    ram_cell[   21739] = 32'h3ce35dbe;
    ram_cell[   21740] = 32'h3f6e837d;
    ram_cell[   21741] = 32'h9c5b642d;
    ram_cell[   21742] = 32'h16d11af9;
    ram_cell[   21743] = 32'h1073f435;
    ram_cell[   21744] = 32'he2cae853;
    ram_cell[   21745] = 32'h4078da7d;
    ram_cell[   21746] = 32'h5b2f9b7b;
    ram_cell[   21747] = 32'ha15c4fa1;
    ram_cell[   21748] = 32'h614f8a55;
    ram_cell[   21749] = 32'h97647fb1;
    ram_cell[   21750] = 32'h79bae8f9;
    ram_cell[   21751] = 32'ha7d48c9b;
    ram_cell[   21752] = 32'h44d7685b;
    ram_cell[   21753] = 32'h0a8e54d7;
    ram_cell[   21754] = 32'h5ea65cc0;
    ram_cell[   21755] = 32'h755c4405;
    ram_cell[   21756] = 32'h4de5e836;
    ram_cell[   21757] = 32'h6b3533a9;
    ram_cell[   21758] = 32'h80f14bce;
    ram_cell[   21759] = 32'h2526b7d8;
    ram_cell[   21760] = 32'h0e6ac78b;
    ram_cell[   21761] = 32'h1e9a00c2;
    ram_cell[   21762] = 32'h09fb8608;
    ram_cell[   21763] = 32'ha8a38f87;
    ram_cell[   21764] = 32'h39659ac2;
    ram_cell[   21765] = 32'hd0a422ed;
    ram_cell[   21766] = 32'h567a9688;
    ram_cell[   21767] = 32'heb3f0516;
    ram_cell[   21768] = 32'h34b20cb9;
    ram_cell[   21769] = 32'h902d08c5;
    ram_cell[   21770] = 32'h591e58e7;
    ram_cell[   21771] = 32'h19305e6f;
    ram_cell[   21772] = 32'hc8d26a93;
    ram_cell[   21773] = 32'hde9ded55;
    ram_cell[   21774] = 32'h9be15cb9;
    ram_cell[   21775] = 32'h51124db1;
    ram_cell[   21776] = 32'h4f2d453a;
    ram_cell[   21777] = 32'h8a9906f3;
    ram_cell[   21778] = 32'h828533dc;
    ram_cell[   21779] = 32'h1e967785;
    ram_cell[   21780] = 32'hcc981c52;
    ram_cell[   21781] = 32'hedd73852;
    ram_cell[   21782] = 32'h4bf732c2;
    ram_cell[   21783] = 32'hf0020a26;
    ram_cell[   21784] = 32'hd7d88ceb;
    ram_cell[   21785] = 32'he132b342;
    ram_cell[   21786] = 32'hc056afc6;
    ram_cell[   21787] = 32'hc017095e;
    ram_cell[   21788] = 32'h8d6f4058;
    ram_cell[   21789] = 32'h81579158;
    ram_cell[   21790] = 32'h738ca4c1;
    ram_cell[   21791] = 32'h5ee83a52;
    ram_cell[   21792] = 32'h763d76aa;
    ram_cell[   21793] = 32'ha0e9dae8;
    ram_cell[   21794] = 32'hf0f129e0;
    ram_cell[   21795] = 32'hb824d3a4;
    ram_cell[   21796] = 32'hc07dd5df;
    ram_cell[   21797] = 32'hf9366466;
    ram_cell[   21798] = 32'h6aa4e09b;
    ram_cell[   21799] = 32'h06e5d5e2;
    ram_cell[   21800] = 32'hc7679d37;
    ram_cell[   21801] = 32'hf44b8349;
    ram_cell[   21802] = 32'h96a6917b;
    ram_cell[   21803] = 32'h7fc31c28;
    ram_cell[   21804] = 32'h0b7c092d;
    ram_cell[   21805] = 32'hce4e7d8e;
    ram_cell[   21806] = 32'hb493f6c4;
    ram_cell[   21807] = 32'h53edb578;
    ram_cell[   21808] = 32'h6647e4f1;
    ram_cell[   21809] = 32'hf6a7b23e;
    ram_cell[   21810] = 32'h3a38aaac;
    ram_cell[   21811] = 32'h01491834;
    ram_cell[   21812] = 32'h1557e635;
    ram_cell[   21813] = 32'h45f7bfc0;
    ram_cell[   21814] = 32'h37258fde;
    ram_cell[   21815] = 32'h08b71f49;
    ram_cell[   21816] = 32'h799cb2d0;
    ram_cell[   21817] = 32'h32515a3b;
    ram_cell[   21818] = 32'h3ae0ad85;
    ram_cell[   21819] = 32'h1d645950;
    ram_cell[   21820] = 32'h7178903c;
    ram_cell[   21821] = 32'hb775038c;
    ram_cell[   21822] = 32'he38cf46a;
    ram_cell[   21823] = 32'hbd1f0dbf;
    ram_cell[   21824] = 32'hd790ab90;
    ram_cell[   21825] = 32'h2dea1835;
    ram_cell[   21826] = 32'h2da833ef;
    ram_cell[   21827] = 32'ha6ec3e04;
    ram_cell[   21828] = 32'hc351bb35;
    ram_cell[   21829] = 32'h513b802a;
    ram_cell[   21830] = 32'hcb9f524a;
    ram_cell[   21831] = 32'h9a6bdbd1;
    ram_cell[   21832] = 32'hbe1dfdd7;
    ram_cell[   21833] = 32'hbf04c4f6;
    ram_cell[   21834] = 32'hc25224d0;
    ram_cell[   21835] = 32'h0da6438d;
    ram_cell[   21836] = 32'h53e47f53;
    ram_cell[   21837] = 32'h34db31be;
    ram_cell[   21838] = 32'he64e3ba5;
    ram_cell[   21839] = 32'h364c4dad;
    ram_cell[   21840] = 32'hdfc00ab1;
    ram_cell[   21841] = 32'hfcfc0687;
    ram_cell[   21842] = 32'h3cd5fc54;
    ram_cell[   21843] = 32'h2898664a;
    ram_cell[   21844] = 32'hd4653083;
    ram_cell[   21845] = 32'h42c94004;
    ram_cell[   21846] = 32'h8385a9ec;
    ram_cell[   21847] = 32'hd9d171df;
    ram_cell[   21848] = 32'hb2069b6d;
    ram_cell[   21849] = 32'h2b77b35a;
    ram_cell[   21850] = 32'h2a26b2ce;
    ram_cell[   21851] = 32'hf50b1134;
    ram_cell[   21852] = 32'h2da460a0;
    ram_cell[   21853] = 32'h70888186;
    ram_cell[   21854] = 32'h1c1cc2bd;
    ram_cell[   21855] = 32'ha59151ef;
    ram_cell[   21856] = 32'h94e7c953;
    ram_cell[   21857] = 32'h052da0de;
    ram_cell[   21858] = 32'h3ac8c689;
    ram_cell[   21859] = 32'h4aaeef6a;
    ram_cell[   21860] = 32'h8c873674;
    ram_cell[   21861] = 32'h6b5b2dac;
    ram_cell[   21862] = 32'h4aa2504c;
    ram_cell[   21863] = 32'h9dbe1d31;
    ram_cell[   21864] = 32'h025054b1;
    ram_cell[   21865] = 32'h9302c260;
    ram_cell[   21866] = 32'h3dbe65e8;
    ram_cell[   21867] = 32'hf0a84146;
    ram_cell[   21868] = 32'h116e4acf;
    ram_cell[   21869] = 32'h6cd6f666;
    ram_cell[   21870] = 32'h1db5c3f9;
    ram_cell[   21871] = 32'hdf32e932;
    ram_cell[   21872] = 32'h740b8d41;
    ram_cell[   21873] = 32'hc70bc307;
    ram_cell[   21874] = 32'h77f40748;
    ram_cell[   21875] = 32'hd88524f7;
    ram_cell[   21876] = 32'h5ae801d9;
    ram_cell[   21877] = 32'hed64cee3;
    ram_cell[   21878] = 32'h78143095;
    ram_cell[   21879] = 32'hd73901bb;
    ram_cell[   21880] = 32'haaf42404;
    ram_cell[   21881] = 32'he97987b7;
    ram_cell[   21882] = 32'h0dd1f5fb;
    ram_cell[   21883] = 32'h8ebde3e3;
    ram_cell[   21884] = 32'h34061c51;
    ram_cell[   21885] = 32'h10b9ec57;
    ram_cell[   21886] = 32'hded54ab2;
    ram_cell[   21887] = 32'h1854f3ae;
    ram_cell[   21888] = 32'h874a48a9;
    ram_cell[   21889] = 32'h8cd9cedd;
    ram_cell[   21890] = 32'h75fc0f5b;
    ram_cell[   21891] = 32'ha3042c00;
    ram_cell[   21892] = 32'h86991756;
    ram_cell[   21893] = 32'hfdfe1b7c;
    ram_cell[   21894] = 32'h3a84c56e;
    ram_cell[   21895] = 32'hd7457789;
    ram_cell[   21896] = 32'h8b70f62f;
    ram_cell[   21897] = 32'hd2c4998e;
    ram_cell[   21898] = 32'hed534ec7;
    ram_cell[   21899] = 32'h2cafb860;
    ram_cell[   21900] = 32'h16f31645;
    ram_cell[   21901] = 32'hef07b609;
    ram_cell[   21902] = 32'he6c626f0;
    ram_cell[   21903] = 32'h6a7a6e27;
    ram_cell[   21904] = 32'h9d6e16b0;
    ram_cell[   21905] = 32'hddc820cd;
    ram_cell[   21906] = 32'h2a2033ef;
    ram_cell[   21907] = 32'hba0b40dc;
    ram_cell[   21908] = 32'h40e86966;
    ram_cell[   21909] = 32'h8ed87491;
    ram_cell[   21910] = 32'h7f320b3e;
    ram_cell[   21911] = 32'h6a883820;
    ram_cell[   21912] = 32'h7d931f8c;
    ram_cell[   21913] = 32'h2677e556;
    ram_cell[   21914] = 32'h9818f335;
    ram_cell[   21915] = 32'h14719d32;
    ram_cell[   21916] = 32'hb8dd28f9;
    ram_cell[   21917] = 32'h9f98d57e;
    ram_cell[   21918] = 32'h7ba66774;
    ram_cell[   21919] = 32'h7d59a353;
    ram_cell[   21920] = 32'h6ef993d2;
    ram_cell[   21921] = 32'h47eefa5c;
    ram_cell[   21922] = 32'h07cda280;
    ram_cell[   21923] = 32'h1a8bab41;
    ram_cell[   21924] = 32'h5440f6fa;
    ram_cell[   21925] = 32'h69885c2c;
    ram_cell[   21926] = 32'h4391ea21;
    ram_cell[   21927] = 32'hc2d91c45;
    ram_cell[   21928] = 32'h2fe3aedd;
    ram_cell[   21929] = 32'hd61a1503;
    ram_cell[   21930] = 32'hb048ecb8;
    ram_cell[   21931] = 32'h828b71a2;
    ram_cell[   21932] = 32'h5916ad35;
    ram_cell[   21933] = 32'h2af5adab;
    ram_cell[   21934] = 32'h4d535388;
    ram_cell[   21935] = 32'h431a0037;
    ram_cell[   21936] = 32'h03e5a4be;
    ram_cell[   21937] = 32'h2c7cb3f3;
    ram_cell[   21938] = 32'h86e118b4;
    ram_cell[   21939] = 32'he67a4506;
    ram_cell[   21940] = 32'h44a13d6c;
    ram_cell[   21941] = 32'he53cbd4a;
    ram_cell[   21942] = 32'h516100dd;
    ram_cell[   21943] = 32'ha778bd66;
    ram_cell[   21944] = 32'h5bd123c3;
    ram_cell[   21945] = 32'hc94450af;
    ram_cell[   21946] = 32'h04a49306;
    ram_cell[   21947] = 32'h0b0ec9e0;
    ram_cell[   21948] = 32'hd80f14ba;
    ram_cell[   21949] = 32'he99b7d4d;
    ram_cell[   21950] = 32'h0d3ef261;
    ram_cell[   21951] = 32'h85827488;
    ram_cell[   21952] = 32'h071d3d6b;
    ram_cell[   21953] = 32'h25aadbac;
    ram_cell[   21954] = 32'h856dd3b6;
    ram_cell[   21955] = 32'h30893e2a;
    ram_cell[   21956] = 32'h7fabc011;
    ram_cell[   21957] = 32'h15020f7f;
    ram_cell[   21958] = 32'h927cdf43;
    ram_cell[   21959] = 32'h30849b01;
    ram_cell[   21960] = 32'h18ac00d0;
    ram_cell[   21961] = 32'h93a87546;
    ram_cell[   21962] = 32'h24493200;
    ram_cell[   21963] = 32'h70bf59e4;
    ram_cell[   21964] = 32'h11aade16;
    ram_cell[   21965] = 32'h8a3f4f30;
    ram_cell[   21966] = 32'h4bff65eb;
    ram_cell[   21967] = 32'h0979aa3f;
    ram_cell[   21968] = 32'hbf126463;
    ram_cell[   21969] = 32'h2f3fc525;
    ram_cell[   21970] = 32'h549e86ad;
    ram_cell[   21971] = 32'h760e8bf6;
    ram_cell[   21972] = 32'h073d035b;
    ram_cell[   21973] = 32'hd7b37e1d;
    ram_cell[   21974] = 32'hf78b0ab0;
    ram_cell[   21975] = 32'h0ce0de33;
    ram_cell[   21976] = 32'hba8faef6;
    ram_cell[   21977] = 32'hbe60dc96;
    ram_cell[   21978] = 32'h73b5d737;
    ram_cell[   21979] = 32'h77e93ec7;
    ram_cell[   21980] = 32'hf1e07468;
    ram_cell[   21981] = 32'h1f43f4eb;
    ram_cell[   21982] = 32'h759886e5;
    ram_cell[   21983] = 32'h8ecfc992;
    ram_cell[   21984] = 32'h32589e56;
    ram_cell[   21985] = 32'h13ac1a84;
    ram_cell[   21986] = 32'hdbd50bcd;
    ram_cell[   21987] = 32'hb4950e46;
    ram_cell[   21988] = 32'hf91083cd;
    ram_cell[   21989] = 32'hebc938a3;
    ram_cell[   21990] = 32'he7e53572;
    ram_cell[   21991] = 32'h1812c44d;
    ram_cell[   21992] = 32'ha2598d39;
    ram_cell[   21993] = 32'h93d2a736;
    ram_cell[   21994] = 32'h600a70c5;
    ram_cell[   21995] = 32'h120af498;
    ram_cell[   21996] = 32'hc3b416ab;
    ram_cell[   21997] = 32'h891a4270;
    ram_cell[   21998] = 32'h56b4085f;
    ram_cell[   21999] = 32'hffa686a6;
    ram_cell[   22000] = 32'h4e67416c;
    ram_cell[   22001] = 32'h99d82b35;
    ram_cell[   22002] = 32'h7d1b4d0b;
    ram_cell[   22003] = 32'hacc13da9;
    ram_cell[   22004] = 32'h807544c4;
    ram_cell[   22005] = 32'h3a6fbeeb;
    ram_cell[   22006] = 32'hd55bc80d;
    ram_cell[   22007] = 32'h356fd303;
    ram_cell[   22008] = 32'hf17f4176;
    ram_cell[   22009] = 32'h6a8ccad6;
    ram_cell[   22010] = 32'h6e99d8bb;
    ram_cell[   22011] = 32'hac4c15c8;
    ram_cell[   22012] = 32'h20f78808;
    ram_cell[   22013] = 32'h2cfe54c5;
    ram_cell[   22014] = 32'h19a7f432;
    ram_cell[   22015] = 32'h5777a580;
    ram_cell[   22016] = 32'hdd5a2282;
    ram_cell[   22017] = 32'hc212ed51;
    ram_cell[   22018] = 32'h04977ced;
    ram_cell[   22019] = 32'hd3df5b2e;
    ram_cell[   22020] = 32'h7274dc1d;
    ram_cell[   22021] = 32'hfe393a34;
    ram_cell[   22022] = 32'h15eed566;
    ram_cell[   22023] = 32'h25a96fcc;
    ram_cell[   22024] = 32'h2b0b4134;
    ram_cell[   22025] = 32'hc438e60e;
    ram_cell[   22026] = 32'h8256a1cf;
    ram_cell[   22027] = 32'h4a09c86e;
    ram_cell[   22028] = 32'h1f67dee0;
    ram_cell[   22029] = 32'hb91b5d79;
    ram_cell[   22030] = 32'hd66fcdfb;
    ram_cell[   22031] = 32'hf6f81866;
    ram_cell[   22032] = 32'h60857ede;
    ram_cell[   22033] = 32'h744ed60b;
    ram_cell[   22034] = 32'hceea01b3;
    ram_cell[   22035] = 32'h296677e7;
    ram_cell[   22036] = 32'h4288b68d;
    ram_cell[   22037] = 32'h77a8c002;
    ram_cell[   22038] = 32'h8b599573;
    ram_cell[   22039] = 32'hb9466780;
    ram_cell[   22040] = 32'h204412ce;
    ram_cell[   22041] = 32'h47301c57;
    ram_cell[   22042] = 32'h3f5a8635;
    ram_cell[   22043] = 32'h5dd00be0;
    ram_cell[   22044] = 32'h2ae49b81;
    ram_cell[   22045] = 32'ha01741ca;
    ram_cell[   22046] = 32'h9e9f4d28;
    ram_cell[   22047] = 32'h158b6807;
    ram_cell[   22048] = 32'h04ae16b6;
    ram_cell[   22049] = 32'hfbe18b42;
    ram_cell[   22050] = 32'h334c4fe7;
    ram_cell[   22051] = 32'h49829009;
    ram_cell[   22052] = 32'h92d5ebab;
    ram_cell[   22053] = 32'h782319e3;
    ram_cell[   22054] = 32'h4575b373;
    ram_cell[   22055] = 32'h6579ea01;
    ram_cell[   22056] = 32'hf9d8db9e;
    ram_cell[   22057] = 32'h870718ed;
    ram_cell[   22058] = 32'h98052930;
    ram_cell[   22059] = 32'h4ba8b036;
    ram_cell[   22060] = 32'he585898d;
    ram_cell[   22061] = 32'h04aa7d5d;
    ram_cell[   22062] = 32'h4d02ba09;
    ram_cell[   22063] = 32'h5cb5a8e1;
    ram_cell[   22064] = 32'h17aa6278;
    ram_cell[   22065] = 32'h9f1445af;
    ram_cell[   22066] = 32'h61d7b730;
    ram_cell[   22067] = 32'hbc693115;
    ram_cell[   22068] = 32'h66fc91e5;
    ram_cell[   22069] = 32'h14c60588;
    ram_cell[   22070] = 32'hdfc1baad;
    ram_cell[   22071] = 32'h7d3e8b6d;
    ram_cell[   22072] = 32'h8d89ad44;
    ram_cell[   22073] = 32'hb4d84f2f;
    ram_cell[   22074] = 32'hf517e6fb;
    ram_cell[   22075] = 32'h31949afd;
    ram_cell[   22076] = 32'h3d990e75;
    ram_cell[   22077] = 32'h5655573f;
    ram_cell[   22078] = 32'h9074a6f0;
    ram_cell[   22079] = 32'h88f865a5;
    ram_cell[   22080] = 32'h61853034;
    ram_cell[   22081] = 32'he514251d;
    ram_cell[   22082] = 32'h7601c9a4;
    ram_cell[   22083] = 32'h1f04ead8;
    ram_cell[   22084] = 32'h35c36f97;
    ram_cell[   22085] = 32'hce637ed2;
    ram_cell[   22086] = 32'he6829aa2;
    ram_cell[   22087] = 32'hebaf7b29;
    ram_cell[   22088] = 32'hf9170fbe;
    ram_cell[   22089] = 32'h95b4de6c;
    ram_cell[   22090] = 32'hbd77a401;
    ram_cell[   22091] = 32'h3379deb4;
    ram_cell[   22092] = 32'h3a724c09;
    ram_cell[   22093] = 32'h30cc1cff;
    ram_cell[   22094] = 32'h557131d5;
    ram_cell[   22095] = 32'h8ffb372b;
    ram_cell[   22096] = 32'h25eb8b9b;
    ram_cell[   22097] = 32'hc9cc90f9;
    ram_cell[   22098] = 32'h9e60851d;
    ram_cell[   22099] = 32'hef24dc2d;
    ram_cell[   22100] = 32'h5cb65009;
    ram_cell[   22101] = 32'h7e5bd54e;
    ram_cell[   22102] = 32'h7786a9c1;
    ram_cell[   22103] = 32'h97212886;
    ram_cell[   22104] = 32'h4bc7289f;
    ram_cell[   22105] = 32'ha7475328;
    ram_cell[   22106] = 32'hcc686345;
    ram_cell[   22107] = 32'he2423d1b;
    ram_cell[   22108] = 32'h0403340e;
    ram_cell[   22109] = 32'h29fcdc0e;
    ram_cell[   22110] = 32'h08307133;
    ram_cell[   22111] = 32'h5eb83cd4;
    ram_cell[   22112] = 32'h39793c19;
    ram_cell[   22113] = 32'h327d7a43;
    ram_cell[   22114] = 32'h5bb4f2e7;
    ram_cell[   22115] = 32'hed749576;
    ram_cell[   22116] = 32'h63a8f817;
    ram_cell[   22117] = 32'h1792e433;
    ram_cell[   22118] = 32'ha0f1e785;
    ram_cell[   22119] = 32'h0b1ff938;
    ram_cell[   22120] = 32'h3a2c2dc6;
    ram_cell[   22121] = 32'hf28e5c14;
    ram_cell[   22122] = 32'h8191738c;
    ram_cell[   22123] = 32'hc430ca9b;
    ram_cell[   22124] = 32'h19658add;
    ram_cell[   22125] = 32'h0c555068;
    ram_cell[   22126] = 32'h96b256e5;
    ram_cell[   22127] = 32'h11a331e4;
    ram_cell[   22128] = 32'h62498a8a;
    ram_cell[   22129] = 32'hb44c8703;
    ram_cell[   22130] = 32'h52d4a135;
    ram_cell[   22131] = 32'he27e430d;
    ram_cell[   22132] = 32'hbe0947e8;
    ram_cell[   22133] = 32'hafb5e248;
    ram_cell[   22134] = 32'h602de2d4;
    ram_cell[   22135] = 32'h852c56e8;
    ram_cell[   22136] = 32'h1e74ee03;
    ram_cell[   22137] = 32'hf949b9cf;
    ram_cell[   22138] = 32'he40d126a;
    ram_cell[   22139] = 32'h7060569e;
    ram_cell[   22140] = 32'hea098d79;
    ram_cell[   22141] = 32'h1daa890e;
    ram_cell[   22142] = 32'h14114c35;
    ram_cell[   22143] = 32'h8eec9e02;
    ram_cell[   22144] = 32'hc6913d8d;
    ram_cell[   22145] = 32'h20ee0d77;
    ram_cell[   22146] = 32'h98c5aad6;
    ram_cell[   22147] = 32'h8f3ac301;
    ram_cell[   22148] = 32'h8b6147ba;
    ram_cell[   22149] = 32'ha4c4d03f;
    ram_cell[   22150] = 32'h4590687f;
    ram_cell[   22151] = 32'he2ede9c3;
    ram_cell[   22152] = 32'h3fda5ccd;
    ram_cell[   22153] = 32'h8bfefdf0;
    ram_cell[   22154] = 32'h608d00a7;
    ram_cell[   22155] = 32'ha8f17bdf;
    ram_cell[   22156] = 32'h02b9f69e;
    ram_cell[   22157] = 32'h7f5fbdde;
    ram_cell[   22158] = 32'hfea6a214;
    ram_cell[   22159] = 32'h9bba532c;
    ram_cell[   22160] = 32'h71228119;
    ram_cell[   22161] = 32'h867876b6;
    ram_cell[   22162] = 32'hf18d6158;
    ram_cell[   22163] = 32'hbce4cd04;
    ram_cell[   22164] = 32'h80e3a885;
    ram_cell[   22165] = 32'hfee7d5ca;
    ram_cell[   22166] = 32'h49e603b7;
    ram_cell[   22167] = 32'h0bf7dea1;
    ram_cell[   22168] = 32'h9b409226;
    ram_cell[   22169] = 32'hf5924385;
    ram_cell[   22170] = 32'h199b5233;
    ram_cell[   22171] = 32'h0afddb6f;
    ram_cell[   22172] = 32'h4b1739f0;
    ram_cell[   22173] = 32'h688c4d87;
    ram_cell[   22174] = 32'h82ec8115;
    ram_cell[   22175] = 32'h94a53644;
    ram_cell[   22176] = 32'hcdf53231;
    ram_cell[   22177] = 32'hc546d12e;
    ram_cell[   22178] = 32'h6d9b6b46;
    ram_cell[   22179] = 32'h36531674;
    ram_cell[   22180] = 32'h3f8bb772;
    ram_cell[   22181] = 32'hfea1e93b;
    ram_cell[   22182] = 32'h53d54254;
    ram_cell[   22183] = 32'hb1cabca3;
    ram_cell[   22184] = 32'hb840c4b3;
    ram_cell[   22185] = 32'h2ea5fc08;
    ram_cell[   22186] = 32'h5076392e;
    ram_cell[   22187] = 32'h21c40750;
    ram_cell[   22188] = 32'h4aded64b;
    ram_cell[   22189] = 32'hbaf6abbc;
    ram_cell[   22190] = 32'h74a98f81;
    ram_cell[   22191] = 32'h89ce8605;
    ram_cell[   22192] = 32'h456a2b53;
    ram_cell[   22193] = 32'hec6120d9;
    ram_cell[   22194] = 32'h6226a700;
    ram_cell[   22195] = 32'hff6a9f78;
    ram_cell[   22196] = 32'h288dac93;
    ram_cell[   22197] = 32'h2e9cf2d2;
    ram_cell[   22198] = 32'h7f72661c;
    ram_cell[   22199] = 32'hb1e5aa4c;
    ram_cell[   22200] = 32'h035dbf12;
    ram_cell[   22201] = 32'h5f18dcba;
    ram_cell[   22202] = 32'hcbb9a229;
    ram_cell[   22203] = 32'hd40f7677;
    ram_cell[   22204] = 32'hec1441af;
    ram_cell[   22205] = 32'h49bdd14a;
    ram_cell[   22206] = 32'h0bf6fad3;
    ram_cell[   22207] = 32'hf88cb2d0;
    ram_cell[   22208] = 32'h3a395674;
    ram_cell[   22209] = 32'hd0b70866;
    ram_cell[   22210] = 32'h7ac7d2d5;
    ram_cell[   22211] = 32'h49b76acf;
    ram_cell[   22212] = 32'h933f5cbf;
    ram_cell[   22213] = 32'h2a97e69a;
    ram_cell[   22214] = 32'haf12bd57;
    ram_cell[   22215] = 32'h09928295;
    ram_cell[   22216] = 32'h94e30497;
    ram_cell[   22217] = 32'hb28b84c3;
    ram_cell[   22218] = 32'h98228c9e;
    ram_cell[   22219] = 32'ha93d5492;
    ram_cell[   22220] = 32'h75808d24;
    ram_cell[   22221] = 32'hdd54cb9a;
    ram_cell[   22222] = 32'h677141cd;
    ram_cell[   22223] = 32'h5cace93f;
    ram_cell[   22224] = 32'hdec0ee92;
    ram_cell[   22225] = 32'hc72e6fde;
    ram_cell[   22226] = 32'hdfcf417d;
    ram_cell[   22227] = 32'h855254bc;
    ram_cell[   22228] = 32'hfc847a0e;
    ram_cell[   22229] = 32'h40115de0;
    ram_cell[   22230] = 32'h55803ca3;
    ram_cell[   22231] = 32'h80d20aa4;
    ram_cell[   22232] = 32'hd2a5611c;
    ram_cell[   22233] = 32'hd2855cf3;
    ram_cell[   22234] = 32'h90118a9e;
    ram_cell[   22235] = 32'h4e8b77ba;
    ram_cell[   22236] = 32'hb421ca05;
    ram_cell[   22237] = 32'hd26b3903;
    ram_cell[   22238] = 32'h3c8f8387;
    ram_cell[   22239] = 32'h8c57c997;
    ram_cell[   22240] = 32'h55e4fb74;
    ram_cell[   22241] = 32'hbee36061;
    ram_cell[   22242] = 32'he5f9c544;
    ram_cell[   22243] = 32'he32e5f6c;
    ram_cell[   22244] = 32'h4052d06b;
    ram_cell[   22245] = 32'h71eab676;
    ram_cell[   22246] = 32'h38cd5fdd;
    ram_cell[   22247] = 32'h2e9f05db;
    ram_cell[   22248] = 32'h1ef2b7a0;
    ram_cell[   22249] = 32'h9ec21ec6;
    ram_cell[   22250] = 32'h890a0c08;
    ram_cell[   22251] = 32'h312432cd;
    ram_cell[   22252] = 32'h25a94feb;
    ram_cell[   22253] = 32'h52923cc6;
    ram_cell[   22254] = 32'haa8bd806;
    ram_cell[   22255] = 32'h123de58f;
    ram_cell[   22256] = 32'h93ceba1f;
    ram_cell[   22257] = 32'h616bdfbc;
    ram_cell[   22258] = 32'hc09bffd1;
    ram_cell[   22259] = 32'hf3711f0e;
    ram_cell[   22260] = 32'h9ce80e59;
    ram_cell[   22261] = 32'h3dd4076d;
    ram_cell[   22262] = 32'h2bffe5cc;
    ram_cell[   22263] = 32'hadc1445b;
    ram_cell[   22264] = 32'hbc4104fd;
    ram_cell[   22265] = 32'hb3351ba7;
    ram_cell[   22266] = 32'h1a28ea83;
    ram_cell[   22267] = 32'h80757984;
    ram_cell[   22268] = 32'h7f80530b;
    ram_cell[   22269] = 32'h77d6021a;
    ram_cell[   22270] = 32'hdf38e045;
    ram_cell[   22271] = 32'h72b8dfcc;
    ram_cell[   22272] = 32'h43386a1c;
    ram_cell[   22273] = 32'h609233e6;
    ram_cell[   22274] = 32'h1206da27;
    ram_cell[   22275] = 32'hd4ec6f26;
    ram_cell[   22276] = 32'h09c93f42;
    ram_cell[   22277] = 32'h15354e20;
    ram_cell[   22278] = 32'h49f75192;
    ram_cell[   22279] = 32'h47b123ce;
    ram_cell[   22280] = 32'h1ef7b205;
    ram_cell[   22281] = 32'h463e8f53;
    ram_cell[   22282] = 32'h27b20c92;
    ram_cell[   22283] = 32'h9589b6fc;
    ram_cell[   22284] = 32'h3cdfc9eb;
    ram_cell[   22285] = 32'hc955b250;
    ram_cell[   22286] = 32'h376c294f;
    ram_cell[   22287] = 32'h78e4ab2c;
    ram_cell[   22288] = 32'h140ede45;
    ram_cell[   22289] = 32'h78560430;
    ram_cell[   22290] = 32'he0da5d79;
    ram_cell[   22291] = 32'h72dbc759;
    ram_cell[   22292] = 32'hd3f00d2c;
    ram_cell[   22293] = 32'h3c1cf99b;
    ram_cell[   22294] = 32'h19851445;
    ram_cell[   22295] = 32'hbb3ba5d6;
    ram_cell[   22296] = 32'h6313666e;
    ram_cell[   22297] = 32'h07edbf9a;
    ram_cell[   22298] = 32'he697a3c5;
    ram_cell[   22299] = 32'h87056b5d;
    ram_cell[   22300] = 32'hd3e73be2;
    ram_cell[   22301] = 32'h33507aa1;
    ram_cell[   22302] = 32'h6e80ef1c;
    ram_cell[   22303] = 32'h2f2d4494;
    ram_cell[   22304] = 32'he0d0c4c7;
    ram_cell[   22305] = 32'h64499e07;
    ram_cell[   22306] = 32'h447aa10d;
    ram_cell[   22307] = 32'h07edda75;
    ram_cell[   22308] = 32'h1b117d01;
    ram_cell[   22309] = 32'hecc8891c;
    ram_cell[   22310] = 32'h7ccfaf4c;
    ram_cell[   22311] = 32'hf8f99afd;
    ram_cell[   22312] = 32'h277eaab0;
    ram_cell[   22313] = 32'h5d40e978;
    ram_cell[   22314] = 32'hfa115cc6;
    ram_cell[   22315] = 32'h94a24d05;
    ram_cell[   22316] = 32'h9dfab981;
    ram_cell[   22317] = 32'hbd43a954;
    ram_cell[   22318] = 32'hae981eed;
    ram_cell[   22319] = 32'h9070b193;
    ram_cell[   22320] = 32'h75bfe54c;
    ram_cell[   22321] = 32'h8c700050;
    ram_cell[   22322] = 32'ha8784021;
    ram_cell[   22323] = 32'hf77a3d32;
    ram_cell[   22324] = 32'h4611bf01;
    ram_cell[   22325] = 32'h38299f4b;
    ram_cell[   22326] = 32'hb0c23bd1;
    ram_cell[   22327] = 32'hc4e7e813;
    ram_cell[   22328] = 32'h2b5ba1a1;
    ram_cell[   22329] = 32'h5376df98;
    ram_cell[   22330] = 32'haf3fa6de;
    ram_cell[   22331] = 32'h6b7b1840;
    ram_cell[   22332] = 32'h5e1a88ed;
    ram_cell[   22333] = 32'h96723a3e;
    ram_cell[   22334] = 32'hbd6a87b6;
    ram_cell[   22335] = 32'h4ce050a2;
    ram_cell[   22336] = 32'h3bd42a75;
    ram_cell[   22337] = 32'h54b615d5;
    ram_cell[   22338] = 32'h28975c87;
    ram_cell[   22339] = 32'hb0430399;
    ram_cell[   22340] = 32'hb10f0052;
    ram_cell[   22341] = 32'hb0f49089;
    ram_cell[   22342] = 32'h39ac0d01;
    ram_cell[   22343] = 32'h81e75703;
    ram_cell[   22344] = 32'h38dea85d;
    ram_cell[   22345] = 32'hda6db326;
    ram_cell[   22346] = 32'h67761046;
    ram_cell[   22347] = 32'h3595af52;
    ram_cell[   22348] = 32'h8f96a342;
    ram_cell[   22349] = 32'h305740ac;
    ram_cell[   22350] = 32'haa5a169d;
    ram_cell[   22351] = 32'hb4d3dea8;
    ram_cell[   22352] = 32'h64c1dd79;
    ram_cell[   22353] = 32'h992cb5f2;
    ram_cell[   22354] = 32'hafcdd1d0;
    ram_cell[   22355] = 32'hc6568fa8;
    ram_cell[   22356] = 32'hc6f3a8da;
    ram_cell[   22357] = 32'he17dc11b;
    ram_cell[   22358] = 32'h14057836;
    ram_cell[   22359] = 32'h777a7277;
    ram_cell[   22360] = 32'h6a75e5ef;
    ram_cell[   22361] = 32'ha8dde984;
    ram_cell[   22362] = 32'h9862530c;
    ram_cell[   22363] = 32'h505ae439;
    ram_cell[   22364] = 32'hbd248a1a;
    ram_cell[   22365] = 32'h6ca12300;
    ram_cell[   22366] = 32'h363e8b4f;
    ram_cell[   22367] = 32'h45bcf000;
    ram_cell[   22368] = 32'hab1cbf88;
    ram_cell[   22369] = 32'h85847add;
    ram_cell[   22370] = 32'h0e785cef;
    ram_cell[   22371] = 32'h748adbd2;
    ram_cell[   22372] = 32'h4f83b3e1;
    ram_cell[   22373] = 32'h05bcfc12;
    ram_cell[   22374] = 32'hfe31db2a;
    ram_cell[   22375] = 32'h774e7c53;
    ram_cell[   22376] = 32'h9c071c69;
    ram_cell[   22377] = 32'ha678ca73;
    ram_cell[   22378] = 32'ha747c52a;
    ram_cell[   22379] = 32'h49db0518;
    ram_cell[   22380] = 32'hfbd164f7;
    ram_cell[   22381] = 32'h27fea5c2;
    ram_cell[   22382] = 32'h2ab0cabd;
    ram_cell[   22383] = 32'h7712b1ab;
    ram_cell[   22384] = 32'hb0135e86;
    ram_cell[   22385] = 32'h4e0f8809;
    ram_cell[   22386] = 32'h06e08c4c;
    ram_cell[   22387] = 32'h15094b2d;
    ram_cell[   22388] = 32'h5e5ffe51;
    ram_cell[   22389] = 32'ha2ff1650;
    ram_cell[   22390] = 32'h238e0c24;
    ram_cell[   22391] = 32'h114ee9ac;
    ram_cell[   22392] = 32'h8455d7dd;
    ram_cell[   22393] = 32'hf8bb0d34;
    ram_cell[   22394] = 32'h3c30fca2;
    ram_cell[   22395] = 32'hf31c9534;
    ram_cell[   22396] = 32'h835a4788;
    ram_cell[   22397] = 32'hbf5f093a;
    ram_cell[   22398] = 32'h559ba400;
    ram_cell[   22399] = 32'h2ae26686;
    ram_cell[   22400] = 32'hfd6a79d0;
    ram_cell[   22401] = 32'h4ad1382a;
    ram_cell[   22402] = 32'h37c6c88c;
    ram_cell[   22403] = 32'ha847cba1;
    ram_cell[   22404] = 32'hf421f94d;
    ram_cell[   22405] = 32'h64f702b8;
    ram_cell[   22406] = 32'hedf3377d;
    ram_cell[   22407] = 32'h4c328d33;
    ram_cell[   22408] = 32'h837f67c2;
    ram_cell[   22409] = 32'h4e5d94cc;
    ram_cell[   22410] = 32'h51ab4272;
    ram_cell[   22411] = 32'h56a9f753;
    ram_cell[   22412] = 32'h033a8d83;
    ram_cell[   22413] = 32'hc0a4bc8d;
    ram_cell[   22414] = 32'h49cd8010;
    ram_cell[   22415] = 32'hc7111400;
    ram_cell[   22416] = 32'h4b6f840d;
    ram_cell[   22417] = 32'h87dd2d6d;
    ram_cell[   22418] = 32'h771e9239;
    ram_cell[   22419] = 32'h27ab1780;
    ram_cell[   22420] = 32'hc956623a;
    ram_cell[   22421] = 32'h3f10c8ad;
    ram_cell[   22422] = 32'hda0c7386;
    ram_cell[   22423] = 32'ha15773d4;
    ram_cell[   22424] = 32'h1fede7ca;
    ram_cell[   22425] = 32'h558c0a9a;
    ram_cell[   22426] = 32'h6f81ba4f;
    ram_cell[   22427] = 32'h1f4af481;
    ram_cell[   22428] = 32'h9c1b9f36;
    ram_cell[   22429] = 32'he7db029b;
    ram_cell[   22430] = 32'hbe7564fd;
    ram_cell[   22431] = 32'h1c62666f;
    ram_cell[   22432] = 32'h4838fe00;
    ram_cell[   22433] = 32'hbe4b0899;
    ram_cell[   22434] = 32'hf6f44481;
    ram_cell[   22435] = 32'hba412621;
    ram_cell[   22436] = 32'hbebe16b7;
    ram_cell[   22437] = 32'h0ae6535d;
    ram_cell[   22438] = 32'hb9e65b34;
    ram_cell[   22439] = 32'h6686097a;
    ram_cell[   22440] = 32'hee962a78;
    ram_cell[   22441] = 32'heac62d62;
    ram_cell[   22442] = 32'h31ef5a75;
    ram_cell[   22443] = 32'h30598f33;
    ram_cell[   22444] = 32'hdbaafa2a;
    ram_cell[   22445] = 32'h616aa1ea;
    ram_cell[   22446] = 32'h80852535;
    ram_cell[   22447] = 32'h4701c4e1;
    ram_cell[   22448] = 32'h4d3208c7;
    ram_cell[   22449] = 32'h1b1ae9f6;
    ram_cell[   22450] = 32'hb934b51a;
    ram_cell[   22451] = 32'hc44ac609;
    ram_cell[   22452] = 32'h7d4824c8;
    ram_cell[   22453] = 32'h8342e9bc;
    ram_cell[   22454] = 32'he224a8a2;
    ram_cell[   22455] = 32'h99c847fc;
    ram_cell[   22456] = 32'hf03278ea;
    ram_cell[   22457] = 32'h01f19b26;
    ram_cell[   22458] = 32'h90338c43;
    ram_cell[   22459] = 32'h3edfe26a;
    ram_cell[   22460] = 32'h8e9135bf;
    ram_cell[   22461] = 32'h6f628bfe;
    ram_cell[   22462] = 32'hfe0d3fb8;
    ram_cell[   22463] = 32'h10f86a22;
    ram_cell[   22464] = 32'h2d943565;
    ram_cell[   22465] = 32'h41a08656;
    ram_cell[   22466] = 32'h96d9eacd;
    ram_cell[   22467] = 32'h8acdce77;
    ram_cell[   22468] = 32'h99bed7d0;
    ram_cell[   22469] = 32'h344c2bc6;
    ram_cell[   22470] = 32'h958d4630;
    ram_cell[   22471] = 32'hda49e141;
    ram_cell[   22472] = 32'had1e19b3;
    ram_cell[   22473] = 32'h14ff83ab;
    ram_cell[   22474] = 32'ha9ba1dc3;
    ram_cell[   22475] = 32'h17884504;
    ram_cell[   22476] = 32'h58c35214;
    ram_cell[   22477] = 32'ha32822e2;
    ram_cell[   22478] = 32'he1eb3762;
    ram_cell[   22479] = 32'heb177fb7;
    ram_cell[   22480] = 32'h1e247776;
    ram_cell[   22481] = 32'h8759cd38;
    ram_cell[   22482] = 32'h7dd72530;
    ram_cell[   22483] = 32'hcc32f455;
    ram_cell[   22484] = 32'h7cc8f282;
    ram_cell[   22485] = 32'hcdf17f8f;
    ram_cell[   22486] = 32'he01d9867;
    ram_cell[   22487] = 32'h03351072;
    ram_cell[   22488] = 32'h2e98dc81;
    ram_cell[   22489] = 32'h6c913a5e;
    ram_cell[   22490] = 32'h314ea400;
    ram_cell[   22491] = 32'hef226627;
    ram_cell[   22492] = 32'ha94b5146;
    ram_cell[   22493] = 32'hd86eadb7;
    ram_cell[   22494] = 32'hccf0f7ed;
    ram_cell[   22495] = 32'ha6500c57;
    ram_cell[   22496] = 32'h307b9358;
    ram_cell[   22497] = 32'h314984c9;
    ram_cell[   22498] = 32'hadc593f8;
    ram_cell[   22499] = 32'h0c9ecd64;
    ram_cell[   22500] = 32'h5f9f65b0;
    ram_cell[   22501] = 32'h5e0e6a34;
    ram_cell[   22502] = 32'hdda87b73;
    ram_cell[   22503] = 32'h1a103401;
    ram_cell[   22504] = 32'hb97a9cd4;
    ram_cell[   22505] = 32'hc089e7a9;
    ram_cell[   22506] = 32'h3615bba2;
    ram_cell[   22507] = 32'he067d3ae;
    ram_cell[   22508] = 32'h3ca0d4fe;
    ram_cell[   22509] = 32'hfa0ead53;
    ram_cell[   22510] = 32'h73181c4f;
    ram_cell[   22511] = 32'h7de14cd9;
    ram_cell[   22512] = 32'ha8c1fead;
    ram_cell[   22513] = 32'h440acb59;
    ram_cell[   22514] = 32'h7618b9df;
    ram_cell[   22515] = 32'h6fc3c724;
    ram_cell[   22516] = 32'h6f04b1ca;
    ram_cell[   22517] = 32'hf1b1e734;
    ram_cell[   22518] = 32'ha5d7e076;
    ram_cell[   22519] = 32'h8c12679e;
    ram_cell[   22520] = 32'hc8ab72f9;
    ram_cell[   22521] = 32'hd9ba3595;
    ram_cell[   22522] = 32'hf899f830;
    ram_cell[   22523] = 32'hcf729a10;
    ram_cell[   22524] = 32'h306d301c;
    ram_cell[   22525] = 32'hf9cc4398;
    ram_cell[   22526] = 32'h66029a74;
    ram_cell[   22527] = 32'h2757c6f6;
    ram_cell[   22528] = 32'h4753cec1;
    ram_cell[   22529] = 32'hcbd572f4;
    ram_cell[   22530] = 32'h342331c3;
    ram_cell[   22531] = 32'h66906adf;
    ram_cell[   22532] = 32'h62f959dc;
    ram_cell[   22533] = 32'h7c8cc957;
    ram_cell[   22534] = 32'h55bc63e8;
    ram_cell[   22535] = 32'h3d6db447;
    ram_cell[   22536] = 32'h04caea84;
    ram_cell[   22537] = 32'haa1b6142;
    ram_cell[   22538] = 32'hc633ca1b;
    ram_cell[   22539] = 32'h10c6a936;
    ram_cell[   22540] = 32'h727f096b;
    ram_cell[   22541] = 32'h40553f5c;
    ram_cell[   22542] = 32'hc38aceef;
    ram_cell[   22543] = 32'hcdf1a960;
    ram_cell[   22544] = 32'h6e97aedf;
    ram_cell[   22545] = 32'hf8886fb1;
    ram_cell[   22546] = 32'h1396476f;
    ram_cell[   22547] = 32'h630321ef;
    ram_cell[   22548] = 32'ha6824cc8;
    ram_cell[   22549] = 32'hc0185c03;
    ram_cell[   22550] = 32'hc1a8f8eb;
    ram_cell[   22551] = 32'hbb936ece;
    ram_cell[   22552] = 32'h2026d9ae;
    ram_cell[   22553] = 32'h558e05e0;
    ram_cell[   22554] = 32'he7629ab7;
    ram_cell[   22555] = 32'hec6f4049;
    ram_cell[   22556] = 32'h748c7811;
    ram_cell[   22557] = 32'h307ec623;
    ram_cell[   22558] = 32'hf3731e0a;
    ram_cell[   22559] = 32'h22a02d25;
    ram_cell[   22560] = 32'h5801a2e5;
    ram_cell[   22561] = 32'h49b7295b;
    ram_cell[   22562] = 32'hee026365;
    ram_cell[   22563] = 32'hdb5e4a4c;
    ram_cell[   22564] = 32'h11e7c060;
    ram_cell[   22565] = 32'ha5346d4e;
    ram_cell[   22566] = 32'he708b1aa;
    ram_cell[   22567] = 32'h9f50879f;
    ram_cell[   22568] = 32'h43a64c4e;
    ram_cell[   22569] = 32'hf8ac5a1c;
    ram_cell[   22570] = 32'h21fd7928;
    ram_cell[   22571] = 32'h7c4303f5;
    ram_cell[   22572] = 32'h3b022e0e;
    ram_cell[   22573] = 32'hc82e3c18;
    ram_cell[   22574] = 32'h8abc9882;
    ram_cell[   22575] = 32'h33720079;
    ram_cell[   22576] = 32'h16ceebae;
    ram_cell[   22577] = 32'h2bb0ca66;
    ram_cell[   22578] = 32'h724f7d48;
    ram_cell[   22579] = 32'hb267031c;
    ram_cell[   22580] = 32'h59929cda;
    ram_cell[   22581] = 32'hfbf820fd;
    ram_cell[   22582] = 32'h5ebc0afd;
    ram_cell[   22583] = 32'h3b03bb61;
    ram_cell[   22584] = 32'h65124845;
    ram_cell[   22585] = 32'h8f52a5cb;
    ram_cell[   22586] = 32'hf2838834;
    ram_cell[   22587] = 32'h443456e3;
    ram_cell[   22588] = 32'h2dfbf9f2;
    ram_cell[   22589] = 32'h2f0a5c0b;
    ram_cell[   22590] = 32'h1e217e66;
    ram_cell[   22591] = 32'h41acee3a;
    ram_cell[   22592] = 32'hc2b362f5;
    ram_cell[   22593] = 32'h8d9cdb6d;
    ram_cell[   22594] = 32'h1a4675bc;
    ram_cell[   22595] = 32'h7b8268bc;
    ram_cell[   22596] = 32'hb76be3eb;
    ram_cell[   22597] = 32'h500f4f8d;
    ram_cell[   22598] = 32'hca25b358;
    ram_cell[   22599] = 32'hdca4c0be;
    ram_cell[   22600] = 32'hd5544c88;
    ram_cell[   22601] = 32'h77e67339;
    ram_cell[   22602] = 32'ha9bdea1b;
    ram_cell[   22603] = 32'h84fafd50;
    ram_cell[   22604] = 32'h450e8d9f;
    ram_cell[   22605] = 32'hc3eed472;
    ram_cell[   22606] = 32'hac64b8b7;
    ram_cell[   22607] = 32'h9c288849;
    ram_cell[   22608] = 32'hc27e9138;
    ram_cell[   22609] = 32'h853fdb1e;
    ram_cell[   22610] = 32'h68bce69b;
    ram_cell[   22611] = 32'h555b3f93;
    ram_cell[   22612] = 32'h110729b1;
    ram_cell[   22613] = 32'hf4acb082;
    ram_cell[   22614] = 32'hf352d72e;
    ram_cell[   22615] = 32'h10ecb815;
    ram_cell[   22616] = 32'h4c079212;
    ram_cell[   22617] = 32'he6486f0b;
    ram_cell[   22618] = 32'hbf51f14f;
    ram_cell[   22619] = 32'h454084d7;
    ram_cell[   22620] = 32'h84b4105a;
    ram_cell[   22621] = 32'hcac835fb;
    ram_cell[   22622] = 32'hc454ef94;
    ram_cell[   22623] = 32'h8c2c9c93;
    ram_cell[   22624] = 32'he6c5d87c;
    ram_cell[   22625] = 32'ha75cb584;
    ram_cell[   22626] = 32'h4290d46b;
    ram_cell[   22627] = 32'h3cbf2a7d;
    ram_cell[   22628] = 32'he50bf529;
    ram_cell[   22629] = 32'hfd1c1fa4;
    ram_cell[   22630] = 32'he9ca95ac;
    ram_cell[   22631] = 32'hafc5e8b0;
    ram_cell[   22632] = 32'h848369aa;
    ram_cell[   22633] = 32'he4285b1d;
    ram_cell[   22634] = 32'h2e501bf9;
    ram_cell[   22635] = 32'h19a0d323;
    ram_cell[   22636] = 32'hb5e848ce;
    ram_cell[   22637] = 32'hf6bb9409;
    ram_cell[   22638] = 32'h7347699c;
    ram_cell[   22639] = 32'h6d647def;
    ram_cell[   22640] = 32'h91db5e79;
    ram_cell[   22641] = 32'h3666e1d6;
    ram_cell[   22642] = 32'h370d9150;
    ram_cell[   22643] = 32'h7e3d7618;
    ram_cell[   22644] = 32'hbdf1354f;
    ram_cell[   22645] = 32'h72b25ef7;
    ram_cell[   22646] = 32'h48f3138e;
    ram_cell[   22647] = 32'h3819f31d;
    ram_cell[   22648] = 32'hfe0d7c6c;
    ram_cell[   22649] = 32'h2942b947;
    ram_cell[   22650] = 32'h31bc35b6;
    ram_cell[   22651] = 32'h435fafe4;
    ram_cell[   22652] = 32'h09f2b492;
    ram_cell[   22653] = 32'h9d691b84;
    ram_cell[   22654] = 32'h73dd4a73;
    ram_cell[   22655] = 32'h7403ca9b;
    ram_cell[   22656] = 32'h389d97d3;
    ram_cell[   22657] = 32'hd79cfdfb;
    ram_cell[   22658] = 32'h5e36bcfd;
    ram_cell[   22659] = 32'h3377b690;
    ram_cell[   22660] = 32'h4b7f5c35;
    ram_cell[   22661] = 32'hc046f80d;
    ram_cell[   22662] = 32'h24fef2d4;
    ram_cell[   22663] = 32'ha5f0b096;
    ram_cell[   22664] = 32'h3556b0f4;
    ram_cell[   22665] = 32'h08ed17a2;
    ram_cell[   22666] = 32'h1847426f;
    ram_cell[   22667] = 32'ha0140d85;
    ram_cell[   22668] = 32'h62ed8de9;
    ram_cell[   22669] = 32'h4e6278d7;
    ram_cell[   22670] = 32'h24f9f9a4;
    ram_cell[   22671] = 32'h01dd20a0;
    ram_cell[   22672] = 32'hdb04b0df;
    ram_cell[   22673] = 32'h15c9dd34;
    ram_cell[   22674] = 32'h4aa670cc;
    ram_cell[   22675] = 32'h28df5de4;
    ram_cell[   22676] = 32'h7ef457e9;
    ram_cell[   22677] = 32'h8c521f5a;
    ram_cell[   22678] = 32'hbd5cd896;
    ram_cell[   22679] = 32'h79d2db37;
    ram_cell[   22680] = 32'h8c756cf4;
    ram_cell[   22681] = 32'hab62a179;
    ram_cell[   22682] = 32'h377275ea;
    ram_cell[   22683] = 32'h4fa95b25;
    ram_cell[   22684] = 32'h39341333;
    ram_cell[   22685] = 32'h3837f209;
    ram_cell[   22686] = 32'h31dc6842;
    ram_cell[   22687] = 32'he071c1d4;
    ram_cell[   22688] = 32'h2760ae2b;
    ram_cell[   22689] = 32'hb0600ce3;
    ram_cell[   22690] = 32'h3b78432f;
    ram_cell[   22691] = 32'hb3c01194;
    ram_cell[   22692] = 32'h894b752d;
    ram_cell[   22693] = 32'h158a2fbd;
    ram_cell[   22694] = 32'h4e2e2963;
    ram_cell[   22695] = 32'h92400811;
    ram_cell[   22696] = 32'h3ce41563;
    ram_cell[   22697] = 32'hd46f2aff;
    ram_cell[   22698] = 32'h2e9a8833;
    ram_cell[   22699] = 32'hbbda62b4;
    ram_cell[   22700] = 32'h4d4667cd;
    ram_cell[   22701] = 32'h153387c0;
    ram_cell[   22702] = 32'h2c81cf29;
    ram_cell[   22703] = 32'h62e9cd73;
    ram_cell[   22704] = 32'h9a919e97;
    ram_cell[   22705] = 32'h5782a582;
    ram_cell[   22706] = 32'h63f7625f;
    ram_cell[   22707] = 32'hc54cbc68;
    ram_cell[   22708] = 32'h737f1a62;
    ram_cell[   22709] = 32'hc6388f9a;
    ram_cell[   22710] = 32'h8654edb5;
    ram_cell[   22711] = 32'hcda6b5a9;
    ram_cell[   22712] = 32'h0c18f05f;
    ram_cell[   22713] = 32'hade1727a;
    ram_cell[   22714] = 32'h760343c0;
    ram_cell[   22715] = 32'h8c8a713b;
    ram_cell[   22716] = 32'hbdac8c71;
    ram_cell[   22717] = 32'hedaa7555;
    ram_cell[   22718] = 32'he81d8741;
    ram_cell[   22719] = 32'hf91e78e4;
    ram_cell[   22720] = 32'h311fdfb8;
    ram_cell[   22721] = 32'h939eb433;
    ram_cell[   22722] = 32'h791a1936;
    ram_cell[   22723] = 32'hfdda4267;
    ram_cell[   22724] = 32'hacf95b08;
    ram_cell[   22725] = 32'h94e8d8ba;
    ram_cell[   22726] = 32'h3da64135;
    ram_cell[   22727] = 32'hc79128a1;
    ram_cell[   22728] = 32'h257a1013;
    ram_cell[   22729] = 32'hab75eaf5;
    ram_cell[   22730] = 32'h29d08d73;
    ram_cell[   22731] = 32'hcb34dced;
    ram_cell[   22732] = 32'h2d860443;
    ram_cell[   22733] = 32'hd3a3779b;
    ram_cell[   22734] = 32'h7aba9f71;
    ram_cell[   22735] = 32'h69a3b2e2;
    ram_cell[   22736] = 32'hde7a985c;
    ram_cell[   22737] = 32'had9b58b0;
    ram_cell[   22738] = 32'hf817c3cd;
    ram_cell[   22739] = 32'hfffc6f8b;
    ram_cell[   22740] = 32'he122224d;
    ram_cell[   22741] = 32'h6206a5db;
    ram_cell[   22742] = 32'h1703d658;
    ram_cell[   22743] = 32'h9621f02d;
    ram_cell[   22744] = 32'hb993eac9;
    ram_cell[   22745] = 32'h6da8fbd7;
    ram_cell[   22746] = 32'hde41bbf0;
    ram_cell[   22747] = 32'h5eaf9cea;
    ram_cell[   22748] = 32'h6086f8d4;
    ram_cell[   22749] = 32'hc8f350e0;
    ram_cell[   22750] = 32'h406f99b5;
    ram_cell[   22751] = 32'h1e5c9735;
    ram_cell[   22752] = 32'h5c50bc98;
    ram_cell[   22753] = 32'h3b93d63c;
    ram_cell[   22754] = 32'heb6acf01;
    ram_cell[   22755] = 32'h3293c685;
    ram_cell[   22756] = 32'ha9ffc44b;
    ram_cell[   22757] = 32'h1b172624;
    ram_cell[   22758] = 32'hc40f4df4;
    ram_cell[   22759] = 32'hb400b617;
    ram_cell[   22760] = 32'he0e1a3e0;
    ram_cell[   22761] = 32'h77e6c484;
    ram_cell[   22762] = 32'h746117d1;
    ram_cell[   22763] = 32'h638955f9;
    ram_cell[   22764] = 32'h75ffc5d6;
    ram_cell[   22765] = 32'h2e509ae9;
    ram_cell[   22766] = 32'h89284685;
    ram_cell[   22767] = 32'hd5779875;
    ram_cell[   22768] = 32'h8d84780b;
    ram_cell[   22769] = 32'h7f97d034;
    ram_cell[   22770] = 32'h8ff6f6e5;
    ram_cell[   22771] = 32'h4014bf66;
    ram_cell[   22772] = 32'h5319fb9f;
    ram_cell[   22773] = 32'hdad31c3a;
    ram_cell[   22774] = 32'hfcc29f8f;
    ram_cell[   22775] = 32'h254524da;
    ram_cell[   22776] = 32'hd9c75123;
    ram_cell[   22777] = 32'hc852b288;
    ram_cell[   22778] = 32'h860adb26;
    ram_cell[   22779] = 32'h3a7db91e;
    ram_cell[   22780] = 32'h8d231a9b;
    ram_cell[   22781] = 32'hed82b6b1;
    ram_cell[   22782] = 32'h8780fe4a;
    ram_cell[   22783] = 32'hee48d55c;
    ram_cell[   22784] = 32'h1a28b44f;
    ram_cell[   22785] = 32'h81f63735;
    ram_cell[   22786] = 32'h207f892e;
    ram_cell[   22787] = 32'hdd6a6ec2;
    ram_cell[   22788] = 32'hb0a85aef;
    ram_cell[   22789] = 32'h8532d938;
    ram_cell[   22790] = 32'he85f171e;
    ram_cell[   22791] = 32'h1303f7f7;
    ram_cell[   22792] = 32'h3ca84699;
    ram_cell[   22793] = 32'hfecbe70c;
    ram_cell[   22794] = 32'h954c0561;
    ram_cell[   22795] = 32'hf1aad91a;
    ram_cell[   22796] = 32'h1e98c2ce;
    ram_cell[   22797] = 32'h0e7a3abc;
    ram_cell[   22798] = 32'h6e25ad18;
    ram_cell[   22799] = 32'h3ac49795;
    ram_cell[   22800] = 32'h300f263f;
    ram_cell[   22801] = 32'he0cb67f3;
    ram_cell[   22802] = 32'hb3a1b04b;
    ram_cell[   22803] = 32'h392ab14d;
    ram_cell[   22804] = 32'h9fa3d9a5;
    ram_cell[   22805] = 32'hc23b90bc;
    ram_cell[   22806] = 32'h61d5cedf;
    ram_cell[   22807] = 32'h609b13ef;
    ram_cell[   22808] = 32'h59911534;
    ram_cell[   22809] = 32'hbde7e044;
    ram_cell[   22810] = 32'h8cdf4b7c;
    ram_cell[   22811] = 32'h90ddc9c3;
    ram_cell[   22812] = 32'h4808cc4c;
    ram_cell[   22813] = 32'h7af7d030;
    ram_cell[   22814] = 32'hd4ec7f2b;
    ram_cell[   22815] = 32'h8268a724;
    ram_cell[   22816] = 32'h8d7ec980;
    ram_cell[   22817] = 32'hc84264e0;
    ram_cell[   22818] = 32'hf86d6bbc;
    ram_cell[   22819] = 32'hfb5efe8a;
    ram_cell[   22820] = 32'h40a2e4cc;
    ram_cell[   22821] = 32'h81f6c6ed;
    ram_cell[   22822] = 32'hbcb42f25;
    ram_cell[   22823] = 32'h3db657ed;
    ram_cell[   22824] = 32'he1599921;
    ram_cell[   22825] = 32'hb8adc137;
    ram_cell[   22826] = 32'h7819b299;
    ram_cell[   22827] = 32'h3bd31008;
    ram_cell[   22828] = 32'hf225be85;
    ram_cell[   22829] = 32'h9db7f82e;
    ram_cell[   22830] = 32'h5f0332e0;
    ram_cell[   22831] = 32'h38a545dd;
    ram_cell[   22832] = 32'hb2247ac4;
    ram_cell[   22833] = 32'hc3d8e0ff;
    ram_cell[   22834] = 32'h44a9405a;
    ram_cell[   22835] = 32'h8aa0d856;
    ram_cell[   22836] = 32'h6a3a1a12;
    ram_cell[   22837] = 32'h643c6795;
    ram_cell[   22838] = 32'h4a52f152;
    ram_cell[   22839] = 32'h5331cfee;
    ram_cell[   22840] = 32'h00bfa915;
    ram_cell[   22841] = 32'h3828465d;
    ram_cell[   22842] = 32'h5d1113a8;
    ram_cell[   22843] = 32'hbcef8097;
    ram_cell[   22844] = 32'h866c1c46;
    ram_cell[   22845] = 32'h9e02d5a0;
    ram_cell[   22846] = 32'hf720c96b;
    ram_cell[   22847] = 32'h694459f6;
    ram_cell[   22848] = 32'ha34fb378;
    ram_cell[   22849] = 32'he1f35b27;
    ram_cell[   22850] = 32'had4ab221;
    ram_cell[   22851] = 32'h1282719d;
    ram_cell[   22852] = 32'h83f61730;
    ram_cell[   22853] = 32'he9b3a673;
    ram_cell[   22854] = 32'h7e5bfca4;
    ram_cell[   22855] = 32'h597fe511;
    ram_cell[   22856] = 32'he4f997ed;
    ram_cell[   22857] = 32'h2b9f11ec;
    ram_cell[   22858] = 32'h390df0d5;
    ram_cell[   22859] = 32'h14b8af6d;
    ram_cell[   22860] = 32'h761f80d5;
    ram_cell[   22861] = 32'ha11bbf15;
    ram_cell[   22862] = 32'hc6b1efab;
    ram_cell[   22863] = 32'h059aecee;
    ram_cell[   22864] = 32'hbe6f11b3;
    ram_cell[   22865] = 32'h04c8c383;
    ram_cell[   22866] = 32'h29c1003f;
    ram_cell[   22867] = 32'h0a50e5dd;
    ram_cell[   22868] = 32'h7b517df9;
    ram_cell[   22869] = 32'h74de5c0c;
    ram_cell[   22870] = 32'h267734cf;
    ram_cell[   22871] = 32'hb41e6e16;
    ram_cell[   22872] = 32'h2ea45682;
    ram_cell[   22873] = 32'h4f9232cb;
    ram_cell[   22874] = 32'hf8667c9a;
    ram_cell[   22875] = 32'hb25cc9f3;
    ram_cell[   22876] = 32'h4e991f62;
    ram_cell[   22877] = 32'ha9f6c9b4;
    ram_cell[   22878] = 32'hdd0fa6cc;
    ram_cell[   22879] = 32'hc357e166;
    ram_cell[   22880] = 32'h7a9fd035;
    ram_cell[   22881] = 32'h8b82bca1;
    ram_cell[   22882] = 32'h0912adfb;
    ram_cell[   22883] = 32'h321701ac;
    ram_cell[   22884] = 32'h9a5bd8af;
    ram_cell[   22885] = 32'h6a9919af;
    ram_cell[   22886] = 32'h98b4b14a;
    ram_cell[   22887] = 32'h89798383;
    ram_cell[   22888] = 32'h1a0d0d4a;
    ram_cell[   22889] = 32'h0ce2d04c;
    ram_cell[   22890] = 32'h24416506;
    ram_cell[   22891] = 32'h18877fc5;
    ram_cell[   22892] = 32'hf0437fbb;
    ram_cell[   22893] = 32'hc9dd572a;
    ram_cell[   22894] = 32'heef507be;
    ram_cell[   22895] = 32'h92e58862;
    ram_cell[   22896] = 32'hcc3b97d8;
    ram_cell[   22897] = 32'h2b92c9a2;
    ram_cell[   22898] = 32'hdbb15223;
    ram_cell[   22899] = 32'hf8ed88af;
    ram_cell[   22900] = 32'h8197ca4c;
    ram_cell[   22901] = 32'hde1a03db;
    ram_cell[   22902] = 32'h160a5904;
    ram_cell[   22903] = 32'h76bea4d4;
    ram_cell[   22904] = 32'h3eb237f7;
    ram_cell[   22905] = 32'hb7640446;
    ram_cell[   22906] = 32'h7a1d19b3;
    ram_cell[   22907] = 32'h760fc2fc;
    ram_cell[   22908] = 32'he3780726;
    ram_cell[   22909] = 32'h12578c0f;
    ram_cell[   22910] = 32'h271e651e;
    ram_cell[   22911] = 32'hddf72407;
    ram_cell[   22912] = 32'he4679cc5;
    ram_cell[   22913] = 32'h9b8a8b6a;
    ram_cell[   22914] = 32'hde832213;
    ram_cell[   22915] = 32'hfc252358;
    ram_cell[   22916] = 32'h76ed15d0;
    ram_cell[   22917] = 32'h8ea43827;
    ram_cell[   22918] = 32'h721290b3;
    ram_cell[   22919] = 32'hbfac9041;
    ram_cell[   22920] = 32'hd6836718;
    ram_cell[   22921] = 32'h87661e05;
    ram_cell[   22922] = 32'h60234c1a;
    ram_cell[   22923] = 32'h9768dd34;
    ram_cell[   22924] = 32'h13de1fbe;
    ram_cell[   22925] = 32'hf6cd78c4;
    ram_cell[   22926] = 32'h3397ccc4;
    ram_cell[   22927] = 32'hcd22537f;
    ram_cell[   22928] = 32'hb4ed189c;
    ram_cell[   22929] = 32'h1702791b;
    ram_cell[   22930] = 32'h93c23675;
    ram_cell[   22931] = 32'h711a6852;
    ram_cell[   22932] = 32'h60740588;
    ram_cell[   22933] = 32'h5068845e;
    ram_cell[   22934] = 32'h18ec74d0;
    ram_cell[   22935] = 32'hff08dea2;
    ram_cell[   22936] = 32'h4daaabba;
    ram_cell[   22937] = 32'h5f2ecd23;
    ram_cell[   22938] = 32'he00d4a9a;
    ram_cell[   22939] = 32'h32e8edc9;
    ram_cell[   22940] = 32'h8f6fa85a;
    ram_cell[   22941] = 32'h3c9e405a;
    ram_cell[   22942] = 32'h7a964c39;
    ram_cell[   22943] = 32'h6524f1cd;
    ram_cell[   22944] = 32'hdea5d97d;
    ram_cell[   22945] = 32'ha9a526cf;
    ram_cell[   22946] = 32'h5bd90aec;
    ram_cell[   22947] = 32'h0197c181;
    ram_cell[   22948] = 32'h2f1f9c3c;
    ram_cell[   22949] = 32'h09581875;
    ram_cell[   22950] = 32'hcc5f007a;
    ram_cell[   22951] = 32'h42a91195;
    ram_cell[   22952] = 32'hd2b59c64;
    ram_cell[   22953] = 32'h4eba6711;
    ram_cell[   22954] = 32'hb0469837;
    ram_cell[   22955] = 32'h9568b15e;
    ram_cell[   22956] = 32'h07f71038;
    ram_cell[   22957] = 32'h06ec8f96;
    ram_cell[   22958] = 32'h08a81feb;
    ram_cell[   22959] = 32'he47087ae;
    ram_cell[   22960] = 32'hbd3187f9;
    ram_cell[   22961] = 32'he8d6887b;
    ram_cell[   22962] = 32'hc45cdf1e;
    ram_cell[   22963] = 32'h7a28cbf9;
    ram_cell[   22964] = 32'hae552000;
    ram_cell[   22965] = 32'hd6f41de7;
    ram_cell[   22966] = 32'h1c734168;
    ram_cell[   22967] = 32'h4f5329fd;
    ram_cell[   22968] = 32'h1b47db1e;
    ram_cell[   22969] = 32'h9f6b035d;
    ram_cell[   22970] = 32'h557e5280;
    ram_cell[   22971] = 32'hbd58eaf4;
    ram_cell[   22972] = 32'h37054ab3;
    ram_cell[   22973] = 32'h76070a74;
    ram_cell[   22974] = 32'h809aea6d;
    ram_cell[   22975] = 32'h3cb2c3c2;
    ram_cell[   22976] = 32'hc32e0f31;
    ram_cell[   22977] = 32'hdea32ae9;
    ram_cell[   22978] = 32'h26f612a6;
    ram_cell[   22979] = 32'hb9f538cc;
    ram_cell[   22980] = 32'hc02a152e;
    ram_cell[   22981] = 32'hdf77cf6e;
    ram_cell[   22982] = 32'h7cfaca58;
    ram_cell[   22983] = 32'h36ba49ec;
    ram_cell[   22984] = 32'haf84df54;
    ram_cell[   22985] = 32'hf5ce17f2;
    ram_cell[   22986] = 32'ha0e2fa65;
    ram_cell[   22987] = 32'h07244d66;
    ram_cell[   22988] = 32'hf397a057;
    ram_cell[   22989] = 32'h1f4fd1ad;
    ram_cell[   22990] = 32'heeb4793c;
    ram_cell[   22991] = 32'h331a3d41;
    ram_cell[   22992] = 32'h706ea2d5;
    ram_cell[   22993] = 32'hf0ea18f6;
    ram_cell[   22994] = 32'h3909e114;
    ram_cell[   22995] = 32'h1556ba26;
    ram_cell[   22996] = 32'h698425ff;
    ram_cell[   22997] = 32'hedc50c41;
    ram_cell[   22998] = 32'h361bf268;
    ram_cell[   22999] = 32'hae2ebae5;
    ram_cell[   23000] = 32'h7a329994;
    ram_cell[   23001] = 32'hc886a607;
    ram_cell[   23002] = 32'hc4a0fc26;
    ram_cell[   23003] = 32'h9edff478;
    ram_cell[   23004] = 32'h95d18f70;
    ram_cell[   23005] = 32'he97abbf0;
    ram_cell[   23006] = 32'heedcfc65;
    ram_cell[   23007] = 32'h493c5119;
    ram_cell[   23008] = 32'hf9d79cbd;
    ram_cell[   23009] = 32'hafd1a8d9;
    ram_cell[   23010] = 32'h3a840df2;
    ram_cell[   23011] = 32'ha43a2b0e;
    ram_cell[   23012] = 32'ha015b339;
    ram_cell[   23013] = 32'h2b9326f6;
    ram_cell[   23014] = 32'hb0eca27b;
    ram_cell[   23015] = 32'haaea6d04;
    ram_cell[   23016] = 32'h9fdad56d;
    ram_cell[   23017] = 32'h4b452f69;
    ram_cell[   23018] = 32'h940b3889;
    ram_cell[   23019] = 32'hd1f18a30;
    ram_cell[   23020] = 32'hb6e3dc09;
    ram_cell[   23021] = 32'h9a66ddd7;
    ram_cell[   23022] = 32'hc92a7a8b;
    ram_cell[   23023] = 32'h2203b0ca;
    ram_cell[   23024] = 32'hc346b9b2;
    ram_cell[   23025] = 32'hae8fac2d;
    ram_cell[   23026] = 32'h163b897c;
    ram_cell[   23027] = 32'h88ba56ce;
    ram_cell[   23028] = 32'h49c7c41c;
    ram_cell[   23029] = 32'h272fedc6;
    ram_cell[   23030] = 32'h7d7439e1;
    ram_cell[   23031] = 32'hedbb436e;
    ram_cell[   23032] = 32'ha8e71fff;
    ram_cell[   23033] = 32'h9e9149df;
    ram_cell[   23034] = 32'hb048d848;
    ram_cell[   23035] = 32'h82634411;
    ram_cell[   23036] = 32'hf791f9ab;
    ram_cell[   23037] = 32'h23912151;
    ram_cell[   23038] = 32'h20870680;
    ram_cell[   23039] = 32'h5c4350b7;
    ram_cell[   23040] = 32'h0b822f31;
    ram_cell[   23041] = 32'h27cdc143;
    ram_cell[   23042] = 32'h2b85eca6;
    ram_cell[   23043] = 32'h044b3de8;
    ram_cell[   23044] = 32'hdeb78bde;
    ram_cell[   23045] = 32'h094b0df0;
    ram_cell[   23046] = 32'h55069069;
    ram_cell[   23047] = 32'h3c3a0af0;
    ram_cell[   23048] = 32'hd8e5585a;
    ram_cell[   23049] = 32'h3f53b072;
    ram_cell[   23050] = 32'h217e4055;
    ram_cell[   23051] = 32'h17ceb8e3;
    ram_cell[   23052] = 32'hfaa12e93;
    ram_cell[   23053] = 32'h20db804e;
    ram_cell[   23054] = 32'h0416ecbd;
    ram_cell[   23055] = 32'h488ffde1;
    ram_cell[   23056] = 32'hd470f070;
    ram_cell[   23057] = 32'hd3643f30;
    ram_cell[   23058] = 32'hc1519fa9;
    ram_cell[   23059] = 32'haae0d597;
    ram_cell[   23060] = 32'hd54838e8;
    ram_cell[   23061] = 32'ha12c6524;
    ram_cell[   23062] = 32'he6e56401;
    ram_cell[   23063] = 32'h038f65c2;
    ram_cell[   23064] = 32'he0f3b8a7;
    ram_cell[   23065] = 32'hdaba928d;
    ram_cell[   23066] = 32'h6fc486c5;
    ram_cell[   23067] = 32'hcc27c159;
    ram_cell[   23068] = 32'h188cf9d1;
    ram_cell[   23069] = 32'ha1bc05ad;
    ram_cell[   23070] = 32'h1727b34d;
    ram_cell[   23071] = 32'hd8f09088;
    ram_cell[   23072] = 32'he4d057fc;
    ram_cell[   23073] = 32'h0e79d9f6;
    ram_cell[   23074] = 32'hef177dfd;
    ram_cell[   23075] = 32'h999280cb;
    ram_cell[   23076] = 32'h2394e9db;
    ram_cell[   23077] = 32'h7c82af7c;
    ram_cell[   23078] = 32'hc2a8e90c;
    ram_cell[   23079] = 32'h93b60eb1;
    ram_cell[   23080] = 32'hbe40992e;
    ram_cell[   23081] = 32'h1b515d69;
    ram_cell[   23082] = 32'h07b7b0dd;
    ram_cell[   23083] = 32'hdda7e4e4;
    ram_cell[   23084] = 32'h7edaae22;
    ram_cell[   23085] = 32'hf37b9ed1;
    ram_cell[   23086] = 32'h7f5e7c1a;
    ram_cell[   23087] = 32'h5b40f2e7;
    ram_cell[   23088] = 32'h79f4a3c0;
    ram_cell[   23089] = 32'h189f0157;
    ram_cell[   23090] = 32'h5e96cb85;
    ram_cell[   23091] = 32'hf878e707;
    ram_cell[   23092] = 32'h3019cef4;
    ram_cell[   23093] = 32'h8035a1de;
    ram_cell[   23094] = 32'h24cc5a74;
    ram_cell[   23095] = 32'h0e8a7e92;
    ram_cell[   23096] = 32'h8e8ad5ea;
    ram_cell[   23097] = 32'ha895f047;
    ram_cell[   23098] = 32'h7ba510d7;
    ram_cell[   23099] = 32'h97631e02;
    ram_cell[   23100] = 32'h90cbd426;
    ram_cell[   23101] = 32'he398cd68;
    ram_cell[   23102] = 32'h10a38364;
    ram_cell[   23103] = 32'hcf3bae82;
    ram_cell[   23104] = 32'h4ce7b383;
    ram_cell[   23105] = 32'hbc133ca8;
    ram_cell[   23106] = 32'h5a2f2682;
    ram_cell[   23107] = 32'h5141449d;
    ram_cell[   23108] = 32'hf4d6ada5;
    ram_cell[   23109] = 32'hb470c38f;
    ram_cell[   23110] = 32'h85b05bbb;
    ram_cell[   23111] = 32'hb3741b00;
    ram_cell[   23112] = 32'h8c722dfe;
    ram_cell[   23113] = 32'h43b39d08;
    ram_cell[   23114] = 32'hb1cb5412;
    ram_cell[   23115] = 32'h86bf0ed7;
    ram_cell[   23116] = 32'h1a61de8a;
    ram_cell[   23117] = 32'hbe217792;
    ram_cell[   23118] = 32'h4ce15128;
    ram_cell[   23119] = 32'h06ca813a;
    ram_cell[   23120] = 32'h94780d2a;
    ram_cell[   23121] = 32'h430e9299;
    ram_cell[   23122] = 32'h7a00b80f;
    ram_cell[   23123] = 32'ha40f7402;
    ram_cell[   23124] = 32'h5d3e27c0;
    ram_cell[   23125] = 32'he7d13832;
    ram_cell[   23126] = 32'h6de5b94f;
    ram_cell[   23127] = 32'h54fb4c1b;
    ram_cell[   23128] = 32'hf7f13c05;
    ram_cell[   23129] = 32'h1b307a9a;
    ram_cell[   23130] = 32'hfb20c7ea;
    ram_cell[   23131] = 32'h81823435;
    ram_cell[   23132] = 32'h716673fb;
    ram_cell[   23133] = 32'had3de595;
    ram_cell[   23134] = 32'h26252383;
    ram_cell[   23135] = 32'h913d6908;
    ram_cell[   23136] = 32'he7789661;
    ram_cell[   23137] = 32'h859e5816;
    ram_cell[   23138] = 32'hfc1adb3c;
    ram_cell[   23139] = 32'h1aeff135;
    ram_cell[   23140] = 32'h768a67cd;
    ram_cell[   23141] = 32'hcb8cf68d;
    ram_cell[   23142] = 32'h3bdaba11;
    ram_cell[   23143] = 32'h2b97a770;
    ram_cell[   23144] = 32'hbff5cd4b;
    ram_cell[   23145] = 32'h1f1182c9;
    ram_cell[   23146] = 32'h96fceb82;
    ram_cell[   23147] = 32'h9952e642;
    ram_cell[   23148] = 32'hfc02888f;
    ram_cell[   23149] = 32'h4181da45;
    ram_cell[   23150] = 32'h6f8a180a;
    ram_cell[   23151] = 32'h9263e114;
    ram_cell[   23152] = 32'h34ad6ac5;
    ram_cell[   23153] = 32'hd0dd8d18;
    ram_cell[   23154] = 32'h78f0f205;
    ram_cell[   23155] = 32'h5dc3df15;
    ram_cell[   23156] = 32'hbb9a785b;
    ram_cell[   23157] = 32'hff84dfdd;
    ram_cell[   23158] = 32'hc7676381;
    ram_cell[   23159] = 32'h479a2b2a;
    ram_cell[   23160] = 32'hb0ee7ad9;
    ram_cell[   23161] = 32'h0cdc8f4b;
    ram_cell[   23162] = 32'ha0d79d9e;
    ram_cell[   23163] = 32'h84d823c1;
    ram_cell[   23164] = 32'hca467a00;
    ram_cell[   23165] = 32'hdaa94947;
    ram_cell[   23166] = 32'h867fc919;
    ram_cell[   23167] = 32'hc4612272;
    ram_cell[   23168] = 32'h437fc6ae;
    ram_cell[   23169] = 32'h0e1803bf;
    ram_cell[   23170] = 32'hce11face;
    ram_cell[   23171] = 32'hec2b9b18;
    ram_cell[   23172] = 32'hf2003814;
    ram_cell[   23173] = 32'hb21d2017;
    ram_cell[   23174] = 32'h5baab06e;
    ram_cell[   23175] = 32'h602eba43;
    ram_cell[   23176] = 32'h1dbd4cd7;
    ram_cell[   23177] = 32'h17783f95;
    ram_cell[   23178] = 32'hc86877db;
    ram_cell[   23179] = 32'h661c1b60;
    ram_cell[   23180] = 32'h0219a616;
    ram_cell[   23181] = 32'h0469de48;
    ram_cell[   23182] = 32'hd3b1878e;
    ram_cell[   23183] = 32'hb501a7d9;
    ram_cell[   23184] = 32'h45a2a30c;
    ram_cell[   23185] = 32'h99d307e9;
    ram_cell[   23186] = 32'ha083a425;
    ram_cell[   23187] = 32'he4bfd1e5;
    ram_cell[   23188] = 32'h38d3fcb2;
    ram_cell[   23189] = 32'h41226914;
    ram_cell[   23190] = 32'ha2d94ec6;
    ram_cell[   23191] = 32'h75fb7302;
    ram_cell[   23192] = 32'h9596a807;
    ram_cell[   23193] = 32'h36d21e2c;
    ram_cell[   23194] = 32'h401a3fe2;
    ram_cell[   23195] = 32'hf779a5dd;
    ram_cell[   23196] = 32'h7004f3a0;
    ram_cell[   23197] = 32'had01e640;
    ram_cell[   23198] = 32'h55ad032a;
    ram_cell[   23199] = 32'h079d488b;
    ram_cell[   23200] = 32'h602c49a5;
    ram_cell[   23201] = 32'hb0df4227;
    ram_cell[   23202] = 32'hfa884c46;
    ram_cell[   23203] = 32'ha75dd2d7;
    ram_cell[   23204] = 32'hd77af055;
    ram_cell[   23205] = 32'hfaed2a89;
    ram_cell[   23206] = 32'h9020da8b;
    ram_cell[   23207] = 32'h038596fe;
    ram_cell[   23208] = 32'hcfe0023e;
    ram_cell[   23209] = 32'h641ccf22;
    ram_cell[   23210] = 32'h2cff9296;
    ram_cell[   23211] = 32'h8c644bdc;
    ram_cell[   23212] = 32'h4c43ae2c;
    ram_cell[   23213] = 32'hdad42384;
    ram_cell[   23214] = 32'hdfb93999;
    ram_cell[   23215] = 32'hf9b509ff;
    ram_cell[   23216] = 32'h49b3d895;
    ram_cell[   23217] = 32'h949fabd9;
    ram_cell[   23218] = 32'hc8d73842;
    ram_cell[   23219] = 32'h0f0db497;
    ram_cell[   23220] = 32'hf38331b9;
    ram_cell[   23221] = 32'h78f997c9;
    ram_cell[   23222] = 32'h00542572;
    ram_cell[   23223] = 32'haf7c1354;
    ram_cell[   23224] = 32'h79ee9e6c;
    ram_cell[   23225] = 32'h26da5d1b;
    ram_cell[   23226] = 32'h6e8e7ded;
    ram_cell[   23227] = 32'hacc3eef9;
    ram_cell[   23228] = 32'hfb672c09;
    ram_cell[   23229] = 32'h92f7bcf5;
    ram_cell[   23230] = 32'h172ef4ec;
    ram_cell[   23231] = 32'h2b302899;
    ram_cell[   23232] = 32'h074e2e8e;
    ram_cell[   23233] = 32'hd202b669;
    ram_cell[   23234] = 32'h9936b2e7;
    ram_cell[   23235] = 32'h4b12b730;
    ram_cell[   23236] = 32'h32b0455b;
    ram_cell[   23237] = 32'h04870f6f;
    ram_cell[   23238] = 32'hf7f9a7ab;
    ram_cell[   23239] = 32'h6236f19f;
    ram_cell[   23240] = 32'h80922be7;
    ram_cell[   23241] = 32'h1f290c27;
    ram_cell[   23242] = 32'hf1183d47;
    ram_cell[   23243] = 32'hb2358c07;
    ram_cell[   23244] = 32'hbb22cc5c;
    ram_cell[   23245] = 32'h2e8fce3a;
    ram_cell[   23246] = 32'h4bf7cc1c;
    ram_cell[   23247] = 32'h2aa956ea;
    ram_cell[   23248] = 32'h4b3ec79d;
    ram_cell[   23249] = 32'h326e6e7a;
    ram_cell[   23250] = 32'h779f9eed;
    ram_cell[   23251] = 32'h11ea6261;
    ram_cell[   23252] = 32'hea278dd6;
    ram_cell[   23253] = 32'h987cf96a;
    ram_cell[   23254] = 32'hf9584386;
    ram_cell[   23255] = 32'h71a73d84;
    ram_cell[   23256] = 32'h08c48082;
    ram_cell[   23257] = 32'hd3d1bf4b;
    ram_cell[   23258] = 32'h7731ce92;
    ram_cell[   23259] = 32'h82c55df5;
    ram_cell[   23260] = 32'h29b96e36;
    ram_cell[   23261] = 32'h6c2d23c7;
    ram_cell[   23262] = 32'h4712f9da;
    ram_cell[   23263] = 32'ha938e56c;
    ram_cell[   23264] = 32'h868cd568;
    ram_cell[   23265] = 32'hdde0a70a;
    ram_cell[   23266] = 32'hd4c5ca16;
    ram_cell[   23267] = 32'haa7442a2;
    ram_cell[   23268] = 32'hc738d174;
    ram_cell[   23269] = 32'hdb4b8d06;
    ram_cell[   23270] = 32'hd6ffe151;
    ram_cell[   23271] = 32'ha9988999;
    ram_cell[   23272] = 32'h50348035;
    ram_cell[   23273] = 32'h58c16110;
    ram_cell[   23274] = 32'h04cad09e;
    ram_cell[   23275] = 32'hfe0dfcfd;
    ram_cell[   23276] = 32'h14913220;
    ram_cell[   23277] = 32'h3b1dd30b;
    ram_cell[   23278] = 32'ha4bd9b54;
    ram_cell[   23279] = 32'h631d57b8;
    ram_cell[   23280] = 32'h440b6b12;
    ram_cell[   23281] = 32'h39ef5839;
    ram_cell[   23282] = 32'h79509343;
    ram_cell[   23283] = 32'h2e9179ad;
    ram_cell[   23284] = 32'ha4851339;
    ram_cell[   23285] = 32'h07797975;
    ram_cell[   23286] = 32'h11efa595;
    ram_cell[   23287] = 32'h6987d138;
    ram_cell[   23288] = 32'h9de78962;
    ram_cell[   23289] = 32'h716d2c6b;
    ram_cell[   23290] = 32'h20c501ef;
    ram_cell[   23291] = 32'h0104129c;
    ram_cell[   23292] = 32'h6c024b1b;
    ram_cell[   23293] = 32'haa1928e5;
    ram_cell[   23294] = 32'hb8ed3e53;
    ram_cell[   23295] = 32'h0dc91853;
    ram_cell[   23296] = 32'hc3041e7f;
    ram_cell[   23297] = 32'h06369b3b;
    ram_cell[   23298] = 32'h2f2f1f3d;
    ram_cell[   23299] = 32'h3e94c68e;
    ram_cell[   23300] = 32'heea9783c;
    ram_cell[   23301] = 32'h9e2eab58;
    ram_cell[   23302] = 32'h8fa24b43;
    ram_cell[   23303] = 32'h7f067611;
    ram_cell[   23304] = 32'h2385ad2b;
    ram_cell[   23305] = 32'hfd696ad5;
    ram_cell[   23306] = 32'h71b8ad68;
    ram_cell[   23307] = 32'h24def7a6;
    ram_cell[   23308] = 32'h0372683a;
    ram_cell[   23309] = 32'hc46e0290;
    ram_cell[   23310] = 32'hdd7ea260;
    ram_cell[   23311] = 32'h2aca5e3a;
    ram_cell[   23312] = 32'h5cbc985c;
    ram_cell[   23313] = 32'h7229d7f5;
    ram_cell[   23314] = 32'h37135ab4;
    ram_cell[   23315] = 32'h1df7e666;
    ram_cell[   23316] = 32'h33e94651;
    ram_cell[   23317] = 32'h424589e1;
    ram_cell[   23318] = 32'h3c49579c;
    ram_cell[   23319] = 32'ha6aa94a5;
    ram_cell[   23320] = 32'he006519c;
    ram_cell[   23321] = 32'h20c4c17a;
    ram_cell[   23322] = 32'hef20ec0a;
    ram_cell[   23323] = 32'h99e0d789;
    ram_cell[   23324] = 32'h84272688;
    ram_cell[   23325] = 32'h5de30c73;
    ram_cell[   23326] = 32'h1dba0815;
    ram_cell[   23327] = 32'h4094fad2;
    ram_cell[   23328] = 32'h5a5701de;
    ram_cell[   23329] = 32'h9c7dd80b;
    ram_cell[   23330] = 32'h16047fc0;
    ram_cell[   23331] = 32'hb11c11c4;
    ram_cell[   23332] = 32'h01f32d5e;
    ram_cell[   23333] = 32'h24c98450;
    ram_cell[   23334] = 32'hc380d772;
    ram_cell[   23335] = 32'h6954763b;
    ram_cell[   23336] = 32'h3d56840b;
    ram_cell[   23337] = 32'h2c65afd8;
    ram_cell[   23338] = 32'h5685455d;
    ram_cell[   23339] = 32'h9ae93d55;
    ram_cell[   23340] = 32'h9a652eb1;
    ram_cell[   23341] = 32'h895b6e76;
    ram_cell[   23342] = 32'hddfa8ca8;
    ram_cell[   23343] = 32'h166f8b93;
    ram_cell[   23344] = 32'h5fe738a2;
    ram_cell[   23345] = 32'h29610819;
    ram_cell[   23346] = 32'h434218ce;
    ram_cell[   23347] = 32'h0ae82b80;
    ram_cell[   23348] = 32'h9460d5c8;
    ram_cell[   23349] = 32'hceb5a853;
    ram_cell[   23350] = 32'ha61bc29e;
    ram_cell[   23351] = 32'hc107716c;
    ram_cell[   23352] = 32'h9c975dd7;
    ram_cell[   23353] = 32'hee170f35;
    ram_cell[   23354] = 32'hf7927de4;
    ram_cell[   23355] = 32'h3cbf8f1d;
    ram_cell[   23356] = 32'h5eb2862e;
    ram_cell[   23357] = 32'h87221e21;
    ram_cell[   23358] = 32'hb8abb2cc;
    ram_cell[   23359] = 32'h4843950f;
    ram_cell[   23360] = 32'hdadc4217;
    ram_cell[   23361] = 32'hc2dd0cc3;
    ram_cell[   23362] = 32'h10b72997;
    ram_cell[   23363] = 32'ha924e660;
    ram_cell[   23364] = 32'h49c15d92;
    ram_cell[   23365] = 32'h8acdb68e;
    ram_cell[   23366] = 32'h85d1686a;
    ram_cell[   23367] = 32'hb90fdd3e;
    ram_cell[   23368] = 32'hcc335989;
    ram_cell[   23369] = 32'h8a4579bc;
    ram_cell[   23370] = 32'h8357b7c0;
    ram_cell[   23371] = 32'h74f83d3f;
    ram_cell[   23372] = 32'hd439e31f;
    ram_cell[   23373] = 32'h7856f60e;
    ram_cell[   23374] = 32'h50b0c3e0;
    ram_cell[   23375] = 32'h023cacbb;
    ram_cell[   23376] = 32'hd6ae3d52;
    ram_cell[   23377] = 32'h6d2663da;
    ram_cell[   23378] = 32'hddeb9e66;
    ram_cell[   23379] = 32'h2c2327cc;
    ram_cell[   23380] = 32'h6d50bf19;
    ram_cell[   23381] = 32'h64902dc5;
    ram_cell[   23382] = 32'he864de6a;
    ram_cell[   23383] = 32'h2687a2c6;
    ram_cell[   23384] = 32'h1324f7cc;
    ram_cell[   23385] = 32'h570471a5;
    ram_cell[   23386] = 32'h968cfde1;
    ram_cell[   23387] = 32'h475e2a14;
    ram_cell[   23388] = 32'hd960c5a6;
    ram_cell[   23389] = 32'h921c946f;
    ram_cell[   23390] = 32'h541705a4;
    ram_cell[   23391] = 32'h2580c7ce;
    ram_cell[   23392] = 32'h5aecbdc7;
    ram_cell[   23393] = 32'haffd1644;
    ram_cell[   23394] = 32'h6f8e57b8;
    ram_cell[   23395] = 32'ha3b1eb02;
    ram_cell[   23396] = 32'hf152b5a6;
    ram_cell[   23397] = 32'haf6e8619;
    ram_cell[   23398] = 32'h4e4c6f63;
    ram_cell[   23399] = 32'h5935486e;
    ram_cell[   23400] = 32'hf5e4afd5;
    ram_cell[   23401] = 32'hdec25c68;
    ram_cell[   23402] = 32'h9ac11385;
    ram_cell[   23403] = 32'h67bdafd2;
    ram_cell[   23404] = 32'h5efc984e;
    ram_cell[   23405] = 32'h22b7180e;
    ram_cell[   23406] = 32'hd0840e7a;
    ram_cell[   23407] = 32'hc6e3484c;
    ram_cell[   23408] = 32'h39114f7a;
    ram_cell[   23409] = 32'h286d8cea;
    ram_cell[   23410] = 32'h168efb33;
    ram_cell[   23411] = 32'h3037f041;
    ram_cell[   23412] = 32'h6a2e2072;
    ram_cell[   23413] = 32'hfae57152;
    ram_cell[   23414] = 32'h7d9e6f2a;
    ram_cell[   23415] = 32'hd85caedc;
    ram_cell[   23416] = 32'h382a96df;
    ram_cell[   23417] = 32'h5a5e2105;
    ram_cell[   23418] = 32'ha424026e;
    ram_cell[   23419] = 32'hd92ec1bc;
    ram_cell[   23420] = 32'h5684ae54;
    ram_cell[   23421] = 32'h49c70d68;
    ram_cell[   23422] = 32'h34958b28;
    ram_cell[   23423] = 32'h14123af7;
    ram_cell[   23424] = 32'h82473beb;
    ram_cell[   23425] = 32'hf3023f6a;
    ram_cell[   23426] = 32'h54b68fa0;
    ram_cell[   23427] = 32'h44e0d825;
    ram_cell[   23428] = 32'h2602cec1;
    ram_cell[   23429] = 32'hd6678d53;
    ram_cell[   23430] = 32'h311be3b2;
    ram_cell[   23431] = 32'h9336a948;
    ram_cell[   23432] = 32'h623a9dc4;
    ram_cell[   23433] = 32'h5241c844;
    ram_cell[   23434] = 32'h3f58a464;
    ram_cell[   23435] = 32'h65c32825;
    ram_cell[   23436] = 32'h31b4412b;
    ram_cell[   23437] = 32'h1798fabe;
    ram_cell[   23438] = 32'h962396a2;
    ram_cell[   23439] = 32'h7ae11291;
    ram_cell[   23440] = 32'h0c159624;
    ram_cell[   23441] = 32'heb7b0de7;
    ram_cell[   23442] = 32'h52f76fc7;
    ram_cell[   23443] = 32'h1c8a4101;
    ram_cell[   23444] = 32'hc0bba836;
    ram_cell[   23445] = 32'hfd5bb0d9;
    ram_cell[   23446] = 32'h20555f33;
    ram_cell[   23447] = 32'h67b053b6;
    ram_cell[   23448] = 32'h77f6ee42;
    ram_cell[   23449] = 32'h0dd2a39d;
    ram_cell[   23450] = 32'h5c315e74;
    ram_cell[   23451] = 32'hc82b4166;
    ram_cell[   23452] = 32'h2ae3abcf;
    ram_cell[   23453] = 32'h9744424e;
    ram_cell[   23454] = 32'h3492eec5;
    ram_cell[   23455] = 32'h9c1eb125;
    ram_cell[   23456] = 32'hf6e9bb69;
    ram_cell[   23457] = 32'h284e8d64;
    ram_cell[   23458] = 32'h0d7cc3c1;
    ram_cell[   23459] = 32'h78ca6f36;
    ram_cell[   23460] = 32'h7681ac9f;
    ram_cell[   23461] = 32'h4177b94f;
    ram_cell[   23462] = 32'h1c9a3a85;
    ram_cell[   23463] = 32'ha57cf7e6;
    ram_cell[   23464] = 32'h6e1863f1;
    ram_cell[   23465] = 32'h3965ab5c;
    ram_cell[   23466] = 32'h3650d174;
    ram_cell[   23467] = 32'hf9bf0c7c;
    ram_cell[   23468] = 32'h84ded4ee;
    ram_cell[   23469] = 32'hfffdf9ba;
    ram_cell[   23470] = 32'hd3910ca9;
    ram_cell[   23471] = 32'h832f9b76;
    ram_cell[   23472] = 32'ha0ffe309;
    ram_cell[   23473] = 32'h9b4fa1a8;
    ram_cell[   23474] = 32'h628b0403;
    ram_cell[   23475] = 32'h5050ee63;
    ram_cell[   23476] = 32'h73f89239;
    ram_cell[   23477] = 32'h5f1dd393;
    ram_cell[   23478] = 32'hfe0ec2bb;
    ram_cell[   23479] = 32'hadfcfa18;
    ram_cell[   23480] = 32'hd6c7afd5;
    ram_cell[   23481] = 32'hbe3b6502;
    ram_cell[   23482] = 32'h01234327;
    ram_cell[   23483] = 32'hda9e7c90;
    ram_cell[   23484] = 32'hd07466df;
    ram_cell[   23485] = 32'hcde7303e;
    ram_cell[   23486] = 32'h4c5594a0;
    ram_cell[   23487] = 32'h664617e4;
    ram_cell[   23488] = 32'h971ef66f;
    ram_cell[   23489] = 32'h7b435630;
    ram_cell[   23490] = 32'hcc6fc229;
    ram_cell[   23491] = 32'h74ad2805;
    ram_cell[   23492] = 32'hfade6457;
    ram_cell[   23493] = 32'h9dc10b77;
    ram_cell[   23494] = 32'hab02cb32;
    ram_cell[   23495] = 32'h42155514;
    ram_cell[   23496] = 32'h122d6f5c;
    ram_cell[   23497] = 32'h27924f9a;
    ram_cell[   23498] = 32'hab3c6324;
    ram_cell[   23499] = 32'hf3b262c6;
    ram_cell[   23500] = 32'h5785dfdc;
    ram_cell[   23501] = 32'h17b2817d;
    ram_cell[   23502] = 32'hcf6becf0;
    ram_cell[   23503] = 32'he3070e0d;
    ram_cell[   23504] = 32'h478674c4;
    ram_cell[   23505] = 32'h0359d43b;
    ram_cell[   23506] = 32'h8933b065;
    ram_cell[   23507] = 32'hdf997949;
    ram_cell[   23508] = 32'hdbaa5919;
    ram_cell[   23509] = 32'h5ff8cac8;
    ram_cell[   23510] = 32'hc6297354;
    ram_cell[   23511] = 32'h93e57e9a;
    ram_cell[   23512] = 32'h8971b599;
    ram_cell[   23513] = 32'h2782e49d;
    ram_cell[   23514] = 32'hf2f1a6ee;
    ram_cell[   23515] = 32'h3961065b;
    ram_cell[   23516] = 32'h873ec9f5;
    ram_cell[   23517] = 32'hba3130b2;
    ram_cell[   23518] = 32'hc05ed70d;
    ram_cell[   23519] = 32'hb8ccdb75;
    ram_cell[   23520] = 32'hc8ae745c;
    ram_cell[   23521] = 32'h3ed7b0b8;
    ram_cell[   23522] = 32'h4b764e1e;
    ram_cell[   23523] = 32'he3016784;
    ram_cell[   23524] = 32'hea979d3a;
    ram_cell[   23525] = 32'h699e02b1;
    ram_cell[   23526] = 32'h824764f9;
    ram_cell[   23527] = 32'h63f9b72d;
    ram_cell[   23528] = 32'h4f872c62;
    ram_cell[   23529] = 32'hed14a418;
    ram_cell[   23530] = 32'h375c653a;
    ram_cell[   23531] = 32'hde9b36ac;
    ram_cell[   23532] = 32'hd1a6e36e;
    ram_cell[   23533] = 32'he88be08a;
    ram_cell[   23534] = 32'hb19e3a6d;
    ram_cell[   23535] = 32'hd34f61e0;
    ram_cell[   23536] = 32'hc69a0033;
    ram_cell[   23537] = 32'h8c758a58;
    ram_cell[   23538] = 32'h79729816;
    ram_cell[   23539] = 32'h79931bf7;
    ram_cell[   23540] = 32'hb5b4f3e5;
    ram_cell[   23541] = 32'hb01acbfb;
    ram_cell[   23542] = 32'haf0a02a3;
    ram_cell[   23543] = 32'h47246a3e;
    ram_cell[   23544] = 32'hd376532e;
    ram_cell[   23545] = 32'h2ef3df23;
    ram_cell[   23546] = 32'ha38a4d66;
    ram_cell[   23547] = 32'ha01986c9;
    ram_cell[   23548] = 32'he12f0d92;
    ram_cell[   23549] = 32'h920c0334;
    ram_cell[   23550] = 32'h42389da5;
    ram_cell[   23551] = 32'h5985a02d;
    ram_cell[   23552] = 32'h18071612;
    ram_cell[   23553] = 32'hfe849f35;
    ram_cell[   23554] = 32'h82e06b5d;
    ram_cell[   23555] = 32'h30a4d68d;
    ram_cell[   23556] = 32'hdc9f0cd7;
    ram_cell[   23557] = 32'hf0d015ca;
    ram_cell[   23558] = 32'h8bbcf339;
    ram_cell[   23559] = 32'h5596daba;
    ram_cell[   23560] = 32'h7cfa0d3a;
    ram_cell[   23561] = 32'h59666808;
    ram_cell[   23562] = 32'h21be1822;
    ram_cell[   23563] = 32'hf3fcf0b8;
    ram_cell[   23564] = 32'h68312f74;
    ram_cell[   23565] = 32'h23b3f877;
    ram_cell[   23566] = 32'hd30d97ff;
    ram_cell[   23567] = 32'h31286cac;
    ram_cell[   23568] = 32'h4c5ca59a;
    ram_cell[   23569] = 32'hfefc6861;
    ram_cell[   23570] = 32'h77005032;
    ram_cell[   23571] = 32'hd604796d;
    ram_cell[   23572] = 32'h27d1c949;
    ram_cell[   23573] = 32'hd14b290d;
    ram_cell[   23574] = 32'h5cd36e0f;
    ram_cell[   23575] = 32'h6c7f7e36;
    ram_cell[   23576] = 32'h8aa8cf8e;
    ram_cell[   23577] = 32'hf3f609ee;
    ram_cell[   23578] = 32'hfaf78001;
    ram_cell[   23579] = 32'h0c7087bb;
    ram_cell[   23580] = 32'haa1c8445;
    ram_cell[   23581] = 32'hca18e908;
    ram_cell[   23582] = 32'h70918094;
    ram_cell[   23583] = 32'hae088856;
    ram_cell[   23584] = 32'h32275f58;
    ram_cell[   23585] = 32'h6df1d3b0;
    ram_cell[   23586] = 32'hecfdf801;
    ram_cell[   23587] = 32'h0936830e;
    ram_cell[   23588] = 32'h94cd8594;
    ram_cell[   23589] = 32'ha10986b2;
    ram_cell[   23590] = 32'h6993212c;
    ram_cell[   23591] = 32'h80bf5ffb;
    ram_cell[   23592] = 32'h47633990;
    ram_cell[   23593] = 32'h0bd10e72;
    ram_cell[   23594] = 32'hf9198e94;
    ram_cell[   23595] = 32'h7a1a55fb;
    ram_cell[   23596] = 32'hdc78bf4b;
    ram_cell[   23597] = 32'hb1d058a2;
    ram_cell[   23598] = 32'hcc37f355;
    ram_cell[   23599] = 32'h38a7c17a;
    ram_cell[   23600] = 32'he0557faf;
    ram_cell[   23601] = 32'h5c38b553;
    ram_cell[   23602] = 32'h45492690;
    ram_cell[   23603] = 32'h760bf575;
    ram_cell[   23604] = 32'h61f9fe26;
    ram_cell[   23605] = 32'h9bacdac8;
    ram_cell[   23606] = 32'h2845081b;
    ram_cell[   23607] = 32'haa97373a;
    ram_cell[   23608] = 32'h273ddb82;
    ram_cell[   23609] = 32'h89cee46e;
    ram_cell[   23610] = 32'ha3e18ec2;
    ram_cell[   23611] = 32'h844b2b42;
    ram_cell[   23612] = 32'hda99f30e;
    ram_cell[   23613] = 32'hb7f4cdc7;
    ram_cell[   23614] = 32'h7fe500f0;
    ram_cell[   23615] = 32'hd6fe0436;
    ram_cell[   23616] = 32'h39b9b96b;
    ram_cell[   23617] = 32'hd66adb8b;
    ram_cell[   23618] = 32'h9f82467c;
    ram_cell[   23619] = 32'h3934c852;
    ram_cell[   23620] = 32'h81d5629b;
    ram_cell[   23621] = 32'he1121705;
    ram_cell[   23622] = 32'h4b5abb69;
    ram_cell[   23623] = 32'h05ce0dfa;
    ram_cell[   23624] = 32'h306dadbb;
    ram_cell[   23625] = 32'hc94ef2cd;
    ram_cell[   23626] = 32'hdfdb4b03;
    ram_cell[   23627] = 32'hd614761b;
    ram_cell[   23628] = 32'h17565a70;
    ram_cell[   23629] = 32'hde33f204;
    ram_cell[   23630] = 32'hdeb5ab33;
    ram_cell[   23631] = 32'h5be7a01b;
    ram_cell[   23632] = 32'hf07f93a8;
    ram_cell[   23633] = 32'h533ae1a6;
    ram_cell[   23634] = 32'hb7e27dec;
    ram_cell[   23635] = 32'h780bf316;
    ram_cell[   23636] = 32'h2078dd04;
    ram_cell[   23637] = 32'h3534581b;
    ram_cell[   23638] = 32'h009ca276;
    ram_cell[   23639] = 32'h6e404aef;
    ram_cell[   23640] = 32'h844f15bb;
    ram_cell[   23641] = 32'h912d6d0a;
    ram_cell[   23642] = 32'hd39e6165;
    ram_cell[   23643] = 32'hfdd6f0e8;
    ram_cell[   23644] = 32'hcafa49a2;
    ram_cell[   23645] = 32'h7945e978;
    ram_cell[   23646] = 32'h3dd10755;
    ram_cell[   23647] = 32'hd38e6925;
    ram_cell[   23648] = 32'h45847f88;
    ram_cell[   23649] = 32'h88252335;
    ram_cell[   23650] = 32'hb8cd78d0;
    ram_cell[   23651] = 32'ha84d8cf7;
    ram_cell[   23652] = 32'h190e1528;
    ram_cell[   23653] = 32'h69a49aee;
    ram_cell[   23654] = 32'h5c155bdc;
    ram_cell[   23655] = 32'h4c2365a2;
    ram_cell[   23656] = 32'h097d235e;
    ram_cell[   23657] = 32'h02fa24ae;
    ram_cell[   23658] = 32'hf25945fb;
    ram_cell[   23659] = 32'haa3100f8;
    ram_cell[   23660] = 32'h9c972876;
    ram_cell[   23661] = 32'h5e53b5f6;
    ram_cell[   23662] = 32'h4a6e3b60;
    ram_cell[   23663] = 32'h5a64eb30;
    ram_cell[   23664] = 32'h3fb508ab;
    ram_cell[   23665] = 32'h2f443ca1;
    ram_cell[   23666] = 32'ha28a234a;
    ram_cell[   23667] = 32'ha53c5054;
    ram_cell[   23668] = 32'h3458b439;
    ram_cell[   23669] = 32'hf3db4787;
    ram_cell[   23670] = 32'hb0661618;
    ram_cell[   23671] = 32'h97b21501;
    ram_cell[   23672] = 32'hf4f2f59f;
    ram_cell[   23673] = 32'hf20fb44f;
    ram_cell[   23674] = 32'h9c799cd5;
    ram_cell[   23675] = 32'h55e76207;
    ram_cell[   23676] = 32'h33bb0eb4;
    ram_cell[   23677] = 32'h57505c3b;
    ram_cell[   23678] = 32'hfd1cf457;
    ram_cell[   23679] = 32'h37a7d418;
    ram_cell[   23680] = 32'h22ad6757;
    ram_cell[   23681] = 32'h5f04fb60;
    ram_cell[   23682] = 32'h205ffc22;
    ram_cell[   23683] = 32'h4ba9f3a9;
    ram_cell[   23684] = 32'h268b3dee;
    ram_cell[   23685] = 32'hc265f762;
    ram_cell[   23686] = 32'h6de20617;
    ram_cell[   23687] = 32'ha5a2f126;
    ram_cell[   23688] = 32'hadeee78b;
    ram_cell[   23689] = 32'hbeef81a2;
    ram_cell[   23690] = 32'h37b161c8;
    ram_cell[   23691] = 32'hc6571275;
    ram_cell[   23692] = 32'hba34a0cd;
    ram_cell[   23693] = 32'h1f98a49c;
    ram_cell[   23694] = 32'hf7a136c0;
    ram_cell[   23695] = 32'h31623454;
    ram_cell[   23696] = 32'hdb459abf;
    ram_cell[   23697] = 32'he18fa987;
    ram_cell[   23698] = 32'hc4afa6ec;
    ram_cell[   23699] = 32'h3b984ca5;
    ram_cell[   23700] = 32'h89c57754;
    ram_cell[   23701] = 32'h56256078;
    ram_cell[   23702] = 32'h068bff62;
    ram_cell[   23703] = 32'hf88da6ee;
    ram_cell[   23704] = 32'h3392972a;
    ram_cell[   23705] = 32'ha718a6bb;
    ram_cell[   23706] = 32'hda68bd0c;
    ram_cell[   23707] = 32'hface69be;
    ram_cell[   23708] = 32'h624913db;
    ram_cell[   23709] = 32'h3afbbea9;
    ram_cell[   23710] = 32'h579011ca;
    ram_cell[   23711] = 32'hb5238e5d;
    ram_cell[   23712] = 32'hd6cf21ec;
    ram_cell[   23713] = 32'h98b6c996;
    ram_cell[   23714] = 32'h7bfd2a19;
    ram_cell[   23715] = 32'hf23c5ecb;
    ram_cell[   23716] = 32'h146a529e;
    ram_cell[   23717] = 32'h1216550a;
    ram_cell[   23718] = 32'h71b02dca;
    ram_cell[   23719] = 32'h916790dd;
    ram_cell[   23720] = 32'hc6805bf2;
    ram_cell[   23721] = 32'h723ffe3c;
    ram_cell[   23722] = 32'h54592f66;
    ram_cell[   23723] = 32'hfdcfd972;
    ram_cell[   23724] = 32'h8307b389;
    ram_cell[   23725] = 32'h4bed61f7;
    ram_cell[   23726] = 32'hb297643a;
    ram_cell[   23727] = 32'he292a15c;
    ram_cell[   23728] = 32'he8cd6922;
    ram_cell[   23729] = 32'hfa3228d3;
    ram_cell[   23730] = 32'h974c7715;
    ram_cell[   23731] = 32'h1e1432a5;
    ram_cell[   23732] = 32'h1991aab1;
    ram_cell[   23733] = 32'h75ea8d71;
    ram_cell[   23734] = 32'he7ea6134;
    ram_cell[   23735] = 32'h6741936a;
    ram_cell[   23736] = 32'h93f7d9ce;
    ram_cell[   23737] = 32'h4ba15cda;
    ram_cell[   23738] = 32'hf9f90aed;
    ram_cell[   23739] = 32'hfc3ce2ed;
    ram_cell[   23740] = 32'h5cd1cb1c;
    ram_cell[   23741] = 32'hbd0da76d;
    ram_cell[   23742] = 32'h8812b785;
    ram_cell[   23743] = 32'h44d2ffd7;
    ram_cell[   23744] = 32'hd0044f40;
    ram_cell[   23745] = 32'hdf978d23;
    ram_cell[   23746] = 32'h9eb67c49;
    ram_cell[   23747] = 32'h5572bf73;
    ram_cell[   23748] = 32'h8746a3a3;
    ram_cell[   23749] = 32'h909d7764;
    ram_cell[   23750] = 32'ha94d42eb;
    ram_cell[   23751] = 32'h345c6927;
    ram_cell[   23752] = 32'h74974194;
    ram_cell[   23753] = 32'h78a42177;
    ram_cell[   23754] = 32'ha8c91e94;
    ram_cell[   23755] = 32'haffbba9a;
    ram_cell[   23756] = 32'h5c41195d;
    ram_cell[   23757] = 32'hdf2c58d6;
    ram_cell[   23758] = 32'h7e4294e7;
    ram_cell[   23759] = 32'hc39c1728;
    ram_cell[   23760] = 32'h39615916;
    ram_cell[   23761] = 32'h562a32b4;
    ram_cell[   23762] = 32'h072a1f74;
    ram_cell[   23763] = 32'h66f5659d;
    ram_cell[   23764] = 32'h6ab5e358;
    ram_cell[   23765] = 32'h1b10a31c;
    ram_cell[   23766] = 32'h826e166b;
    ram_cell[   23767] = 32'hea3deaad;
    ram_cell[   23768] = 32'hffc0500b;
    ram_cell[   23769] = 32'h1feb149d;
    ram_cell[   23770] = 32'hb9ad4b70;
    ram_cell[   23771] = 32'h91466b7e;
    ram_cell[   23772] = 32'hb3bc072e;
    ram_cell[   23773] = 32'h1f26bee9;
    ram_cell[   23774] = 32'h9b4495e2;
    ram_cell[   23775] = 32'h224a1b2c;
    ram_cell[   23776] = 32'hc6efadfd;
    ram_cell[   23777] = 32'h5a83844a;
    ram_cell[   23778] = 32'h5ea40de0;
    ram_cell[   23779] = 32'h5a1233ae;
    ram_cell[   23780] = 32'h489a5acd;
    ram_cell[   23781] = 32'h0be55981;
    ram_cell[   23782] = 32'h9deb1272;
    ram_cell[   23783] = 32'h2166d132;
    ram_cell[   23784] = 32'h3f93bcdf;
    ram_cell[   23785] = 32'hca1a3c59;
    ram_cell[   23786] = 32'h314cbbe9;
    ram_cell[   23787] = 32'hd0b309b8;
    ram_cell[   23788] = 32'he7115344;
    ram_cell[   23789] = 32'h6a53eaa6;
    ram_cell[   23790] = 32'he876c6ee;
    ram_cell[   23791] = 32'hbbb3545b;
    ram_cell[   23792] = 32'hc828d8b8;
    ram_cell[   23793] = 32'haa44be6e;
    ram_cell[   23794] = 32'hbe5ecbb5;
    ram_cell[   23795] = 32'hd326b162;
    ram_cell[   23796] = 32'h14c6c7c1;
    ram_cell[   23797] = 32'h451bc841;
    ram_cell[   23798] = 32'hcf504691;
    ram_cell[   23799] = 32'hd09fc04c;
    ram_cell[   23800] = 32'hde8d53c5;
    ram_cell[   23801] = 32'hf3e7e59a;
    ram_cell[   23802] = 32'hca143b48;
    ram_cell[   23803] = 32'hb301dfba;
    ram_cell[   23804] = 32'h592a81ba;
    ram_cell[   23805] = 32'ha30c73e3;
    ram_cell[   23806] = 32'h033fadfd;
    ram_cell[   23807] = 32'h2ed235d7;
    ram_cell[   23808] = 32'h4f886fa8;
    ram_cell[   23809] = 32'hf6000a1e;
    ram_cell[   23810] = 32'hbcdca263;
    ram_cell[   23811] = 32'ha6ce073a;
    ram_cell[   23812] = 32'h625a073b;
    ram_cell[   23813] = 32'h7c9975a4;
    ram_cell[   23814] = 32'h3aacf891;
    ram_cell[   23815] = 32'h5d8e5e9c;
    ram_cell[   23816] = 32'h3cad9017;
    ram_cell[   23817] = 32'hb52d7021;
    ram_cell[   23818] = 32'ha40481c7;
    ram_cell[   23819] = 32'he69a774d;
    ram_cell[   23820] = 32'h19e353ef;
    ram_cell[   23821] = 32'hc7efc219;
    ram_cell[   23822] = 32'hd69fbfff;
    ram_cell[   23823] = 32'hc2cf3dfb;
    ram_cell[   23824] = 32'ha22bf9a4;
    ram_cell[   23825] = 32'h5e300406;
    ram_cell[   23826] = 32'h3c155844;
    ram_cell[   23827] = 32'h85b75593;
    ram_cell[   23828] = 32'hb657bdd7;
    ram_cell[   23829] = 32'h465bcc73;
    ram_cell[   23830] = 32'h0919680e;
    ram_cell[   23831] = 32'h2de3db46;
    ram_cell[   23832] = 32'hce896c88;
    ram_cell[   23833] = 32'h45f8bd7d;
    ram_cell[   23834] = 32'hc3ba19ef;
    ram_cell[   23835] = 32'h4d2ee2a7;
    ram_cell[   23836] = 32'h4cecaad7;
    ram_cell[   23837] = 32'hfca526ea;
    ram_cell[   23838] = 32'h3b02c37c;
    ram_cell[   23839] = 32'h9df3c2a0;
    ram_cell[   23840] = 32'h92f5e787;
    ram_cell[   23841] = 32'hc9fbde06;
    ram_cell[   23842] = 32'hc0e5ec43;
    ram_cell[   23843] = 32'h1d0e76df;
    ram_cell[   23844] = 32'h9ad99a8b;
    ram_cell[   23845] = 32'h5add42b5;
    ram_cell[   23846] = 32'h99289116;
    ram_cell[   23847] = 32'h5df91579;
    ram_cell[   23848] = 32'h812a9ebe;
    ram_cell[   23849] = 32'hecb56791;
    ram_cell[   23850] = 32'h53d68072;
    ram_cell[   23851] = 32'h91b46274;
    ram_cell[   23852] = 32'ha7c61c3b;
    ram_cell[   23853] = 32'h8d3d8f9c;
    ram_cell[   23854] = 32'hc41dc15f;
    ram_cell[   23855] = 32'hfcf5e34a;
    ram_cell[   23856] = 32'h5112726f;
    ram_cell[   23857] = 32'hacb2673d;
    ram_cell[   23858] = 32'h2ce5e9d9;
    ram_cell[   23859] = 32'h5fe67f19;
    ram_cell[   23860] = 32'h180a1865;
    ram_cell[   23861] = 32'hfd121815;
    ram_cell[   23862] = 32'hcc15429d;
    ram_cell[   23863] = 32'h80e36b83;
    ram_cell[   23864] = 32'h438b66ad;
    ram_cell[   23865] = 32'h865451f6;
    ram_cell[   23866] = 32'hcb8cd138;
    ram_cell[   23867] = 32'h52738812;
    ram_cell[   23868] = 32'h28c5f11c;
    ram_cell[   23869] = 32'h32deeb51;
    ram_cell[   23870] = 32'hc1842c68;
    ram_cell[   23871] = 32'h061742be;
    ram_cell[   23872] = 32'h83b43484;
    ram_cell[   23873] = 32'h68f63854;
    ram_cell[   23874] = 32'h9ff42082;
    ram_cell[   23875] = 32'h1823d48a;
    ram_cell[   23876] = 32'h51c53b57;
    ram_cell[   23877] = 32'hffbaaf9f;
    ram_cell[   23878] = 32'h2bbf6811;
    ram_cell[   23879] = 32'hcc4150f6;
    ram_cell[   23880] = 32'h65397685;
    ram_cell[   23881] = 32'ha9429809;
    ram_cell[   23882] = 32'hc21c739d;
    ram_cell[   23883] = 32'h5d9e4111;
    ram_cell[   23884] = 32'hf99870ba;
    ram_cell[   23885] = 32'h86cd81e6;
    ram_cell[   23886] = 32'h049a2a3c;
    ram_cell[   23887] = 32'h0f963910;
    ram_cell[   23888] = 32'hb8f87e68;
    ram_cell[   23889] = 32'hb781dd7e;
    ram_cell[   23890] = 32'h0ef7ae20;
    ram_cell[   23891] = 32'hca95721b;
    ram_cell[   23892] = 32'h8fef3954;
    ram_cell[   23893] = 32'hf1acb7ac;
    ram_cell[   23894] = 32'h6d5e19ef;
    ram_cell[   23895] = 32'he2ffbf4c;
    ram_cell[   23896] = 32'hb44a7e97;
    ram_cell[   23897] = 32'hab37ef8d;
    ram_cell[   23898] = 32'h8de7b487;
    ram_cell[   23899] = 32'hf684aa84;
    ram_cell[   23900] = 32'hfdf95551;
    ram_cell[   23901] = 32'h77a728a1;
    ram_cell[   23902] = 32'hfcceb93d;
    ram_cell[   23903] = 32'hc109edea;
    ram_cell[   23904] = 32'h939d5090;
    ram_cell[   23905] = 32'h5ae69329;
    ram_cell[   23906] = 32'h89031072;
    ram_cell[   23907] = 32'h80014221;
    ram_cell[   23908] = 32'h4f01accf;
    ram_cell[   23909] = 32'h2b429997;
    ram_cell[   23910] = 32'h418407c7;
    ram_cell[   23911] = 32'hb9a0b12d;
    ram_cell[   23912] = 32'h40362a39;
    ram_cell[   23913] = 32'hd0ae11b2;
    ram_cell[   23914] = 32'hfefdfa50;
    ram_cell[   23915] = 32'h709493f6;
    ram_cell[   23916] = 32'h2b1605ac;
    ram_cell[   23917] = 32'hb67f2ad3;
    ram_cell[   23918] = 32'hdd734da4;
    ram_cell[   23919] = 32'hd681d7de;
    ram_cell[   23920] = 32'hb67717df;
    ram_cell[   23921] = 32'h9aad1e46;
    ram_cell[   23922] = 32'h17b155b0;
    ram_cell[   23923] = 32'hf50dc11b;
    ram_cell[   23924] = 32'hf241cf90;
    ram_cell[   23925] = 32'h74c54e5d;
    ram_cell[   23926] = 32'he71a1a13;
    ram_cell[   23927] = 32'h1f68bab6;
    ram_cell[   23928] = 32'h1de144c7;
    ram_cell[   23929] = 32'h13acb3c3;
    ram_cell[   23930] = 32'h5d2fec1a;
    ram_cell[   23931] = 32'h4182503e;
    ram_cell[   23932] = 32'hfb7f9b9b;
    ram_cell[   23933] = 32'h679526aa;
    ram_cell[   23934] = 32'hbdb4c579;
    ram_cell[   23935] = 32'hf2dd27d3;
    ram_cell[   23936] = 32'hdf41f994;
    ram_cell[   23937] = 32'h748e9a70;
    ram_cell[   23938] = 32'he6f2ad4a;
    ram_cell[   23939] = 32'h29fb562e;
    ram_cell[   23940] = 32'h7cf7fc6b;
    ram_cell[   23941] = 32'h213bc0fc;
    ram_cell[   23942] = 32'h15c54d70;
    ram_cell[   23943] = 32'ha685bc5f;
    ram_cell[   23944] = 32'hdc3ea1e2;
    ram_cell[   23945] = 32'h06fa16b8;
    ram_cell[   23946] = 32'h0e5beea1;
    ram_cell[   23947] = 32'hed087744;
    ram_cell[   23948] = 32'hfcf304f8;
    ram_cell[   23949] = 32'h3ab434db;
    ram_cell[   23950] = 32'hbdc5f263;
    ram_cell[   23951] = 32'hb6d93a3d;
    ram_cell[   23952] = 32'h838f20dc;
    ram_cell[   23953] = 32'h85a1387a;
    ram_cell[   23954] = 32'h1561c987;
    ram_cell[   23955] = 32'h42b1d61c;
    ram_cell[   23956] = 32'h0eaede3d;
    ram_cell[   23957] = 32'hb2bf047b;
    ram_cell[   23958] = 32'hc93f59b5;
    ram_cell[   23959] = 32'h88f32cb9;
    ram_cell[   23960] = 32'h3055db92;
    ram_cell[   23961] = 32'hfdb7ae7b;
    ram_cell[   23962] = 32'h9b4bd2ff;
    ram_cell[   23963] = 32'ha615c33a;
    ram_cell[   23964] = 32'h1b337860;
    ram_cell[   23965] = 32'hed246b29;
    ram_cell[   23966] = 32'h13e52d84;
    ram_cell[   23967] = 32'h7e39e63a;
    ram_cell[   23968] = 32'h131848ec;
    ram_cell[   23969] = 32'h8e8b64dc;
    ram_cell[   23970] = 32'h1d580f2e;
    ram_cell[   23971] = 32'h45e3d90a;
    ram_cell[   23972] = 32'h9a2abdf6;
    ram_cell[   23973] = 32'hf06ee739;
    ram_cell[   23974] = 32'hf8472c3c;
    ram_cell[   23975] = 32'h3d4c9c2b;
    ram_cell[   23976] = 32'ha962ca5b;
    ram_cell[   23977] = 32'h46d921ef;
    ram_cell[   23978] = 32'hdf508ef1;
    ram_cell[   23979] = 32'h87d86fbe;
    ram_cell[   23980] = 32'h396d14ea;
    ram_cell[   23981] = 32'hecfb5115;
    ram_cell[   23982] = 32'hc15490f2;
    ram_cell[   23983] = 32'h6e04c4c8;
    ram_cell[   23984] = 32'h6b21b8f4;
    ram_cell[   23985] = 32'h48fe4c86;
    ram_cell[   23986] = 32'h932811cc;
    ram_cell[   23987] = 32'h006dbd3f;
    ram_cell[   23988] = 32'ha02adf71;
    ram_cell[   23989] = 32'h109516a7;
    ram_cell[   23990] = 32'he3f95b06;
    ram_cell[   23991] = 32'h97c72f4b;
    ram_cell[   23992] = 32'hb33ae1b0;
    ram_cell[   23993] = 32'h07114b79;
    ram_cell[   23994] = 32'h91cc21bd;
    ram_cell[   23995] = 32'haa877e1d;
    ram_cell[   23996] = 32'h5cafbec6;
    ram_cell[   23997] = 32'h906608b6;
    ram_cell[   23998] = 32'hc29056c1;
    ram_cell[   23999] = 32'h4545facb;
    ram_cell[   24000] = 32'h69756c83;
    ram_cell[   24001] = 32'h9506389c;
    ram_cell[   24002] = 32'h2db8305c;
    ram_cell[   24003] = 32'h91048423;
    ram_cell[   24004] = 32'haf2c0e90;
    ram_cell[   24005] = 32'hfa4e7755;
    ram_cell[   24006] = 32'h65285e63;
    ram_cell[   24007] = 32'hf640dfd8;
    ram_cell[   24008] = 32'h13e00c96;
    ram_cell[   24009] = 32'h514e729e;
    ram_cell[   24010] = 32'haa189c31;
    ram_cell[   24011] = 32'h5c1308c1;
    ram_cell[   24012] = 32'hf258d47a;
    ram_cell[   24013] = 32'h255b4bc0;
    ram_cell[   24014] = 32'h67522a93;
    ram_cell[   24015] = 32'ha4a4e234;
    ram_cell[   24016] = 32'h5b9eeb33;
    ram_cell[   24017] = 32'h9b8f0b38;
    ram_cell[   24018] = 32'hb67d18af;
    ram_cell[   24019] = 32'h99e00e21;
    ram_cell[   24020] = 32'h6c411403;
    ram_cell[   24021] = 32'he15726a3;
    ram_cell[   24022] = 32'h8a7f7d5d;
    ram_cell[   24023] = 32'h3982d692;
    ram_cell[   24024] = 32'h94b2dd32;
    ram_cell[   24025] = 32'h81b26739;
    ram_cell[   24026] = 32'h25e83c9d;
    ram_cell[   24027] = 32'h4437a87b;
    ram_cell[   24028] = 32'h49a8ce5e;
    ram_cell[   24029] = 32'h089b49c7;
    ram_cell[   24030] = 32'ha1c8400a;
    ram_cell[   24031] = 32'hd9a81924;
    ram_cell[   24032] = 32'h78f9b38f;
    ram_cell[   24033] = 32'h734b15a8;
    ram_cell[   24034] = 32'h69bbccfc;
    ram_cell[   24035] = 32'h74ac073a;
    ram_cell[   24036] = 32'h3bc5ff14;
    ram_cell[   24037] = 32'haae9940b;
    ram_cell[   24038] = 32'he2deea25;
    ram_cell[   24039] = 32'h4d2c8ca3;
    ram_cell[   24040] = 32'h56ffbaa9;
    ram_cell[   24041] = 32'hc4f72c57;
    ram_cell[   24042] = 32'hd25c58a7;
    ram_cell[   24043] = 32'h7d49628b;
    ram_cell[   24044] = 32'h44000c9a;
    ram_cell[   24045] = 32'h2fb5c937;
    ram_cell[   24046] = 32'h9ba3cda3;
    ram_cell[   24047] = 32'h86ad9e8a;
    ram_cell[   24048] = 32'h7542c0f5;
    ram_cell[   24049] = 32'h4eef5be5;
    ram_cell[   24050] = 32'h8b88e795;
    ram_cell[   24051] = 32'hd58434d6;
    ram_cell[   24052] = 32'h129ffe39;
    ram_cell[   24053] = 32'hd248ccf1;
    ram_cell[   24054] = 32'h2575db82;
    ram_cell[   24055] = 32'h0a572d75;
    ram_cell[   24056] = 32'h50985ac5;
    ram_cell[   24057] = 32'hea0b3698;
    ram_cell[   24058] = 32'hb0691ddc;
    ram_cell[   24059] = 32'h85159d77;
    ram_cell[   24060] = 32'h08dcd207;
    ram_cell[   24061] = 32'hdf9e32cc;
    ram_cell[   24062] = 32'h9ecdd3cf;
    ram_cell[   24063] = 32'hb5a62115;
    ram_cell[   24064] = 32'h0f13b18d;
    ram_cell[   24065] = 32'heab5bd65;
    ram_cell[   24066] = 32'h666c8af8;
    ram_cell[   24067] = 32'hbfe1c547;
    ram_cell[   24068] = 32'hd5b59e41;
    ram_cell[   24069] = 32'h0e530bb3;
    ram_cell[   24070] = 32'h1a7c05d2;
    ram_cell[   24071] = 32'hcc01f1e3;
    ram_cell[   24072] = 32'h4528b331;
    ram_cell[   24073] = 32'h058ff6a6;
    ram_cell[   24074] = 32'hff35f334;
    ram_cell[   24075] = 32'h74fe4b3a;
    ram_cell[   24076] = 32'h15ddaf90;
    ram_cell[   24077] = 32'hb1c3556c;
    ram_cell[   24078] = 32'h07f648e4;
    ram_cell[   24079] = 32'h3aff3a21;
    ram_cell[   24080] = 32'h273680e8;
    ram_cell[   24081] = 32'h5fa95451;
    ram_cell[   24082] = 32'h31080c9f;
    ram_cell[   24083] = 32'h4fa396b3;
    ram_cell[   24084] = 32'h3b147940;
    ram_cell[   24085] = 32'h4b2f5a9a;
    ram_cell[   24086] = 32'h6015542e;
    ram_cell[   24087] = 32'hdd2624a8;
    ram_cell[   24088] = 32'hc6f5aa09;
    ram_cell[   24089] = 32'h65f28abf;
    ram_cell[   24090] = 32'h7fd5f9df;
    ram_cell[   24091] = 32'h29a3f11d;
    ram_cell[   24092] = 32'h09b34483;
    ram_cell[   24093] = 32'h3b4c1808;
    ram_cell[   24094] = 32'hf2445128;
    ram_cell[   24095] = 32'ha3b51886;
    ram_cell[   24096] = 32'h1cba0e43;
    ram_cell[   24097] = 32'hf873ce23;
    ram_cell[   24098] = 32'hf7a0cebe;
    ram_cell[   24099] = 32'h7ae66fce;
    ram_cell[   24100] = 32'hbdd2cd06;
    ram_cell[   24101] = 32'he5544c9e;
    ram_cell[   24102] = 32'hfcbbea70;
    ram_cell[   24103] = 32'hfe65ac83;
    ram_cell[   24104] = 32'h1cd4fe0b;
    ram_cell[   24105] = 32'had903db5;
    ram_cell[   24106] = 32'h11a22808;
    ram_cell[   24107] = 32'h688a948a;
    ram_cell[   24108] = 32'h553f7320;
    ram_cell[   24109] = 32'h30024908;
    ram_cell[   24110] = 32'h4c9a6009;
    ram_cell[   24111] = 32'h5ce92056;
    ram_cell[   24112] = 32'hb3148e8e;
    ram_cell[   24113] = 32'ha42ddcc6;
    ram_cell[   24114] = 32'h5154a34c;
    ram_cell[   24115] = 32'h3557a1b9;
    ram_cell[   24116] = 32'hd1554df4;
    ram_cell[   24117] = 32'h6c9252b8;
    ram_cell[   24118] = 32'h1adc7b1e;
    ram_cell[   24119] = 32'h863f0d86;
    ram_cell[   24120] = 32'h93bb3369;
    ram_cell[   24121] = 32'h8ac13213;
    ram_cell[   24122] = 32'hcc75fdab;
    ram_cell[   24123] = 32'h620baddd;
    ram_cell[   24124] = 32'h9baa9e58;
    ram_cell[   24125] = 32'h5b1decdd;
    ram_cell[   24126] = 32'h5309239f;
    ram_cell[   24127] = 32'hdc8dd006;
    ram_cell[   24128] = 32'h6929f378;
    ram_cell[   24129] = 32'heda07780;
    ram_cell[   24130] = 32'h4a8ff515;
    ram_cell[   24131] = 32'hfc4d2c67;
    ram_cell[   24132] = 32'h635361b8;
    ram_cell[   24133] = 32'h5a943707;
    ram_cell[   24134] = 32'h2bd7ec08;
    ram_cell[   24135] = 32'h646f1141;
    ram_cell[   24136] = 32'h8f56b100;
    ram_cell[   24137] = 32'h4ba1bc08;
    ram_cell[   24138] = 32'h727b12aa;
    ram_cell[   24139] = 32'h60cf99e4;
    ram_cell[   24140] = 32'hff1ecb0d;
    ram_cell[   24141] = 32'hba4e545d;
    ram_cell[   24142] = 32'h902f71f3;
    ram_cell[   24143] = 32'h5cd31ccf;
    ram_cell[   24144] = 32'h27758c90;
    ram_cell[   24145] = 32'hea5e5e61;
    ram_cell[   24146] = 32'habe825fd;
    ram_cell[   24147] = 32'h0b24f0f1;
    ram_cell[   24148] = 32'h8142014e;
    ram_cell[   24149] = 32'h9eaf04fe;
    ram_cell[   24150] = 32'h1d2d47a3;
    ram_cell[   24151] = 32'ha211a9ac;
    ram_cell[   24152] = 32'h80803686;
    ram_cell[   24153] = 32'hf35cb0be;
    ram_cell[   24154] = 32'h624aff7c;
    ram_cell[   24155] = 32'h1c8dae72;
    ram_cell[   24156] = 32'hd432c600;
    ram_cell[   24157] = 32'h67c1545d;
    ram_cell[   24158] = 32'h9ff386df;
    ram_cell[   24159] = 32'h9d8ec5b9;
    ram_cell[   24160] = 32'h6ed22d6e;
    ram_cell[   24161] = 32'h6a71fedf;
    ram_cell[   24162] = 32'h83f70b3b;
    ram_cell[   24163] = 32'hc99925ae;
    ram_cell[   24164] = 32'ha152571f;
    ram_cell[   24165] = 32'h2bc4aa97;
    ram_cell[   24166] = 32'hfa36000d;
    ram_cell[   24167] = 32'h242dade3;
    ram_cell[   24168] = 32'h84642508;
    ram_cell[   24169] = 32'h6fe2a1bc;
    ram_cell[   24170] = 32'h261d8e06;
    ram_cell[   24171] = 32'h97e2caf8;
    ram_cell[   24172] = 32'h3c66a2ca;
    ram_cell[   24173] = 32'hf25fe9ad;
    ram_cell[   24174] = 32'habb7ec34;
    ram_cell[   24175] = 32'h8ada663b;
    ram_cell[   24176] = 32'h77c38a80;
    ram_cell[   24177] = 32'h70eb1d32;
    ram_cell[   24178] = 32'h89af2cd9;
    ram_cell[   24179] = 32'he5180175;
    ram_cell[   24180] = 32'hc0a8c462;
    ram_cell[   24181] = 32'h07d42aa0;
    ram_cell[   24182] = 32'h9430ab6c;
    ram_cell[   24183] = 32'h1fd29fb6;
    ram_cell[   24184] = 32'hb91aeaa7;
    ram_cell[   24185] = 32'ha9e500fe;
    ram_cell[   24186] = 32'h5039d893;
    ram_cell[   24187] = 32'h75ee8a5e;
    ram_cell[   24188] = 32'h017a84e6;
    ram_cell[   24189] = 32'hf43ab05a;
    ram_cell[   24190] = 32'hff7128ef;
    ram_cell[   24191] = 32'haddc7c65;
    ram_cell[   24192] = 32'h0987c8e5;
    ram_cell[   24193] = 32'he3f74b84;
    ram_cell[   24194] = 32'ha98a9494;
    ram_cell[   24195] = 32'h4b29b89a;
    ram_cell[   24196] = 32'h6e053bf4;
    ram_cell[   24197] = 32'hcd63211a;
    ram_cell[   24198] = 32'hc886ad3e;
    ram_cell[   24199] = 32'hb245b3e1;
    ram_cell[   24200] = 32'h0af0d868;
    ram_cell[   24201] = 32'ha84e6edf;
    ram_cell[   24202] = 32'hbc43eb33;
    ram_cell[   24203] = 32'hc5bd418f;
    ram_cell[   24204] = 32'h33ee44a1;
    ram_cell[   24205] = 32'hfaa70d68;
    ram_cell[   24206] = 32'hf3a268a1;
    ram_cell[   24207] = 32'hcec58c4f;
    ram_cell[   24208] = 32'hb0aaddab;
    ram_cell[   24209] = 32'hf7f4e9a9;
    ram_cell[   24210] = 32'h75e59b66;
    ram_cell[   24211] = 32'h0439e893;
    ram_cell[   24212] = 32'h07e3614f;
    ram_cell[   24213] = 32'h4cb02ebb;
    ram_cell[   24214] = 32'h38e01271;
    ram_cell[   24215] = 32'he74106fe;
    ram_cell[   24216] = 32'hae57afc2;
    ram_cell[   24217] = 32'hea2a334e;
    ram_cell[   24218] = 32'h0086ee8d;
    ram_cell[   24219] = 32'hfee89ec8;
    ram_cell[   24220] = 32'h4c250369;
    ram_cell[   24221] = 32'h98d4a25c;
    ram_cell[   24222] = 32'h01effb30;
    ram_cell[   24223] = 32'h3aab1aa7;
    ram_cell[   24224] = 32'hd4a0fc32;
    ram_cell[   24225] = 32'hbdf86194;
    ram_cell[   24226] = 32'ha2611a27;
    ram_cell[   24227] = 32'h5cc33c8f;
    ram_cell[   24228] = 32'h037192f0;
    ram_cell[   24229] = 32'h82aa6c86;
    ram_cell[   24230] = 32'h0bc42e81;
    ram_cell[   24231] = 32'hd9001fee;
    ram_cell[   24232] = 32'h28ce1262;
    ram_cell[   24233] = 32'h18760966;
    ram_cell[   24234] = 32'ha33357f2;
    ram_cell[   24235] = 32'h36a51928;
    ram_cell[   24236] = 32'h2919f565;
    ram_cell[   24237] = 32'h33111c23;
    ram_cell[   24238] = 32'h2d94c90d;
    ram_cell[   24239] = 32'h7ae66e26;
    ram_cell[   24240] = 32'h14f7465a;
    ram_cell[   24241] = 32'ha9bd5424;
    ram_cell[   24242] = 32'h5099cc87;
    ram_cell[   24243] = 32'h370730f9;
    ram_cell[   24244] = 32'h77d61ec7;
    ram_cell[   24245] = 32'h0ac52b35;
    ram_cell[   24246] = 32'h6d1d170a;
    ram_cell[   24247] = 32'h538192db;
    ram_cell[   24248] = 32'hfd9af19b;
    ram_cell[   24249] = 32'h7fc0a912;
    ram_cell[   24250] = 32'h6ff74ba3;
    ram_cell[   24251] = 32'h555a022f;
    ram_cell[   24252] = 32'h31c8a9ca;
    ram_cell[   24253] = 32'h170135f5;
    ram_cell[   24254] = 32'h07e7f2ef;
    ram_cell[   24255] = 32'hd5e64856;
    ram_cell[   24256] = 32'hbc61f725;
    ram_cell[   24257] = 32'h111e4159;
    ram_cell[   24258] = 32'h9ab20ec0;
    ram_cell[   24259] = 32'h480bf58e;
    ram_cell[   24260] = 32'hd441bebc;
    ram_cell[   24261] = 32'hf2fe34d9;
    ram_cell[   24262] = 32'h60689420;
    ram_cell[   24263] = 32'h7086dde0;
    ram_cell[   24264] = 32'hb87cb87b;
    ram_cell[   24265] = 32'h69111556;
    ram_cell[   24266] = 32'hadfeab43;
    ram_cell[   24267] = 32'h88180408;
    ram_cell[   24268] = 32'h49d8c606;
    ram_cell[   24269] = 32'hd6d0813e;
    ram_cell[   24270] = 32'hd95dc8d4;
    ram_cell[   24271] = 32'h79eea2e8;
    ram_cell[   24272] = 32'h7b027b73;
    ram_cell[   24273] = 32'h487fd201;
    ram_cell[   24274] = 32'h029d83da;
    ram_cell[   24275] = 32'h41df947c;
    ram_cell[   24276] = 32'h8e1d1649;
    ram_cell[   24277] = 32'h2f2a944b;
    ram_cell[   24278] = 32'h607eb011;
    ram_cell[   24279] = 32'h8de5c06f;
    ram_cell[   24280] = 32'h0bb1bb6a;
    ram_cell[   24281] = 32'hfba38705;
    ram_cell[   24282] = 32'h187bb709;
    ram_cell[   24283] = 32'hdec0d252;
    ram_cell[   24284] = 32'h73fd3820;
    ram_cell[   24285] = 32'h4aeaccc3;
    ram_cell[   24286] = 32'hcd0a8b51;
    ram_cell[   24287] = 32'ha3531b65;
    ram_cell[   24288] = 32'h4333c086;
    ram_cell[   24289] = 32'h8eb45ba7;
    ram_cell[   24290] = 32'h91bf8945;
    ram_cell[   24291] = 32'h5b865c42;
    ram_cell[   24292] = 32'h05f09226;
    ram_cell[   24293] = 32'he2966387;
    ram_cell[   24294] = 32'ha21701e0;
    ram_cell[   24295] = 32'hc6a1eb9e;
    ram_cell[   24296] = 32'h4c0c91a4;
    ram_cell[   24297] = 32'hd4f731a9;
    ram_cell[   24298] = 32'h6641cd18;
    ram_cell[   24299] = 32'h9126c22d;
    ram_cell[   24300] = 32'h48016fa8;
    ram_cell[   24301] = 32'h40fb3af8;
    ram_cell[   24302] = 32'hd618b79b;
    ram_cell[   24303] = 32'hee42c889;
    ram_cell[   24304] = 32'h7c898b5a;
    ram_cell[   24305] = 32'hbbaed1cd;
    ram_cell[   24306] = 32'hb379d30c;
    ram_cell[   24307] = 32'h85a9a30d;
    ram_cell[   24308] = 32'h1a3c9441;
    ram_cell[   24309] = 32'hc0c87e9b;
    ram_cell[   24310] = 32'h412fc74f;
    ram_cell[   24311] = 32'h2be5baa7;
    ram_cell[   24312] = 32'h5dc7f34d;
    ram_cell[   24313] = 32'h375d9960;
    ram_cell[   24314] = 32'h72185624;
    ram_cell[   24315] = 32'h7ce713ad;
    ram_cell[   24316] = 32'ha8310eb5;
    ram_cell[   24317] = 32'ha844d633;
    ram_cell[   24318] = 32'h42560b12;
    ram_cell[   24319] = 32'hb575aa75;
    ram_cell[   24320] = 32'h7f797217;
    ram_cell[   24321] = 32'hfce1ee2e;
    ram_cell[   24322] = 32'h594d18f0;
    ram_cell[   24323] = 32'h8e075134;
    ram_cell[   24324] = 32'hf5c1e447;
    ram_cell[   24325] = 32'h539a077b;
    ram_cell[   24326] = 32'h119ae5d9;
    ram_cell[   24327] = 32'he249b356;
    ram_cell[   24328] = 32'h78f7a0c4;
    ram_cell[   24329] = 32'h814149da;
    ram_cell[   24330] = 32'h86940368;
    ram_cell[   24331] = 32'h623e8972;
    ram_cell[   24332] = 32'h71b5cb87;
    ram_cell[   24333] = 32'h79de35c5;
    ram_cell[   24334] = 32'hb21b215d;
    ram_cell[   24335] = 32'h655aa08c;
    ram_cell[   24336] = 32'hd305279f;
    ram_cell[   24337] = 32'h7ab823b9;
    ram_cell[   24338] = 32'h22e96b60;
    ram_cell[   24339] = 32'h36266681;
    ram_cell[   24340] = 32'h4c7b005b;
    ram_cell[   24341] = 32'hf9708eb2;
    ram_cell[   24342] = 32'h510ab628;
    ram_cell[   24343] = 32'hbb36d6cf;
    ram_cell[   24344] = 32'hb981d369;
    ram_cell[   24345] = 32'h993678d0;
    ram_cell[   24346] = 32'h5095b89a;
    ram_cell[   24347] = 32'hef05d13e;
    ram_cell[   24348] = 32'hec33f7a2;
    ram_cell[   24349] = 32'h8a127b08;
    ram_cell[   24350] = 32'h004a324a;
    ram_cell[   24351] = 32'h0789eb36;
    ram_cell[   24352] = 32'h2c4d6ddf;
    ram_cell[   24353] = 32'h0818eece;
    ram_cell[   24354] = 32'h4d49a9df;
    ram_cell[   24355] = 32'h19d964ac;
    ram_cell[   24356] = 32'he03c0f36;
    ram_cell[   24357] = 32'hebaef238;
    ram_cell[   24358] = 32'h099a5541;
    ram_cell[   24359] = 32'hd5226eff;
    ram_cell[   24360] = 32'h36878427;
    ram_cell[   24361] = 32'ha7ef4008;
    ram_cell[   24362] = 32'h88c22b1e;
    ram_cell[   24363] = 32'h2a8def87;
    ram_cell[   24364] = 32'h40ef12a0;
    ram_cell[   24365] = 32'h438f9442;
    ram_cell[   24366] = 32'h31fef427;
    ram_cell[   24367] = 32'hb56b1773;
    ram_cell[   24368] = 32'hed896a42;
    ram_cell[   24369] = 32'h5d425802;
    ram_cell[   24370] = 32'hb313b426;
    ram_cell[   24371] = 32'h9453bca3;
    ram_cell[   24372] = 32'h59bd098d;
    ram_cell[   24373] = 32'h1dcc33f9;
    ram_cell[   24374] = 32'h73bb7d19;
    ram_cell[   24375] = 32'h8cf7df50;
    ram_cell[   24376] = 32'hfddc0457;
    ram_cell[   24377] = 32'h07f47193;
    ram_cell[   24378] = 32'h6caa32b7;
    ram_cell[   24379] = 32'hbd452a33;
    ram_cell[   24380] = 32'h116e3032;
    ram_cell[   24381] = 32'h484d723c;
    ram_cell[   24382] = 32'h9c983a2e;
    ram_cell[   24383] = 32'h5b98faa7;
    ram_cell[   24384] = 32'hbc910447;
    ram_cell[   24385] = 32'hf63b2215;
    ram_cell[   24386] = 32'h3b0b25bc;
    ram_cell[   24387] = 32'h02a36cbc;
    ram_cell[   24388] = 32'hcdc2cab5;
    ram_cell[   24389] = 32'hb2ac30a4;
    ram_cell[   24390] = 32'hfe4df3b1;
    ram_cell[   24391] = 32'h8a185520;
    ram_cell[   24392] = 32'h109294e9;
    ram_cell[   24393] = 32'hfd5cc39c;
    ram_cell[   24394] = 32'hd27f37c7;
    ram_cell[   24395] = 32'h1d7be080;
    ram_cell[   24396] = 32'ha8a6b40e;
    ram_cell[   24397] = 32'hbe10b626;
    ram_cell[   24398] = 32'h73184168;
    ram_cell[   24399] = 32'h5226d260;
    ram_cell[   24400] = 32'h731cef2e;
    ram_cell[   24401] = 32'h29127468;
    ram_cell[   24402] = 32'h3ed635eb;
    ram_cell[   24403] = 32'ha61cd024;
    ram_cell[   24404] = 32'h975beb89;
    ram_cell[   24405] = 32'h94a46d11;
    ram_cell[   24406] = 32'h42ae0029;
    ram_cell[   24407] = 32'h5ca9f205;
    ram_cell[   24408] = 32'h50ce57e8;
    ram_cell[   24409] = 32'hd8d6f89d;
    ram_cell[   24410] = 32'h4c282316;
    ram_cell[   24411] = 32'h4073ef78;
    ram_cell[   24412] = 32'ha8c57f6d;
    ram_cell[   24413] = 32'hf0deb14a;
    ram_cell[   24414] = 32'ha7dd68ab;
    ram_cell[   24415] = 32'hc767cfef;
    ram_cell[   24416] = 32'h246734d8;
    ram_cell[   24417] = 32'h9a3fab1d;
    ram_cell[   24418] = 32'h606ef248;
    ram_cell[   24419] = 32'hf5a36ac3;
    ram_cell[   24420] = 32'h7efd0ff9;
    ram_cell[   24421] = 32'h121d5355;
    ram_cell[   24422] = 32'h22340531;
    ram_cell[   24423] = 32'h16d31fa0;
    ram_cell[   24424] = 32'h3b13365d;
    ram_cell[   24425] = 32'hb3eaeb36;
    ram_cell[   24426] = 32'he66cee45;
    ram_cell[   24427] = 32'h4f519651;
    ram_cell[   24428] = 32'h3e22f027;
    ram_cell[   24429] = 32'h2bf83be3;
    ram_cell[   24430] = 32'h1628eb15;
    ram_cell[   24431] = 32'hc9eb0e47;
    ram_cell[   24432] = 32'h90b6afef;
    ram_cell[   24433] = 32'h7b774fa5;
    ram_cell[   24434] = 32'h00f313d8;
    ram_cell[   24435] = 32'h23bada8c;
    ram_cell[   24436] = 32'h45092b3d;
    ram_cell[   24437] = 32'h976572bc;
    ram_cell[   24438] = 32'hcac3a163;
    ram_cell[   24439] = 32'he212e03c;
    ram_cell[   24440] = 32'h5e44d89a;
    ram_cell[   24441] = 32'h0deb7cc0;
    ram_cell[   24442] = 32'hd3bcb4d2;
    ram_cell[   24443] = 32'h4c0d9859;
    ram_cell[   24444] = 32'hd10b5154;
    ram_cell[   24445] = 32'h87e95136;
    ram_cell[   24446] = 32'h0bd4bc2c;
    ram_cell[   24447] = 32'hb7fdc839;
    ram_cell[   24448] = 32'hdb806af7;
    ram_cell[   24449] = 32'h04f88970;
    ram_cell[   24450] = 32'h50995e51;
    ram_cell[   24451] = 32'h5bbe695a;
    ram_cell[   24452] = 32'h80f1be30;
    ram_cell[   24453] = 32'he9587522;
    ram_cell[   24454] = 32'h2471d615;
    ram_cell[   24455] = 32'h9cccc9b9;
    ram_cell[   24456] = 32'h31beef62;
    ram_cell[   24457] = 32'h5b0d2e99;
    ram_cell[   24458] = 32'ha1159f49;
    ram_cell[   24459] = 32'h149a28ef;
    ram_cell[   24460] = 32'h6b49ae0e;
    ram_cell[   24461] = 32'ha7a916a8;
    ram_cell[   24462] = 32'hf8ae71e0;
    ram_cell[   24463] = 32'h26b7aa50;
    ram_cell[   24464] = 32'h16369fa8;
    ram_cell[   24465] = 32'h27cb37cc;
    ram_cell[   24466] = 32'hfec6a01f;
    ram_cell[   24467] = 32'hf9eeba75;
    ram_cell[   24468] = 32'hf7d7ea91;
    ram_cell[   24469] = 32'h4a72a215;
    ram_cell[   24470] = 32'h97776e78;
    ram_cell[   24471] = 32'h6c6d1ccd;
    ram_cell[   24472] = 32'h12a00941;
    ram_cell[   24473] = 32'h1b436103;
    ram_cell[   24474] = 32'h95340257;
    ram_cell[   24475] = 32'haa48b11d;
    ram_cell[   24476] = 32'h9f50d0bf;
    ram_cell[   24477] = 32'hcf80e39c;
    ram_cell[   24478] = 32'hbff7739d;
    ram_cell[   24479] = 32'h3e2ca88b;
    ram_cell[   24480] = 32'h2417206c;
    ram_cell[   24481] = 32'hba4c91ac;
    ram_cell[   24482] = 32'h6ecbd683;
    ram_cell[   24483] = 32'h4c393edc;
    ram_cell[   24484] = 32'h9592c026;
    ram_cell[   24485] = 32'he6aee81f;
    ram_cell[   24486] = 32'hd955af14;
    ram_cell[   24487] = 32'h9529cf86;
    ram_cell[   24488] = 32'hcefe40a7;
    ram_cell[   24489] = 32'h5ecbdbfa;
    ram_cell[   24490] = 32'hc5f661d1;
    ram_cell[   24491] = 32'h6fe94af2;
    ram_cell[   24492] = 32'he150fb6e;
    ram_cell[   24493] = 32'hd32dcedd;
    ram_cell[   24494] = 32'h97b99978;
    ram_cell[   24495] = 32'h6edfa897;
    ram_cell[   24496] = 32'h36b62635;
    ram_cell[   24497] = 32'h6b3ba7bb;
    ram_cell[   24498] = 32'h0b984140;
    ram_cell[   24499] = 32'hd851cb5b;
    ram_cell[   24500] = 32'hfc40e529;
    ram_cell[   24501] = 32'hd4144eda;
    ram_cell[   24502] = 32'h41862caf;
    ram_cell[   24503] = 32'h6dc98d3a;
    ram_cell[   24504] = 32'hfaaebc84;
    ram_cell[   24505] = 32'habc48a8b;
    ram_cell[   24506] = 32'h0ca162c5;
    ram_cell[   24507] = 32'h7a5436d0;
    ram_cell[   24508] = 32'hd9b96709;
    ram_cell[   24509] = 32'hea979d7f;
    ram_cell[   24510] = 32'he306c66e;
    ram_cell[   24511] = 32'h6b98d70c;
    ram_cell[   24512] = 32'h2b1c64db;
    ram_cell[   24513] = 32'he802593a;
    ram_cell[   24514] = 32'he2f2dfdc;
    ram_cell[   24515] = 32'hd5979774;
    ram_cell[   24516] = 32'hd2af5254;
    ram_cell[   24517] = 32'h7d8bb847;
    ram_cell[   24518] = 32'h5fc3ff2d;
    ram_cell[   24519] = 32'hce3fe54e;
    ram_cell[   24520] = 32'h8160ab71;
    ram_cell[   24521] = 32'h12c633ab;
    ram_cell[   24522] = 32'h6d7e52aa;
    ram_cell[   24523] = 32'hc0058371;
    ram_cell[   24524] = 32'hb79eba9b;
    ram_cell[   24525] = 32'h95e6039c;
    ram_cell[   24526] = 32'h33bbceb1;
    ram_cell[   24527] = 32'h7c765743;
    ram_cell[   24528] = 32'hbc4bd163;
    ram_cell[   24529] = 32'hd2196b3e;
    ram_cell[   24530] = 32'h9d777347;
    ram_cell[   24531] = 32'hfdf3c299;
    ram_cell[   24532] = 32'hdf4e14be;
    ram_cell[   24533] = 32'h2fcc4939;
    ram_cell[   24534] = 32'h34485e48;
    ram_cell[   24535] = 32'h4e51c7a3;
    ram_cell[   24536] = 32'hfb6e95c3;
    ram_cell[   24537] = 32'ha0b40e39;
    ram_cell[   24538] = 32'hb0a7c343;
    ram_cell[   24539] = 32'h2cca937b;
    ram_cell[   24540] = 32'hdbb56754;
    ram_cell[   24541] = 32'hfe5eee7b;
    ram_cell[   24542] = 32'h58008dc6;
    ram_cell[   24543] = 32'hea39ed0d;
    ram_cell[   24544] = 32'h3e6bddc4;
    ram_cell[   24545] = 32'h063b46ce;
    ram_cell[   24546] = 32'hb9ac5f76;
    ram_cell[   24547] = 32'h4dcc096f;
    ram_cell[   24548] = 32'h98bc02d9;
    ram_cell[   24549] = 32'ha31e6540;
    ram_cell[   24550] = 32'he28d3e2c;
    ram_cell[   24551] = 32'h24b157b3;
    ram_cell[   24552] = 32'h007209e4;
    ram_cell[   24553] = 32'hedc5f2b1;
    ram_cell[   24554] = 32'hf5237626;
    ram_cell[   24555] = 32'h75554970;
    ram_cell[   24556] = 32'h0db831d5;
    ram_cell[   24557] = 32'h10b15666;
    ram_cell[   24558] = 32'h83c616b7;
    ram_cell[   24559] = 32'h901a88d0;
    ram_cell[   24560] = 32'h0445eba8;
    ram_cell[   24561] = 32'h395ede54;
    ram_cell[   24562] = 32'h8b2314a4;
    ram_cell[   24563] = 32'h84fa45eb;
    ram_cell[   24564] = 32'hb6a662df;
    ram_cell[   24565] = 32'h984e073d;
    ram_cell[   24566] = 32'h3437fbb3;
    ram_cell[   24567] = 32'ha1685548;
    ram_cell[   24568] = 32'h476811de;
    ram_cell[   24569] = 32'h4da3b62c;
    ram_cell[   24570] = 32'hcdcbfe89;
    ram_cell[   24571] = 32'hfa648850;
    ram_cell[   24572] = 32'h0d8cf452;
    ram_cell[   24573] = 32'h89ffeb12;
    ram_cell[   24574] = 32'h235d26e3;
    ram_cell[   24575] = 32'h4eca2abe;
    ram_cell[   24576] = 32'hf930fb39;
    ram_cell[   24577] = 32'h98e2816b;
    ram_cell[   24578] = 32'h9c814012;
    ram_cell[   24579] = 32'haf5282fe;
    ram_cell[   24580] = 32'h699ea38e;
    ram_cell[   24581] = 32'h56254472;
    ram_cell[   24582] = 32'h474cc932;
    ram_cell[   24583] = 32'h1b196c7b;
    ram_cell[   24584] = 32'h2cd161dd;
    ram_cell[   24585] = 32'h37eb7294;
    ram_cell[   24586] = 32'hb0a145e1;
    ram_cell[   24587] = 32'h0b38e7d5;
    ram_cell[   24588] = 32'hced7bb5a;
    ram_cell[   24589] = 32'h45359276;
    ram_cell[   24590] = 32'he6fc9e55;
    ram_cell[   24591] = 32'h0ab14a68;
    ram_cell[   24592] = 32'h22f78ed1;
    ram_cell[   24593] = 32'hd05e4527;
    ram_cell[   24594] = 32'h19abbe14;
    ram_cell[   24595] = 32'h58dc5321;
    ram_cell[   24596] = 32'h57af3574;
    ram_cell[   24597] = 32'hc553fa20;
    ram_cell[   24598] = 32'h784a7411;
    ram_cell[   24599] = 32'h5a601439;
    ram_cell[   24600] = 32'h0f6a4cb7;
    ram_cell[   24601] = 32'h4ec112b5;
    ram_cell[   24602] = 32'h0465bbe1;
    ram_cell[   24603] = 32'h3145db34;
    ram_cell[   24604] = 32'h8dcd437e;
    ram_cell[   24605] = 32'hf87968c3;
    ram_cell[   24606] = 32'hab31e0f5;
    ram_cell[   24607] = 32'hffe4af6a;
    ram_cell[   24608] = 32'h9118fa2f;
    ram_cell[   24609] = 32'h322a8cb5;
    ram_cell[   24610] = 32'hc09471a9;
    ram_cell[   24611] = 32'ha737e9dc;
    ram_cell[   24612] = 32'hbfff2a25;
    ram_cell[   24613] = 32'hc4cd8cd4;
    ram_cell[   24614] = 32'h764eb229;
    ram_cell[   24615] = 32'h22fe4d6d;
    ram_cell[   24616] = 32'h32a5f016;
    ram_cell[   24617] = 32'h9cc0b82e;
    ram_cell[   24618] = 32'hea713f4a;
    ram_cell[   24619] = 32'h0cd76c23;
    ram_cell[   24620] = 32'h58c83d34;
    ram_cell[   24621] = 32'h25d58f5e;
    ram_cell[   24622] = 32'hfbd793f9;
    ram_cell[   24623] = 32'h2a317fb5;
    ram_cell[   24624] = 32'hbc48dc6b;
    ram_cell[   24625] = 32'h332a2120;
    ram_cell[   24626] = 32'h4fe81769;
    ram_cell[   24627] = 32'hc7080c0b;
    ram_cell[   24628] = 32'h277846ec;
    ram_cell[   24629] = 32'hd94a60ef;
    ram_cell[   24630] = 32'h13266cc0;
    ram_cell[   24631] = 32'h052e847d;
    ram_cell[   24632] = 32'h597d9146;
    ram_cell[   24633] = 32'ha954a716;
    ram_cell[   24634] = 32'hf821c70a;
    ram_cell[   24635] = 32'h9c2d06ec;
    ram_cell[   24636] = 32'h99027c0f;
    ram_cell[   24637] = 32'h86592ad7;
    ram_cell[   24638] = 32'hbd5da56a;
    ram_cell[   24639] = 32'ha369b80a;
    ram_cell[   24640] = 32'h10423d84;
    ram_cell[   24641] = 32'he59859d9;
    ram_cell[   24642] = 32'ha8f7a46f;
    ram_cell[   24643] = 32'h77de5bf8;
    ram_cell[   24644] = 32'h38fa12ab;
    ram_cell[   24645] = 32'h078b1485;
    ram_cell[   24646] = 32'h10d6f328;
    ram_cell[   24647] = 32'h74d156f9;
    ram_cell[   24648] = 32'ha55fb2d7;
    ram_cell[   24649] = 32'h8f1d8706;
    ram_cell[   24650] = 32'hdd1fbc65;
    ram_cell[   24651] = 32'had80e942;
    ram_cell[   24652] = 32'h98904438;
    ram_cell[   24653] = 32'h182612cb;
    ram_cell[   24654] = 32'h16494ac8;
    ram_cell[   24655] = 32'hd2f678b4;
    ram_cell[   24656] = 32'h2ffadb7c;
    ram_cell[   24657] = 32'h5b1410b7;
    ram_cell[   24658] = 32'hff5392f0;
    ram_cell[   24659] = 32'h7f8ea2c1;
    ram_cell[   24660] = 32'h02c8d457;
    ram_cell[   24661] = 32'h082dd638;
    ram_cell[   24662] = 32'haebe3e60;
    ram_cell[   24663] = 32'ha4786140;
    ram_cell[   24664] = 32'hf0691097;
    ram_cell[   24665] = 32'hbc9cf878;
    ram_cell[   24666] = 32'h790be829;
    ram_cell[   24667] = 32'hc0bd41fe;
    ram_cell[   24668] = 32'hb2b6b02d;
    ram_cell[   24669] = 32'hc12cf82e;
    ram_cell[   24670] = 32'ha81c3ee0;
    ram_cell[   24671] = 32'h703ec207;
    ram_cell[   24672] = 32'hd9b8619f;
    ram_cell[   24673] = 32'h2d106963;
    ram_cell[   24674] = 32'h6e4b2307;
    ram_cell[   24675] = 32'h514e46a3;
    ram_cell[   24676] = 32'he6e9197d;
    ram_cell[   24677] = 32'hb956f3cb;
    ram_cell[   24678] = 32'hdff5cbdf;
    ram_cell[   24679] = 32'h599123f2;
    ram_cell[   24680] = 32'hb7175c7c;
    ram_cell[   24681] = 32'hf8cc44fd;
    ram_cell[   24682] = 32'hc152fbf7;
    ram_cell[   24683] = 32'h3a0f3bad;
    ram_cell[   24684] = 32'h5db3a00b;
    ram_cell[   24685] = 32'hffac16f0;
    ram_cell[   24686] = 32'h863a24b2;
    ram_cell[   24687] = 32'h57862386;
    ram_cell[   24688] = 32'hd7ceba67;
    ram_cell[   24689] = 32'h844b73de;
    ram_cell[   24690] = 32'hc2cda05a;
    ram_cell[   24691] = 32'h0d6c407d;
    ram_cell[   24692] = 32'hde9ba67a;
    ram_cell[   24693] = 32'h3e7dad18;
    ram_cell[   24694] = 32'hca9bd5ed;
    ram_cell[   24695] = 32'h46bcbd50;
    ram_cell[   24696] = 32'h20ec4238;
    ram_cell[   24697] = 32'hd501b557;
    ram_cell[   24698] = 32'h7c6611d4;
    ram_cell[   24699] = 32'h982999a8;
    ram_cell[   24700] = 32'h886758b2;
    ram_cell[   24701] = 32'hb31bb99b;
    ram_cell[   24702] = 32'he510e8fe;
    ram_cell[   24703] = 32'h28b40aac;
    ram_cell[   24704] = 32'h4dfbd9b6;
    ram_cell[   24705] = 32'hca8efd40;
    ram_cell[   24706] = 32'h882db125;
    ram_cell[   24707] = 32'h73a4124c;
    ram_cell[   24708] = 32'h4296ad0a;
    ram_cell[   24709] = 32'hd5b40513;
    ram_cell[   24710] = 32'h74cffe7b;
    ram_cell[   24711] = 32'h974908f6;
    ram_cell[   24712] = 32'h7519c5ba;
    ram_cell[   24713] = 32'hc03a3158;
    ram_cell[   24714] = 32'h3a6311ad;
    ram_cell[   24715] = 32'h0b622cc7;
    ram_cell[   24716] = 32'he7190492;
    ram_cell[   24717] = 32'hcf9a7a78;
    ram_cell[   24718] = 32'hcf97a920;
    ram_cell[   24719] = 32'h00260b90;
    ram_cell[   24720] = 32'h3ccb2ef4;
    ram_cell[   24721] = 32'hf2dfdf89;
    ram_cell[   24722] = 32'h2d79b0a6;
    ram_cell[   24723] = 32'h491515cc;
    ram_cell[   24724] = 32'h1bf2db4d;
    ram_cell[   24725] = 32'h78ca11a5;
    ram_cell[   24726] = 32'h488a97fc;
    ram_cell[   24727] = 32'h8586585a;
    ram_cell[   24728] = 32'h00676147;
    ram_cell[   24729] = 32'he3207d7e;
    ram_cell[   24730] = 32'h25c929b7;
    ram_cell[   24731] = 32'hdac2c200;
    ram_cell[   24732] = 32'h1020e184;
    ram_cell[   24733] = 32'h92f8155b;
    ram_cell[   24734] = 32'hddd2df5b;
    ram_cell[   24735] = 32'hc1984fb5;
    ram_cell[   24736] = 32'h4bfdc676;
    ram_cell[   24737] = 32'h4827358c;
    ram_cell[   24738] = 32'h7b33cfbe;
    ram_cell[   24739] = 32'h95d124b9;
    ram_cell[   24740] = 32'h664f81c7;
    ram_cell[   24741] = 32'hfa28e46e;
    ram_cell[   24742] = 32'h1c28b266;
    ram_cell[   24743] = 32'hfd8da858;
    ram_cell[   24744] = 32'hc42405b3;
    ram_cell[   24745] = 32'hcde55e17;
    ram_cell[   24746] = 32'hf053fa08;
    ram_cell[   24747] = 32'h81b19614;
    ram_cell[   24748] = 32'hb48abfa2;
    ram_cell[   24749] = 32'h65b3677d;
    ram_cell[   24750] = 32'h792270f9;
    ram_cell[   24751] = 32'hb933ffef;
    ram_cell[   24752] = 32'he9789287;
    ram_cell[   24753] = 32'h331a6870;
    ram_cell[   24754] = 32'hc0f5ac85;
    ram_cell[   24755] = 32'hf47bc676;
    ram_cell[   24756] = 32'h7a0b5f14;
    ram_cell[   24757] = 32'h93637f61;
    ram_cell[   24758] = 32'h669d3c16;
    ram_cell[   24759] = 32'h2b0eaa09;
    ram_cell[   24760] = 32'ha3869d72;
    ram_cell[   24761] = 32'haeafa8fa;
    ram_cell[   24762] = 32'h90c68e70;
    ram_cell[   24763] = 32'h2be2d2ed;
    ram_cell[   24764] = 32'hf7f1984f;
    ram_cell[   24765] = 32'h811aae12;
    ram_cell[   24766] = 32'hbb79b4af;
    ram_cell[   24767] = 32'hb7a70a77;
    ram_cell[   24768] = 32'ha5e1e908;
    ram_cell[   24769] = 32'h6ba19f19;
    ram_cell[   24770] = 32'h7935b93b;
    ram_cell[   24771] = 32'haf314dbd;
    ram_cell[   24772] = 32'hc167090b;
    ram_cell[   24773] = 32'h7296e4ae;
    ram_cell[   24774] = 32'hdc3ba13e;
    ram_cell[   24775] = 32'h3faeae44;
    ram_cell[   24776] = 32'h55eb2f7b;
    ram_cell[   24777] = 32'ha55d3c26;
    ram_cell[   24778] = 32'hedf314ed;
    ram_cell[   24779] = 32'h8466e090;
    ram_cell[   24780] = 32'h4dafc079;
    ram_cell[   24781] = 32'hd897f890;
    ram_cell[   24782] = 32'h4a0bdf9c;
    ram_cell[   24783] = 32'hd2015efa;
    ram_cell[   24784] = 32'h906b5149;
    ram_cell[   24785] = 32'ha7a025f9;
    ram_cell[   24786] = 32'hc0196448;
    ram_cell[   24787] = 32'h134caef7;
    ram_cell[   24788] = 32'hc88236ca;
    ram_cell[   24789] = 32'h673e3efb;
    ram_cell[   24790] = 32'h02ff9290;
    ram_cell[   24791] = 32'h11b761c4;
    ram_cell[   24792] = 32'hed2465ea;
    ram_cell[   24793] = 32'h916e54fc;
    ram_cell[   24794] = 32'h26da8d44;
    ram_cell[   24795] = 32'h465673d6;
    ram_cell[   24796] = 32'h6c4f7194;
    ram_cell[   24797] = 32'h1e06923b;
    ram_cell[   24798] = 32'h92fd8125;
    ram_cell[   24799] = 32'h4c92a7e6;
    ram_cell[   24800] = 32'hcdfc3518;
    ram_cell[   24801] = 32'h59afebe4;
    ram_cell[   24802] = 32'he96620cb;
    ram_cell[   24803] = 32'hddaf0831;
    ram_cell[   24804] = 32'h2a544a88;
    ram_cell[   24805] = 32'hc10df9be;
    ram_cell[   24806] = 32'h63126ea3;
    ram_cell[   24807] = 32'hf5f21d8f;
    ram_cell[   24808] = 32'h03a9a89d;
    ram_cell[   24809] = 32'hdd41f1d3;
    ram_cell[   24810] = 32'h07d52cd5;
    ram_cell[   24811] = 32'h66dead19;
    ram_cell[   24812] = 32'hc0473692;
    ram_cell[   24813] = 32'h27c9ca5a;
    ram_cell[   24814] = 32'h6bc340d9;
    ram_cell[   24815] = 32'h5bb1482c;
    ram_cell[   24816] = 32'hfb9403f8;
    ram_cell[   24817] = 32'h4c31671e;
    ram_cell[   24818] = 32'haec694c8;
    ram_cell[   24819] = 32'h80758ef3;
    ram_cell[   24820] = 32'h7fc88cd0;
    ram_cell[   24821] = 32'h33aa5a54;
    ram_cell[   24822] = 32'h0b9c9f16;
    ram_cell[   24823] = 32'he4aac761;
    ram_cell[   24824] = 32'hea5dac45;
    ram_cell[   24825] = 32'h53fb3c7d;
    ram_cell[   24826] = 32'h4632095c;
    ram_cell[   24827] = 32'ha97720a6;
    ram_cell[   24828] = 32'h5f67fba4;
    ram_cell[   24829] = 32'hff5698ef;
    ram_cell[   24830] = 32'ha6f8af7e;
    ram_cell[   24831] = 32'ha147c526;
    ram_cell[   24832] = 32'hf62fc435;
    ram_cell[   24833] = 32'h76023f1c;
    ram_cell[   24834] = 32'h70ff04a3;
    ram_cell[   24835] = 32'hd6e4195b;
    ram_cell[   24836] = 32'h4f79f8dd;
    ram_cell[   24837] = 32'h0823a66c;
    ram_cell[   24838] = 32'h2086012b;
    ram_cell[   24839] = 32'h7cb660e9;
    ram_cell[   24840] = 32'h09c30b2a;
    ram_cell[   24841] = 32'hea1530cc;
    ram_cell[   24842] = 32'h3655242d;
    ram_cell[   24843] = 32'h3cfd023a;
    ram_cell[   24844] = 32'h80619a4f;
    ram_cell[   24845] = 32'hde4f8370;
    ram_cell[   24846] = 32'h5f832ea4;
    ram_cell[   24847] = 32'hde597567;
    ram_cell[   24848] = 32'he400d33d;
    ram_cell[   24849] = 32'h3ae56967;
    ram_cell[   24850] = 32'h2ee988c2;
    ram_cell[   24851] = 32'h665f5e1a;
    ram_cell[   24852] = 32'ha1d3698e;
    ram_cell[   24853] = 32'hb7e53a96;
    ram_cell[   24854] = 32'hb5e685d3;
    ram_cell[   24855] = 32'h6b4d537c;
    ram_cell[   24856] = 32'ha1373079;
    ram_cell[   24857] = 32'hbfefbb26;
    ram_cell[   24858] = 32'h6f8fb782;
    ram_cell[   24859] = 32'hd18d4451;
    ram_cell[   24860] = 32'h53b34c85;
    ram_cell[   24861] = 32'h34999859;
    ram_cell[   24862] = 32'ha83a94e5;
    ram_cell[   24863] = 32'h56fb67f3;
    ram_cell[   24864] = 32'h90ba96d5;
    ram_cell[   24865] = 32'h879a20b0;
    ram_cell[   24866] = 32'h7c545dc4;
    ram_cell[   24867] = 32'h30578acf;
    ram_cell[   24868] = 32'h2dce542a;
    ram_cell[   24869] = 32'hbb81a077;
    ram_cell[   24870] = 32'hef9ef767;
    ram_cell[   24871] = 32'hb63fbfe5;
    ram_cell[   24872] = 32'ha246a982;
    ram_cell[   24873] = 32'hcbdfec48;
    ram_cell[   24874] = 32'hd01322d2;
    ram_cell[   24875] = 32'h801ada7e;
    ram_cell[   24876] = 32'hd8838bfe;
    ram_cell[   24877] = 32'h93936bf1;
    ram_cell[   24878] = 32'h7ac0fa50;
    ram_cell[   24879] = 32'hdf628990;
    ram_cell[   24880] = 32'h569a82e7;
    ram_cell[   24881] = 32'h9786c7db;
    ram_cell[   24882] = 32'had68246a;
    ram_cell[   24883] = 32'hd31055ff;
    ram_cell[   24884] = 32'h1ab37a06;
    ram_cell[   24885] = 32'ha5f7cb27;
    ram_cell[   24886] = 32'hc3ee7ca5;
    ram_cell[   24887] = 32'hef0ceb02;
    ram_cell[   24888] = 32'hfd2910ce;
    ram_cell[   24889] = 32'h279a7859;
    ram_cell[   24890] = 32'h02c54584;
    ram_cell[   24891] = 32'h04e841fe;
    ram_cell[   24892] = 32'hc9c422e8;
    ram_cell[   24893] = 32'ha5ee9a91;
    ram_cell[   24894] = 32'h07642588;
    ram_cell[   24895] = 32'hb788f8a8;
    ram_cell[   24896] = 32'h86bcd5b5;
    ram_cell[   24897] = 32'h986f87b3;
    ram_cell[   24898] = 32'h010a36c4;
    ram_cell[   24899] = 32'h930c374e;
    ram_cell[   24900] = 32'hf8cf5d39;
    ram_cell[   24901] = 32'h6e59c9df;
    ram_cell[   24902] = 32'hab900278;
    ram_cell[   24903] = 32'hfa09cf19;
    ram_cell[   24904] = 32'h2ba6556a;
    ram_cell[   24905] = 32'hb3563dd4;
    ram_cell[   24906] = 32'h29c2da39;
    ram_cell[   24907] = 32'h78ac210c;
    ram_cell[   24908] = 32'h2e090b7b;
    ram_cell[   24909] = 32'hba075320;
    ram_cell[   24910] = 32'h051da227;
    ram_cell[   24911] = 32'h9b700862;
    ram_cell[   24912] = 32'h070fc8d6;
    ram_cell[   24913] = 32'h8888d389;
    ram_cell[   24914] = 32'h959244c0;
    ram_cell[   24915] = 32'h5cef8ec6;
    ram_cell[   24916] = 32'hff537f8f;
    ram_cell[   24917] = 32'h64f286c7;
    ram_cell[   24918] = 32'he2ba362d;
    ram_cell[   24919] = 32'h3c004aff;
    ram_cell[   24920] = 32'h0edda6c3;
    ram_cell[   24921] = 32'h2e1d8fb3;
    ram_cell[   24922] = 32'h9a23c74b;
    ram_cell[   24923] = 32'hc53c4af6;
    ram_cell[   24924] = 32'h40c01151;
    ram_cell[   24925] = 32'h04ab39d2;
    ram_cell[   24926] = 32'h12383c08;
    ram_cell[   24927] = 32'h755b318c;
    ram_cell[   24928] = 32'ha67a6545;
    ram_cell[   24929] = 32'h2fd7df60;
    ram_cell[   24930] = 32'hb799e030;
    ram_cell[   24931] = 32'h4548d0ab;
    ram_cell[   24932] = 32'h0f74dd04;
    ram_cell[   24933] = 32'h1cc902e5;
    ram_cell[   24934] = 32'he49fec77;
    ram_cell[   24935] = 32'hc8b6e9b1;
    ram_cell[   24936] = 32'hff602109;
    ram_cell[   24937] = 32'h0fb3c245;
    ram_cell[   24938] = 32'h43011050;
    ram_cell[   24939] = 32'h5fd6f68f;
    ram_cell[   24940] = 32'h0816901c;
    ram_cell[   24941] = 32'ha049a898;
    ram_cell[   24942] = 32'hf0cffb79;
    ram_cell[   24943] = 32'h88ff7263;
    ram_cell[   24944] = 32'h8b00632e;
    ram_cell[   24945] = 32'h1e6cc151;
    ram_cell[   24946] = 32'h248ffe70;
    ram_cell[   24947] = 32'h41899b25;
    ram_cell[   24948] = 32'hdb9521f4;
    ram_cell[   24949] = 32'he2ad2660;
    ram_cell[   24950] = 32'h89abf345;
    ram_cell[   24951] = 32'h7b4420bc;
    ram_cell[   24952] = 32'h5114f016;
    ram_cell[   24953] = 32'h6f279131;
    ram_cell[   24954] = 32'hcfa08585;
    ram_cell[   24955] = 32'hcac2c90b;
    ram_cell[   24956] = 32'hef36fea6;
    ram_cell[   24957] = 32'heefc5380;
    ram_cell[   24958] = 32'h7c416dcb;
    ram_cell[   24959] = 32'h0b2b1798;
    ram_cell[   24960] = 32'h68372874;
    ram_cell[   24961] = 32'h9685338a;
    ram_cell[   24962] = 32'h7471784b;
    ram_cell[   24963] = 32'h6d05c710;
    ram_cell[   24964] = 32'hef8d5d26;
    ram_cell[   24965] = 32'h24bf27a3;
    ram_cell[   24966] = 32'h2ffdcc72;
    ram_cell[   24967] = 32'hd7c23ec0;
    ram_cell[   24968] = 32'ha9afc4ca;
    ram_cell[   24969] = 32'h588e8cc2;
    ram_cell[   24970] = 32'h8733ff2c;
    ram_cell[   24971] = 32'h99e657af;
    ram_cell[   24972] = 32'hc8e121f4;
    ram_cell[   24973] = 32'he6cb5865;
    ram_cell[   24974] = 32'ha52900e7;
    ram_cell[   24975] = 32'h07c5c397;
    ram_cell[   24976] = 32'h3dcc618f;
    ram_cell[   24977] = 32'h9ad171b5;
    ram_cell[   24978] = 32'h97c8aeb3;
    ram_cell[   24979] = 32'hc6a56ff5;
    ram_cell[   24980] = 32'h00c0143a;
    ram_cell[   24981] = 32'h469fa369;
    ram_cell[   24982] = 32'h357712aa;
    ram_cell[   24983] = 32'h33072928;
    ram_cell[   24984] = 32'hcaf10866;
    ram_cell[   24985] = 32'h419339a4;
    ram_cell[   24986] = 32'h91857ccc;
    ram_cell[   24987] = 32'hfff79c19;
    ram_cell[   24988] = 32'ha3fe7e72;
    ram_cell[   24989] = 32'h5a5684f7;
    ram_cell[   24990] = 32'h6248f2c0;
    ram_cell[   24991] = 32'h2d02d800;
    ram_cell[   24992] = 32'h81f81f5b;
    ram_cell[   24993] = 32'h3b4fe7b7;
    ram_cell[   24994] = 32'h19ae2bc6;
    ram_cell[   24995] = 32'hae2136a4;
    ram_cell[   24996] = 32'h51bcf263;
    ram_cell[   24997] = 32'h4e86bff6;
    ram_cell[   24998] = 32'hd5c35e17;
    ram_cell[   24999] = 32'had14f498;
    ram_cell[   25000] = 32'hea5e57c8;
    ram_cell[   25001] = 32'h93085a04;
    ram_cell[   25002] = 32'h9acc7e81;
    ram_cell[   25003] = 32'h396127ac;
    ram_cell[   25004] = 32'h487b1212;
    ram_cell[   25005] = 32'h9ba22803;
    ram_cell[   25006] = 32'h70e870b5;
    ram_cell[   25007] = 32'hc722abfe;
    ram_cell[   25008] = 32'h2e0115c9;
    ram_cell[   25009] = 32'hcf4bfbee;
    ram_cell[   25010] = 32'h43475e91;
    ram_cell[   25011] = 32'hecc30faf;
    ram_cell[   25012] = 32'h8ff5104a;
    ram_cell[   25013] = 32'hb7dbca70;
    ram_cell[   25014] = 32'h41957594;
    ram_cell[   25015] = 32'hb974d7e8;
    ram_cell[   25016] = 32'h8826d042;
    ram_cell[   25017] = 32'h8f4ed6a0;
    ram_cell[   25018] = 32'he29f22d7;
    ram_cell[   25019] = 32'h7dfdbfc6;
    ram_cell[   25020] = 32'h173e79f5;
    ram_cell[   25021] = 32'hdf30203d;
    ram_cell[   25022] = 32'hae8d1414;
    ram_cell[   25023] = 32'h986280bd;
    ram_cell[   25024] = 32'h889e0c61;
    ram_cell[   25025] = 32'h5674c82c;
    ram_cell[   25026] = 32'hb1ba7294;
    ram_cell[   25027] = 32'h5ced6e73;
    ram_cell[   25028] = 32'hebc4ea28;
    ram_cell[   25029] = 32'ha1066d49;
    ram_cell[   25030] = 32'hbbd73b8f;
    ram_cell[   25031] = 32'h5c4964ba;
    ram_cell[   25032] = 32'h36a7fea1;
    ram_cell[   25033] = 32'h652bae5b;
    ram_cell[   25034] = 32'h8fb70cdd;
    ram_cell[   25035] = 32'he344de37;
    ram_cell[   25036] = 32'hb08694e0;
    ram_cell[   25037] = 32'h0bd00cbf;
    ram_cell[   25038] = 32'hcbdc8008;
    ram_cell[   25039] = 32'hcfffd859;
    ram_cell[   25040] = 32'h4630fcf3;
    ram_cell[   25041] = 32'h95f1d196;
    ram_cell[   25042] = 32'h2752a31e;
    ram_cell[   25043] = 32'h067f86e1;
    ram_cell[   25044] = 32'h93b4a6a0;
    ram_cell[   25045] = 32'h0ef1080a;
    ram_cell[   25046] = 32'h8a685f75;
    ram_cell[   25047] = 32'hc07b1812;
    ram_cell[   25048] = 32'hc564422b;
    ram_cell[   25049] = 32'h5098a3b3;
    ram_cell[   25050] = 32'h8aacaa83;
    ram_cell[   25051] = 32'h68458b30;
    ram_cell[   25052] = 32'hdf5da4a6;
    ram_cell[   25053] = 32'h07b5692e;
    ram_cell[   25054] = 32'h6f1d2c1f;
    ram_cell[   25055] = 32'h5afa5d4a;
    ram_cell[   25056] = 32'ha82dd901;
    ram_cell[   25057] = 32'hbe3de26e;
    ram_cell[   25058] = 32'h3aa9395d;
    ram_cell[   25059] = 32'ha4b22b82;
    ram_cell[   25060] = 32'h91feaa54;
    ram_cell[   25061] = 32'h8733a79a;
    ram_cell[   25062] = 32'h04417a6d;
    ram_cell[   25063] = 32'h606660fa;
    ram_cell[   25064] = 32'h092678ce;
    ram_cell[   25065] = 32'haec77024;
    ram_cell[   25066] = 32'ha945db00;
    ram_cell[   25067] = 32'h3fb41514;
    ram_cell[   25068] = 32'h19094ff4;
    ram_cell[   25069] = 32'h2ca353ed;
    ram_cell[   25070] = 32'h3f609958;
    ram_cell[   25071] = 32'h135190b3;
    ram_cell[   25072] = 32'h3b7c7581;
    ram_cell[   25073] = 32'h3e352642;
    ram_cell[   25074] = 32'h17b6644c;
    ram_cell[   25075] = 32'h713edfbd;
    ram_cell[   25076] = 32'h399aca16;
    ram_cell[   25077] = 32'h861c5f8d;
    ram_cell[   25078] = 32'h13244345;
    ram_cell[   25079] = 32'h77d8a1a6;
    ram_cell[   25080] = 32'h85613afd;
    ram_cell[   25081] = 32'h4d0b9017;
    ram_cell[   25082] = 32'h4b1320f6;
    ram_cell[   25083] = 32'h5c75bf6c;
    ram_cell[   25084] = 32'h781992bc;
    ram_cell[   25085] = 32'h0f47953e;
    ram_cell[   25086] = 32'h9df7a36d;
    ram_cell[   25087] = 32'h27efb6ae;
    ram_cell[   25088] = 32'hddf450c5;
    ram_cell[   25089] = 32'h5b2918c5;
    ram_cell[   25090] = 32'h6525b461;
    ram_cell[   25091] = 32'hfdcc4e8e;
    ram_cell[   25092] = 32'h41e87309;
    ram_cell[   25093] = 32'h8786d9c2;
    ram_cell[   25094] = 32'hda8001d9;
    ram_cell[   25095] = 32'h28e941d6;
    ram_cell[   25096] = 32'hfce6334e;
    ram_cell[   25097] = 32'h8167a1ec;
    ram_cell[   25098] = 32'hbc5bace3;
    ram_cell[   25099] = 32'h1a66e676;
    ram_cell[   25100] = 32'h7b26c8e4;
    ram_cell[   25101] = 32'h5c475de9;
    ram_cell[   25102] = 32'hf2c03c83;
    ram_cell[   25103] = 32'h6ee92b4b;
    ram_cell[   25104] = 32'hf9fa0311;
    ram_cell[   25105] = 32'h5a6c56df;
    ram_cell[   25106] = 32'hecec3939;
    ram_cell[   25107] = 32'h2b80de78;
    ram_cell[   25108] = 32'he5e14e96;
    ram_cell[   25109] = 32'h39dc95a7;
    ram_cell[   25110] = 32'h443019dc;
    ram_cell[   25111] = 32'hbbbf9fb0;
    ram_cell[   25112] = 32'hc61bd18e;
    ram_cell[   25113] = 32'h46efe4aa;
    ram_cell[   25114] = 32'h39efa7b2;
    ram_cell[   25115] = 32'h68d1d85c;
    ram_cell[   25116] = 32'h9e1e3a33;
    ram_cell[   25117] = 32'h7981cd39;
    ram_cell[   25118] = 32'h4f4bf706;
    ram_cell[   25119] = 32'hf771ef31;
    ram_cell[   25120] = 32'h973fca8d;
    ram_cell[   25121] = 32'h2865b70a;
    ram_cell[   25122] = 32'hd2416f04;
    ram_cell[   25123] = 32'he9cf8d90;
    ram_cell[   25124] = 32'h10a39908;
    ram_cell[   25125] = 32'h7bbb57b8;
    ram_cell[   25126] = 32'hdfbc9158;
    ram_cell[   25127] = 32'h1af678f5;
    ram_cell[   25128] = 32'hefee39c1;
    ram_cell[   25129] = 32'h3bdd230b;
    ram_cell[   25130] = 32'h573f2456;
    ram_cell[   25131] = 32'heccd2fbb;
    ram_cell[   25132] = 32'hdb96da17;
    ram_cell[   25133] = 32'h19ebfd5e;
    ram_cell[   25134] = 32'h2084e8a8;
    ram_cell[   25135] = 32'h2275e00e;
    ram_cell[   25136] = 32'hb839cb94;
    ram_cell[   25137] = 32'h3306f898;
    ram_cell[   25138] = 32'hafb228a6;
    ram_cell[   25139] = 32'h00ff1f54;
    ram_cell[   25140] = 32'hd983b7cc;
    ram_cell[   25141] = 32'h6dd115cd;
    ram_cell[   25142] = 32'h0ca0a595;
    ram_cell[   25143] = 32'h26aa710b;
    ram_cell[   25144] = 32'h25f4501b;
    ram_cell[   25145] = 32'h6d1a286f;
    ram_cell[   25146] = 32'h8d35ec8e;
    ram_cell[   25147] = 32'h7074a919;
    ram_cell[   25148] = 32'hfc53b507;
    ram_cell[   25149] = 32'h9be2d932;
    ram_cell[   25150] = 32'hbd8d423a;
    ram_cell[   25151] = 32'h4256aa9e;
    ram_cell[   25152] = 32'ha39d68de;
    ram_cell[   25153] = 32'h8d6bef81;
    ram_cell[   25154] = 32'h32d48143;
    ram_cell[   25155] = 32'haa5cfda8;
    ram_cell[   25156] = 32'h467d2c25;
    ram_cell[   25157] = 32'h8bb4bf41;
    ram_cell[   25158] = 32'h3fafd6e3;
    ram_cell[   25159] = 32'h8573c035;
    ram_cell[   25160] = 32'h9dbc4d1b;
    ram_cell[   25161] = 32'h8c06bb5a;
    ram_cell[   25162] = 32'h6ba948fd;
    ram_cell[   25163] = 32'he63cbdac;
    ram_cell[   25164] = 32'h55e7f342;
    ram_cell[   25165] = 32'hdfe9a253;
    ram_cell[   25166] = 32'hab63cc13;
    ram_cell[   25167] = 32'h71aa4a80;
    ram_cell[   25168] = 32'hbc17f10c;
    ram_cell[   25169] = 32'hc7a52b1e;
    ram_cell[   25170] = 32'h01ef6594;
    ram_cell[   25171] = 32'h231ba902;
    ram_cell[   25172] = 32'he7d9a7f5;
    ram_cell[   25173] = 32'h6de307eb;
    ram_cell[   25174] = 32'h0d4d709a;
    ram_cell[   25175] = 32'h6c11efe4;
    ram_cell[   25176] = 32'h06920a1c;
    ram_cell[   25177] = 32'hca50c380;
    ram_cell[   25178] = 32'h332b3932;
    ram_cell[   25179] = 32'h9cd907d5;
    ram_cell[   25180] = 32'hcb9f1b0b;
    ram_cell[   25181] = 32'h8148e2a2;
    ram_cell[   25182] = 32'hba002d4c;
    ram_cell[   25183] = 32'h04891c39;
    ram_cell[   25184] = 32'h2337904e;
    ram_cell[   25185] = 32'h85017f2e;
    ram_cell[   25186] = 32'h27728f94;
    ram_cell[   25187] = 32'h68e51952;
    ram_cell[   25188] = 32'h75c72a64;
    ram_cell[   25189] = 32'hd00564c8;
    ram_cell[   25190] = 32'hb040f2bf;
    ram_cell[   25191] = 32'h08304cd6;
    ram_cell[   25192] = 32'h7c6bcb2e;
    ram_cell[   25193] = 32'h40d91efc;
    ram_cell[   25194] = 32'h5c6b07a5;
    ram_cell[   25195] = 32'ha264f71c;
    ram_cell[   25196] = 32'hbf903162;
    ram_cell[   25197] = 32'h098c6fdd;
    ram_cell[   25198] = 32'h79ab3f3f;
    ram_cell[   25199] = 32'hbd8ea0f1;
    ram_cell[   25200] = 32'hf9863b75;
    ram_cell[   25201] = 32'h77e5d954;
    ram_cell[   25202] = 32'h8108006d;
    ram_cell[   25203] = 32'h00d95b0b;
    ram_cell[   25204] = 32'hd367affc;
    ram_cell[   25205] = 32'hdbe82631;
    ram_cell[   25206] = 32'hd9d4d207;
    ram_cell[   25207] = 32'hd98bcd16;
    ram_cell[   25208] = 32'h90161d2f;
    ram_cell[   25209] = 32'h333f8aab;
    ram_cell[   25210] = 32'h5149f34f;
    ram_cell[   25211] = 32'heecbaf56;
    ram_cell[   25212] = 32'hb82dacc6;
    ram_cell[   25213] = 32'h08943d70;
    ram_cell[   25214] = 32'hb52204ec;
    ram_cell[   25215] = 32'h32b5e2c5;
    ram_cell[   25216] = 32'hdffa37d9;
    ram_cell[   25217] = 32'he7bda99a;
    ram_cell[   25218] = 32'h9e6fd8e2;
    ram_cell[   25219] = 32'h23030c2b;
    ram_cell[   25220] = 32'h180d5d62;
    ram_cell[   25221] = 32'h84d88571;
    ram_cell[   25222] = 32'h14851257;
    ram_cell[   25223] = 32'hf90c4c65;
    ram_cell[   25224] = 32'ha78e6654;
    ram_cell[   25225] = 32'h344f773e;
    ram_cell[   25226] = 32'hfdd71ff7;
    ram_cell[   25227] = 32'hcfd37a90;
    ram_cell[   25228] = 32'h381d558c;
    ram_cell[   25229] = 32'h1684dd91;
    ram_cell[   25230] = 32'h096406fb;
    ram_cell[   25231] = 32'h0214b8d7;
    ram_cell[   25232] = 32'h89333d07;
    ram_cell[   25233] = 32'hc5d37b2c;
    ram_cell[   25234] = 32'hb064b7a9;
    ram_cell[   25235] = 32'h5644f60c;
    ram_cell[   25236] = 32'hbc12b708;
    ram_cell[   25237] = 32'h3a7671f2;
    ram_cell[   25238] = 32'hc10ccaac;
    ram_cell[   25239] = 32'h483496cb;
    ram_cell[   25240] = 32'h9fcf95b5;
    ram_cell[   25241] = 32'h712f3fdb;
    ram_cell[   25242] = 32'hae73c563;
    ram_cell[   25243] = 32'h98e502f4;
    ram_cell[   25244] = 32'he2fc0470;
    ram_cell[   25245] = 32'h6602d6af;
    ram_cell[   25246] = 32'h29eb1797;
    ram_cell[   25247] = 32'h43bace5f;
    ram_cell[   25248] = 32'h52894d92;
    ram_cell[   25249] = 32'h4401f157;
    ram_cell[   25250] = 32'h803f2c66;
    ram_cell[   25251] = 32'hbf1dc52d;
    ram_cell[   25252] = 32'h5d5bddba;
    ram_cell[   25253] = 32'h2f9078ea;
    ram_cell[   25254] = 32'h57a270a2;
    ram_cell[   25255] = 32'h31a6bca3;
    ram_cell[   25256] = 32'h2d251ca4;
    ram_cell[   25257] = 32'h32df3198;
    ram_cell[   25258] = 32'h467c0cd0;
    ram_cell[   25259] = 32'hffa454b9;
    ram_cell[   25260] = 32'h1ab54a76;
    ram_cell[   25261] = 32'h7caaf785;
    ram_cell[   25262] = 32'hef18f99c;
    ram_cell[   25263] = 32'hfbb1c105;
    ram_cell[   25264] = 32'ha1279881;
    ram_cell[   25265] = 32'haa7d5abf;
    ram_cell[   25266] = 32'h3a113b56;
    ram_cell[   25267] = 32'h940c093a;
    ram_cell[   25268] = 32'h60d0dcdb;
    ram_cell[   25269] = 32'h5323cf86;
    ram_cell[   25270] = 32'h82105a61;
    ram_cell[   25271] = 32'hff6ac825;
    ram_cell[   25272] = 32'hd2fe678f;
    ram_cell[   25273] = 32'h79d8162c;
    ram_cell[   25274] = 32'h44f0482d;
    ram_cell[   25275] = 32'h3303996c;
    ram_cell[   25276] = 32'h29cdf992;
    ram_cell[   25277] = 32'he4feda6b;
    ram_cell[   25278] = 32'h772b4f48;
    ram_cell[   25279] = 32'h74bd4dd4;
    ram_cell[   25280] = 32'hc23e874f;
    ram_cell[   25281] = 32'hb50068b6;
    ram_cell[   25282] = 32'h156a7cd6;
    ram_cell[   25283] = 32'ha9653b75;
    ram_cell[   25284] = 32'h8f1418c7;
    ram_cell[   25285] = 32'h58885c70;
    ram_cell[   25286] = 32'h4044d4e2;
    ram_cell[   25287] = 32'h52494a51;
    ram_cell[   25288] = 32'h19258405;
    ram_cell[   25289] = 32'hb5cabe2b;
    ram_cell[   25290] = 32'h278520b3;
    ram_cell[   25291] = 32'hfbb93dbc;
    ram_cell[   25292] = 32'h2936a665;
    ram_cell[   25293] = 32'h12b64109;
    ram_cell[   25294] = 32'h11e883f9;
    ram_cell[   25295] = 32'h411a20fa;
    ram_cell[   25296] = 32'h02bb9fe7;
    ram_cell[   25297] = 32'h99211dab;
    ram_cell[   25298] = 32'he57aa158;
    ram_cell[   25299] = 32'hac114fbd;
    ram_cell[   25300] = 32'hfe13a510;
    ram_cell[   25301] = 32'ha8cfd1df;
    ram_cell[   25302] = 32'h41d828c4;
    ram_cell[   25303] = 32'h76f26147;
    ram_cell[   25304] = 32'hea32b02b;
    ram_cell[   25305] = 32'hcd15aa3a;
    ram_cell[   25306] = 32'h7efee3ae;
    ram_cell[   25307] = 32'hdf9f7dc3;
    ram_cell[   25308] = 32'hf8b9f518;
    ram_cell[   25309] = 32'h432331bd;
    ram_cell[   25310] = 32'h6de0eaba;
    ram_cell[   25311] = 32'h10b1a2ca;
    ram_cell[   25312] = 32'hf8dd9940;
    ram_cell[   25313] = 32'h13708d28;
    ram_cell[   25314] = 32'h1e4fd745;
    ram_cell[   25315] = 32'h7a0e50f5;
    ram_cell[   25316] = 32'hd3df8655;
    ram_cell[   25317] = 32'h417d65b0;
    ram_cell[   25318] = 32'he2ace59f;
    ram_cell[   25319] = 32'he481f885;
    ram_cell[   25320] = 32'h2b88012f;
    ram_cell[   25321] = 32'h8c5b57cf;
    ram_cell[   25322] = 32'h9c0eb8c5;
    ram_cell[   25323] = 32'h3136eaae;
    ram_cell[   25324] = 32'hefc32b7c;
    ram_cell[   25325] = 32'h07a5e8d5;
    ram_cell[   25326] = 32'h2d662f8f;
    ram_cell[   25327] = 32'h8621b7b0;
    ram_cell[   25328] = 32'hb283a93e;
    ram_cell[   25329] = 32'h4a8126e9;
    ram_cell[   25330] = 32'h652edc21;
    ram_cell[   25331] = 32'h1a7bea1e;
    ram_cell[   25332] = 32'h101e8ed1;
    ram_cell[   25333] = 32'h6e762f71;
    ram_cell[   25334] = 32'hbbc96bac;
    ram_cell[   25335] = 32'h6cc40496;
    ram_cell[   25336] = 32'h4ce318d7;
    ram_cell[   25337] = 32'h45173766;
    ram_cell[   25338] = 32'h713ae750;
    ram_cell[   25339] = 32'hb81bb3c5;
    ram_cell[   25340] = 32'h9d61cd91;
    ram_cell[   25341] = 32'h02d5cc7e;
    ram_cell[   25342] = 32'h38a46d02;
    ram_cell[   25343] = 32'h6d6b3d2b;
    ram_cell[   25344] = 32'hfa7756e9;
    ram_cell[   25345] = 32'h2c1cb1cf;
    ram_cell[   25346] = 32'h229b2625;
    ram_cell[   25347] = 32'h3d9c4bcb;
    ram_cell[   25348] = 32'h1910a84e;
    ram_cell[   25349] = 32'he219c433;
    ram_cell[   25350] = 32'h7ebb8a0a;
    ram_cell[   25351] = 32'h4a8afda8;
    ram_cell[   25352] = 32'h0d12f31e;
    ram_cell[   25353] = 32'haf35e1dd;
    ram_cell[   25354] = 32'h9bdcb68e;
    ram_cell[   25355] = 32'hc9fa4a98;
    ram_cell[   25356] = 32'h8a102cd8;
    ram_cell[   25357] = 32'h25c90a23;
    ram_cell[   25358] = 32'h6d524a6a;
    ram_cell[   25359] = 32'h852db1e4;
    ram_cell[   25360] = 32'h12fc146e;
    ram_cell[   25361] = 32'h998a01d9;
    ram_cell[   25362] = 32'ha49819ad;
    ram_cell[   25363] = 32'h63da39fe;
    ram_cell[   25364] = 32'hfa6c1e18;
    ram_cell[   25365] = 32'h4dbd394d;
    ram_cell[   25366] = 32'h73688ddf;
    ram_cell[   25367] = 32'hfcfaf2ae;
    ram_cell[   25368] = 32'h0ec3c675;
    ram_cell[   25369] = 32'hddf46713;
    ram_cell[   25370] = 32'hc207cc42;
    ram_cell[   25371] = 32'ha13c1521;
    ram_cell[   25372] = 32'hdfbd3b17;
    ram_cell[   25373] = 32'h707a64d9;
    ram_cell[   25374] = 32'h813e8630;
    ram_cell[   25375] = 32'h5da3800e;
    ram_cell[   25376] = 32'h6404800a;
    ram_cell[   25377] = 32'hff729794;
    ram_cell[   25378] = 32'he6c5b671;
    ram_cell[   25379] = 32'h63b940c1;
    ram_cell[   25380] = 32'h64ca4825;
    ram_cell[   25381] = 32'h0bb4457d;
    ram_cell[   25382] = 32'h7659bc19;
    ram_cell[   25383] = 32'hcc0e18ee;
    ram_cell[   25384] = 32'h412ec739;
    ram_cell[   25385] = 32'hdbd71ad7;
    ram_cell[   25386] = 32'hcef6bf90;
    ram_cell[   25387] = 32'h53ab50e1;
    ram_cell[   25388] = 32'h7f601edb;
    ram_cell[   25389] = 32'h219fa392;
    ram_cell[   25390] = 32'h8983cc6a;
    ram_cell[   25391] = 32'hae89cb5c;
    ram_cell[   25392] = 32'hc6e0b2e3;
    ram_cell[   25393] = 32'haf3bffe2;
    ram_cell[   25394] = 32'h66fb44ac;
    ram_cell[   25395] = 32'h7c3ff582;
    ram_cell[   25396] = 32'h0b42e3aa;
    ram_cell[   25397] = 32'h9e5a36e8;
    ram_cell[   25398] = 32'hbb5d1252;
    ram_cell[   25399] = 32'h101615c5;
    ram_cell[   25400] = 32'hc5d349b4;
    ram_cell[   25401] = 32'h6e5e816d;
    ram_cell[   25402] = 32'hc8c31a36;
    ram_cell[   25403] = 32'h9d28c1b8;
    ram_cell[   25404] = 32'hb4df9c72;
    ram_cell[   25405] = 32'h8a0c9704;
    ram_cell[   25406] = 32'hdd37780e;
    ram_cell[   25407] = 32'heba75b54;
    ram_cell[   25408] = 32'h3d76cf30;
    ram_cell[   25409] = 32'h4c847352;
    ram_cell[   25410] = 32'h841d4c9e;
    ram_cell[   25411] = 32'h9c49f3dc;
    ram_cell[   25412] = 32'h6f1f90b5;
    ram_cell[   25413] = 32'h1d834f6d;
    ram_cell[   25414] = 32'hdaeb8ab0;
    ram_cell[   25415] = 32'h74a352d3;
    ram_cell[   25416] = 32'he1e2cb01;
    ram_cell[   25417] = 32'hd71a24e7;
    ram_cell[   25418] = 32'h41245350;
    ram_cell[   25419] = 32'h074fc742;
    ram_cell[   25420] = 32'hc7e2648f;
    ram_cell[   25421] = 32'h8a0d4082;
    ram_cell[   25422] = 32'h2966c22b;
    ram_cell[   25423] = 32'h5ea16d43;
    ram_cell[   25424] = 32'h2ce23b0b;
    ram_cell[   25425] = 32'h935b1fc8;
    ram_cell[   25426] = 32'h2937ef34;
    ram_cell[   25427] = 32'hee39f839;
    ram_cell[   25428] = 32'he859bb4c;
    ram_cell[   25429] = 32'h25c6faed;
    ram_cell[   25430] = 32'h6cbc8ec3;
    ram_cell[   25431] = 32'h0de67246;
    ram_cell[   25432] = 32'hdfb097b9;
    ram_cell[   25433] = 32'h78578865;
    ram_cell[   25434] = 32'hf3a3ea47;
    ram_cell[   25435] = 32'h41502f1f;
    ram_cell[   25436] = 32'h366e2b02;
    ram_cell[   25437] = 32'hb4092ffb;
    ram_cell[   25438] = 32'ha34de2a0;
    ram_cell[   25439] = 32'h485f4943;
    ram_cell[   25440] = 32'h5ef4f240;
    ram_cell[   25441] = 32'h01926a92;
    ram_cell[   25442] = 32'hf4febd41;
    ram_cell[   25443] = 32'h8584e6a7;
    ram_cell[   25444] = 32'hd8f01e00;
    ram_cell[   25445] = 32'h7d4736cc;
    ram_cell[   25446] = 32'hd56006e4;
    ram_cell[   25447] = 32'ha77ebbf6;
    ram_cell[   25448] = 32'h217422ee;
    ram_cell[   25449] = 32'h2cc58eb3;
    ram_cell[   25450] = 32'ha59b7da0;
    ram_cell[   25451] = 32'h62298867;
    ram_cell[   25452] = 32'hf74b1cd2;
    ram_cell[   25453] = 32'h68e2f9bc;
    ram_cell[   25454] = 32'h50981090;
    ram_cell[   25455] = 32'h6e6cf0a2;
    ram_cell[   25456] = 32'h797acbca;
    ram_cell[   25457] = 32'hbba83108;
    ram_cell[   25458] = 32'h2c81dfb4;
    ram_cell[   25459] = 32'hb2a92178;
    ram_cell[   25460] = 32'h2c2b9191;
    ram_cell[   25461] = 32'hbdef6a7e;
    ram_cell[   25462] = 32'hb3daca19;
    ram_cell[   25463] = 32'h45b2b045;
    ram_cell[   25464] = 32'h5b9f0420;
    ram_cell[   25465] = 32'h9ae83866;
    ram_cell[   25466] = 32'h3ba48c85;
    ram_cell[   25467] = 32'h8ca8a8ea;
    ram_cell[   25468] = 32'hf70fd57d;
    ram_cell[   25469] = 32'hd2815786;
    ram_cell[   25470] = 32'h67ce2cc1;
    ram_cell[   25471] = 32'h4b828451;
    ram_cell[   25472] = 32'hf50b8cf3;
    ram_cell[   25473] = 32'h562ce865;
    ram_cell[   25474] = 32'h381c54ac;
    ram_cell[   25475] = 32'hd4631a32;
    ram_cell[   25476] = 32'h5cad8da9;
    ram_cell[   25477] = 32'h676263fa;
    ram_cell[   25478] = 32'h4fa7692c;
    ram_cell[   25479] = 32'h6c08ad14;
    ram_cell[   25480] = 32'h99b0f803;
    ram_cell[   25481] = 32'hdad181b5;
    ram_cell[   25482] = 32'h2dbbc49b;
    ram_cell[   25483] = 32'h23ac6709;
    ram_cell[   25484] = 32'hc313acb3;
    ram_cell[   25485] = 32'h40fb4a6f;
    ram_cell[   25486] = 32'h75cb8b01;
    ram_cell[   25487] = 32'hca48fc77;
    ram_cell[   25488] = 32'hf1a8c4b3;
    ram_cell[   25489] = 32'hba8060d6;
    ram_cell[   25490] = 32'h251484c6;
    ram_cell[   25491] = 32'hdcb07967;
    ram_cell[   25492] = 32'h3877f42e;
    ram_cell[   25493] = 32'h925141d7;
    ram_cell[   25494] = 32'he387c87c;
    ram_cell[   25495] = 32'hff55a3a0;
    ram_cell[   25496] = 32'h87311721;
    ram_cell[   25497] = 32'h5c2d90a6;
    ram_cell[   25498] = 32'h15e834e2;
    ram_cell[   25499] = 32'haaec1770;
    ram_cell[   25500] = 32'hd81982d4;
    ram_cell[   25501] = 32'h9c83a735;
    ram_cell[   25502] = 32'h727e645b;
    ram_cell[   25503] = 32'h9990da60;
    ram_cell[   25504] = 32'he913080f;
    ram_cell[   25505] = 32'h53fdc6be;
    ram_cell[   25506] = 32'h5dd1534c;
    ram_cell[   25507] = 32'h2d329529;
    ram_cell[   25508] = 32'h79a75eb1;
    ram_cell[   25509] = 32'h07feeada;
    ram_cell[   25510] = 32'h51c89ca1;
    ram_cell[   25511] = 32'ha0977815;
    ram_cell[   25512] = 32'h7d178d62;
    ram_cell[   25513] = 32'had52f443;
    ram_cell[   25514] = 32'hf392f9e4;
    ram_cell[   25515] = 32'h4c9fd1cf;
    ram_cell[   25516] = 32'hd968d62e;
    ram_cell[   25517] = 32'hac67c502;
    ram_cell[   25518] = 32'h728d3df6;
    ram_cell[   25519] = 32'h19796d32;
    ram_cell[   25520] = 32'hc48b3a87;
    ram_cell[   25521] = 32'h5d087b66;
    ram_cell[   25522] = 32'h957976c4;
    ram_cell[   25523] = 32'hba0519a6;
    ram_cell[   25524] = 32'hbfe73ff6;
    ram_cell[   25525] = 32'h2a2438e0;
    ram_cell[   25526] = 32'hbaa58b68;
    ram_cell[   25527] = 32'h0ffa4b2b;
    ram_cell[   25528] = 32'h339b226d;
    ram_cell[   25529] = 32'h2a5a6929;
    ram_cell[   25530] = 32'h7687855c;
    ram_cell[   25531] = 32'h3a3ae661;
    ram_cell[   25532] = 32'h9ffe20b6;
    ram_cell[   25533] = 32'h7fa53715;
    ram_cell[   25534] = 32'h891d5236;
    ram_cell[   25535] = 32'h71472504;
    ram_cell[   25536] = 32'ha0962b4b;
    ram_cell[   25537] = 32'h620e39be;
    ram_cell[   25538] = 32'hf6c9c69b;
    ram_cell[   25539] = 32'h44e56790;
    ram_cell[   25540] = 32'h783d79a6;
    ram_cell[   25541] = 32'h674f23de;
    ram_cell[   25542] = 32'h26cd9d19;
    ram_cell[   25543] = 32'h7287fab1;
    ram_cell[   25544] = 32'h562870eb;
    ram_cell[   25545] = 32'h4e398d45;
    ram_cell[   25546] = 32'h98d30225;
    ram_cell[   25547] = 32'hff1b8a7e;
    ram_cell[   25548] = 32'he50c54c0;
    ram_cell[   25549] = 32'haffac245;
    ram_cell[   25550] = 32'haf2cf27a;
    ram_cell[   25551] = 32'hd4090d8d;
    ram_cell[   25552] = 32'hf1aa9f1a;
    ram_cell[   25553] = 32'hb28b068b;
    ram_cell[   25554] = 32'h11782187;
    ram_cell[   25555] = 32'h1ba6f800;
    ram_cell[   25556] = 32'hb2ab6516;
    ram_cell[   25557] = 32'ha814eda1;
    ram_cell[   25558] = 32'hdc3c3fbe;
    ram_cell[   25559] = 32'h47148380;
    ram_cell[   25560] = 32'h4a3ca2b6;
    ram_cell[   25561] = 32'h38c751e9;
    ram_cell[   25562] = 32'h62b893aa;
    ram_cell[   25563] = 32'ha54e8b73;
    ram_cell[   25564] = 32'hd85e1bcf;
    ram_cell[   25565] = 32'h941b66a3;
    ram_cell[   25566] = 32'h36f14c0d;
    ram_cell[   25567] = 32'h1981b030;
    ram_cell[   25568] = 32'h9eaa97b0;
    ram_cell[   25569] = 32'hc75704ed;
    ram_cell[   25570] = 32'hbf7a423c;
    ram_cell[   25571] = 32'h19f26c74;
    ram_cell[   25572] = 32'he8407e63;
    ram_cell[   25573] = 32'hf9ef49b7;
    ram_cell[   25574] = 32'h47c9af3c;
    ram_cell[   25575] = 32'he9365a15;
    ram_cell[   25576] = 32'hd4826953;
    ram_cell[   25577] = 32'hf2593e00;
    ram_cell[   25578] = 32'h640dcb30;
    ram_cell[   25579] = 32'h03110c47;
    ram_cell[   25580] = 32'h0564852d;
    ram_cell[   25581] = 32'h8b76c0d5;
    ram_cell[   25582] = 32'h2d794764;
    ram_cell[   25583] = 32'h913e7f5f;
    ram_cell[   25584] = 32'h295a7b7d;
    ram_cell[   25585] = 32'hcfa1e9a3;
    ram_cell[   25586] = 32'h7b5a0cb5;
    ram_cell[   25587] = 32'hb04d8a43;
    ram_cell[   25588] = 32'hd65a53df;
    ram_cell[   25589] = 32'h3200f5ee;
    ram_cell[   25590] = 32'h77c854bd;
    ram_cell[   25591] = 32'h32fa1a09;
    ram_cell[   25592] = 32'h4ebc3d4a;
    ram_cell[   25593] = 32'hb02c1b04;
    ram_cell[   25594] = 32'h067bbde0;
    ram_cell[   25595] = 32'h813d74a3;
    ram_cell[   25596] = 32'h65c4db35;
    ram_cell[   25597] = 32'h387ec10a;
    ram_cell[   25598] = 32'h5c0f53aa;
    ram_cell[   25599] = 32'h7e0a22f7;
    ram_cell[   25600] = 32'hea75f798;
    ram_cell[   25601] = 32'hb36eb245;
    ram_cell[   25602] = 32'hc32032fb;
    ram_cell[   25603] = 32'h1938fa80;
    ram_cell[   25604] = 32'h542274e0;
    ram_cell[   25605] = 32'hd21ebcae;
    ram_cell[   25606] = 32'h5653350c;
    ram_cell[   25607] = 32'h45c0a36e;
    ram_cell[   25608] = 32'h530f0d3a;
    ram_cell[   25609] = 32'h1650b763;
    ram_cell[   25610] = 32'h70c3edef;
    ram_cell[   25611] = 32'hae8d44fc;
    ram_cell[   25612] = 32'h9bd78ab8;
    ram_cell[   25613] = 32'h4a22cbea;
    ram_cell[   25614] = 32'h4553e0b3;
    ram_cell[   25615] = 32'hc078aa1e;
    ram_cell[   25616] = 32'h34507d6c;
    ram_cell[   25617] = 32'hcb62e9b1;
    ram_cell[   25618] = 32'h55f23d25;
    ram_cell[   25619] = 32'h2a4ad06d;
    ram_cell[   25620] = 32'h629b1be0;
    ram_cell[   25621] = 32'h8326b167;
    ram_cell[   25622] = 32'h82a84902;
    ram_cell[   25623] = 32'hd4232133;
    ram_cell[   25624] = 32'h347cf154;
    ram_cell[   25625] = 32'h9709d9a5;
    ram_cell[   25626] = 32'h6e7dacba;
    ram_cell[   25627] = 32'h99d2ef66;
    ram_cell[   25628] = 32'h36ec4cf3;
    ram_cell[   25629] = 32'h9faaf5a6;
    ram_cell[   25630] = 32'hc2352418;
    ram_cell[   25631] = 32'h5a1cbd6e;
    ram_cell[   25632] = 32'hb876f957;
    ram_cell[   25633] = 32'h200b9e08;
    ram_cell[   25634] = 32'h4b6e93ab;
    ram_cell[   25635] = 32'he4744364;
    ram_cell[   25636] = 32'hbbea4b4c;
    ram_cell[   25637] = 32'h28ae9854;
    ram_cell[   25638] = 32'ha6f51a4e;
    ram_cell[   25639] = 32'hc8dbfcd8;
    ram_cell[   25640] = 32'h7c337416;
    ram_cell[   25641] = 32'heb261138;
    ram_cell[   25642] = 32'h061a975a;
    ram_cell[   25643] = 32'h0bd65646;
    ram_cell[   25644] = 32'h9515631e;
    ram_cell[   25645] = 32'hc3e89bfa;
    ram_cell[   25646] = 32'hf8e5bf88;
    ram_cell[   25647] = 32'h4e6ba980;
    ram_cell[   25648] = 32'ha1b4ce58;
    ram_cell[   25649] = 32'hebe26f42;
    ram_cell[   25650] = 32'hb01b85ad;
    ram_cell[   25651] = 32'h57863cf8;
    ram_cell[   25652] = 32'hf3ff4d18;
    ram_cell[   25653] = 32'h0cc0f0b7;
    ram_cell[   25654] = 32'h97b435ed;
    ram_cell[   25655] = 32'ha204a631;
    ram_cell[   25656] = 32'h4dda4f3c;
    ram_cell[   25657] = 32'h03238086;
    ram_cell[   25658] = 32'h8dc42f78;
    ram_cell[   25659] = 32'ha4048b7a;
    ram_cell[   25660] = 32'h90549b2e;
    ram_cell[   25661] = 32'h64084198;
    ram_cell[   25662] = 32'hc61db7f8;
    ram_cell[   25663] = 32'hf8f113ea;
    ram_cell[   25664] = 32'h793f5d8f;
    ram_cell[   25665] = 32'h562051da;
    ram_cell[   25666] = 32'h7f86679d;
    ram_cell[   25667] = 32'h68043490;
    ram_cell[   25668] = 32'h7c0ff6c5;
    ram_cell[   25669] = 32'h7918d1a5;
    ram_cell[   25670] = 32'h5b87a980;
    ram_cell[   25671] = 32'hfda19ddc;
    ram_cell[   25672] = 32'h0c0f03e8;
    ram_cell[   25673] = 32'h087c5ec1;
    ram_cell[   25674] = 32'h6c08fac3;
    ram_cell[   25675] = 32'h194c152a;
    ram_cell[   25676] = 32'h476a7943;
    ram_cell[   25677] = 32'hbf6c053f;
    ram_cell[   25678] = 32'he59d15c4;
    ram_cell[   25679] = 32'he7d81292;
    ram_cell[   25680] = 32'hc077bffa;
    ram_cell[   25681] = 32'h1edcc68f;
    ram_cell[   25682] = 32'h14d798fc;
    ram_cell[   25683] = 32'h1514c778;
    ram_cell[   25684] = 32'h18efb073;
    ram_cell[   25685] = 32'hc2d1d479;
    ram_cell[   25686] = 32'h13fd332e;
    ram_cell[   25687] = 32'h467ec654;
    ram_cell[   25688] = 32'hdba3696d;
    ram_cell[   25689] = 32'h17b7e12a;
    ram_cell[   25690] = 32'hcbc160e2;
    ram_cell[   25691] = 32'h2c33d20a;
    ram_cell[   25692] = 32'hc4ed080a;
    ram_cell[   25693] = 32'h005cea88;
    ram_cell[   25694] = 32'h720d5f2e;
    ram_cell[   25695] = 32'h19f6df2c;
    ram_cell[   25696] = 32'h12028492;
    ram_cell[   25697] = 32'h77404c4f;
    ram_cell[   25698] = 32'he24d8deb;
    ram_cell[   25699] = 32'h1f3f8611;
    ram_cell[   25700] = 32'hf4a0115a;
    ram_cell[   25701] = 32'hcc6eadcd;
    ram_cell[   25702] = 32'he73a9855;
    ram_cell[   25703] = 32'h42f200a9;
    ram_cell[   25704] = 32'hf9658481;
    ram_cell[   25705] = 32'hbd78006d;
    ram_cell[   25706] = 32'h3c9c605d;
    ram_cell[   25707] = 32'h4186b065;
    ram_cell[   25708] = 32'hd196b5ed;
    ram_cell[   25709] = 32'h63e10b3a;
    ram_cell[   25710] = 32'h5d6ac6ab;
    ram_cell[   25711] = 32'ha6e77a11;
    ram_cell[   25712] = 32'h67a7a944;
    ram_cell[   25713] = 32'h3333d240;
    ram_cell[   25714] = 32'ha81170cd;
    ram_cell[   25715] = 32'h1a071470;
    ram_cell[   25716] = 32'h706b49b0;
    ram_cell[   25717] = 32'h76e84d19;
    ram_cell[   25718] = 32'hb3bf6efe;
    ram_cell[   25719] = 32'h3fecfdc9;
    ram_cell[   25720] = 32'h7c3fa77b;
    ram_cell[   25721] = 32'hc67680db;
    ram_cell[   25722] = 32'ha57f02b2;
    ram_cell[   25723] = 32'hf0701d86;
    ram_cell[   25724] = 32'h71d707c0;
    ram_cell[   25725] = 32'h1312c535;
    ram_cell[   25726] = 32'heab2630b;
    ram_cell[   25727] = 32'h36ea5f61;
    ram_cell[   25728] = 32'h7774803b;
    ram_cell[   25729] = 32'ha1afbc06;
    ram_cell[   25730] = 32'h19bebd2a;
    ram_cell[   25731] = 32'h9def9486;
    ram_cell[   25732] = 32'h34a5e268;
    ram_cell[   25733] = 32'hf03e7f5d;
    ram_cell[   25734] = 32'h20ba060d;
    ram_cell[   25735] = 32'hc0855ab2;
    ram_cell[   25736] = 32'h1621e698;
    ram_cell[   25737] = 32'h7f36d4a9;
    ram_cell[   25738] = 32'h65653407;
    ram_cell[   25739] = 32'hc001876a;
    ram_cell[   25740] = 32'he638c9dd;
    ram_cell[   25741] = 32'h6d72994a;
    ram_cell[   25742] = 32'hbb5d38b0;
    ram_cell[   25743] = 32'h0ae1233d;
    ram_cell[   25744] = 32'h3a995c12;
    ram_cell[   25745] = 32'h9a53fe50;
    ram_cell[   25746] = 32'h2c07c1d1;
    ram_cell[   25747] = 32'h20c8a340;
    ram_cell[   25748] = 32'hec85fc14;
    ram_cell[   25749] = 32'h8c271221;
    ram_cell[   25750] = 32'h2293d603;
    ram_cell[   25751] = 32'h4ab0423f;
    ram_cell[   25752] = 32'h37b5e6f9;
    ram_cell[   25753] = 32'h84fb3023;
    ram_cell[   25754] = 32'h7d7066b7;
    ram_cell[   25755] = 32'h4e257328;
    ram_cell[   25756] = 32'hcd22f875;
    ram_cell[   25757] = 32'h60df0cb7;
    ram_cell[   25758] = 32'hbc4feb68;
    ram_cell[   25759] = 32'h91899bda;
    ram_cell[   25760] = 32'h36fb326c;
    ram_cell[   25761] = 32'h00c5ff10;
    ram_cell[   25762] = 32'h85b2be30;
    ram_cell[   25763] = 32'hfc865180;
    ram_cell[   25764] = 32'hf2478c32;
    ram_cell[   25765] = 32'h7adb588f;
    ram_cell[   25766] = 32'h62b92b5a;
    ram_cell[   25767] = 32'h6f0a6506;
    ram_cell[   25768] = 32'h03669071;
    ram_cell[   25769] = 32'hedb277c2;
    ram_cell[   25770] = 32'h8ad29048;
    ram_cell[   25771] = 32'hf0b62eb3;
    ram_cell[   25772] = 32'he3a5fed7;
    ram_cell[   25773] = 32'hf911db22;
    ram_cell[   25774] = 32'h6752d829;
    ram_cell[   25775] = 32'ha5322e5f;
    ram_cell[   25776] = 32'hb52b9b5a;
    ram_cell[   25777] = 32'h9b23aa20;
    ram_cell[   25778] = 32'h9e9c591f;
    ram_cell[   25779] = 32'h99b6550c;
    ram_cell[   25780] = 32'h4fca8c53;
    ram_cell[   25781] = 32'h0aff4efc;
    ram_cell[   25782] = 32'h7ff978b1;
    ram_cell[   25783] = 32'he55c8b70;
    ram_cell[   25784] = 32'h13e6175e;
    ram_cell[   25785] = 32'h0f58bd14;
    ram_cell[   25786] = 32'hda6ae61e;
    ram_cell[   25787] = 32'hcb21e8eb;
    ram_cell[   25788] = 32'hc59835c3;
    ram_cell[   25789] = 32'haac86d20;
    ram_cell[   25790] = 32'hc1773c0a;
    ram_cell[   25791] = 32'h13df9fc5;
    ram_cell[   25792] = 32'heff06439;
    ram_cell[   25793] = 32'hbda2c56c;
    ram_cell[   25794] = 32'h5f061a43;
    ram_cell[   25795] = 32'h44f76bbb;
    ram_cell[   25796] = 32'h38488ae4;
    ram_cell[   25797] = 32'hfe88b200;
    ram_cell[   25798] = 32'h0a7bb9d8;
    ram_cell[   25799] = 32'h2cae9f15;
    ram_cell[   25800] = 32'h911237dd;
    ram_cell[   25801] = 32'hc8de6f6d;
    ram_cell[   25802] = 32'haf03042b;
    ram_cell[   25803] = 32'hcde8e486;
    ram_cell[   25804] = 32'h6731b628;
    ram_cell[   25805] = 32'h38bce4f6;
    ram_cell[   25806] = 32'ha0ac18d9;
    ram_cell[   25807] = 32'hd7e4929b;
    ram_cell[   25808] = 32'h58bd9de5;
    ram_cell[   25809] = 32'hf01d6181;
    ram_cell[   25810] = 32'h1570be47;
    ram_cell[   25811] = 32'h1771d1f9;
    ram_cell[   25812] = 32'he184bcab;
    ram_cell[   25813] = 32'hb0bd3acb;
    ram_cell[   25814] = 32'h510e5db6;
    ram_cell[   25815] = 32'h49967394;
    ram_cell[   25816] = 32'h7d68aaba;
    ram_cell[   25817] = 32'he38fd45b;
    ram_cell[   25818] = 32'hb97c1350;
    ram_cell[   25819] = 32'hd56a9871;
    ram_cell[   25820] = 32'hde265805;
    ram_cell[   25821] = 32'h251c4dfc;
    ram_cell[   25822] = 32'he89a412c;
    ram_cell[   25823] = 32'h2d5dfe40;
    ram_cell[   25824] = 32'he70fb7ce;
    ram_cell[   25825] = 32'h45a3b4bb;
    ram_cell[   25826] = 32'h158c5695;
    ram_cell[   25827] = 32'hb26cc3a0;
    ram_cell[   25828] = 32'hbe61bb71;
    ram_cell[   25829] = 32'h90d6f0fb;
    ram_cell[   25830] = 32'hf11cffa6;
    ram_cell[   25831] = 32'hcb58eef0;
    ram_cell[   25832] = 32'ha70e6741;
    ram_cell[   25833] = 32'hd09053a9;
    ram_cell[   25834] = 32'h92c9e60b;
    ram_cell[   25835] = 32'hf8e0978e;
    ram_cell[   25836] = 32'hb0e81892;
    ram_cell[   25837] = 32'h8d00af80;
    ram_cell[   25838] = 32'h9ae26786;
    ram_cell[   25839] = 32'hd9c9ba6a;
    ram_cell[   25840] = 32'h14a2ab38;
    ram_cell[   25841] = 32'hdee76a01;
    ram_cell[   25842] = 32'hbc4c947d;
    ram_cell[   25843] = 32'hd2da6f3d;
    ram_cell[   25844] = 32'hb2b5de3a;
    ram_cell[   25845] = 32'h12f159df;
    ram_cell[   25846] = 32'hb0ad91f4;
    ram_cell[   25847] = 32'h5df2b9a8;
    ram_cell[   25848] = 32'h19e33110;
    ram_cell[   25849] = 32'hc35569ae;
    ram_cell[   25850] = 32'h5c48355c;
    ram_cell[   25851] = 32'h0506031a;
    ram_cell[   25852] = 32'h38760151;
    ram_cell[   25853] = 32'h6dcda48b;
    ram_cell[   25854] = 32'h178a5738;
    ram_cell[   25855] = 32'h371374f6;
    ram_cell[   25856] = 32'h62fe90fc;
    ram_cell[   25857] = 32'h07596b27;
    ram_cell[   25858] = 32'hb7116644;
    ram_cell[   25859] = 32'h3c78759d;
    ram_cell[   25860] = 32'h3d8e797e;
    ram_cell[   25861] = 32'h53730647;
    ram_cell[   25862] = 32'h7864f8da;
    ram_cell[   25863] = 32'h74b1a05f;
    ram_cell[   25864] = 32'h4ac9d618;
    ram_cell[   25865] = 32'h013a21b8;
    ram_cell[   25866] = 32'hba2c2af0;
    ram_cell[   25867] = 32'h47b30c2f;
    ram_cell[   25868] = 32'h2778942d;
    ram_cell[   25869] = 32'h2e6303bf;
    ram_cell[   25870] = 32'hd487dc7c;
    ram_cell[   25871] = 32'h9a78a448;
    ram_cell[   25872] = 32'h3fca03c4;
    ram_cell[   25873] = 32'h27e57cad;
    ram_cell[   25874] = 32'hd2168972;
    ram_cell[   25875] = 32'hc977faae;
    ram_cell[   25876] = 32'h727095ee;
    ram_cell[   25877] = 32'h4abb11b0;
    ram_cell[   25878] = 32'h3bee188a;
    ram_cell[   25879] = 32'hbca661a1;
    ram_cell[   25880] = 32'h2ad1edd2;
    ram_cell[   25881] = 32'h6f713ebc;
    ram_cell[   25882] = 32'h9ce400b2;
    ram_cell[   25883] = 32'h11b4227b;
    ram_cell[   25884] = 32'ha4df84b8;
    ram_cell[   25885] = 32'he98e47a3;
    ram_cell[   25886] = 32'h04ce2d35;
    ram_cell[   25887] = 32'h2b3b6aa8;
    ram_cell[   25888] = 32'h189a1657;
    ram_cell[   25889] = 32'ha4745279;
    ram_cell[   25890] = 32'h6c4fb344;
    ram_cell[   25891] = 32'h1d25d17b;
    ram_cell[   25892] = 32'he176b580;
    ram_cell[   25893] = 32'h0f8491e0;
    ram_cell[   25894] = 32'h7b3d13c6;
    ram_cell[   25895] = 32'hc9cf89cf;
    ram_cell[   25896] = 32'he2b11dcd;
    ram_cell[   25897] = 32'h44e6e0c8;
    ram_cell[   25898] = 32'h07ff6834;
    ram_cell[   25899] = 32'h60e67720;
    ram_cell[   25900] = 32'hf95a5a04;
    ram_cell[   25901] = 32'he6cf45bb;
    ram_cell[   25902] = 32'h0896605b;
    ram_cell[   25903] = 32'hfb28237f;
    ram_cell[   25904] = 32'h5badf238;
    ram_cell[   25905] = 32'h430321c8;
    ram_cell[   25906] = 32'hde17c5c8;
    ram_cell[   25907] = 32'h2e2cc021;
    ram_cell[   25908] = 32'he523808b;
    ram_cell[   25909] = 32'hccc37efd;
    ram_cell[   25910] = 32'haac28764;
    ram_cell[   25911] = 32'hd374a806;
    ram_cell[   25912] = 32'hc86a9624;
    ram_cell[   25913] = 32'h990c4b84;
    ram_cell[   25914] = 32'hcf940a34;
    ram_cell[   25915] = 32'he2b03ebe;
    ram_cell[   25916] = 32'hde13c1c6;
    ram_cell[   25917] = 32'h1e8251c2;
    ram_cell[   25918] = 32'hecea4e61;
    ram_cell[   25919] = 32'h33259a52;
    ram_cell[   25920] = 32'h868a71c5;
    ram_cell[   25921] = 32'h583a51ea;
    ram_cell[   25922] = 32'h1ab7220a;
    ram_cell[   25923] = 32'hd9c057a5;
    ram_cell[   25924] = 32'h3a5ba802;
    ram_cell[   25925] = 32'hc43ba1d1;
    ram_cell[   25926] = 32'h580ff136;
    ram_cell[   25927] = 32'hb494679c;
    ram_cell[   25928] = 32'h3d73c4d9;
    ram_cell[   25929] = 32'h5971e78e;
    ram_cell[   25930] = 32'h7c5d34e7;
    ram_cell[   25931] = 32'h3610ee3c;
    ram_cell[   25932] = 32'h7fef6c5d;
    ram_cell[   25933] = 32'h17da9e55;
    ram_cell[   25934] = 32'h8398bdf1;
    ram_cell[   25935] = 32'hc2f5db9e;
    ram_cell[   25936] = 32'hae1e1fea;
    ram_cell[   25937] = 32'h8e91f4a7;
    ram_cell[   25938] = 32'hc7902c9b;
    ram_cell[   25939] = 32'h5402a5d2;
    ram_cell[   25940] = 32'h0c23fde0;
    ram_cell[   25941] = 32'h7a6a05f2;
    ram_cell[   25942] = 32'hd5578296;
    ram_cell[   25943] = 32'hb7cb56d2;
    ram_cell[   25944] = 32'h6a25acd4;
    ram_cell[   25945] = 32'hec43a9d3;
    ram_cell[   25946] = 32'hdbdc1473;
    ram_cell[   25947] = 32'he653ef69;
    ram_cell[   25948] = 32'h095f0a01;
    ram_cell[   25949] = 32'h844b3008;
    ram_cell[   25950] = 32'hdd56ca78;
    ram_cell[   25951] = 32'h8547b0cd;
    ram_cell[   25952] = 32'h8048747b;
    ram_cell[   25953] = 32'h08ef1a87;
    ram_cell[   25954] = 32'h9df3e120;
    ram_cell[   25955] = 32'h877ff346;
    ram_cell[   25956] = 32'h5be7ad37;
    ram_cell[   25957] = 32'hee20246e;
    ram_cell[   25958] = 32'hba77366e;
    ram_cell[   25959] = 32'h6fc65b99;
    ram_cell[   25960] = 32'h99341503;
    ram_cell[   25961] = 32'h0b4c989a;
    ram_cell[   25962] = 32'hacd1cd0f;
    ram_cell[   25963] = 32'ha34d9805;
    ram_cell[   25964] = 32'hd53a6e49;
    ram_cell[   25965] = 32'h2b18e30b;
    ram_cell[   25966] = 32'h3714a254;
    ram_cell[   25967] = 32'hdf106546;
    ram_cell[   25968] = 32'he054086c;
    ram_cell[   25969] = 32'h6dfa660f;
    ram_cell[   25970] = 32'hd92abffb;
    ram_cell[   25971] = 32'h68d14959;
    ram_cell[   25972] = 32'hf0401065;
    ram_cell[   25973] = 32'h3476057a;
    ram_cell[   25974] = 32'h60f5f5a0;
    ram_cell[   25975] = 32'hf39994af;
    ram_cell[   25976] = 32'h45affcad;
    ram_cell[   25977] = 32'h3af6fe0f;
    ram_cell[   25978] = 32'h1b6db4e7;
    ram_cell[   25979] = 32'hb7b44ca1;
    ram_cell[   25980] = 32'h1a64ef01;
    ram_cell[   25981] = 32'h11914a79;
    ram_cell[   25982] = 32'h84ef7875;
    ram_cell[   25983] = 32'h5394f5bb;
    ram_cell[   25984] = 32'h630f453f;
    ram_cell[   25985] = 32'h1f9786f0;
    ram_cell[   25986] = 32'hee659997;
    ram_cell[   25987] = 32'h0a15f2a3;
    ram_cell[   25988] = 32'haf2787ae;
    ram_cell[   25989] = 32'h06daaef4;
    ram_cell[   25990] = 32'hbac464e8;
    ram_cell[   25991] = 32'hde2aa542;
    ram_cell[   25992] = 32'h1f70c3ab;
    ram_cell[   25993] = 32'hee7d9f42;
    ram_cell[   25994] = 32'h1b6da8f4;
    ram_cell[   25995] = 32'hd60a98fc;
    ram_cell[   25996] = 32'hc453ac8a;
    ram_cell[   25997] = 32'h91d8e840;
    ram_cell[   25998] = 32'h67c949bd;
    ram_cell[   25999] = 32'hbb27b654;
    ram_cell[   26000] = 32'h1b122203;
    ram_cell[   26001] = 32'h242ab169;
    ram_cell[   26002] = 32'h10dcc9ce;
    ram_cell[   26003] = 32'hd777a7e3;
    ram_cell[   26004] = 32'h7108d816;
    ram_cell[   26005] = 32'h6caab5f3;
    ram_cell[   26006] = 32'hd5bd3adb;
    ram_cell[   26007] = 32'he1f125a3;
    ram_cell[   26008] = 32'h71b5a792;
    ram_cell[   26009] = 32'hb6803f58;
    ram_cell[   26010] = 32'he1b95792;
    ram_cell[   26011] = 32'h521d5444;
    ram_cell[   26012] = 32'h742915cb;
    ram_cell[   26013] = 32'hca9ae46c;
    ram_cell[   26014] = 32'h84f9f01c;
    ram_cell[   26015] = 32'h7dc2b83f;
    ram_cell[   26016] = 32'he0465891;
    ram_cell[   26017] = 32'h0c3e7b42;
    ram_cell[   26018] = 32'h81c4a8fb;
    ram_cell[   26019] = 32'h1cd12b27;
    ram_cell[   26020] = 32'h7b9f632c;
    ram_cell[   26021] = 32'hed24a9d3;
    ram_cell[   26022] = 32'h4ee3cb84;
    ram_cell[   26023] = 32'h56a98213;
    ram_cell[   26024] = 32'h48e12ac7;
    ram_cell[   26025] = 32'h6dd00c83;
    ram_cell[   26026] = 32'hb89753d8;
    ram_cell[   26027] = 32'h1b73fdd8;
    ram_cell[   26028] = 32'he7c933ac;
    ram_cell[   26029] = 32'h0d61e188;
    ram_cell[   26030] = 32'h04e8dbfc;
    ram_cell[   26031] = 32'hc82eb35c;
    ram_cell[   26032] = 32'h301471cc;
    ram_cell[   26033] = 32'h36aff25b;
    ram_cell[   26034] = 32'he13c544c;
    ram_cell[   26035] = 32'h55c92fc3;
    ram_cell[   26036] = 32'h6c3dff07;
    ram_cell[   26037] = 32'h8e9d2609;
    ram_cell[   26038] = 32'h9219c7fb;
    ram_cell[   26039] = 32'h0dcf482c;
    ram_cell[   26040] = 32'h11c16c66;
    ram_cell[   26041] = 32'h0115d5b1;
    ram_cell[   26042] = 32'h37159627;
    ram_cell[   26043] = 32'h3d58e0a5;
    ram_cell[   26044] = 32'haf35cf1f;
    ram_cell[   26045] = 32'h0113bac9;
    ram_cell[   26046] = 32'hccf21a25;
    ram_cell[   26047] = 32'h58c22608;
    ram_cell[   26048] = 32'hd7881350;
    ram_cell[   26049] = 32'ha80a3749;
    ram_cell[   26050] = 32'hed925248;
    ram_cell[   26051] = 32'he85dc5ae;
    ram_cell[   26052] = 32'h1cf2a682;
    ram_cell[   26053] = 32'hd8eb1320;
    ram_cell[   26054] = 32'hdf2a9c6d;
    ram_cell[   26055] = 32'hef16ae19;
    ram_cell[   26056] = 32'h3e00744d;
    ram_cell[   26057] = 32'he4d48f5a;
    ram_cell[   26058] = 32'hcfebdc33;
    ram_cell[   26059] = 32'hb76a7999;
    ram_cell[   26060] = 32'h4ecf509d;
    ram_cell[   26061] = 32'heb6984b0;
    ram_cell[   26062] = 32'h1fc19f41;
    ram_cell[   26063] = 32'h77586a6c;
    ram_cell[   26064] = 32'ha1268044;
    ram_cell[   26065] = 32'h9209c606;
    ram_cell[   26066] = 32'hbe4fb045;
    ram_cell[   26067] = 32'hbe800083;
    ram_cell[   26068] = 32'h06ec506d;
    ram_cell[   26069] = 32'h40dad373;
    ram_cell[   26070] = 32'h2e42718e;
    ram_cell[   26071] = 32'h78a7a113;
    ram_cell[   26072] = 32'hfc4f26d9;
    ram_cell[   26073] = 32'hc6cb88a5;
    ram_cell[   26074] = 32'h3482fee1;
    ram_cell[   26075] = 32'h5be110da;
    ram_cell[   26076] = 32'h4c461b91;
    ram_cell[   26077] = 32'hc9e191d0;
    ram_cell[   26078] = 32'h85e9eea5;
    ram_cell[   26079] = 32'h5c68e2c1;
    ram_cell[   26080] = 32'h1627ea1c;
    ram_cell[   26081] = 32'h889fb235;
    ram_cell[   26082] = 32'h84bc4ddc;
    ram_cell[   26083] = 32'hd5bb3d62;
    ram_cell[   26084] = 32'h71588d23;
    ram_cell[   26085] = 32'h408fe2c1;
    ram_cell[   26086] = 32'hf976cf20;
    ram_cell[   26087] = 32'hd191f1cd;
    ram_cell[   26088] = 32'ha4a4dc17;
    ram_cell[   26089] = 32'h6998bde3;
    ram_cell[   26090] = 32'hba5b6552;
    ram_cell[   26091] = 32'h58c0d086;
    ram_cell[   26092] = 32'h42218103;
    ram_cell[   26093] = 32'h1e30c110;
    ram_cell[   26094] = 32'h971ba55a;
    ram_cell[   26095] = 32'h0f9aa241;
    ram_cell[   26096] = 32'hee4f48a6;
    ram_cell[   26097] = 32'he50d396f;
    ram_cell[   26098] = 32'hf6a02c94;
    ram_cell[   26099] = 32'hb74850fc;
    ram_cell[   26100] = 32'haf9ee9da;
    ram_cell[   26101] = 32'he272d80f;
    ram_cell[   26102] = 32'h6cfc897e;
    ram_cell[   26103] = 32'h46366c0e;
    ram_cell[   26104] = 32'hc70b80f9;
    ram_cell[   26105] = 32'h4b282fe2;
    ram_cell[   26106] = 32'h2f3f8713;
    ram_cell[   26107] = 32'h6e5666e9;
    ram_cell[   26108] = 32'hac73adf7;
    ram_cell[   26109] = 32'h71c64c7b;
    ram_cell[   26110] = 32'hcb6435e4;
    ram_cell[   26111] = 32'h5769e769;
    ram_cell[   26112] = 32'h6b72b288;
    ram_cell[   26113] = 32'h1d00f2c9;
    ram_cell[   26114] = 32'h896499fd;
    ram_cell[   26115] = 32'hc275cd14;
    ram_cell[   26116] = 32'hb04b3a92;
    ram_cell[   26117] = 32'hc5c2bfbf;
    ram_cell[   26118] = 32'h42550930;
    ram_cell[   26119] = 32'h16e5cf3e;
    ram_cell[   26120] = 32'h71c484db;
    ram_cell[   26121] = 32'h87f35c24;
    ram_cell[   26122] = 32'h9daa5e97;
    ram_cell[   26123] = 32'hd61db1aa;
    ram_cell[   26124] = 32'hbe736444;
    ram_cell[   26125] = 32'haa7a32aa;
    ram_cell[   26126] = 32'he093b3f7;
    ram_cell[   26127] = 32'hf7ac9c66;
    ram_cell[   26128] = 32'h9f656f28;
    ram_cell[   26129] = 32'hab9be800;
    ram_cell[   26130] = 32'h9e50590f;
    ram_cell[   26131] = 32'h859951f6;
    ram_cell[   26132] = 32'h65a656c5;
    ram_cell[   26133] = 32'hb2b53a6f;
    ram_cell[   26134] = 32'h6a2ad3c6;
    ram_cell[   26135] = 32'h69cdb0ab;
    ram_cell[   26136] = 32'ha4008988;
    ram_cell[   26137] = 32'h81e77cf8;
    ram_cell[   26138] = 32'hd983d74e;
    ram_cell[   26139] = 32'he45f34fb;
    ram_cell[   26140] = 32'hb3c568e7;
    ram_cell[   26141] = 32'h47cd3cc6;
    ram_cell[   26142] = 32'h65d52ed5;
    ram_cell[   26143] = 32'h315139e2;
    ram_cell[   26144] = 32'hb0d7e61b;
    ram_cell[   26145] = 32'h7f1ea9b4;
    ram_cell[   26146] = 32'h8f4c1188;
    ram_cell[   26147] = 32'h0fca9085;
    ram_cell[   26148] = 32'hfc516a2a;
    ram_cell[   26149] = 32'h096ab4e0;
    ram_cell[   26150] = 32'h89b6f768;
    ram_cell[   26151] = 32'h608a65aa;
    ram_cell[   26152] = 32'hc50e8489;
    ram_cell[   26153] = 32'h5cc43714;
    ram_cell[   26154] = 32'hc45bbb9b;
    ram_cell[   26155] = 32'h078fbe69;
    ram_cell[   26156] = 32'h2e6a9706;
    ram_cell[   26157] = 32'hef7cb6a7;
    ram_cell[   26158] = 32'h90c47591;
    ram_cell[   26159] = 32'hd81578db;
    ram_cell[   26160] = 32'h9550f85d;
    ram_cell[   26161] = 32'h6b3fcc56;
    ram_cell[   26162] = 32'hf3456b2e;
    ram_cell[   26163] = 32'hcba2c74e;
    ram_cell[   26164] = 32'h3f2e42a4;
    ram_cell[   26165] = 32'he1d0dc99;
    ram_cell[   26166] = 32'hc8602f4a;
    ram_cell[   26167] = 32'he2c7a5a9;
    ram_cell[   26168] = 32'h65f73f6c;
    ram_cell[   26169] = 32'hb2a69a7b;
    ram_cell[   26170] = 32'h6e24e6a6;
    ram_cell[   26171] = 32'ha4477e19;
    ram_cell[   26172] = 32'h2a0f27a3;
    ram_cell[   26173] = 32'hab5fc883;
    ram_cell[   26174] = 32'heefadbd4;
    ram_cell[   26175] = 32'h534fad7d;
    ram_cell[   26176] = 32'h1f1eb915;
    ram_cell[   26177] = 32'h0e04e68b;
    ram_cell[   26178] = 32'hcc746a1b;
    ram_cell[   26179] = 32'hf7c3a325;
    ram_cell[   26180] = 32'ha251ca96;
    ram_cell[   26181] = 32'hd55e9e1a;
    ram_cell[   26182] = 32'hf2828f92;
    ram_cell[   26183] = 32'h6a31948a;
    ram_cell[   26184] = 32'hcd55ee6a;
    ram_cell[   26185] = 32'hcd6db28f;
    ram_cell[   26186] = 32'hf517a6a3;
    ram_cell[   26187] = 32'hbb0908f6;
    ram_cell[   26188] = 32'hf1d0a1be;
    ram_cell[   26189] = 32'h5b6369c2;
    ram_cell[   26190] = 32'hbd58597e;
    ram_cell[   26191] = 32'h28f39d12;
    ram_cell[   26192] = 32'h336eaf4b;
    ram_cell[   26193] = 32'hc168c8a3;
    ram_cell[   26194] = 32'h45cc7c72;
    ram_cell[   26195] = 32'hfc0aaeda;
    ram_cell[   26196] = 32'h74d62fe8;
    ram_cell[   26197] = 32'h67f9a1db;
    ram_cell[   26198] = 32'h92ae6ef2;
    ram_cell[   26199] = 32'hac7b0c00;
    ram_cell[   26200] = 32'hd5312918;
    ram_cell[   26201] = 32'h14cbdd2c;
    ram_cell[   26202] = 32'hd1be8480;
    ram_cell[   26203] = 32'h95756005;
    ram_cell[   26204] = 32'h3a905c1b;
    ram_cell[   26205] = 32'h1f84d83a;
    ram_cell[   26206] = 32'h1eb97bf4;
    ram_cell[   26207] = 32'h333dfaa8;
    ram_cell[   26208] = 32'h65efc790;
    ram_cell[   26209] = 32'hdbccd418;
    ram_cell[   26210] = 32'h4b278bd2;
    ram_cell[   26211] = 32'h479485ea;
    ram_cell[   26212] = 32'h2282fafc;
    ram_cell[   26213] = 32'h1b584b78;
    ram_cell[   26214] = 32'h62d688bd;
    ram_cell[   26215] = 32'h8abced93;
    ram_cell[   26216] = 32'h7f7dab5c;
    ram_cell[   26217] = 32'ha136f032;
    ram_cell[   26218] = 32'he40f9b9d;
    ram_cell[   26219] = 32'h67f559ba;
    ram_cell[   26220] = 32'hc0b155d0;
    ram_cell[   26221] = 32'h815ac62a;
    ram_cell[   26222] = 32'h3fb14235;
    ram_cell[   26223] = 32'h904e12e5;
    ram_cell[   26224] = 32'he6839822;
    ram_cell[   26225] = 32'h16898445;
    ram_cell[   26226] = 32'he51dd504;
    ram_cell[   26227] = 32'h385e9265;
    ram_cell[   26228] = 32'hb6654d3e;
    ram_cell[   26229] = 32'hbe890727;
    ram_cell[   26230] = 32'h1185dc6a;
    ram_cell[   26231] = 32'h4cd4dcc6;
    ram_cell[   26232] = 32'he56452d1;
    ram_cell[   26233] = 32'h491efb36;
    ram_cell[   26234] = 32'hf71d6dba;
    ram_cell[   26235] = 32'h2bd62812;
    ram_cell[   26236] = 32'h19b32585;
    ram_cell[   26237] = 32'hc9ac2be3;
    ram_cell[   26238] = 32'h2572b8c9;
    ram_cell[   26239] = 32'hd7fac6d7;
    ram_cell[   26240] = 32'hb568f80c;
    ram_cell[   26241] = 32'h23950dbd;
    ram_cell[   26242] = 32'he6077b91;
    ram_cell[   26243] = 32'h1b88866c;
    ram_cell[   26244] = 32'h4888aa32;
    ram_cell[   26245] = 32'h08bce455;
    ram_cell[   26246] = 32'h2dd18394;
    ram_cell[   26247] = 32'hc7704fac;
    ram_cell[   26248] = 32'h1f9c0198;
    ram_cell[   26249] = 32'h2030b87d;
    ram_cell[   26250] = 32'h79df3e27;
    ram_cell[   26251] = 32'h52738a03;
    ram_cell[   26252] = 32'h462f10cf;
    ram_cell[   26253] = 32'hd267a8ad;
    ram_cell[   26254] = 32'h83aab4aa;
    ram_cell[   26255] = 32'h69eea37b;
    ram_cell[   26256] = 32'h3df738b6;
    ram_cell[   26257] = 32'hd7a6b862;
    ram_cell[   26258] = 32'h1db9e797;
    ram_cell[   26259] = 32'h269c413b;
    ram_cell[   26260] = 32'hbb85bfea;
    ram_cell[   26261] = 32'h38a83955;
    ram_cell[   26262] = 32'h53f6eff8;
    ram_cell[   26263] = 32'hc4361808;
    ram_cell[   26264] = 32'hde40c365;
    ram_cell[   26265] = 32'h53101d5c;
    ram_cell[   26266] = 32'h21a9f82a;
    ram_cell[   26267] = 32'h8109d319;
    ram_cell[   26268] = 32'h827a4b0a;
    ram_cell[   26269] = 32'hdcdb243a;
    ram_cell[   26270] = 32'h82bb2696;
    ram_cell[   26271] = 32'h90137ce8;
    ram_cell[   26272] = 32'h0444ffef;
    ram_cell[   26273] = 32'h8d26b97a;
    ram_cell[   26274] = 32'h3c24756b;
    ram_cell[   26275] = 32'h1ce8332a;
    ram_cell[   26276] = 32'hb2dc6714;
    ram_cell[   26277] = 32'hf7952034;
    ram_cell[   26278] = 32'h80126c55;
    ram_cell[   26279] = 32'hd878978a;
    ram_cell[   26280] = 32'h9486a230;
    ram_cell[   26281] = 32'hf3df6c9d;
    ram_cell[   26282] = 32'h0a6d2600;
    ram_cell[   26283] = 32'he42a2aa8;
    ram_cell[   26284] = 32'ha247f72c;
    ram_cell[   26285] = 32'he24012f1;
    ram_cell[   26286] = 32'hdd787480;
    ram_cell[   26287] = 32'hf8568f59;
    ram_cell[   26288] = 32'h277fca74;
    ram_cell[   26289] = 32'h045780c0;
    ram_cell[   26290] = 32'hc12bb068;
    ram_cell[   26291] = 32'h8b68a3f9;
    ram_cell[   26292] = 32'hd955e53a;
    ram_cell[   26293] = 32'hf0855f53;
    ram_cell[   26294] = 32'hce286380;
    ram_cell[   26295] = 32'h0f32ef0a;
    ram_cell[   26296] = 32'h4a483670;
    ram_cell[   26297] = 32'h0b6e5e9b;
    ram_cell[   26298] = 32'h17657999;
    ram_cell[   26299] = 32'hc0201e09;
    ram_cell[   26300] = 32'h2bca122b;
    ram_cell[   26301] = 32'h0b72223f;
    ram_cell[   26302] = 32'hf6156fc2;
    ram_cell[   26303] = 32'h007054fc;
    ram_cell[   26304] = 32'had702ad0;
    ram_cell[   26305] = 32'hca6acd5d;
    ram_cell[   26306] = 32'h54d28009;
    ram_cell[   26307] = 32'hb9e74e5c;
    ram_cell[   26308] = 32'he2d229d3;
    ram_cell[   26309] = 32'hcf546602;
    ram_cell[   26310] = 32'hc04285fe;
    ram_cell[   26311] = 32'h887e9b94;
    ram_cell[   26312] = 32'h7348c06d;
    ram_cell[   26313] = 32'h37ecb100;
    ram_cell[   26314] = 32'h6f2c0249;
    ram_cell[   26315] = 32'h9600ccff;
    ram_cell[   26316] = 32'he9cefad4;
    ram_cell[   26317] = 32'h9d4453fa;
    ram_cell[   26318] = 32'h735a832b;
    ram_cell[   26319] = 32'h60b4f6c3;
    ram_cell[   26320] = 32'h1fc7dd7c;
    ram_cell[   26321] = 32'hdcc6c264;
    ram_cell[   26322] = 32'h5224c696;
    ram_cell[   26323] = 32'h491f08a0;
    ram_cell[   26324] = 32'h1aa5fa2d;
    ram_cell[   26325] = 32'h4317650d;
    ram_cell[   26326] = 32'h1bb78515;
    ram_cell[   26327] = 32'h645754f4;
    ram_cell[   26328] = 32'h45326d67;
    ram_cell[   26329] = 32'hf31788b8;
    ram_cell[   26330] = 32'hc6e598b1;
    ram_cell[   26331] = 32'hbab298fa;
    ram_cell[   26332] = 32'hc4f1e597;
    ram_cell[   26333] = 32'hfc51418f;
    ram_cell[   26334] = 32'h535b7a08;
    ram_cell[   26335] = 32'h9daa1c23;
    ram_cell[   26336] = 32'h10213c71;
    ram_cell[   26337] = 32'hcc6088db;
    ram_cell[   26338] = 32'hb534ac70;
    ram_cell[   26339] = 32'hf834d2f0;
    ram_cell[   26340] = 32'h99efc53d;
    ram_cell[   26341] = 32'hf7e9c629;
    ram_cell[   26342] = 32'ha87c2f89;
    ram_cell[   26343] = 32'hdeaac3f2;
    ram_cell[   26344] = 32'h3b6b6c47;
    ram_cell[   26345] = 32'hafb99710;
    ram_cell[   26346] = 32'h38335227;
    ram_cell[   26347] = 32'h81423e5d;
    ram_cell[   26348] = 32'h0fc1a3b3;
    ram_cell[   26349] = 32'h70c4a15f;
    ram_cell[   26350] = 32'h0c1e2504;
    ram_cell[   26351] = 32'he0228e54;
    ram_cell[   26352] = 32'h4eae0c37;
    ram_cell[   26353] = 32'hf7e48f88;
    ram_cell[   26354] = 32'haff8a5a5;
    ram_cell[   26355] = 32'hea331aba;
    ram_cell[   26356] = 32'h2420b2ad;
    ram_cell[   26357] = 32'hde113ce6;
    ram_cell[   26358] = 32'h3e6a6705;
    ram_cell[   26359] = 32'h51cbe377;
    ram_cell[   26360] = 32'hc21d8919;
    ram_cell[   26361] = 32'h19246f5c;
    ram_cell[   26362] = 32'hdbbc393e;
    ram_cell[   26363] = 32'h802cc54b;
    ram_cell[   26364] = 32'h9f8f9493;
    ram_cell[   26365] = 32'h0a19045a;
    ram_cell[   26366] = 32'h79fe83b5;
    ram_cell[   26367] = 32'h28a72b84;
    ram_cell[   26368] = 32'h2334c34b;
    ram_cell[   26369] = 32'h78a82eb6;
    ram_cell[   26370] = 32'h99e15aa7;
    ram_cell[   26371] = 32'h561fae87;
    ram_cell[   26372] = 32'h31db7bd1;
    ram_cell[   26373] = 32'hbe9ee044;
    ram_cell[   26374] = 32'h03475e4f;
    ram_cell[   26375] = 32'hca428585;
    ram_cell[   26376] = 32'hc68f5751;
    ram_cell[   26377] = 32'h3c40ca64;
    ram_cell[   26378] = 32'hdd066436;
    ram_cell[   26379] = 32'he7556508;
    ram_cell[   26380] = 32'hafd72124;
    ram_cell[   26381] = 32'h40e28769;
    ram_cell[   26382] = 32'h08fb4f9e;
    ram_cell[   26383] = 32'hcb0c8a85;
    ram_cell[   26384] = 32'ha40e1186;
    ram_cell[   26385] = 32'hb788d029;
    ram_cell[   26386] = 32'h525db7cc;
    ram_cell[   26387] = 32'hb6352230;
    ram_cell[   26388] = 32'h5fcb8740;
    ram_cell[   26389] = 32'hd28053bc;
    ram_cell[   26390] = 32'h85aa1896;
    ram_cell[   26391] = 32'h045a3dfc;
    ram_cell[   26392] = 32'h1318f2b4;
    ram_cell[   26393] = 32'hbe94331c;
    ram_cell[   26394] = 32'hd9d2652b;
    ram_cell[   26395] = 32'hbc32a1fb;
    ram_cell[   26396] = 32'h5f3f4070;
    ram_cell[   26397] = 32'ha64d4f4f;
    ram_cell[   26398] = 32'h3f0f8b12;
    ram_cell[   26399] = 32'h12e6133c;
    ram_cell[   26400] = 32'hfb113cc2;
    ram_cell[   26401] = 32'h12b7cc5b;
    ram_cell[   26402] = 32'h2208d79d;
    ram_cell[   26403] = 32'h97c2abcb;
    ram_cell[   26404] = 32'h0208885a;
    ram_cell[   26405] = 32'h92b159c7;
    ram_cell[   26406] = 32'hbc6e214c;
    ram_cell[   26407] = 32'hf93b02e9;
    ram_cell[   26408] = 32'h2cae213d;
    ram_cell[   26409] = 32'he87233da;
    ram_cell[   26410] = 32'h64ac6172;
    ram_cell[   26411] = 32'h82c13820;
    ram_cell[   26412] = 32'hf95f3a45;
    ram_cell[   26413] = 32'h36c0f711;
    ram_cell[   26414] = 32'h15aa66fa;
    ram_cell[   26415] = 32'h1f114222;
    ram_cell[   26416] = 32'hb6794fda;
    ram_cell[   26417] = 32'h11b26b66;
    ram_cell[   26418] = 32'ha806f2b6;
    ram_cell[   26419] = 32'h7978c1fd;
    ram_cell[   26420] = 32'h58d41653;
    ram_cell[   26421] = 32'h6d02d37f;
    ram_cell[   26422] = 32'h44b49e2d;
    ram_cell[   26423] = 32'heeba033f;
    ram_cell[   26424] = 32'h06019d1f;
    ram_cell[   26425] = 32'h369f2392;
    ram_cell[   26426] = 32'h3706b562;
    ram_cell[   26427] = 32'hc6f2d934;
    ram_cell[   26428] = 32'hc62743b1;
    ram_cell[   26429] = 32'h035a27fd;
    ram_cell[   26430] = 32'h28c86983;
    ram_cell[   26431] = 32'h0519ddfb;
    ram_cell[   26432] = 32'h330cc0dc;
    ram_cell[   26433] = 32'hf239c3b0;
    ram_cell[   26434] = 32'h03c63883;
    ram_cell[   26435] = 32'h0f1d2d69;
    ram_cell[   26436] = 32'h0b574625;
    ram_cell[   26437] = 32'ha8c4836d;
    ram_cell[   26438] = 32'h07ee24a2;
    ram_cell[   26439] = 32'h3bc87c03;
    ram_cell[   26440] = 32'h9627fdc5;
    ram_cell[   26441] = 32'hed2413cb;
    ram_cell[   26442] = 32'h1422a9df;
    ram_cell[   26443] = 32'hf75af9ac;
    ram_cell[   26444] = 32'he2480d93;
    ram_cell[   26445] = 32'h580a57c7;
    ram_cell[   26446] = 32'h2c4b1961;
    ram_cell[   26447] = 32'hb721fe34;
    ram_cell[   26448] = 32'hab12b776;
    ram_cell[   26449] = 32'h369565ac;
    ram_cell[   26450] = 32'ha6990d04;
    ram_cell[   26451] = 32'hff0f2b90;
    ram_cell[   26452] = 32'h739f376a;
    ram_cell[   26453] = 32'h0f3c1629;
    ram_cell[   26454] = 32'h122bc055;
    ram_cell[   26455] = 32'h5309f4b7;
    ram_cell[   26456] = 32'h08dca9b5;
    ram_cell[   26457] = 32'h489b7d6e;
    ram_cell[   26458] = 32'hdd991ccc;
    ram_cell[   26459] = 32'h4b2d29c5;
    ram_cell[   26460] = 32'h683a5f93;
    ram_cell[   26461] = 32'h05ee7b89;
    ram_cell[   26462] = 32'hf82a250e;
    ram_cell[   26463] = 32'hf037b719;
    ram_cell[   26464] = 32'hfb56d5d8;
    ram_cell[   26465] = 32'hcea0a82e;
    ram_cell[   26466] = 32'h8a2e63a2;
    ram_cell[   26467] = 32'hb7e62ece;
    ram_cell[   26468] = 32'h8f1f6f7b;
    ram_cell[   26469] = 32'h3172df7e;
    ram_cell[   26470] = 32'h4c9f7e25;
    ram_cell[   26471] = 32'h6e006914;
    ram_cell[   26472] = 32'hbca1b8b7;
    ram_cell[   26473] = 32'hb4d7686c;
    ram_cell[   26474] = 32'hbd9d1d0d;
    ram_cell[   26475] = 32'h71bb060c;
    ram_cell[   26476] = 32'hf236d49b;
    ram_cell[   26477] = 32'hd1e73a73;
    ram_cell[   26478] = 32'h5562aeaa;
    ram_cell[   26479] = 32'hab8ad0d2;
    ram_cell[   26480] = 32'h8ff27fa4;
    ram_cell[   26481] = 32'hbf71e04c;
    ram_cell[   26482] = 32'hbf35aa3e;
    ram_cell[   26483] = 32'h8e479a3f;
    ram_cell[   26484] = 32'h7e7a449f;
    ram_cell[   26485] = 32'h87717aaa;
    ram_cell[   26486] = 32'h99953942;
    ram_cell[   26487] = 32'hc3e5a647;
    ram_cell[   26488] = 32'haa070a96;
    ram_cell[   26489] = 32'h3dcda4d1;
    ram_cell[   26490] = 32'he888568d;
    ram_cell[   26491] = 32'h43908f35;
    ram_cell[   26492] = 32'hce662628;
    ram_cell[   26493] = 32'h04875b09;
    ram_cell[   26494] = 32'hb919ab8a;
    ram_cell[   26495] = 32'h19abdc74;
    ram_cell[   26496] = 32'hf37b6154;
    ram_cell[   26497] = 32'h2a777c66;
    ram_cell[   26498] = 32'hcf468927;
    ram_cell[   26499] = 32'hc6e1c8dd;
    ram_cell[   26500] = 32'h708d4bcc;
    ram_cell[   26501] = 32'hfb801207;
    ram_cell[   26502] = 32'h02239df1;
    ram_cell[   26503] = 32'h9d6a5913;
    ram_cell[   26504] = 32'h6a7ea219;
    ram_cell[   26505] = 32'h9045d940;
    ram_cell[   26506] = 32'h9c66c9f1;
    ram_cell[   26507] = 32'h0bc95d3f;
    ram_cell[   26508] = 32'hdf41db55;
    ram_cell[   26509] = 32'h1772a41b;
    ram_cell[   26510] = 32'ha60d8cd7;
    ram_cell[   26511] = 32'h672c9042;
    ram_cell[   26512] = 32'h83af174d;
    ram_cell[   26513] = 32'hed22f75d;
    ram_cell[   26514] = 32'h428851af;
    ram_cell[   26515] = 32'hc50f52c7;
    ram_cell[   26516] = 32'h74d62035;
    ram_cell[   26517] = 32'h19fdb5e9;
    ram_cell[   26518] = 32'h275381be;
    ram_cell[   26519] = 32'had0fe604;
    ram_cell[   26520] = 32'h8df21ecf;
    ram_cell[   26521] = 32'h1705a54d;
    ram_cell[   26522] = 32'hf1b198df;
    ram_cell[   26523] = 32'hab376d24;
    ram_cell[   26524] = 32'h7a79e044;
    ram_cell[   26525] = 32'hdf50db69;
    ram_cell[   26526] = 32'h5c000591;
    ram_cell[   26527] = 32'h5f596ae1;
    ram_cell[   26528] = 32'h19bf1caa;
    ram_cell[   26529] = 32'h898d2718;
    ram_cell[   26530] = 32'he675b42e;
    ram_cell[   26531] = 32'h1519662b;
    ram_cell[   26532] = 32'h29f78f20;
    ram_cell[   26533] = 32'h5628b794;
    ram_cell[   26534] = 32'h3e50438f;
    ram_cell[   26535] = 32'hac505827;
    ram_cell[   26536] = 32'h73f9837e;
    ram_cell[   26537] = 32'h8eb22058;
    ram_cell[   26538] = 32'hd05d7451;
    ram_cell[   26539] = 32'h74a52e1b;
    ram_cell[   26540] = 32'h6bd03e0f;
    ram_cell[   26541] = 32'h6c32354e;
    ram_cell[   26542] = 32'hf2b0c2b5;
    ram_cell[   26543] = 32'hbe574602;
    ram_cell[   26544] = 32'h635a14fb;
    ram_cell[   26545] = 32'hf2284384;
    ram_cell[   26546] = 32'h244d5ba5;
    ram_cell[   26547] = 32'hfe399124;
    ram_cell[   26548] = 32'h61f0f4a4;
    ram_cell[   26549] = 32'h08fb6e5e;
    ram_cell[   26550] = 32'hd6609f52;
    ram_cell[   26551] = 32'h5632276d;
    ram_cell[   26552] = 32'hb3e6f7d7;
    ram_cell[   26553] = 32'h525c3ced;
    ram_cell[   26554] = 32'h82211990;
    ram_cell[   26555] = 32'h0fbc7864;
    ram_cell[   26556] = 32'h18b94879;
    ram_cell[   26557] = 32'hd416302d;
    ram_cell[   26558] = 32'h3e19eef3;
    ram_cell[   26559] = 32'h686b956f;
    ram_cell[   26560] = 32'h09e87534;
    ram_cell[   26561] = 32'h5a72861e;
    ram_cell[   26562] = 32'h4ee8e0a0;
    ram_cell[   26563] = 32'h263241cb;
    ram_cell[   26564] = 32'h4a51f702;
    ram_cell[   26565] = 32'had57070a;
    ram_cell[   26566] = 32'hebde7d47;
    ram_cell[   26567] = 32'ha8f25c5e;
    ram_cell[   26568] = 32'h6f571e06;
    ram_cell[   26569] = 32'h442cc645;
    ram_cell[   26570] = 32'hf7b9cbfd;
    ram_cell[   26571] = 32'hd9d7fb1d;
    ram_cell[   26572] = 32'hf6c35fbd;
    ram_cell[   26573] = 32'h285d5df2;
    ram_cell[   26574] = 32'h72539a15;
    ram_cell[   26575] = 32'hd6b15279;
    ram_cell[   26576] = 32'h1d23716c;
    ram_cell[   26577] = 32'h4bc72148;
    ram_cell[   26578] = 32'h8f874a0b;
    ram_cell[   26579] = 32'h88a2a126;
    ram_cell[   26580] = 32'h56fee837;
    ram_cell[   26581] = 32'hbe6389a9;
    ram_cell[   26582] = 32'h0b418ed9;
    ram_cell[   26583] = 32'h295db9d2;
    ram_cell[   26584] = 32'he3bb6b34;
    ram_cell[   26585] = 32'hd44385bb;
    ram_cell[   26586] = 32'h2aa5d784;
    ram_cell[   26587] = 32'hab6c4adf;
    ram_cell[   26588] = 32'h80ba1016;
    ram_cell[   26589] = 32'haf726945;
    ram_cell[   26590] = 32'h5d9fb3e1;
    ram_cell[   26591] = 32'hed47eb35;
    ram_cell[   26592] = 32'ha1793910;
    ram_cell[   26593] = 32'h080e9f23;
    ram_cell[   26594] = 32'hee3aa304;
    ram_cell[   26595] = 32'h210e5c53;
    ram_cell[   26596] = 32'h74b9136c;
    ram_cell[   26597] = 32'hc934c9dc;
    ram_cell[   26598] = 32'h58a86d61;
    ram_cell[   26599] = 32'h027e3582;
    ram_cell[   26600] = 32'h710783d0;
    ram_cell[   26601] = 32'h4c43f8bc;
    ram_cell[   26602] = 32'h49740de0;
    ram_cell[   26603] = 32'hf2699c55;
    ram_cell[   26604] = 32'h8a46be5d;
    ram_cell[   26605] = 32'hf2798ecb;
    ram_cell[   26606] = 32'h73326a82;
    ram_cell[   26607] = 32'h3570efb1;
    ram_cell[   26608] = 32'h71d98876;
    ram_cell[   26609] = 32'hd07174a8;
    ram_cell[   26610] = 32'hd5b9d064;
    ram_cell[   26611] = 32'h9810d411;
    ram_cell[   26612] = 32'h47f2363d;
    ram_cell[   26613] = 32'h8b5d51d7;
    ram_cell[   26614] = 32'ha0d7fa75;
    ram_cell[   26615] = 32'h84f84d93;
    ram_cell[   26616] = 32'h4ccbb1b2;
    ram_cell[   26617] = 32'h01de1e82;
    ram_cell[   26618] = 32'hb83624ac;
    ram_cell[   26619] = 32'h1584b713;
    ram_cell[   26620] = 32'h22509aa1;
    ram_cell[   26621] = 32'h2078c3b7;
    ram_cell[   26622] = 32'hfac3d891;
    ram_cell[   26623] = 32'hc7b620bc;
    ram_cell[   26624] = 32'hfb3daf95;
    ram_cell[   26625] = 32'h7d29b3fc;
    ram_cell[   26626] = 32'h515a83cc;
    ram_cell[   26627] = 32'h60c8f20f;
    ram_cell[   26628] = 32'h13f6d2df;
    ram_cell[   26629] = 32'h16bc919d;
    ram_cell[   26630] = 32'h6b454db8;
    ram_cell[   26631] = 32'h76047d9f;
    ram_cell[   26632] = 32'hb8fc19c7;
    ram_cell[   26633] = 32'h2ef3386d;
    ram_cell[   26634] = 32'h6e504aec;
    ram_cell[   26635] = 32'hc9670631;
    ram_cell[   26636] = 32'h5858035e;
    ram_cell[   26637] = 32'ha1da76e9;
    ram_cell[   26638] = 32'h4a82a92d;
    ram_cell[   26639] = 32'h91de75ac;
    ram_cell[   26640] = 32'h0bd33da9;
    ram_cell[   26641] = 32'h63ae3c47;
    ram_cell[   26642] = 32'h049da238;
    ram_cell[   26643] = 32'h439fe61c;
    ram_cell[   26644] = 32'h21189918;
    ram_cell[   26645] = 32'hdc5c9e1b;
    ram_cell[   26646] = 32'h1fa86f59;
    ram_cell[   26647] = 32'h45fa391f;
    ram_cell[   26648] = 32'h54e17848;
    ram_cell[   26649] = 32'hf6eb2124;
    ram_cell[   26650] = 32'h2f0f7b06;
    ram_cell[   26651] = 32'hebae7731;
    ram_cell[   26652] = 32'hdbbfdff3;
    ram_cell[   26653] = 32'h0634639d;
    ram_cell[   26654] = 32'hd713e2e3;
    ram_cell[   26655] = 32'h49aefff7;
    ram_cell[   26656] = 32'ha4446c92;
    ram_cell[   26657] = 32'hf02b6049;
    ram_cell[   26658] = 32'hbefb488b;
    ram_cell[   26659] = 32'h8a982c3d;
    ram_cell[   26660] = 32'hf05a1e67;
    ram_cell[   26661] = 32'hfcd2a1cd;
    ram_cell[   26662] = 32'h025d855b;
    ram_cell[   26663] = 32'h222ae2b4;
    ram_cell[   26664] = 32'he06af989;
    ram_cell[   26665] = 32'h16e4891d;
    ram_cell[   26666] = 32'ha350a87c;
    ram_cell[   26667] = 32'h4cd88445;
    ram_cell[   26668] = 32'h6a3cfee9;
    ram_cell[   26669] = 32'hdc2389b1;
    ram_cell[   26670] = 32'hd2c4e089;
    ram_cell[   26671] = 32'hd996e99c;
    ram_cell[   26672] = 32'h6166d01f;
    ram_cell[   26673] = 32'hdd7bf464;
    ram_cell[   26674] = 32'h412d4ce7;
    ram_cell[   26675] = 32'h558096db;
    ram_cell[   26676] = 32'h4d669d74;
    ram_cell[   26677] = 32'hab8896e3;
    ram_cell[   26678] = 32'h35b568c3;
    ram_cell[   26679] = 32'he463a41e;
    ram_cell[   26680] = 32'h7fcaac6b;
    ram_cell[   26681] = 32'hc93ebb88;
    ram_cell[   26682] = 32'h16019373;
    ram_cell[   26683] = 32'hb9187873;
    ram_cell[   26684] = 32'h39bf60a2;
    ram_cell[   26685] = 32'h289a8870;
    ram_cell[   26686] = 32'h50d9597c;
    ram_cell[   26687] = 32'ha09093ca;
    ram_cell[   26688] = 32'hba4aa412;
    ram_cell[   26689] = 32'h6c0b79c4;
    ram_cell[   26690] = 32'he4d7bf76;
    ram_cell[   26691] = 32'hddf6b33e;
    ram_cell[   26692] = 32'h088c3ecb;
    ram_cell[   26693] = 32'h41f83e7c;
    ram_cell[   26694] = 32'h5e6560fe;
    ram_cell[   26695] = 32'h2d400db3;
    ram_cell[   26696] = 32'hc22caca4;
    ram_cell[   26697] = 32'h290214b6;
    ram_cell[   26698] = 32'h4bd7fd18;
    ram_cell[   26699] = 32'h675d484d;
    ram_cell[   26700] = 32'h5fd2d2a1;
    ram_cell[   26701] = 32'hcf892711;
    ram_cell[   26702] = 32'h5c31520b;
    ram_cell[   26703] = 32'h9b123c3e;
    ram_cell[   26704] = 32'h35aabcb1;
    ram_cell[   26705] = 32'h6852cdbb;
    ram_cell[   26706] = 32'h91e64b00;
    ram_cell[   26707] = 32'h5f146546;
    ram_cell[   26708] = 32'h88e9c59c;
    ram_cell[   26709] = 32'h7c25f0d1;
    ram_cell[   26710] = 32'he6f4981e;
    ram_cell[   26711] = 32'h701065df;
    ram_cell[   26712] = 32'h2d9ef214;
    ram_cell[   26713] = 32'he5359638;
    ram_cell[   26714] = 32'ha89ab8fd;
    ram_cell[   26715] = 32'h06924396;
    ram_cell[   26716] = 32'h12184be1;
    ram_cell[   26717] = 32'hb093928c;
    ram_cell[   26718] = 32'hf25babd1;
    ram_cell[   26719] = 32'hc639dace;
    ram_cell[   26720] = 32'h764b9c1c;
    ram_cell[   26721] = 32'h081b3c3e;
    ram_cell[   26722] = 32'h7e86ce73;
    ram_cell[   26723] = 32'h542ac0b5;
    ram_cell[   26724] = 32'hb61e2c08;
    ram_cell[   26725] = 32'h6879294c;
    ram_cell[   26726] = 32'h195b60aa;
    ram_cell[   26727] = 32'h34e83b51;
    ram_cell[   26728] = 32'h298770d3;
    ram_cell[   26729] = 32'hedd55cc6;
    ram_cell[   26730] = 32'h4cfcb90f;
    ram_cell[   26731] = 32'hdb0d0ba4;
    ram_cell[   26732] = 32'h17017e7f;
    ram_cell[   26733] = 32'hadcabf5a;
    ram_cell[   26734] = 32'h800742d7;
    ram_cell[   26735] = 32'hf58555eb;
    ram_cell[   26736] = 32'h973958b5;
    ram_cell[   26737] = 32'h9d9ea9f5;
    ram_cell[   26738] = 32'he9386e2c;
    ram_cell[   26739] = 32'h21250f9f;
    ram_cell[   26740] = 32'hffb40b12;
    ram_cell[   26741] = 32'h910e86fc;
    ram_cell[   26742] = 32'h23b8f57b;
    ram_cell[   26743] = 32'h8a09cf54;
    ram_cell[   26744] = 32'h1f1a1d5c;
    ram_cell[   26745] = 32'h601ea5d7;
    ram_cell[   26746] = 32'h5c0e15c2;
    ram_cell[   26747] = 32'h1f8a051f;
    ram_cell[   26748] = 32'h2f882351;
    ram_cell[   26749] = 32'h248f26e6;
    ram_cell[   26750] = 32'h03f3b42e;
    ram_cell[   26751] = 32'hfbddaf39;
    ram_cell[   26752] = 32'h81ff910a;
    ram_cell[   26753] = 32'h491a8a4f;
    ram_cell[   26754] = 32'h44454b03;
    ram_cell[   26755] = 32'h21138bc7;
    ram_cell[   26756] = 32'h464bb2b5;
    ram_cell[   26757] = 32'hdaaeba59;
    ram_cell[   26758] = 32'hcaeadbdb;
    ram_cell[   26759] = 32'h054fa57d;
    ram_cell[   26760] = 32'h7b798930;
    ram_cell[   26761] = 32'hb329706d;
    ram_cell[   26762] = 32'hc103cf0a;
    ram_cell[   26763] = 32'h7dcd5095;
    ram_cell[   26764] = 32'h495a4bfd;
    ram_cell[   26765] = 32'he587632a;
    ram_cell[   26766] = 32'h10ce8ef2;
    ram_cell[   26767] = 32'h4f749464;
    ram_cell[   26768] = 32'h1f546567;
    ram_cell[   26769] = 32'hb8aa742e;
    ram_cell[   26770] = 32'hb6eaf7a9;
    ram_cell[   26771] = 32'h7aa3862a;
    ram_cell[   26772] = 32'h66847e5c;
    ram_cell[   26773] = 32'h056c52da;
    ram_cell[   26774] = 32'h32e57908;
    ram_cell[   26775] = 32'h71dcfcbe;
    ram_cell[   26776] = 32'h0473c2c0;
    ram_cell[   26777] = 32'h385f01d0;
    ram_cell[   26778] = 32'hc44ddb4f;
    ram_cell[   26779] = 32'h2296e939;
    ram_cell[   26780] = 32'hf4e78efb;
    ram_cell[   26781] = 32'h6d72ed92;
    ram_cell[   26782] = 32'h04f18fc9;
    ram_cell[   26783] = 32'hf8c1a751;
    ram_cell[   26784] = 32'h4fef54b8;
    ram_cell[   26785] = 32'h708744d6;
    ram_cell[   26786] = 32'hdd8282bf;
    ram_cell[   26787] = 32'h8bd5045d;
    ram_cell[   26788] = 32'h674a19d6;
    ram_cell[   26789] = 32'h4db75558;
    ram_cell[   26790] = 32'h14bffb44;
    ram_cell[   26791] = 32'haabdead6;
    ram_cell[   26792] = 32'hf6344607;
    ram_cell[   26793] = 32'h9c0891e1;
    ram_cell[   26794] = 32'hc2b86d63;
    ram_cell[   26795] = 32'h9bdc525c;
    ram_cell[   26796] = 32'hb066c623;
    ram_cell[   26797] = 32'hff23cfce;
    ram_cell[   26798] = 32'hb519e30a;
    ram_cell[   26799] = 32'h5f685a87;
    ram_cell[   26800] = 32'hf1cd089f;
    ram_cell[   26801] = 32'ha7972ef7;
    ram_cell[   26802] = 32'h5d56c1aa;
    ram_cell[   26803] = 32'hb4779ac7;
    ram_cell[   26804] = 32'h577ee597;
    ram_cell[   26805] = 32'he81cc3d1;
    ram_cell[   26806] = 32'h9149d295;
    ram_cell[   26807] = 32'h8eb4981f;
    ram_cell[   26808] = 32'ha02feb03;
    ram_cell[   26809] = 32'he5e2bfe8;
    ram_cell[   26810] = 32'h9404ec92;
    ram_cell[   26811] = 32'h59f72cf9;
    ram_cell[   26812] = 32'ha4595a61;
    ram_cell[   26813] = 32'h4aeec764;
    ram_cell[   26814] = 32'h5d2dca58;
    ram_cell[   26815] = 32'h8d2633d7;
    ram_cell[   26816] = 32'hfd449500;
    ram_cell[   26817] = 32'h88c33cc5;
    ram_cell[   26818] = 32'h3384ac68;
    ram_cell[   26819] = 32'h7c8f8755;
    ram_cell[   26820] = 32'h516aeb2c;
    ram_cell[   26821] = 32'h319450c4;
    ram_cell[   26822] = 32'h3548fe6c;
    ram_cell[   26823] = 32'h69d6355a;
    ram_cell[   26824] = 32'hcc504d69;
    ram_cell[   26825] = 32'h6234ee0d;
    ram_cell[   26826] = 32'h72dd1c18;
    ram_cell[   26827] = 32'h969baa5f;
    ram_cell[   26828] = 32'hbdb1d007;
    ram_cell[   26829] = 32'h26ea5bb4;
    ram_cell[   26830] = 32'ha9675cbb;
    ram_cell[   26831] = 32'h948a492b;
    ram_cell[   26832] = 32'habc2ecf8;
    ram_cell[   26833] = 32'h677b0aa9;
    ram_cell[   26834] = 32'hb340be23;
    ram_cell[   26835] = 32'hb0435133;
    ram_cell[   26836] = 32'h728e210f;
    ram_cell[   26837] = 32'hd3311fcf;
    ram_cell[   26838] = 32'h4ab11a14;
    ram_cell[   26839] = 32'hda3c675d;
    ram_cell[   26840] = 32'h71ef3d9b;
    ram_cell[   26841] = 32'h5fc53abb;
    ram_cell[   26842] = 32'h32cff843;
    ram_cell[   26843] = 32'h8e355cd7;
    ram_cell[   26844] = 32'hac755a41;
    ram_cell[   26845] = 32'h742a7ad8;
    ram_cell[   26846] = 32'heeb0d204;
    ram_cell[   26847] = 32'h5dfa425e;
    ram_cell[   26848] = 32'h20e5b1e6;
    ram_cell[   26849] = 32'h7c8bd134;
    ram_cell[   26850] = 32'hbf85d31c;
    ram_cell[   26851] = 32'h394c97c0;
    ram_cell[   26852] = 32'h49b91917;
    ram_cell[   26853] = 32'h33887122;
    ram_cell[   26854] = 32'h106b6f85;
    ram_cell[   26855] = 32'h7aca733d;
    ram_cell[   26856] = 32'h219311d2;
    ram_cell[   26857] = 32'h11124883;
    ram_cell[   26858] = 32'he8262758;
    ram_cell[   26859] = 32'h138dbbd7;
    ram_cell[   26860] = 32'h6f0275bc;
    ram_cell[   26861] = 32'h5219e0b0;
    ram_cell[   26862] = 32'h831168ca;
    ram_cell[   26863] = 32'h598d6ce9;
    ram_cell[   26864] = 32'h050c463a;
    ram_cell[   26865] = 32'ha9b56ea9;
    ram_cell[   26866] = 32'h71215a5e;
    ram_cell[   26867] = 32'h59020921;
    ram_cell[   26868] = 32'h5c31cd1c;
    ram_cell[   26869] = 32'hf51d0e18;
    ram_cell[   26870] = 32'h12dad382;
    ram_cell[   26871] = 32'h9df9e292;
    ram_cell[   26872] = 32'h58ed95f0;
    ram_cell[   26873] = 32'h924206d1;
    ram_cell[   26874] = 32'h414825e0;
    ram_cell[   26875] = 32'h3c4df626;
    ram_cell[   26876] = 32'h5548cd9e;
    ram_cell[   26877] = 32'h182fb29b;
    ram_cell[   26878] = 32'h4ae491fb;
    ram_cell[   26879] = 32'hec69e50f;
    ram_cell[   26880] = 32'ha8e520de;
    ram_cell[   26881] = 32'h56b60321;
    ram_cell[   26882] = 32'h16122f44;
    ram_cell[   26883] = 32'h8799cf6c;
    ram_cell[   26884] = 32'hf1fd163d;
    ram_cell[   26885] = 32'hfc607164;
    ram_cell[   26886] = 32'hd4811a80;
    ram_cell[   26887] = 32'haa6ef348;
    ram_cell[   26888] = 32'hf259b873;
    ram_cell[   26889] = 32'h6512ba87;
    ram_cell[   26890] = 32'h5dd1e965;
    ram_cell[   26891] = 32'h8a8f8699;
    ram_cell[   26892] = 32'h3ed17f90;
    ram_cell[   26893] = 32'h792d4a9b;
    ram_cell[   26894] = 32'h2eb2ea6e;
    ram_cell[   26895] = 32'h48ad9d08;
    ram_cell[   26896] = 32'h3ffb160b;
    ram_cell[   26897] = 32'h46131741;
    ram_cell[   26898] = 32'h1c0325eb;
    ram_cell[   26899] = 32'h1f0fdbeb;
    ram_cell[   26900] = 32'h7afcb5ed;
    ram_cell[   26901] = 32'h99a05d28;
    ram_cell[   26902] = 32'h738c3a66;
    ram_cell[   26903] = 32'hd8c6e2dc;
    ram_cell[   26904] = 32'hbddac5e8;
    ram_cell[   26905] = 32'h4014fb46;
    ram_cell[   26906] = 32'h257114d0;
    ram_cell[   26907] = 32'h14359fd1;
    ram_cell[   26908] = 32'he1fa9916;
    ram_cell[   26909] = 32'h614bd087;
    ram_cell[   26910] = 32'h59825ef0;
    ram_cell[   26911] = 32'h7738f434;
    ram_cell[   26912] = 32'h5629f100;
    ram_cell[   26913] = 32'hbeceb92b;
    ram_cell[   26914] = 32'h2ddb8309;
    ram_cell[   26915] = 32'hcdd7bcca;
    ram_cell[   26916] = 32'hbe13ef6a;
    ram_cell[   26917] = 32'h609bd325;
    ram_cell[   26918] = 32'h211ceea6;
    ram_cell[   26919] = 32'hb2dd0ee1;
    ram_cell[   26920] = 32'hebf19353;
    ram_cell[   26921] = 32'h87adf68f;
    ram_cell[   26922] = 32'h6e3a86ad;
    ram_cell[   26923] = 32'h4fad4ad4;
    ram_cell[   26924] = 32'hc3a16fb0;
    ram_cell[   26925] = 32'he9fce1db;
    ram_cell[   26926] = 32'h80d003d2;
    ram_cell[   26927] = 32'h40d1d037;
    ram_cell[   26928] = 32'hd4ec43f1;
    ram_cell[   26929] = 32'hf421a7cb;
    ram_cell[   26930] = 32'hb5fdb0f7;
    ram_cell[   26931] = 32'h421d6a52;
    ram_cell[   26932] = 32'haac1ec47;
    ram_cell[   26933] = 32'h7f7f045f;
    ram_cell[   26934] = 32'h13c80cf8;
    ram_cell[   26935] = 32'h0cbc2308;
    ram_cell[   26936] = 32'haa34611f;
    ram_cell[   26937] = 32'h745b30e4;
    ram_cell[   26938] = 32'h9725ba5d;
    ram_cell[   26939] = 32'h76b13d87;
    ram_cell[   26940] = 32'h2ff4144d;
    ram_cell[   26941] = 32'hea073c19;
    ram_cell[   26942] = 32'h4cddc775;
    ram_cell[   26943] = 32'h49b46613;
    ram_cell[   26944] = 32'ha54ea85c;
    ram_cell[   26945] = 32'h2b7978bb;
    ram_cell[   26946] = 32'h4ecd8d0f;
    ram_cell[   26947] = 32'h8f9a60b8;
    ram_cell[   26948] = 32'hdf36fbc5;
    ram_cell[   26949] = 32'he3caefb1;
    ram_cell[   26950] = 32'hfa57b01e;
    ram_cell[   26951] = 32'h763b2892;
    ram_cell[   26952] = 32'h4f53c650;
    ram_cell[   26953] = 32'hb21c5861;
    ram_cell[   26954] = 32'h430a6eb0;
    ram_cell[   26955] = 32'h69168b60;
    ram_cell[   26956] = 32'hc3119e41;
    ram_cell[   26957] = 32'haf67d051;
    ram_cell[   26958] = 32'h801dca43;
    ram_cell[   26959] = 32'hbdd2bf44;
    ram_cell[   26960] = 32'hce0f8f42;
    ram_cell[   26961] = 32'h68f6241f;
    ram_cell[   26962] = 32'he40b4a78;
    ram_cell[   26963] = 32'h9c643e08;
    ram_cell[   26964] = 32'hc61845dc;
    ram_cell[   26965] = 32'h59dc8b6c;
    ram_cell[   26966] = 32'h67741eb1;
    ram_cell[   26967] = 32'h4806510e;
    ram_cell[   26968] = 32'h3bb17fec;
    ram_cell[   26969] = 32'hc065c098;
    ram_cell[   26970] = 32'hdb68dfba;
    ram_cell[   26971] = 32'h1786dea5;
    ram_cell[   26972] = 32'hc4602334;
    ram_cell[   26973] = 32'h53325f63;
    ram_cell[   26974] = 32'h39499e84;
    ram_cell[   26975] = 32'h1a8774bd;
    ram_cell[   26976] = 32'hbb4bea64;
    ram_cell[   26977] = 32'hde7dbd91;
    ram_cell[   26978] = 32'h08b988f2;
    ram_cell[   26979] = 32'hf2465998;
    ram_cell[   26980] = 32'h0a1631a3;
    ram_cell[   26981] = 32'h6ba2bee8;
    ram_cell[   26982] = 32'h0432f8a1;
    ram_cell[   26983] = 32'hcd695763;
    ram_cell[   26984] = 32'hd6d256f8;
    ram_cell[   26985] = 32'h9a1f9d1b;
    ram_cell[   26986] = 32'ha1e87e48;
    ram_cell[   26987] = 32'h1d2770e7;
    ram_cell[   26988] = 32'h20ccae8f;
    ram_cell[   26989] = 32'h74794a5c;
    ram_cell[   26990] = 32'h565137f5;
    ram_cell[   26991] = 32'he2bdd9ad;
    ram_cell[   26992] = 32'h8441d7d5;
    ram_cell[   26993] = 32'h566fb97d;
    ram_cell[   26994] = 32'hcf6ab89e;
    ram_cell[   26995] = 32'hef3d7878;
    ram_cell[   26996] = 32'h27f81e4b;
    ram_cell[   26997] = 32'he9c8113c;
    ram_cell[   26998] = 32'h4436b8fc;
    ram_cell[   26999] = 32'h98256c1a;
    ram_cell[   27000] = 32'h215b8c69;
    ram_cell[   27001] = 32'h8faa2d5d;
    ram_cell[   27002] = 32'hde5d00c4;
    ram_cell[   27003] = 32'hc5e3e178;
    ram_cell[   27004] = 32'hacb728d9;
    ram_cell[   27005] = 32'he3389b4b;
    ram_cell[   27006] = 32'h33d692cb;
    ram_cell[   27007] = 32'h7f71431a;
    ram_cell[   27008] = 32'h0557d87b;
    ram_cell[   27009] = 32'he97b7e60;
    ram_cell[   27010] = 32'h8bb9213d;
    ram_cell[   27011] = 32'h39fce200;
    ram_cell[   27012] = 32'he8728cd1;
    ram_cell[   27013] = 32'h15f97fef;
    ram_cell[   27014] = 32'h7253a62b;
    ram_cell[   27015] = 32'h21679aec;
    ram_cell[   27016] = 32'h9f1a7e12;
    ram_cell[   27017] = 32'hc72276c4;
    ram_cell[   27018] = 32'hbf521b3a;
    ram_cell[   27019] = 32'h74e5b0ca;
    ram_cell[   27020] = 32'ha84a51bf;
    ram_cell[   27021] = 32'h3a3caecd;
    ram_cell[   27022] = 32'h8088fb4d;
    ram_cell[   27023] = 32'h8f71888f;
    ram_cell[   27024] = 32'ha0662f0d;
    ram_cell[   27025] = 32'hec4e594d;
    ram_cell[   27026] = 32'hf2b3ea40;
    ram_cell[   27027] = 32'hb00de623;
    ram_cell[   27028] = 32'h63f0e1ba;
    ram_cell[   27029] = 32'haa773ffe;
    ram_cell[   27030] = 32'h1436bc18;
    ram_cell[   27031] = 32'h50ae30c5;
    ram_cell[   27032] = 32'h039c1d69;
    ram_cell[   27033] = 32'h7b687069;
    ram_cell[   27034] = 32'h8f2cf941;
    ram_cell[   27035] = 32'h63f0e74a;
    ram_cell[   27036] = 32'h6574c372;
    ram_cell[   27037] = 32'he7c635d0;
    ram_cell[   27038] = 32'h7d1440ee;
    ram_cell[   27039] = 32'hb6917215;
    ram_cell[   27040] = 32'h56ab58f9;
    ram_cell[   27041] = 32'h29c4ba1a;
    ram_cell[   27042] = 32'h26ace2da;
    ram_cell[   27043] = 32'hde9da5aa;
    ram_cell[   27044] = 32'h31946585;
    ram_cell[   27045] = 32'hab760924;
    ram_cell[   27046] = 32'hd7ab6849;
    ram_cell[   27047] = 32'hdcd73811;
    ram_cell[   27048] = 32'h6b82dff4;
    ram_cell[   27049] = 32'h6e5245bf;
    ram_cell[   27050] = 32'ha87ab89b;
    ram_cell[   27051] = 32'hfc6182fb;
    ram_cell[   27052] = 32'h68d05fbc;
    ram_cell[   27053] = 32'h5787dc15;
    ram_cell[   27054] = 32'h4f8a2046;
    ram_cell[   27055] = 32'h1b57faa5;
    ram_cell[   27056] = 32'hbcfb8516;
    ram_cell[   27057] = 32'haf0edca0;
    ram_cell[   27058] = 32'h27999f8e;
    ram_cell[   27059] = 32'h78658a3e;
    ram_cell[   27060] = 32'h7ca366de;
    ram_cell[   27061] = 32'h7d3b7ee7;
    ram_cell[   27062] = 32'h1ae53fb9;
    ram_cell[   27063] = 32'hc6f0b384;
    ram_cell[   27064] = 32'hbb217c84;
    ram_cell[   27065] = 32'ha5abf2a2;
    ram_cell[   27066] = 32'hae191c81;
    ram_cell[   27067] = 32'h360f4ee2;
    ram_cell[   27068] = 32'h7eeb7481;
    ram_cell[   27069] = 32'h90e367b9;
    ram_cell[   27070] = 32'hb29238ac;
    ram_cell[   27071] = 32'h476ac1d0;
    ram_cell[   27072] = 32'h69f5c6e1;
    ram_cell[   27073] = 32'hb17e7844;
    ram_cell[   27074] = 32'h09693bc0;
    ram_cell[   27075] = 32'h5dd70f86;
    ram_cell[   27076] = 32'hc9e99227;
    ram_cell[   27077] = 32'h513fbcef;
    ram_cell[   27078] = 32'h632fb8fc;
    ram_cell[   27079] = 32'h7441724d;
    ram_cell[   27080] = 32'h899655b9;
    ram_cell[   27081] = 32'h9a2c30e8;
    ram_cell[   27082] = 32'hec9a4f20;
    ram_cell[   27083] = 32'h33456f73;
    ram_cell[   27084] = 32'h445d47c3;
    ram_cell[   27085] = 32'h4d8738c3;
    ram_cell[   27086] = 32'h2e319c37;
    ram_cell[   27087] = 32'h40e4c435;
    ram_cell[   27088] = 32'hfea3db7e;
    ram_cell[   27089] = 32'he9109ce4;
    ram_cell[   27090] = 32'h88d6df9f;
    ram_cell[   27091] = 32'hafe85f19;
    ram_cell[   27092] = 32'h9c780853;
    ram_cell[   27093] = 32'hb5596b8d;
    ram_cell[   27094] = 32'hd0717fa8;
    ram_cell[   27095] = 32'ha5bc26bf;
    ram_cell[   27096] = 32'had64f327;
    ram_cell[   27097] = 32'h794bc912;
    ram_cell[   27098] = 32'h016abc39;
    ram_cell[   27099] = 32'h7a4b7d73;
    ram_cell[   27100] = 32'h62c1eb5c;
    ram_cell[   27101] = 32'h150874f6;
    ram_cell[   27102] = 32'h4fc8ecb2;
    ram_cell[   27103] = 32'h467425fe;
    ram_cell[   27104] = 32'h4f1df167;
    ram_cell[   27105] = 32'he1cc68f3;
    ram_cell[   27106] = 32'hcca5b535;
    ram_cell[   27107] = 32'h8c1bb1c6;
    ram_cell[   27108] = 32'h4023d6b5;
    ram_cell[   27109] = 32'h42407e49;
    ram_cell[   27110] = 32'h67f6962d;
    ram_cell[   27111] = 32'h3e4f981b;
    ram_cell[   27112] = 32'hd7e4f741;
    ram_cell[   27113] = 32'h666d84a9;
    ram_cell[   27114] = 32'h17cf3fbf;
    ram_cell[   27115] = 32'h0e5e77a8;
    ram_cell[   27116] = 32'hf977d287;
    ram_cell[   27117] = 32'h91efc8e5;
    ram_cell[   27118] = 32'h08732573;
    ram_cell[   27119] = 32'h3eb88ddc;
    ram_cell[   27120] = 32'h4b2a002c;
    ram_cell[   27121] = 32'hd47ef001;
    ram_cell[   27122] = 32'h0306b53e;
    ram_cell[   27123] = 32'h316b7129;
    ram_cell[   27124] = 32'h5caa6467;
    ram_cell[   27125] = 32'h2015518c;
    ram_cell[   27126] = 32'h496b4f38;
    ram_cell[   27127] = 32'h5a6ee9e4;
    ram_cell[   27128] = 32'h97ba5528;
    ram_cell[   27129] = 32'hc1f062e8;
    ram_cell[   27130] = 32'h554fce6c;
    ram_cell[   27131] = 32'h4b57bc4b;
    ram_cell[   27132] = 32'h0ff7371a;
    ram_cell[   27133] = 32'hf6003b78;
    ram_cell[   27134] = 32'h7f49a137;
    ram_cell[   27135] = 32'h8b09c716;
    ram_cell[   27136] = 32'h2784409c;
    ram_cell[   27137] = 32'h4e099998;
    ram_cell[   27138] = 32'ha012888d;
    ram_cell[   27139] = 32'hde75c9ce;
    ram_cell[   27140] = 32'h5e36aed2;
    ram_cell[   27141] = 32'hfd4d91d1;
    ram_cell[   27142] = 32'h41ba924a;
    ram_cell[   27143] = 32'hcac704f3;
    ram_cell[   27144] = 32'he536c4bc;
    ram_cell[   27145] = 32'h1094c7d2;
    ram_cell[   27146] = 32'hef51d84c;
    ram_cell[   27147] = 32'h0fb8fb86;
    ram_cell[   27148] = 32'h2e8b5f41;
    ram_cell[   27149] = 32'h5f9e6f69;
    ram_cell[   27150] = 32'hd7b48907;
    ram_cell[   27151] = 32'hc3705c8d;
    ram_cell[   27152] = 32'h0f7ee877;
    ram_cell[   27153] = 32'he7d9b47f;
    ram_cell[   27154] = 32'hc96abbdf;
    ram_cell[   27155] = 32'h5f7021dd;
    ram_cell[   27156] = 32'h0eee3c2a;
    ram_cell[   27157] = 32'h18e6e3e3;
    ram_cell[   27158] = 32'h302781d0;
    ram_cell[   27159] = 32'h98ac705c;
    ram_cell[   27160] = 32'h51e8a109;
    ram_cell[   27161] = 32'h9a1b098e;
    ram_cell[   27162] = 32'hd60b8b60;
    ram_cell[   27163] = 32'hee40741d;
    ram_cell[   27164] = 32'h481a638a;
    ram_cell[   27165] = 32'h192aeb40;
    ram_cell[   27166] = 32'hbddfe3a6;
    ram_cell[   27167] = 32'h865a1122;
    ram_cell[   27168] = 32'h6c14598a;
    ram_cell[   27169] = 32'hc3994abc;
    ram_cell[   27170] = 32'hadf11482;
    ram_cell[   27171] = 32'h8d810f3a;
    ram_cell[   27172] = 32'hf7692449;
    ram_cell[   27173] = 32'h02357561;
    ram_cell[   27174] = 32'h783251af;
    ram_cell[   27175] = 32'hb8a6df0f;
    ram_cell[   27176] = 32'h82f8aa0f;
    ram_cell[   27177] = 32'h29534c28;
    ram_cell[   27178] = 32'h876979b9;
    ram_cell[   27179] = 32'hab07f17a;
    ram_cell[   27180] = 32'h0ff890b3;
    ram_cell[   27181] = 32'h9650620f;
    ram_cell[   27182] = 32'h60f5a6d5;
    ram_cell[   27183] = 32'h7e115647;
    ram_cell[   27184] = 32'h45c0cf14;
    ram_cell[   27185] = 32'h888a3048;
    ram_cell[   27186] = 32'h03bbdf69;
    ram_cell[   27187] = 32'h58836484;
    ram_cell[   27188] = 32'hf86b7c62;
    ram_cell[   27189] = 32'hf240b7f9;
    ram_cell[   27190] = 32'hacf18a88;
    ram_cell[   27191] = 32'hf4ce5dc8;
    ram_cell[   27192] = 32'hbb7ec1a0;
    ram_cell[   27193] = 32'hf3f36249;
    ram_cell[   27194] = 32'h7ed32d59;
    ram_cell[   27195] = 32'hfaf1f6f4;
    ram_cell[   27196] = 32'h70274949;
    ram_cell[   27197] = 32'h9f15af33;
    ram_cell[   27198] = 32'h30758f12;
    ram_cell[   27199] = 32'h7a5de7f3;
    ram_cell[   27200] = 32'ha25ed632;
    ram_cell[   27201] = 32'h7d33f8ca;
    ram_cell[   27202] = 32'hfb24f573;
    ram_cell[   27203] = 32'hf6c971cc;
    ram_cell[   27204] = 32'h58c28255;
    ram_cell[   27205] = 32'h5b5815e1;
    ram_cell[   27206] = 32'hb814a1de;
    ram_cell[   27207] = 32'h1a7dc51b;
    ram_cell[   27208] = 32'h781d2176;
    ram_cell[   27209] = 32'h27290c76;
    ram_cell[   27210] = 32'hb7e19c2a;
    ram_cell[   27211] = 32'h7b7baef6;
    ram_cell[   27212] = 32'h56a3c111;
    ram_cell[   27213] = 32'h45b62ec9;
    ram_cell[   27214] = 32'h47836462;
    ram_cell[   27215] = 32'h782deaed;
    ram_cell[   27216] = 32'he1e3ae89;
    ram_cell[   27217] = 32'h61c3957a;
    ram_cell[   27218] = 32'h177f9f64;
    ram_cell[   27219] = 32'hc88b9ad0;
    ram_cell[   27220] = 32'hcd3f3431;
    ram_cell[   27221] = 32'hc94c220c;
    ram_cell[   27222] = 32'he5af094e;
    ram_cell[   27223] = 32'h59e96c2e;
    ram_cell[   27224] = 32'h9e96c26d;
    ram_cell[   27225] = 32'h43548fa6;
    ram_cell[   27226] = 32'h09b54a5b;
    ram_cell[   27227] = 32'hf858a49b;
    ram_cell[   27228] = 32'hb940ad90;
    ram_cell[   27229] = 32'hcd42fc01;
    ram_cell[   27230] = 32'h93675713;
    ram_cell[   27231] = 32'hde38d879;
    ram_cell[   27232] = 32'h4aa8a51b;
    ram_cell[   27233] = 32'he4a494f8;
    ram_cell[   27234] = 32'hfc42b8b5;
    ram_cell[   27235] = 32'h718f621b;
    ram_cell[   27236] = 32'ha00a032b;
    ram_cell[   27237] = 32'h761fd0c4;
    ram_cell[   27238] = 32'h1ba52524;
    ram_cell[   27239] = 32'hd60252c5;
    ram_cell[   27240] = 32'h5012bfd0;
    ram_cell[   27241] = 32'h7ed0e787;
    ram_cell[   27242] = 32'hb3c41904;
    ram_cell[   27243] = 32'h5049dfad;
    ram_cell[   27244] = 32'hed57814d;
    ram_cell[   27245] = 32'hf4540247;
    ram_cell[   27246] = 32'h0691185e;
    ram_cell[   27247] = 32'h877d8867;
    ram_cell[   27248] = 32'h24198623;
    ram_cell[   27249] = 32'hfb995558;
    ram_cell[   27250] = 32'h508c61d9;
    ram_cell[   27251] = 32'h16e29064;
    ram_cell[   27252] = 32'h1078ec36;
    ram_cell[   27253] = 32'h100bb634;
    ram_cell[   27254] = 32'h44450bd9;
    ram_cell[   27255] = 32'h2fe4e13e;
    ram_cell[   27256] = 32'h32b10bf9;
    ram_cell[   27257] = 32'h0cb64435;
    ram_cell[   27258] = 32'hb7ae052b;
    ram_cell[   27259] = 32'h71b6c652;
    ram_cell[   27260] = 32'hfeec8fcf;
    ram_cell[   27261] = 32'h6a0ff387;
    ram_cell[   27262] = 32'hec8f18a4;
    ram_cell[   27263] = 32'h175a315b;
    ram_cell[   27264] = 32'ha77a9aea;
    ram_cell[   27265] = 32'h271fefb3;
    ram_cell[   27266] = 32'hb8550017;
    ram_cell[   27267] = 32'h575d1944;
    ram_cell[   27268] = 32'he71ad1b9;
    ram_cell[   27269] = 32'h7991cafe;
    ram_cell[   27270] = 32'h3a7679c6;
    ram_cell[   27271] = 32'h8588c8b3;
    ram_cell[   27272] = 32'h8ca8cc8a;
    ram_cell[   27273] = 32'h169ca44c;
    ram_cell[   27274] = 32'hcf5aa588;
    ram_cell[   27275] = 32'haad7d9a3;
    ram_cell[   27276] = 32'hf0521194;
    ram_cell[   27277] = 32'h59e9e317;
    ram_cell[   27278] = 32'h30b82aad;
    ram_cell[   27279] = 32'h65148d6e;
    ram_cell[   27280] = 32'h305abe10;
    ram_cell[   27281] = 32'h990168bd;
    ram_cell[   27282] = 32'hf29307ab;
    ram_cell[   27283] = 32'hebc6f29b;
    ram_cell[   27284] = 32'h756bfad6;
    ram_cell[   27285] = 32'h4264b4d7;
    ram_cell[   27286] = 32'hef83a2b0;
    ram_cell[   27287] = 32'ha33dfdc1;
    ram_cell[   27288] = 32'hafbee80c;
    ram_cell[   27289] = 32'h23829063;
    ram_cell[   27290] = 32'h901f949a;
    ram_cell[   27291] = 32'h9c975074;
    ram_cell[   27292] = 32'h308f7d42;
    ram_cell[   27293] = 32'h557b5546;
    ram_cell[   27294] = 32'h8fb94eb5;
    ram_cell[   27295] = 32'hf5f8ce0d;
    ram_cell[   27296] = 32'h959e6a96;
    ram_cell[   27297] = 32'h05410b5f;
    ram_cell[   27298] = 32'h260a3a93;
    ram_cell[   27299] = 32'hd7f553ed;
    ram_cell[   27300] = 32'h78aa8d0a;
    ram_cell[   27301] = 32'hc957bcd5;
    ram_cell[   27302] = 32'h9bc0169a;
    ram_cell[   27303] = 32'h581e0a40;
    ram_cell[   27304] = 32'hffb36b6a;
    ram_cell[   27305] = 32'h1fb3a573;
    ram_cell[   27306] = 32'ha708af54;
    ram_cell[   27307] = 32'h1acfa8a6;
    ram_cell[   27308] = 32'hf0d5fff0;
    ram_cell[   27309] = 32'h51cd04cd;
    ram_cell[   27310] = 32'hb6eba68a;
    ram_cell[   27311] = 32'h85e4a757;
    ram_cell[   27312] = 32'h518ef049;
    ram_cell[   27313] = 32'hfc02e43b;
    ram_cell[   27314] = 32'h64c0a606;
    ram_cell[   27315] = 32'h30efa065;
    ram_cell[   27316] = 32'h2c267c9c;
    ram_cell[   27317] = 32'h1f93d5c8;
    ram_cell[   27318] = 32'h7a050697;
    ram_cell[   27319] = 32'hd3094a9b;
    ram_cell[   27320] = 32'h1fcbc5ca;
    ram_cell[   27321] = 32'hff3bbd47;
    ram_cell[   27322] = 32'he0b7a4a2;
    ram_cell[   27323] = 32'h45b0fed5;
    ram_cell[   27324] = 32'h31936365;
    ram_cell[   27325] = 32'hb0d53f0c;
    ram_cell[   27326] = 32'he452ee4b;
    ram_cell[   27327] = 32'h774929ef;
    ram_cell[   27328] = 32'hae2c60d2;
    ram_cell[   27329] = 32'hab92fed3;
    ram_cell[   27330] = 32'ha2f03409;
    ram_cell[   27331] = 32'h13c17a08;
    ram_cell[   27332] = 32'hc867db1c;
    ram_cell[   27333] = 32'h9370a8c3;
    ram_cell[   27334] = 32'hc91c2d55;
    ram_cell[   27335] = 32'hb0b90847;
    ram_cell[   27336] = 32'h25658b09;
    ram_cell[   27337] = 32'hc323dce0;
    ram_cell[   27338] = 32'hdfd9c006;
    ram_cell[   27339] = 32'h2809d2ee;
    ram_cell[   27340] = 32'hcbbef7e5;
    ram_cell[   27341] = 32'hff3d7035;
    ram_cell[   27342] = 32'h1dd575f5;
    ram_cell[   27343] = 32'hcccc22b3;
    ram_cell[   27344] = 32'ha5edf54d;
    ram_cell[   27345] = 32'h6d30dbd7;
    ram_cell[   27346] = 32'h6d94ba57;
    ram_cell[   27347] = 32'hbf63e153;
    ram_cell[   27348] = 32'hac1f7def;
    ram_cell[   27349] = 32'h2aa551ea;
    ram_cell[   27350] = 32'h2baebd18;
    ram_cell[   27351] = 32'h2c3eb2be;
    ram_cell[   27352] = 32'he861d1fb;
    ram_cell[   27353] = 32'hcef0942f;
    ram_cell[   27354] = 32'h7d258084;
    ram_cell[   27355] = 32'hbc3f8c89;
    ram_cell[   27356] = 32'h4286b2c9;
    ram_cell[   27357] = 32'h15645431;
    ram_cell[   27358] = 32'h461b0e4e;
    ram_cell[   27359] = 32'h314b53f1;
    ram_cell[   27360] = 32'h3dd02231;
    ram_cell[   27361] = 32'hb1efd7b7;
    ram_cell[   27362] = 32'h15c44497;
    ram_cell[   27363] = 32'h6bb643f9;
    ram_cell[   27364] = 32'h65d55876;
    ram_cell[   27365] = 32'hdb08b151;
    ram_cell[   27366] = 32'hb9b47bb1;
    ram_cell[   27367] = 32'h8e3dcd3d;
    ram_cell[   27368] = 32'he66ed08f;
    ram_cell[   27369] = 32'haff71ee9;
    ram_cell[   27370] = 32'hb49cb443;
    ram_cell[   27371] = 32'hbc13d6b5;
    ram_cell[   27372] = 32'h6e4c60dc;
    ram_cell[   27373] = 32'h3b8f1372;
    ram_cell[   27374] = 32'h3247c00c;
    ram_cell[   27375] = 32'h0da664da;
    ram_cell[   27376] = 32'hadad1665;
    ram_cell[   27377] = 32'h8b8fe3e7;
    ram_cell[   27378] = 32'h40448fe0;
    ram_cell[   27379] = 32'h113b862d;
    ram_cell[   27380] = 32'hbbef8aea;
    ram_cell[   27381] = 32'hd9bf6411;
    ram_cell[   27382] = 32'hda800c00;
    ram_cell[   27383] = 32'hf7649c22;
    ram_cell[   27384] = 32'h9099cf11;
    ram_cell[   27385] = 32'h2823183f;
    ram_cell[   27386] = 32'hf881040a;
    ram_cell[   27387] = 32'he81d857f;
    ram_cell[   27388] = 32'he537ae81;
    ram_cell[   27389] = 32'h66898962;
    ram_cell[   27390] = 32'h051e5e83;
    ram_cell[   27391] = 32'he5663fbe;
    ram_cell[   27392] = 32'h84c583bf;
    ram_cell[   27393] = 32'hc9d33792;
    ram_cell[   27394] = 32'h4d4b1277;
    ram_cell[   27395] = 32'h92a945b2;
    ram_cell[   27396] = 32'h0a1674f7;
    ram_cell[   27397] = 32'h6df6f142;
    ram_cell[   27398] = 32'h58dfce73;
    ram_cell[   27399] = 32'h67d338a1;
    ram_cell[   27400] = 32'he36f6fa2;
    ram_cell[   27401] = 32'ha61f9170;
    ram_cell[   27402] = 32'h16635a5d;
    ram_cell[   27403] = 32'h949d4fdb;
    ram_cell[   27404] = 32'h3a938078;
    ram_cell[   27405] = 32'hb93a220c;
    ram_cell[   27406] = 32'h73e12bf3;
    ram_cell[   27407] = 32'h1b116f3f;
    ram_cell[   27408] = 32'he07225e5;
    ram_cell[   27409] = 32'h4c758416;
    ram_cell[   27410] = 32'h376e1734;
    ram_cell[   27411] = 32'had286e51;
    ram_cell[   27412] = 32'hf6844924;
    ram_cell[   27413] = 32'h85858ca2;
    ram_cell[   27414] = 32'h6fa7be67;
    ram_cell[   27415] = 32'h156f15e1;
    ram_cell[   27416] = 32'h1203e2c3;
    ram_cell[   27417] = 32'h26559188;
    ram_cell[   27418] = 32'h741881ad;
    ram_cell[   27419] = 32'h23b2978d;
    ram_cell[   27420] = 32'habb50d3a;
    ram_cell[   27421] = 32'h5fe1ae30;
    ram_cell[   27422] = 32'h835032ad;
    ram_cell[   27423] = 32'h587490c2;
    ram_cell[   27424] = 32'hcef9fdf6;
    ram_cell[   27425] = 32'h94f46e6c;
    ram_cell[   27426] = 32'hc2c09c66;
    ram_cell[   27427] = 32'h2be8afef;
    ram_cell[   27428] = 32'h451b38cb;
    ram_cell[   27429] = 32'hc055bb15;
    ram_cell[   27430] = 32'h01cfa4f1;
    ram_cell[   27431] = 32'h3d9cfde6;
    ram_cell[   27432] = 32'h6be7bfbe;
    ram_cell[   27433] = 32'h6885e9aa;
    ram_cell[   27434] = 32'h23dfa9a1;
    ram_cell[   27435] = 32'h252a3c22;
    ram_cell[   27436] = 32'hb85fa737;
    ram_cell[   27437] = 32'h546fc3dd;
    ram_cell[   27438] = 32'h0523074a;
    ram_cell[   27439] = 32'h6871ccd1;
    ram_cell[   27440] = 32'hc2366a82;
    ram_cell[   27441] = 32'h784582d5;
    ram_cell[   27442] = 32'h005eecf5;
    ram_cell[   27443] = 32'h8bb15605;
    ram_cell[   27444] = 32'h205ecb03;
    ram_cell[   27445] = 32'h87e0b6da;
    ram_cell[   27446] = 32'h0fe1f014;
    ram_cell[   27447] = 32'hdaf63467;
    ram_cell[   27448] = 32'h5c76a11a;
    ram_cell[   27449] = 32'hec69ffc7;
    ram_cell[   27450] = 32'h72e628db;
    ram_cell[   27451] = 32'h3fa6cb04;
    ram_cell[   27452] = 32'h922ef838;
    ram_cell[   27453] = 32'hdd2258de;
    ram_cell[   27454] = 32'hcb7563d5;
    ram_cell[   27455] = 32'hf7241676;
    ram_cell[   27456] = 32'h5bb4e522;
    ram_cell[   27457] = 32'h66513dd1;
    ram_cell[   27458] = 32'h82fafa8c;
    ram_cell[   27459] = 32'h193628d9;
    ram_cell[   27460] = 32'he730cb50;
    ram_cell[   27461] = 32'heb99690f;
    ram_cell[   27462] = 32'hf8f797f5;
    ram_cell[   27463] = 32'h94415c9c;
    ram_cell[   27464] = 32'hd90539d4;
    ram_cell[   27465] = 32'h2d0c74ee;
    ram_cell[   27466] = 32'h9f9741e6;
    ram_cell[   27467] = 32'h6281f2fd;
    ram_cell[   27468] = 32'h24b0df4f;
    ram_cell[   27469] = 32'h7c32e77f;
    ram_cell[   27470] = 32'hfb1e9de6;
    ram_cell[   27471] = 32'hd4f173fe;
    ram_cell[   27472] = 32'h21accf5c;
    ram_cell[   27473] = 32'h450ca7fe;
    ram_cell[   27474] = 32'h94e7b2ac;
    ram_cell[   27475] = 32'hca596b12;
    ram_cell[   27476] = 32'h7d775670;
    ram_cell[   27477] = 32'h58df6b99;
    ram_cell[   27478] = 32'h55ce7667;
    ram_cell[   27479] = 32'h4e2a7b18;
    ram_cell[   27480] = 32'h06379cde;
    ram_cell[   27481] = 32'h768c9e50;
    ram_cell[   27482] = 32'he928d678;
    ram_cell[   27483] = 32'h2b2e181d;
    ram_cell[   27484] = 32'h465029cf;
    ram_cell[   27485] = 32'h6ddae159;
    ram_cell[   27486] = 32'h11fde3ed;
    ram_cell[   27487] = 32'h7e8947a1;
    ram_cell[   27488] = 32'hbf195d52;
    ram_cell[   27489] = 32'h547779a2;
    ram_cell[   27490] = 32'h43fb13ed;
    ram_cell[   27491] = 32'h1f94777b;
    ram_cell[   27492] = 32'h928211ab;
    ram_cell[   27493] = 32'h58d583c7;
    ram_cell[   27494] = 32'h338b5984;
    ram_cell[   27495] = 32'he3e21a67;
    ram_cell[   27496] = 32'hf4ce8117;
    ram_cell[   27497] = 32'h19a64119;
    ram_cell[   27498] = 32'h6417abb2;
    ram_cell[   27499] = 32'h7bf99419;
    ram_cell[   27500] = 32'h7bf1b385;
    ram_cell[   27501] = 32'h4ee58d13;
    ram_cell[   27502] = 32'h067c3d0c;
    ram_cell[   27503] = 32'h397b83d0;
    ram_cell[   27504] = 32'h0e26e496;
    ram_cell[   27505] = 32'h5c587ced;
    ram_cell[   27506] = 32'h769fc057;
    ram_cell[   27507] = 32'h106d4aeb;
    ram_cell[   27508] = 32'ha8c385c3;
    ram_cell[   27509] = 32'h2fd978db;
    ram_cell[   27510] = 32'h6e9acec3;
    ram_cell[   27511] = 32'hc12e7bcf;
    ram_cell[   27512] = 32'h5d861dbe;
    ram_cell[   27513] = 32'hf75208de;
    ram_cell[   27514] = 32'h5694ed71;
    ram_cell[   27515] = 32'hb9f44c61;
    ram_cell[   27516] = 32'hbdf960a7;
    ram_cell[   27517] = 32'hf11509c9;
    ram_cell[   27518] = 32'h33f67cb9;
    ram_cell[   27519] = 32'h1fb1d818;
    ram_cell[   27520] = 32'hf6f2f873;
    ram_cell[   27521] = 32'he009d15b;
    ram_cell[   27522] = 32'h64a12ffc;
    ram_cell[   27523] = 32'hf710d85e;
    ram_cell[   27524] = 32'hae05c30f;
    ram_cell[   27525] = 32'h8140ef94;
    ram_cell[   27526] = 32'he81e1cd8;
    ram_cell[   27527] = 32'hb4626e52;
    ram_cell[   27528] = 32'h31c125f6;
    ram_cell[   27529] = 32'h9e522381;
    ram_cell[   27530] = 32'hc8f48bc2;
    ram_cell[   27531] = 32'h58cf68ba;
    ram_cell[   27532] = 32'hc69a15c8;
    ram_cell[   27533] = 32'h2041589e;
    ram_cell[   27534] = 32'h20240989;
    ram_cell[   27535] = 32'hd4d7b8cf;
    ram_cell[   27536] = 32'h93f4d46f;
    ram_cell[   27537] = 32'hc327334e;
    ram_cell[   27538] = 32'h6d66ab4b;
    ram_cell[   27539] = 32'hda4c54a0;
    ram_cell[   27540] = 32'hfe9e35b1;
    ram_cell[   27541] = 32'he288bc1f;
    ram_cell[   27542] = 32'hede7c0d4;
    ram_cell[   27543] = 32'hd7e9bf18;
    ram_cell[   27544] = 32'h381c369b;
    ram_cell[   27545] = 32'h2b7dbe49;
    ram_cell[   27546] = 32'hdf77a092;
    ram_cell[   27547] = 32'h51754bec;
    ram_cell[   27548] = 32'h9c6a92ac;
    ram_cell[   27549] = 32'h8f70cbff;
    ram_cell[   27550] = 32'h9c6518c0;
    ram_cell[   27551] = 32'hedfa1984;
    ram_cell[   27552] = 32'h0777fd91;
    ram_cell[   27553] = 32'h851b973b;
    ram_cell[   27554] = 32'he8b7aea6;
    ram_cell[   27555] = 32'hdcd3623b;
    ram_cell[   27556] = 32'h7decc047;
    ram_cell[   27557] = 32'hddb9b96c;
    ram_cell[   27558] = 32'h4c237169;
    ram_cell[   27559] = 32'hcbbaa168;
    ram_cell[   27560] = 32'hc954e501;
    ram_cell[   27561] = 32'h020692ef;
    ram_cell[   27562] = 32'hae6851ec;
    ram_cell[   27563] = 32'h4d875239;
    ram_cell[   27564] = 32'h8aaf1657;
    ram_cell[   27565] = 32'he75ace24;
    ram_cell[   27566] = 32'h52eef99e;
    ram_cell[   27567] = 32'ha776265e;
    ram_cell[   27568] = 32'h1930eefb;
    ram_cell[   27569] = 32'h1785a014;
    ram_cell[   27570] = 32'h652fe9ac;
    ram_cell[   27571] = 32'hb144f546;
    ram_cell[   27572] = 32'hb5b8b9c5;
    ram_cell[   27573] = 32'h3090d832;
    ram_cell[   27574] = 32'hc6b0057f;
    ram_cell[   27575] = 32'h76ad8499;
    ram_cell[   27576] = 32'h5216c223;
    ram_cell[   27577] = 32'h98e2261f;
    ram_cell[   27578] = 32'hf6945a15;
    ram_cell[   27579] = 32'heba30fc7;
    ram_cell[   27580] = 32'he8acc580;
    ram_cell[   27581] = 32'h1dc86468;
    ram_cell[   27582] = 32'h2034891b;
    ram_cell[   27583] = 32'hb1d87f3b;
    ram_cell[   27584] = 32'hb6b30208;
    ram_cell[   27585] = 32'heb6a678d;
    ram_cell[   27586] = 32'h443d2aaf;
    ram_cell[   27587] = 32'h1d6743dd;
    ram_cell[   27588] = 32'h0a1126a2;
    ram_cell[   27589] = 32'h54de3322;
    ram_cell[   27590] = 32'h72fc0dfc;
    ram_cell[   27591] = 32'h6aee7950;
    ram_cell[   27592] = 32'h1cd39dfb;
    ram_cell[   27593] = 32'h8a1a0b93;
    ram_cell[   27594] = 32'ha4d06002;
    ram_cell[   27595] = 32'ha909535d;
    ram_cell[   27596] = 32'h243e3e25;
    ram_cell[   27597] = 32'hd5320d8c;
    ram_cell[   27598] = 32'h65a47480;
    ram_cell[   27599] = 32'h6eb65872;
    ram_cell[   27600] = 32'h9b4191f6;
    ram_cell[   27601] = 32'hee195e5f;
    ram_cell[   27602] = 32'h0925c126;
    ram_cell[   27603] = 32'h05ff5abf;
    ram_cell[   27604] = 32'h13b76448;
    ram_cell[   27605] = 32'h6da65b6b;
    ram_cell[   27606] = 32'h8052e0e1;
    ram_cell[   27607] = 32'hdb8ea188;
    ram_cell[   27608] = 32'ha894cb69;
    ram_cell[   27609] = 32'h118122cb;
    ram_cell[   27610] = 32'hbc2f237e;
    ram_cell[   27611] = 32'hf8cea9c6;
    ram_cell[   27612] = 32'hf67d3433;
    ram_cell[   27613] = 32'h76d1cf3e;
    ram_cell[   27614] = 32'hc4d7cf5c;
    ram_cell[   27615] = 32'hdf873d92;
    ram_cell[   27616] = 32'ha85dcbe1;
    ram_cell[   27617] = 32'hcfe3a03a;
    ram_cell[   27618] = 32'h2abe9d45;
    ram_cell[   27619] = 32'h6a797e85;
    ram_cell[   27620] = 32'h36683cdb;
    ram_cell[   27621] = 32'h69abe5c9;
    ram_cell[   27622] = 32'h8ba0591f;
    ram_cell[   27623] = 32'hfe5f6fc6;
    ram_cell[   27624] = 32'h752a16e6;
    ram_cell[   27625] = 32'hdf0e6ba4;
    ram_cell[   27626] = 32'hbf11bc6a;
    ram_cell[   27627] = 32'he0bafe8d;
    ram_cell[   27628] = 32'h1147ff00;
    ram_cell[   27629] = 32'hd1f6cfca;
    ram_cell[   27630] = 32'h2c562197;
    ram_cell[   27631] = 32'h8f24bbd7;
    ram_cell[   27632] = 32'h7c47899b;
    ram_cell[   27633] = 32'hbadf5609;
    ram_cell[   27634] = 32'he4ff3857;
    ram_cell[   27635] = 32'hb50a93ea;
    ram_cell[   27636] = 32'h4c09c942;
    ram_cell[   27637] = 32'h97be2f57;
    ram_cell[   27638] = 32'h550031b8;
    ram_cell[   27639] = 32'hf2f53780;
    ram_cell[   27640] = 32'h5e8b8a66;
    ram_cell[   27641] = 32'h070e65da;
    ram_cell[   27642] = 32'h6de30a5b;
    ram_cell[   27643] = 32'hd386b685;
    ram_cell[   27644] = 32'h4f8e29bd;
    ram_cell[   27645] = 32'he12812fc;
    ram_cell[   27646] = 32'h0112b0e6;
    ram_cell[   27647] = 32'h77c17126;
    ram_cell[   27648] = 32'h285b8ab0;
    ram_cell[   27649] = 32'h764beaa8;
    ram_cell[   27650] = 32'h1244c671;
    ram_cell[   27651] = 32'h57ac79b4;
    ram_cell[   27652] = 32'hea824175;
    ram_cell[   27653] = 32'hea258bcc;
    ram_cell[   27654] = 32'h11fc0b2f;
    ram_cell[   27655] = 32'h060d7894;
    ram_cell[   27656] = 32'h65752e67;
    ram_cell[   27657] = 32'h172a64ac;
    ram_cell[   27658] = 32'h302ce545;
    ram_cell[   27659] = 32'h6d63d002;
    ram_cell[   27660] = 32'h9553b47f;
    ram_cell[   27661] = 32'hdb3203a1;
    ram_cell[   27662] = 32'h1f317d61;
    ram_cell[   27663] = 32'h584b8460;
    ram_cell[   27664] = 32'hd7e817ba;
    ram_cell[   27665] = 32'h0973e938;
    ram_cell[   27666] = 32'h51b67472;
    ram_cell[   27667] = 32'h339acc03;
    ram_cell[   27668] = 32'h09427839;
    ram_cell[   27669] = 32'h4a7312a5;
    ram_cell[   27670] = 32'hcb929de5;
    ram_cell[   27671] = 32'hd8508baf;
    ram_cell[   27672] = 32'ha53b65f2;
    ram_cell[   27673] = 32'haae00cf0;
    ram_cell[   27674] = 32'h8cc4ea75;
    ram_cell[   27675] = 32'h4c960df1;
    ram_cell[   27676] = 32'he4d5b857;
    ram_cell[   27677] = 32'ha4d3679f;
    ram_cell[   27678] = 32'h89b59105;
    ram_cell[   27679] = 32'h227a1829;
    ram_cell[   27680] = 32'h8b98cf8f;
    ram_cell[   27681] = 32'h04850c30;
    ram_cell[   27682] = 32'hb0c82097;
    ram_cell[   27683] = 32'ha1a12e09;
    ram_cell[   27684] = 32'h7ce7545a;
    ram_cell[   27685] = 32'h604d6835;
    ram_cell[   27686] = 32'h195b5677;
    ram_cell[   27687] = 32'h251c93e3;
    ram_cell[   27688] = 32'hc22c12a3;
    ram_cell[   27689] = 32'hdb09282b;
    ram_cell[   27690] = 32'h68429fb5;
    ram_cell[   27691] = 32'h66f019fa;
    ram_cell[   27692] = 32'hb058a537;
    ram_cell[   27693] = 32'h87e7528f;
    ram_cell[   27694] = 32'h7f95608c;
    ram_cell[   27695] = 32'hf3699028;
    ram_cell[   27696] = 32'h2aa12f30;
    ram_cell[   27697] = 32'h8630e29f;
    ram_cell[   27698] = 32'h57ddcadf;
    ram_cell[   27699] = 32'h5cc52624;
    ram_cell[   27700] = 32'hfb97b1b2;
    ram_cell[   27701] = 32'hdb5122f7;
    ram_cell[   27702] = 32'h361cf944;
    ram_cell[   27703] = 32'ha5044723;
    ram_cell[   27704] = 32'h987aa3c5;
    ram_cell[   27705] = 32'hcc8d9fcd;
    ram_cell[   27706] = 32'hab9b13b8;
    ram_cell[   27707] = 32'he2c1c2ec;
    ram_cell[   27708] = 32'h745a4d42;
    ram_cell[   27709] = 32'hbe2d8641;
    ram_cell[   27710] = 32'h93515b24;
    ram_cell[   27711] = 32'h48caeb15;
    ram_cell[   27712] = 32'h225b4a63;
    ram_cell[   27713] = 32'hd6a153b3;
    ram_cell[   27714] = 32'he9472464;
    ram_cell[   27715] = 32'haff576cc;
    ram_cell[   27716] = 32'h036f6087;
    ram_cell[   27717] = 32'hf2452ccf;
    ram_cell[   27718] = 32'he62a027c;
    ram_cell[   27719] = 32'h2fe23bcd;
    ram_cell[   27720] = 32'h05bbf30f;
    ram_cell[   27721] = 32'h14a70874;
    ram_cell[   27722] = 32'hdb85d233;
    ram_cell[   27723] = 32'hada4ae8c;
    ram_cell[   27724] = 32'h1ceeb2e6;
    ram_cell[   27725] = 32'haa23d6a0;
    ram_cell[   27726] = 32'h907591e9;
    ram_cell[   27727] = 32'hef9b5784;
    ram_cell[   27728] = 32'h0a748eb9;
    ram_cell[   27729] = 32'h98fd0ee4;
    ram_cell[   27730] = 32'he56f312d;
    ram_cell[   27731] = 32'hd8ffd789;
    ram_cell[   27732] = 32'h6e88e71f;
    ram_cell[   27733] = 32'h0a141746;
    ram_cell[   27734] = 32'h41b637ca;
    ram_cell[   27735] = 32'hc24563a2;
    ram_cell[   27736] = 32'hdeb62299;
    ram_cell[   27737] = 32'h5150891c;
    ram_cell[   27738] = 32'hb6f74f99;
    ram_cell[   27739] = 32'hede1848b;
    ram_cell[   27740] = 32'h418e409e;
    ram_cell[   27741] = 32'h5dcd5548;
    ram_cell[   27742] = 32'hfc7967c3;
    ram_cell[   27743] = 32'h47d7381a;
    ram_cell[   27744] = 32'h312cc117;
    ram_cell[   27745] = 32'h379724c2;
    ram_cell[   27746] = 32'h717e8c71;
    ram_cell[   27747] = 32'hf02a333b;
    ram_cell[   27748] = 32'h13d6085f;
    ram_cell[   27749] = 32'h2955ee17;
    ram_cell[   27750] = 32'h0f9c5af3;
    ram_cell[   27751] = 32'h6deaf705;
    ram_cell[   27752] = 32'hb8df6aa2;
    ram_cell[   27753] = 32'ha2c2f402;
    ram_cell[   27754] = 32'hfc1db4e7;
    ram_cell[   27755] = 32'h1e6e2039;
    ram_cell[   27756] = 32'hce5f1142;
    ram_cell[   27757] = 32'ha07608bb;
    ram_cell[   27758] = 32'h7daae026;
    ram_cell[   27759] = 32'he47842d0;
    ram_cell[   27760] = 32'h982084d5;
    ram_cell[   27761] = 32'h6cbfd429;
    ram_cell[   27762] = 32'h5c03133d;
    ram_cell[   27763] = 32'hc4ce2c11;
    ram_cell[   27764] = 32'h257398eb;
    ram_cell[   27765] = 32'hcd76c07f;
    ram_cell[   27766] = 32'heb396449;
    ram_cell[   27767] = 32'hd68053f3;
    ram_cell[   27768] = 32'hf2f8e88a;
    ram_cell[   27769] = 32'h67229578;
    ram_cell[   27770] = 32'hcc7152f0;
    ram_cell[   27771] = 32'h0b278b02;
    ram_cell[   27772] = 32'hda3d5eb3;
    ram_cell[   27773] = 32'hdf939dba;
    ram_cell[   27774] = 32'hbfadba32;
    ram_cell[   27775] = 32'h639e07b0;
    ram_cell[   27776] = 32'h5281be2d;
    ram_cell[   27777] = 32'h4405a05c;
    ram_cell[   27778] = 32'h443e6044;
    ram_cell[   27779] = 32'h037f35a5;
    ram_cell[   27780] = 32'h05efa287;
    ram_cell[   27781] = 32'h6af18646;
    ram_cell[   27782] = 32'h2ee2795d;
    ram_cell[   27783] = 32'hd54ff72c;
    ram_cell[   27784] = 32'h856b17de;
    ram_cell[   27785] = 32'h2d9dfbad;
    ram_cell[   27786] = 32'h7cb62f5f;
    ram_cell[   27787] = 32'hecd65d0d;
    ram_cell[   27788] = 32'h6a5833e4;
    ram_cell[   27789] = 32'he3c7af69;
    ram_cell[   27790] = 32'h219e20e1;
    ram_cell[   27791] = 32'h3ddaf825;
    ram_cell[   27792] = 32'h22af00a3;
    ram_cell[   27793] = 32'h238b5bfe;
    ram_cell[   27794] = 32'hc82128e7;
    ram_cell[   27795] = 32'h172f31fc;
    ram_cell[   27796] = 32'h6a19f585;
    ram_cell[   27797] = 32'h0c66429d;
    ram_cell[   27798] = 32'hb26382a7;
    ram_cell[   27799] = 32'h601a99cd;
    ram_cell[   27800] = 32'heba7cc85;
    ram_cell[   27801] = 32'hda014502;
    ram_cell[   27802] = 32'he1e8f8a6;
    ram_cell[   27803] = 32'hdfffdd76;
    ram_cell[   27804] = 32'hf52949ac;
    ram_cell[   27805] = 32'h564b3bf8;
    ram_cell[   27806] = 32'h44cf9bca;
    ram_cell[   27807] = 32'hf15839fd;
    ram_cell[   27808] = 32'hdaddea4b;
    ram_cell[   27809] = 32'he25123b2;
    ram_cell[   27810] = 32'h6220cd63;
    ram_cell[   27811] = 32'h47b770a1;
    ram_cell[   27812] = 32'h57d1e0ae;
    ram_cell[   27813] = 32'hdb1bb13e;
    ram_cell[   27814] = 32'hc46fa78c;
    ram_cell[   27815] = 32'h77808f70;
    ram_cell[   27816] = 32'h5984fb54;
    ram_cell[   27817] = 32'ha54acabf;
    ram_cell[   27818] = 32'h52cff5d7;
    ram_cell[   27819] = 32'h2727bf14;
    ram_cell[   27820] = 32'he4af5d23;
    ram_cell[   27821] = 32'hf9e5f53c;
    ram_cell[   27822] = 32'hf9ee1e94;
    ram_cell[   27823] = 32'hcd4de527;
    ram_cell[   27824] = 32'hc48a57f3;
    ram_cell[   27825] = 32'ha107d17d;
    ram_cell[   27826] = 32'hd2b7ac14;
    ram_cell[   27827] = 32'h0aba5bf2;
    ram_cell[   27828] = 32'hbf7c4b49;
    ram_cell[   27829] = 32'h74acdfa8;
    ram_cell[   27830] = 32'h7b49f639;
    ram_cell[   27831] = 32'h69dbe3a4;
    ram_cell[   27832] = 32'h8bf957b9;
    ram_cell[   27833] = 32'h2cc3ae1b;
    ram_cell[   27834] = 32'h7b495e08;
    ram_cell[   27835] = 32'hf984b3f8;
    ram_cell[   27836] = 32'hac26be3a;
    ram_cell[   27837] = 32'h6225fec0;
    ram_cell[   27838] = 32'hc84fcd1e;
    ram_cell[   27839] = 32'h285ea627;
    ram_cell[   27840] = 32'hef430b1f;
    ram_cell[   27841] = 32'he423c163;
    ram_cell[   27842] = 32'h94391263;
    ram_cell[   27843] = 32'h746829a7;
    ram_cell[   27844] = 32'h95a3ba41;
    ram_cell[   27845] = 32'h7927da8a;
    ram_cell[   27846] = 32'hef123363;
    ram_cell[   27847] = 32'hb8beef3b;
    ram_cell[   27848] = 32'h567e4b48;
    ram_cell[   27849] = 32'hc74e3655;
    ram_cell[   27850] = 32'hf10807d1;
    ram_cell[   27851] = 32'hf9850636;
    ram_cell[   27852] = 32'hebd6ac17;
    ram_cell[   27853] = 32'hc834a6c6;
    ram_cell[   27854] = 32'h09ae267d;
    ram_cell[   27855] = 32'h3025989e;
    ram_cell[   27856] = 32'h8cd224b1;
    ram_cell[   27857] = 32'h1b82b9eb;
    ram_cell[   27858] = 32'h3317328a;
    ram_cell[   27859] = 32'h93963b4f;
    ram_cell[   27860] = 32'h8f85d52b;
    ram_cell[   27861] = 32'hb0d5cf96;
    ram_cell[   27862] = 32'hadae6311;
    ram_cell[   27863] = 32'h61ecf933;
    ram_cell[   27864] = 32'hfa0ba8c8;
    ram_cell[   27865] = 32'h2fb4b7de;
    ram_cell[   27866] = 32'hf8162e6f;
    ram_cell[   27867] = 32'h9eb47c96;
    ram_cell[   27868] = 32'hd8a277f5;
    ram_cell[   27869] = 32'hacaf3a30;
    ram_cell[   27870] = 32'h956ab02e;
    ram_cell[   27871] = 32'hde945a84;
    ram_cell[   27872] = 32'h84652c79;
    ram_cell[   27873] = 32'hd77504a9;
    ram_cell[   27874] = 32'h729d7a4d;
    ram_cell[   27875] = 32'h33631acb;
    ram_cell[   27876] = 32'h9d59eaab;
    ram_cell[   27877] = 32'hdc5cdb93;
    ram_cell[   27878] = 32'ha80de6e6;
    ram_cell[   27879] = 32'h82995542;
    ram_cell[   27880] = 32'h2cba371f;
    ram_cell[   27881] = 32'h568627ca;
    ram_cell[   27882] = 32'h7e7c6f82;
    ram_cell[   27883] = 32'h0ce3795f;
    ram_cell[   27884] = 32'h607cbaee;
    ram_cell[   27885] = 32'hb655088d;
    ram_cell[   27886] = 32'h26e92fb7;
    ram_cell[   27887] = 32'hd16a24f1;
    ram_cell[   27888] = 32'h6a0ce398;
    ram_cell[   27889] = 32'hd1f1a24a;
    ram_cell[   27890] = 32'hf383d03a;
    ram_cell[   27891] = 32'hce9d9e41;
    ram_cell[   27892] = 32'h7c54ded6;
    ram_cell[   27893] = 32'ha98115fc;
    ram_cell[   27894] = 32'h669e91ea;
    ram_cell[   27895] = 32'h1afed280;
    ram_cell[   27896] = 32'h9372f7e5;
    ram_cell[   27897] = 32'hd035fac9;
    ram_cell[   27898] = 32'hff1e4c28;
    ram_cell[   27899] = 32'h7f3447b9;
    ram_cell[   27900] = 32'h749a6861;
    ram_cell[   27901] = 32'h79c4d33e;
    ram_cell[   27902] = 32'h5bc40f54;
    ram_cell[   27903] = 32'h03adec7a;
    ram_cell[   27904] = 32'h8b519baf;
    ram_cell[   27905] = 32'hb1c0ff97;
    ram_cell[   27906] = 32'hd7ca2e18;
    ram_cell[   27907] = 32'h8b7a6e73;
    ram_cell[   27908] = 32'hc8420b91;
    ram_cell[   27909] = 32'h62e126af;
    ram_cell[   27910] = 32'h9cff87a6;
    ram_cell[   27911] = 32'hd0d5ea44;
    ram_cell[   27912] = 32'h0a38c6c7;
    ram_cell[   27913] = 32'hf12598f7;
    ram_cell[   27914] = 32'hc1545e13;
    ram_cell[   27915] = 32'hde3f98ec;
    ram_cell[   27916] = 32'h030d5e67;
    ram_cell[   27917] = 32'hc5e4b410;
    ram_cell[   27918] = 32'h789194f4;
    ram_cell[   27919] = 32'h55be1f59;
    ram_cell[   27920] = 32'h0b87b0fd;
    ram_cell[   27921] = 32'h0ceb55df;
    ram_cell[   27922] = 32'h283b604c;
    ram_cell[   27923] = 32'h72ef25a0;
    ram_cell[   27924] = 32'hf5945358;
    ram_cell[   27925] = 32'h17aec20b;
    ram_cell[   27926] = 32'hf113f052;
    ram_cell[   27927] = 32'he2151c7b;
    ram_cell[   27928] = 32'hfd01f053;
    ram_cell[   27929] = 32'h2ac297d4;
    ram_cell[   27930] = 32'hc24e34d2;
    ram_cell[   27931] = 32'h6f660251;
    ram_cell[   27932] = 32'h2d68bf4e;
    ram_cell[   27933] = 32'h344c7090;
    ram_cell[   27934] = 32'hb9de946f;
    ram_cell[   27935] = 32'h3ef63a3c;
    ram_cell[   27936] = 32'h6d08dd07;
    ram_cell[   27937] = 32'h77725e76;
    ram_cell[   27938] = 32'hc7999e2c;
    ram_cell[   27939] = 32'h3e41870a;
    ram_cell[   27940] = 32'hf94f3009;
    ram_cell[   27941] = 32'h3c897292;
    ram_cell[   27942] = 32'hadab78b4;
    ram_cell[   27943] = 32'haa5e26ea;
    ram_cell[   27944] = 32'h2bce5129;
    ram_cell[   27945] = 32'h8acb6698;
    ram_cell[   27946] = 32'h13df0e56;
    ram_cell[   27947] = 32'h49aeb7dd;
    ram_cell[   27948] = 32'h544ad152;
    ram_cell[   27949] = 32'h7d07fac8;
    ram_cell[   27950] = 32'hc1ee81fb;
    ram_cell[   27951] = 32'hd569241a;
    ram_cell[   27952] = 32'h6aaa406c;
    ram_cell[   27953] = 32'h41f122dd;
    ram_cell[   27954] = 32'h2453c211;
    ram_cell[   27955] = 32'ha10d8b4a;
    ram_cell[   27956] = 32'hdc572eb1;
    ram_cell[   27957] = 32'h7cc647b7;
    ram_cell[   27958] = 32'hd0f92a81;
    ram_cell[   27959] = 32'h967ab913;
    ram_cell[   27960] = 32'h2e17de3d;
    ram_cell[   27961] = 32'h5ba52117;
    ram_cell[   27962] = 32'h7322ed47;
    ram_cell[   27963] = 32'h37e73f7c;
    ram_cell[   27964] = 32'h3eb89411;
    ram_cell[   27965] = 32'h9edd2ed1;
    ram_cell[   27966] = 32'h71b48ace;
    ram_cell[   27967] = 32'h2a85221b;
    ram_cell[   27968] = 32'h65e53ccb;
    ram_cell[   27969] = 32'hacec3c31;
    ram_cell[   27970] = 32'h61dc801a;
    ram_cell[   27971] = 32'h34fb0eab;
    ram_cell[   27972] = 32'hf436303e;
    ram_cell[   27973] = 32'h4028f0ff;
    ram_cell[   27974] = 32'h743bd3d6;
    ram_cell[   27975] = 32'h7b9f9fc7;
    ram_cell[   27976] = 32'h2565c1a6;
    ram_cell[   27977] = 32'h54dd5e3f;
    ram_cell[   27978] = 32'hc55dda1c;
    ram_cell[   27979] = 32'h58ca9a90;
    ram_cell[   27980] = 32'h513850df;
    ram_cell[   27981] = 32'h07e22e4f;
    ram_cell[   27982] = 32'h899acf7b;
    ram_cell[   27983] = 32'h25d6f9bd;
    ram_cell[   27984] = 32'hc861546c;
    ram_cell[   27985] = 32'hb7aead56;
    ram_cell[   27986] = 32'he4e59bc1;
    ram_cell[   27987] = 32'hd34668b4;
    ram_cell[   27988] = 32'h7b5896cb;
    ram_cell[   27989] = 32'h4c6ae16b;
    ram_cell[   27990] = 32'hb22fb8f6;
    ram_cell[   27991] = 32'h6f49f0ed;
    ram_cell[   27992] = 32'hd77460bb;
    ram_cell[   27993] = 32'hda9401bf;
    ram_cell[   27994] = 32'hc9ba98a3;
    ram_cell[   27995] = 32'hf6988c37;
    ram_cell[   27996] = 32'h7f4c2e54;
    ram_cell[   27997] = 32'h730274bc;
    ram_cell[   27998] = 32'h323e3760;
    ram_cell[   27999] = 32'h96456fc0;
    ram_cell[   28000] = 32'h7b3317c0;
    ram_cell[   28001] = 32'had909475;
    ram_cell[   28002] = 32'h5f3ae22b;
    ram_cell[   28003] = 32'hc833469b;
    ram_cell[   28004] = 32'hf73e9aa9;
    ram_cell[   28005] = 32'h86da32e7;
    ram_cell[   28006] = 32'h355e37bc;
    ram_cell[   28007] = 32'hbdc58b4e;
    ram_cell[   28008] = 32'hd1e54ca7;
    ram_cell[   28009] = 32'he18d4f9d;
    ram_cell[   28010] = 32'h94b978d4;
    ram_cell[   28011] = 32'hba874518;
    ram_cell[   28012] = 32'h5cb01250;
    ram_cell[   28013] = 32'ha6ba3f44;
    ram_cell[   28014] = 32'hf8aaa164;
    ram_cell[   28015] = 32'ha9c57130;
    ram_cell[   28016] = 32'hc8d34346;
    ram_cell[   28017] = 32'hcc2c6c41;
    ram_cell[   28018] = 32'hdb8a0a99;
    ram_cell[   28019] = 32'h1da29e32;
    ram_cell[   28020] = 32'h5bd2c682;
    ram_cell[   28021] = 32'ha3ae085e;
    ram_cell[   28022] = 32'h4fff97fe;
    ram_cell[   28023] = 32'h29f72118;
    ram_cell[   28024] = 32'h1b6f1656;
    ram_cell[   28025] = 32'h3478bc2b;
    ram_cell[   28026] = 32'h946eca74;
    ram_cell[   28027] = 32'hbd3e8ce2;
    ram_cell[   28028] = 32'h68c5485b;
    ram_cell[   28029] = 32'h0218b0ce;
    ram_cell[   28030] = 32'he43e5cba;
    ram_cell[   28031] = 32'h7d0672c4;
    ram_cell[   28032] = 32'h81165e0d;
    ram_cell[   28033] = 32'h21becd3e;
    ram_cell[   28034] = 32'h75a599fd;
    ram_cell[   28035] = 32'h9e7b1e8a;
    ram_cell[   28036] = 32'h628e6ea5;
    ram_cell[   28037] = 32'ha7dced1a;
    ram_cell[   28038] = 32'hce7ef21d;
    ram_cell[   28039] = 32'hc273259a;
    ram_cell[   28040] = 32'h68b53c81;
    ram_cell[   28041] = 32'h0646718b;
    ram_cell[   28042] = 32'h5189a974;
    ram_cell[   28043] = 32'h8789529a;
    ram_cell[   28044] = 32'h0c005951;
    ram_cell[   28045] = 32'h33a727c8;
    ram_cell[   28046] = 32'hefb02981;
    ram_cell[   28047] = 32'h3c8b4548;
    ram_cell[   28048] = 32'h33a44ddc;
    ram_cell[   28049] = 32'hcbece90b;
    ram_cell[   28050] = 32'h83ea48d5;
    ram_cell[   28051] = 32'he3a971f4;
    ram_cell[   28052] = 32'h7ee6aad6;
    ram_cell[   28053] = 32'h15f64bf6;
    ram_cell[   28054] = 32'h29c2a503;
    ram_cell[   28055] = 32'h318af74b;
    ram_cell[   28056] = 32'h788a2664;
    ram_cell[   28057] = 32'h7ed3e563;
    ram_cell[   28058] = 32'h0516ca9e;
    ram_cell[   28059] = 32'hea5efb83;
    ram_cell[   28060] = 32'h1a7bfd1c;
    ram_cell[   28061] = 32'h99ffd501;
    ram_cell[   28062] = 32'h2fb3a95b;
    ram_cell[   28063] = 32'h52e204d1;
    ram_cell[   28064] = 32'hd433c486;
    ram_cell[   28065] = 32'h6885cc41;
    ram_cell[   28066] = 32'h9ccd0bdc;
    ram_cell[   28067] = 32'hd1c9d83d;
    ram_cell[   28068] = 32'h98f92ec4;
    ram_cell[   28069] = 32'h02e09b36;
    ram_cell[   28070] = 32'h73604d3c;
    ram_cell[   28071] = 32'h6be2181f;
    ram_cell[   28072] = 32'h35404ca3;
    ram_cell[   28073] = 32'h2cbc018e;
    ram_cell[   28074] = 32'h3d76cf4b;
    ram_cell[   28075] = 32'hc8bb1d35;
    ram_cell[   28076] = 32'h75986067;
    ram_cell[   28077] = 32'h557ff6ef;
    ram_cell[   28078] = 32'h93e650de;
    ram_cell[   28079] = 32'h2fa6eece;
    ram_cell[   28080] = 32'h32314adc;
    ram_cell[   28081] = 32'h8d6c3163;
    ram_cell[   28082] = 32'h75d1c08f;
    ram_cell[   28083] = 32'h8265f5c2;
    ram_cell[   28084] = 32'hd6d9ca4f;
    ram_cell[   28085] = 32'h2c9ebcf4;
    ram_cell[   28086] = 32'h8e5ddb0f;
    ram_cell[   28087] = 32'h2b238c36;
    ram_cell[   28088] = 32'h75c8fb9c;
    ram_cell[   28089] = 32'h4e6824b0;
    ram_cell[   28090] = 32'h10acdaba;
    ram_cell[   28091] = 32'h72f5f0e0;
    ram_cell[   28092] = 32'hc97de993;
    ram_cell[   28093] = 32'h1e6bc471;
    ram_cell[   28094] = 32'h6f2ce1d1;
    ram_cell[   28095] = 32'he7de895b;
    ram_cell[   28096] = 32'h7bf4754d;
    ram_cell[   28097] = 32'h83fc1f14;
    ram_cell[   28098] = 32'h650b6e18;
    ram_cell[   28099] = 32'h9b780a3e;
    ram_cell[   28100] = 32'hfad90fdc;
    ram_cell[   28101] = 32'h87e28267;
    ram_cell[   28102] = 32'hd4c25a3f;
    ram_cell[   28103] = 32'h4a575b92;
    ram_cell[   28104] = 32'h81a9cae5;
    ram_cell[   28105] = 32'h004d5889;
    ram_cell[   28106] = 32'ha7543d5c;
    ram_cell[   28107] = 32'h5e5043b2;
    ram_cell[   28108] = 32'h8101a211;
    ram_cell[   28109] = 32'hc07e5c0f;
    ram_cell[   28110] = 32'hca28ca9e;
    ram_cell[   28111] = 32'hd85134d2;
    ram_cell[   28112] = 32'hb2946d2a;
    ram_cell[   28113] = 32'h3c150fb0;
    ram_cell[   28114] = 32'h4b3bc992;
    ram_cell[   28115] = 32'h739d817e;
    ram_cell[   28116] = 32'h0b12d2b7;
    ram_cell[   28117] = 32'h5ae111bb;
    ram_cell[   28118] = 32'h1b608ad6;
    ram_cell[   28119] = 32'h79995455;
    ram_cell[   28120] = 32'h8113f521;
    ram_cell[   28121] = 32'h1748d695;
    ram_cell[   28122] = 32'h6fe581a0;
    ram_cell[   28123] = 32'h84d3c0c6;
    ram_cell[   28124] = 32'h125d8f80;
    ram_cell[   28125] = 32'h554819b0;
    ram_cell[   28126] = 32'hc978397b;
    ram_cell[   28127] = 32'h843d5e56;
    ram_cell[   28128] = 32'h968fcfdc;
    ram_cell[   28129] = 32'h60364324;
    ram_cell[   28130] = 32'h0c9a85da;
    ram_cell[   28131] = 32'h97313033;
    ram_cell[   28132] = 32'h4e7dbada;
    ram_cell[   28133] = 32'h09787f4e;
    ram_cell[   28134] = 32'h578af0c7;
    ram_cell[   28135] = 32'h223f4c2e;
    ram_cell[   28136] = 32'he111baf9;
    ram_cell[   28137] = 32'h679eb735;
    ram_cell[   28138] = 32'h52de9738;
    ram_cell[   28139] = 32'h5cab2923;
    ram_cell[   28140] = 32'ha8aeee75;
    ram_cell[   28141] = 32'hc71352fe;
    ram_cell[   28142] = 32'he391c355;
    ram_cell[   28143] = 32'h28c3fcbc;
    ram_cell[   28144] = 32'hdcd16e28;
    ram_cell[   28145] = 32'h5127c22b;
    ram_cell[   28146] = 32'h4cc5e7d8;
    ram_cell[   28147] = 32'h3bf62a4b;
    ram_cell[   28148] = 32'had50d442;
    ram_cell[   28149] = 32'h3c50852e;
    ram_cell[   28150] = 32'hde30403a;
    ram_cell[   28151] = 32'h596cd45e;
    ram_cell[   28152] = 32'h7ef82fc2;
    ram_cell[   28153] = 32'h3f0e5a85;
    ram_cell[   28154] = 32'h1db8d0f5;
    ram_cell[   28155] = 32'h9ced5fa8;
    ram_cell[   28156] = 32'h26efa54e;
    ram_cell[   28157] = 32'h9e972bee;
    ram_cell[   28158] = 32'h618461a4;
    ram_cell[   28159] = 32'hb67bd423;
    ram_cell[   28160] = 32'h55bf1f03;
    ram_cell[   28161] = 32'hc755e564;
    ram_cell[   28162] = 32'h6c60409f;
    ram_cell[   28163] = 32'hc34b6992;
    ram_cell[   28164] = 32'h2052c2e7;
    ram_cell[   28165] = 32'ha505eec0;
    ram_cell[   28166] = 32'h345e84c6;
    ram_cell[   28167] = 32'hc48b74af;
    ram_cell[   28168] = 32'h7186eae0;
    ram_cell[   28169] = 32'h935dd27e;
    ram_cell[   28170] = 32'h2c0facc6;
    ram_cell[   28171] = 32'h5e352e9c;
    ram_cell[   28172] = 32'hda1d849f;
    ram_cell[   28173] = 32'hd61af557;
    ram_cell[   28174] = 32'h12236883;
    ram_cell[   28175] = 32'h7e77664c;
    ram_cell[   28176] = 32'h1a9978fc;
    ram_cell[   28177] = 32'hd2d537ef;
    ram_cell[   28178] = 32'h3872f13f;
    ram_cell[   28179] = 32'hd20eda68;
    ram_cell[   28180] = 32'hdf53d008;
    ram_cell[   28181] = 32'h43fa5ad9;
    ram_cell[   28182] = 32'hd124cfdf;
    ram_cell[   28183] = 32'h44086fa5;
    ram_cell[   28184] = 32'hc01f1e42;
    ram_cell[   28185] = 32'h4f445561;
    ram_cell[   28186] = 32'hf9c4427f;
    ram_cell[   28187] = 32'h7eb1b350;
    ram_cell[   28188] = 32'h5a824cad;
    ram_cell[   28189] = 32'hefe111d1;
    ram_cell[   28190] = 32'hdf63c93d;
    ram_cell[   28191] = 32'h3ff75f7f;
    ram_cell[   28192] = 32'h1fca89cc;
    ram_cell[   28193] = 32'h37518c03;
    ram_cell[   28194] = 32'hc0ba2c23;
    ram_cell[   28195] = 32'h9f46f017;
    ram_cell[   28196] = 32'h6cd45598;
    ram_cell[   28197] = 32'h32c76618;
    ram_cell[   28198] = 32'h83070c8c;
    ram_cell[   28199] = 32'h2f6b0058;
    ram_cell[   28200] = 32'he1f9ae45;
    ram_cell[   28201] = 32'h1dc54516;
    ram_cell[   28202] = 32'h54fe8a86;
    ram_cell[   28203] = 32'heb359694;
    ram_cell[   28204] = 32'h58652f0b;
    ram_cell[   28205] = 32'h359bf9d3;
    ram_cell[   28206] = 32'h25d73a7d;
    ram_cell[   28207] = 32'hae3d612a;
    ram_cell[   28208] = 32'h19da483e;
    ram_cell[   28209] = 32'h4cb0c32b;
    ram_cell[   28210] = 32'h2e4edbda;
    ram_cell[   28211] = 32'h95fa4d5b;
    ram_cell[   28212] = 32'h527d355e;
    ram_cell[   28213] = 32'h03bde512;
    ram_cell[   28214] = 32'h49dd1039;
    ram_cell[   28215] = 32'h071821de;
    ram_cell[   28216] = 32'h5799000c;
    ram_cell[   28217] = 32'h789b04d3;
    ram_cell[   28218] = 32'hc0e92122;
    ram_cell[   28219] = 32'he9caa9e5;
    ram_cell[   28220] = 32'he84ba429;
    ram_cell[   28221] = 32'hcd09a79e;
    ram_cell[   28222] = 32'h9a55a3a9;
    ram_cell[   28223] = 32'he61557e9;
    ram_cell[   28224] = 32'hf69cc56d;
    ram_cell[   28225] = 32'hb75beed6;
    ram_cell[   28226] = 32'h718c55c7;
    ram_cell[   28227] = 32'h39d7ffc2;
    ram_cell[   28228] = 32'h54b04aa8;
    ram_cell[   28229] = 32'h302c605c;
    ram_cell[   28230] = 32'h9b90ee4e;
    ram_cell[   28231] = 32'h84155b38;
    ram_cell[   28232] = 32'h3569376c;
    ram_cell[   28233] = 32'h2026101e;
    ram_cell[   28234] = 32'hf05e74eb;
    ram_cell[   28235] = 32'h58f33074;
    ram_cell[   28236] = 32'hd0bdee2a;
    ram_cell[   28237] = 32'h91f03699;
    ram_cell[   28238] = 32'hc1d192e5;
    ram_cell[   28239] = 32'h6b3964b4;
    ram_cell[   28240] = 32'h230e09f4;
    ram_cell[   28241] = 32'hf28d1feb;
    ram_cell[   28242] = 32'h6a9623ee;
    ram_cell[   28243] = 32'he2a11d3a;
    ram_cell[   28244] = 32'h1ea9f57a;
    ram_cell[   28245] = 32'hcc0b73c0;
    ram_cell[   28246] = 32'h760f6f11;
    ram_cell[   28247] = 32'h2437cd13;
    ram_cell[   28248] = 32'h611cad85;
    ram_cell[   28249] = 32'h3336b23f;
    ram_cell[   28250] = 32'hed375b60;
    ram_cell[   28251] = 32'hebe766fc;
    ram_cell[   28252] = 32'h9530c24b;
    ram_cell[   28253] = 32'hd9c0bf22;
    ram_cell[   28254] = 32'h22efaf3c;
    ram_cell[   28255] = 32'hd8496e92;
    ram_cell[   28256] = 32'h17cf955d;
    ram_cell[   28257] = 32'h270a0ce8;
    ram_cell[   28258] = 32'hfa8bf7b9;
    ram_cell[   28259] = 32'h53ec95fa;
    ram_cell[   28260] = 32'h6dba190d;
    ram_cell[   28261] = 32'h7f8d0d12;
    ram_cell[   28262] = 32'h8001e900;
    ram_cell[   28263] = 32'h55c8a311;
    ram_cell[   28264] = 32'hda51e3e4;
    ram_cell[   28265] = 32'hbd927171;
    ram_cell[   28266] = 32'h004053e6;
    ram_cell[   28267] = 32'ha3ce6b3b;
    ram_cell[   28268] = 32'h1af2eab6;
    ram_cell[   28269] = 32'h6131c917;
    ram_cell[   28270] = 32'hcf3b673a;
    ram_cell[   28271] = 32'h82af75e3;
    ram_cell[   28272] = 32'hcb1ac804;
    ram_cell[   28273] = 32'he08d2388;
    ram_cell[   28274] = 32'h7baa7b53;
    ram_cell[   28275] = 32'h5f58a128;
    ram_cell[   28276] = 32'hb6651c98;
    ram_cell[   28277] = 32'hc74db763;
    ram_cell[   28278] = 32'h487cd866;
    ram_cell[   28279] = 32'h5f88e540;
    ram_cell[   28280] = 32'h81533695;
    ram_cell[   28281] = 32'h77c5229d;
    ram_cell[   28282] = 32'h070a2031;
    ram_cell[   28283] = 32'h94657fd2;
    ram_cell[   28284] = 32'h2aafd370;
    ram_cell[   28285] = 32'h8372afc7;
    ram_cell[   28286] = 32'h1b54fb91;
    ram_cell[   28287] = 32'ha0f88445;
    ram_cell[   28288] = 32'hdbc42467;
    ram_cell[   28289] = 32'hdc26ff8f;
    ram_cell[   28290] = 32'h0fee19ff;
    ram_cell[   28291] = 32'hf75a7e79;
    ram_cell[   28292] = 32'hf74213e4;
    ram_cell[   28293] = 32'hf8d9bbee;
    ram_cell[   28294] = 32'h73492b32;
    ram_cell[   28295] = 32'h190a3829;
    ram_cell[   28296] = 32'hec226239;
    ram_cell[   28297] = 32'h29b65a71;
    ram_cell[   28298] = 32'h5b8d8c5e;
    ram_cell[   28299] = 32'h9db8b488;
    ram_cell[   28300] = 32'h9c18a0d8;
    ram_cell[   28301] = 32'h14adcdb0;
    ram_cell[   28302] = 32'ha994fc1b;
    ram_cell[   28303] = 32'hf5f3e3bf;
    ram_cell[   28304] = 32'h4f34b015;
    ram_cell[   28305] = 32'h412fb935;
    ram_cell[   28306] = 32'hb3ef176e;
    ram_cell[   28307] = 32'h1f136d1c;
    ram_cell[   28308] = 32'hbef01371;
    ram_cell[   28309] = 32'h58a42fee;
    ram_cell[   28310] = 32'h5a4808a1;
    ram_cell[   28311] = 32'h79c90989;
    ram_cell[   28312] = 32'h4a208872;
    ram_cell[   28313] = 32'ha959deb1;
    ram_cell[   28314] = 32'h72aed535;
    ram_cell[   28315] = 32'h6ed381bf;
    ram_cell[   28316] = 32'hb3d1a365;
    ram_cell[   28317] = 32'ha5d8a891;
    ram_cell[   28318] = 32'h866948db;
    ram_cell[   28319] = 32'h10950dc3;
    ram_cell[   28320] = 32'h8984dede;
    ram_cell[   28321] = 32'h63b86051;
    ram_cell[   28322] = 32'h7dfce5e3;
    ram_cell[   28323] = 32'he4fd459e;
    ram_cell[   28324] = 32'hc627bae1;
    ram_cell[   28325] = 32'h15de67f0;
    ram_cell[   28326] = 32'h8d200acb;
    ram_cell[   28327] = 32'h895f0057;
    ram_cell[   28328] = 32'hdff93018;
    ram_cell[   28329] = 32'h721a4bdd;
    ram_cell[   28330] = 32'hc5515ac4;
    ram_cell[   28331] = 32'h68877e53;
    ram_cell[   28332] = 32'h097fe576;
    ram_cell[   28333] = 32'h344bb904;
    ram_cell[   28334] = 32'hf1f8950f;
    ram_cell[   28335] = 32'hec26b7bc;
    ram_cell[   28336] = 32'hb1b80b3c;
    ram_cell[   28337] = 32'hec4dd530;
    ram_cell[   28338] = 32'hda9edcb9;
    ram_cell[   28339] = 32'he022ed71;
    ram_cell[   28340] = 32'h2f8a6dfa;
    ram_cell[   28341] = 32'h52fb74de;
    ram_cell[   28342] = 32'hb9bf0f26;
    ram_cell[   28343] = 32'hb5a3f20f;
    ram_cell[   28344] = 32'h51e63795;
    ram_cell[   28345] = 32'h03b19408;
    ram_cell[   28346] = 32'hf5e2b297;
    ram_cell[   28347] = 32'ha1fd4c9a;
    ram_cell[   28348] = 32'hd63296b8;
    ram_cell[   28349] = 32'h669ae5b4;
    ram_cell[   28350] = 32'h98bbab7d;
    ram_cell[   28351] = 32'h611ee822;
    ram_cell[   28352] = 32'hf14d24d6;
    ram_cell[   28353] = 32'hd778da4e;
    ram_cell[   28354] = 32'hc28f1483;
    ram_cell[   28355] = 32'he8dbf4a7;
    ram_cell[   28356] = 32'h30db0976;
    ram_cell[   28357] = 32'h6d81281d;
    ram_cell[   28358] = 32'h258d5166;
    ram_cell[   28359] = 32'hc4e64e48;
    ram_cell[   28360] = 32'ha2b55a46;
    ram_cell[   28361] = 32'hba64b71c;
    ram_cell[   28362] = 32'hf5e77fa5;
    ram_cell[   28363] = 32'h9ae9147b;
    ram_cell[   28364] = 32'hf8948b21;
    ram_cell[   28365] = 32'h08322465;
    ram_cell[   28366] = 32'hcf43d27b;
    ram_cell[   28367] = 32'h0f1c89e8;
    ram_cell[   28368] = 32'h5abaadc0;
    ram_cell[   28369] = 32'h17695baf;
    ram_cell[   28370] = 32'h9280ee11;
    ram_cell[   28371] = 32'hb880e188;
    ram_cell[   28372] = 32'h2d51c4ba;
    ram_cell[   28373] = 32'haf76e238;
    ram_cell[   28374] = 32'h0b15bd3e;
    ram_cell[   28375] = 32'h6ab226b2;
    ram_cell[   28376] = 32'he70bc25d;
    ram_cell[   28377] = 32'h637190bd;
    ram_cell[   28378] = 32'h219c2a40;
    ram_cell[   28379] = 32'hbe27606b;
    ram_cell[   28380] = 32'h3ad79fb9;
    ram_cell[   28381] = 32'h1ba8d46d;
    ram_cell[   28382] = 32'haa5b757d;
    ram_cell[   28383] = 32'h41f191a8;
    ram_cell[   28384] = 32'h18c1cb4b;
    ram_cell[   28385] = 32'ha1bf2a00;
    ram_cell[   28386] = 32'h3c2abc07;
    ram_cell[   28387] = 32'hdacae04a;
    ram_cell[   28388] = 32'h1b5220da;
    ram_cell[   28389] = 32'h9446534d;
    ram_cell[   28390] = 32'h8dbffbe8;
    ram_cell[   28391] = 32'had02f027;
    ram_cell[   28392] = 32'h780737f5;
    ram_cell[   28393] = 32'he4c512f3;
    ram_cell[   28394] = 32'h57720547;
    ram_cell[   28395] = 32'hcef1214a;
    ram_cell[   28396] = 32'h63f5bda8;
    ram_cell[   28397] = 32'h81fd8792;
    ram_cell[   28398] = 32'he9b7069a;
    ram_cell[   28399] = 32'hea4e34ee;
    ram_cell[   28400] = 32'hea9f7326;
    ram_cell[   28401] = 32'hc20860fe;
    ram_cell[   28402] = 32'hd76c6e91;
    ram_cell[   28403] = 32'h2d032f24;
    ram_cell[   28404] = 32'h55f5ddce;
    ram_cell[   28405] = 32'h81c66fcb;
    ram_cell[   28406] = 32'h395c1310;
    ram_cell[   28407] = 32'h7f4e0034;
    ram_cell[   28408] = 32'hba30f8c5;
    ram_cell[   28409] = 32'h1f94ec3e;
    ram_cell[   28410] = 32'hf371a68c;
    ram_cell[   28411] = 32'hcda71644;
    ram_cell[   28412] = 32'h19e0b7a6;
    ram_cell[   28413] = 32'he8c09313;
    ram_cell[   28414] = 32'h07724984;
    ram_cell[   28415] = 32'hb48f0482;
    ram_cell[   28416] = 32'hc8643675;
    ram_cell[   28417] = 32'h3193071b;
    ram_cell[   28418] = 32'hb85a5eb4;
    ram_cell[   28419] = 32'h3073f85b;
    ram_cell[   28420] = 32'hf10eb7dd;
    ram_cell[   28421] = 32'h558b76ff;
    ram_cell[   28422] = 32'h00e5f25d;
    ram_cell[   28423] = 32'h8c2443cb;
    ram_cell[   28424] = 32'h9ac878fe;
    ram_cell[   28425] = 32'h098e1a30;
    ram_cell[   28426] = 32'h22695522;
    ram_cell[   28427] = 32'hd12c5b89;
    ram_cell[   28428] = 32'h1c3918d7;
    ram_cell[   28429] = 32'hdc630daf;
    ram_cell[   28430] = 32'ha54271d1;
    ram_cell[   28431] = 32'hb6af1210;
    ram_cell[   28432] = 32'h49a0a46d;
    ram_cell[   28433] = 32'h40eeeffb;
    ram_cell[   28434] = 32'h603b2dbb;
    ram_cell[   28435] = 32'h685ad417;
    ram_cell[   28436] = 32'h907c0acd;
    ram_cell[   28437] = 32'h1e61b37d;
    ram_cell[   28438] = 32'h3e41e524;
    ram_cell[   28439] = 32'hc1d84d67;
    ram_cell[   28440] = 32'h8bb2dca5;
    ram_cell[   28441] = 32'h65f142bd;
    ram_cell[   28442] = 32'h3e64c23a;
    ram_cell[   28443] = 32'hb0806b3f;
    ram_cell[   28444] = 32'hff0755dc;
    ram_cell[   28445] = 32'h14ac5a16;
    ram_cell[   28446] = 32'h7429cf5d;
    ram_cell[   28447] = 32'ha8aa67c7;
    ram_cell[   28448] = 32'h3cfd5144;
    ram_cell[   28449] = 32'hd35568cd;
    ram_cell[   28450] = 32'h1917b80f;
    ram_cell[   28451] = 32'had3c9307;
    ram_cell[   28452] = 32'h19257a8c;
    ram_cell[   28453] = 32'h1b4d8cbd;
    ram_cell[   28454] = 32'h9d1442c7;
    ram_cell[   28455] = 32'h6a0b4fde;
    ram_cell[   28456] = 32'h16744f2a;
    ram_cell[   28457] = 32'hed3cba24;
    ram_cell[   28458] = 32'h95b6f14d;
    ram_cell[   28459] = 32'hb43c64cc;
    ram_cell[   28460] = 32'hdceb6551;
    ram_cell[   28461] = 32'h170b1b59;
    ram_cell[   28462] = 32'h923075a6;
    ram_cell[   28463] = 32'hc8aecbdb;
    ram_cell[   28464] = 32'h0a06be41;
    ram_cell[   28465] = 32'h16e77300;
    ram_cell[   28466] = 32'h0b937a84;
    ram_cell[   28467] = 32'h03ff4b67;
    ram_cell[   28468] = 32'h9326ff8d;
    ram_cell[   28469] = 32'h124fc047;
    ram_cell[   28470] = 32'h2e452a65;
    ram_cell[   28471] = 32'h6943edc3;
    ram_cell[   28472] = 32'h0448ab61;
    ram_cell[   28473] = 32'hd723bd2f;
    ram_cell[   28474] = 32'h43d0a3ea;
    ram_cell[   28475] = 32'ha24aa895;
    ram_cell[   28476] = 32'hd7b7af96;
    ram_cell[   28477] = 32'h0c9d5888;
    ram_cell[   28478] = 32'h06831a46;
    ram_cell[   28479] = 32'h062403a2;
    ram_cell[   28480] = 32'ha7e562e5;
    ram_cell[   28481] = 32'hc07732c8;
    ram_cell[   28482] = 32'h0d83ce82;
    ram_cell[   28483] = 32'h947e6b9e;
    ram_cell[   28484] = 32'ha2b32506;
    ram_cell[   28485] = 32'h42ff6d40;
    ram_cell[   28486] = 32'h7bb45350;
    ram_cell[   28487] = 32'hee222b41;
    ram_cell[   28488] = 32'h3c4fd3cd;
    ram_cell[   28489] = 32'h2a0032a9;
    ram_cell[   28490] = 32'hd5349a11;
    ram_cell[   28491] = 32'h392c1cd6;
    ram_cell[   28492] = 32'hc226c820;
    ram_cell[   28493] = 32'h77770ab5;
    ram_cell[   28494] = 32'h455a9731;
    ram_cell[   28495] = 32'h03291a78;
    ram_cell[   28496] = 32'hee8b2347;
    ram_cell[   28497] = 32'h77d71e3d;
    ram_cell[   28498] = 32'h0eed35c6;
    ram_cell[   28499] = 32'h3e70b20f;
    ram_cell[   28500] = 32'h0159edab;
    ram_cell[   28501] = 32'hb0ef0886;
    ram_cell[   28502] = 32'h3a71ac76;
    ram_cell[   28503] = 32'h2d4ffddb;
    ram_cell[   28504] = 32'h631661b8;
    ram_cell[   28505] = 32'h4b697d17;
    ram_cell[   28506] = 32'h22168a7d;
    ram_cell[   28507] = 32'h2bab87aa;
    ram_cell[   28508] = 32'h33034f7e;
    ram_cell[   28509] = 32'h0fe8daad;
    ram_cell[   28510] = 32'he5621c52;
    ram_cell[   28511] = 32'h56936cc9;
    ram_cell[   28512] = 32'h770e6000;
    ram_cell[   28513] = 32'h11a142d6;
    ram_cell[   28514] = 32'h31d68a46;
    ram_cell[   28515] = 32'h3922a416;
    ram_cell[   28516] = 32'h732be58a;
    ram_cell[   28517] = 32'h9818f016;
    ram_cell[   28518] = 32'h7a61796a;
    ram_cell[   28519] = 32'hf337b1f4;
    ram_cell[   28520] = 32'hdedeba91;
    ram_cell[   28521] = 32'hbaba967c;
    ram_cell[   28522] = 32'h874f8ed0;
    ram_cell[   28523] = 32'h3d731492;
    ram_cell[   28524] = 32'h10946e63;
    ram_cell[   28525] = 32'hb271576e;
    ram_cell[   28526] = 32'h67dcb642;
    ram_cell[   28527] = 32'h6d8cf57d;
    ram_cell[   28528] = 32'h56e17b35;
    ram_cell[   28529] = 32'hf63ce21f;
    ram_cell[   28530] = 32'h4e814544;
    ram_cell[   28531] = 32'ha40332ac;
    ram_cell[   28532] = 32'h22f67a27;
    ram_cell[   28533] = 32'hde7ad4d7;
    ram_cell[   28534] = 32'h9b831b1f;
    ram_cell[   28535] = 32'h2ec5bebf;
    ram_cell[   28536] = 32'h0f694740;
    ram_cell[   28537] = 32'hd7a2a841;
    ram_cell[   28538] = 32'h8ed401cd;
    ram_cell[   28539] = 32'h7e933b4b;
    ram_cell[   28540] = 32'hd623c2c2;
    ram_cell[   28541] = 32'h32301d5a;
    ram_cell[   28542] = 32'h958febb2;
    ram_cell[   28543] = 32'h3fdc4525;
    ram_cell[   28544] = 32'h9f3ecb9a;
    ram_cell[   28545] = 32'h0c0c6eaf;
    ram_cell[   28546] = 32'h62328ea2;
    ram_cell[   28547] = 32'hf7b47113;
    ram_cell[   28548] = 32'ha1d02cb8;
    ram_cell[   28549] = 32'h5950fd2d;
    ram_cell[   28550] = 32'hda379718;
    ram_cell[   28551] = 32'h01e63147;
    ram_cell[   28552] = 32'h86bac787;
    ram_cell[   28553] = 32'h1afb1408;
    ram_cell[   28554] = 32'h75d88540;
    ram_cell[   28555] = 32'h0d0ca0f7;
    ram_cell[   28556] = 32'hae94d76d;
    ram_cell[   28557] = 32'h3d88ab7c;
    ram_cell[   28558] = 32'h28ad8565;
    ram_cell[   28559] = 32'h5ed1c29b;
    ram_cell[   28560] = 32'h78df1c2a;
    ram_cell[   28561] = 32'ha73d95e3;
    ram_cell[   28562] = 32'he9d5f7f2;
    ram_cell[   28563] = 32'he8291a46;
    ram_cell[   28564] = 32'hfa000273;
    ram_cell[   28565] = 32'h15962157;
    ram_cell[   28566] = 32'hfb87fb49;
    ram_cell[   28567] = 32'h87265ab0;
    ram_cell[   28568] = 32'hf74f3c2a;
    ram_cell[   28569] = 32'he3b4e586;
    ram_cell[   28570] = 32'h8ecb4fc0;
    ram_cell[   28571] = 32'h82c96713;
    ram_cell[   28572] = 32'h3dcbac9e;
    ram_cell[   28573] = 32'h90d2d88c;
    ram_cell[   28574] = 32'h465d7197;
    ram_cell[   28575] = 32'h2abe3894;
    ram_cell[   28576] = 32'h679ae2ba;
    ram_cell[   28577] = 32'h227657bd;
    ram_cell[   28578] = 32'h2ad70a74;
    ram_cell[   28579] = 32'h3a0ee1d7;
    ram_cell[   28580] = 32'h56b3ad9e;
    ram_cell[   28581] = 32'h01655f08;
    ram_cell[   28582] = 32'h5db497c0;
    ram_cell[   28583] = 32'hb6ed2fff;
    ram_cell[   28584] = 32'hf312c0d0;
    ram_cell[   28585] = 32'h84c69b59;
    ram_cell[   28586] = 32'h92fab2dc;
    ram_cell[   28587] = 32'h1277719b;
    ram_cell[   28588] = 32'h87e5b8f6;
    ram_cell[   28589] = 32'h4a14836b;
    ram_cell[   28590] = 32'h06f91700;
    ram_cell[   28591] = 32'hf950bcf4;
    ram_cell[   28592] = 32'h1a6c19e3;
    ram_cell[   28593] = 32'h9f65c838;
    ram_cell[   28594] = 32'h0fd64bb7;
    ram_cell[   28595] = 32'h42e122df;
    ram_cell[   28596] = 32'h0c09d8a8;
    ram_cell[   28597] = 32'hd70b4d87;
    ram_cell[   28598] = 32'hf6c415a1;
    ram_cell[   28599] = 32'ha05e55b4;
    ram_cell[   28600] = 32'h124fdb3f;
    ram_cell[   28601] = 32'h43ef7708;
    ram_cell[   28602] = 32'h011089a3;
    ram_cell[   28603] = 32'h79f8b498;
    ram_cell[   28604] = 32'h9f9e6a35;
    ram_cell[   28605] = 32'h65cb5768;
    ram_cell[   28606] = 32'hdfffc579;
    ram_cell[   28607] = 32'h20016011;
    ram_cell[   28608] = 32'h10391a48;
    ram_cell[   28609] = 32'he27bb1f4;
    ram_cell[   28610] = 32'ha927cbe1;
    ram_cell[   28611] = 32'h7e8d46df;
    ram_cell[   28612] = 32'h3a5132ae;
    ram_cell[   28613] = 32'h6dc2f65d;
    ram_cell[   28614] = 32'hd441c5ff;
    ram_cell[   28615] = 32'hf5fbecbf;
    ram_cell[   28616] = 32'h8567c12a;
    ram_cell[   28617] = 32'hd546d285;
    ram_cell[   28618] = 32'ha72ac859;
    ram_cell[   28619] = 32'h8db14b6f;
    ram_cell[   28620] = 32'h20ca009c;
    ram_cell[   28621] = 32'hffb5688e;
    ram_cell[   28622] = 32'h86589883;
    ram_cell[   28623] = 32'hf7ade344;
    ram_cell[   28624] = 32'h3a5e889a;
    ram_cell[   28625] = 32'h897a6b78;
    ram_cell[   28626] = 32'had63f9cd;
    ram_cell[   28627] = 32'ha77f005d;
    ram_cell[   28628] = 32'h058e8781;
    ram_cell[   28629] = 32'h8d270e01;
    ram_cell[   28630] = 32'h2d1eac48;
    ram_cell[   28631] = 32'h6af8bf41;
    ram_cell[   28632] = 32'h73cbead1;
    ram_cell[   28633] = 32'h94f576a7;
    ram_cell[   28634] = 32'h2a5491ce;
    ram_cell[   28635] = 32'h173e7c11;
    ram_cell[   28636] = 32'h0317e18c;
    ram_cell[   28637] = 32'hf382b4bb;
    ram_cell[   28638] = 32'h0bf7c651;
    ram_cell[   28639] = 32'hb8729ef3;
    ram_cell[   28640] = 32'hffd46846;
    ram_cell[   28641] = 32'hfebbfdfe;
    ram_cell[   28642] = 32'h624914aa;
    ram_cell[   28643] = 32'h6a8c25d2;
    ram_cell[   28644] = 32'h2a626403;
    ram_cell[   28645] = 32'h067794f0;
    ram_cell[   28646] = 32'h7939a62b;
    ram_cell[   28647] = 32'he837cc30;
    ram_cell[   28648] = 32'h03887cde;
    ram_cell[   28649] = 32'h88b323e7;
    ram_cell[   28650] = 32'h21590c42;
    ram_cell[   28651] = 32'h147c7128;
    ram_cell[   28652] = 32'hd8ab9ff8;
    ram_cell[   28653] = 32'h827efc68;
    ram_cell[   28654] = 32'hce55b40f;
    ram_cell[   28655] = 32'h363f6e38;
    ram_cell[   28656] = 32'h689ef24f;
    ram_cell[   28657] = 32'hafe296a2;
    ram_cell[   28658] = 32'h2351ad35;
    ram_cell[   28659] = 32'hf9c7979d;
    ram_cell[   28660] = 32'h47935f54;
    ram_cell[   28661] = 32'h0e1caeb2;
    ram_cell[   28662] = 32'hbc672d5b;
    ram_cell[   28663] = 32'h0417ce9a;
    ram_cell[   28664] = 32'h9aee2bdd;
    ram_cell[   28665] = 32'h768cf4d0;
    ram_cell[   28666] = 32'h1cd06f8f;
    ram_cell[   28667] = 32'h7304bc72;
    ram_cell[   28668] = 32'h98ea3d97;
    ram_cell[   28669] = 32'h4b3cdb79;
    ram_cell[   28670] = 32'he9dc9249;
    ram_cell[   28671] = 32'hce522f9c;
    ram_cell[   28672] = 32'hb11992e2;
    ram_cell[   28673] = 32'hf0f85e78;
    ram_cell[   28674] = 32'h7dd3865a;
    ram_cell[   28675] = 32'h6acdf37e;
    ram_cell[   28676] = 32'h507dc5ac;
    ram_cell[   28677] = 32'h313c4ec8;
    ram_cell[   28678] = 32'hff40500f;
    ram_cell[   28679] = 32'h1f440718;
    ram_cell[   28680] = 32'h8b3ec336;
    ram_cell[   28681] = 32'h63eca184;
    ram_cell[   28682] = 32'h60ded585;
    ram_cell[   28683] = 32'ha877d3f7;
    ram_cell[   28684] = 32'h2aa224a2;
    ram_cell[   28685] = 32'h79c226d4;
    ram_cell[   28686] = 32'h95d1d246;
    ram_cell[   28687] = 32'h6b0ababd;
    ram_cell[   28688] = 32'hc52faf80;
    ram_cell[   28689] = 32'h870baed4;
    ram_cell[   28690] = 32'hb1ad6d5b;
    ram_cell[   28691] = 32'heed2dacc;
    ram_cell[   28692] = 32'h1381146b;
    ram_cell[   28693] = 32'h945bdb35;
    ram_cell[   28694] = 32'h64043366;
    ram_cell[   28695] = 32'hb13100af;
    ram_cell[   28696] = 32'h141f119b;
    ram_cell[   28697] = 32'h192d6dd7;
    ram_cell[   28698] = 32'h0e414a32;
    ram_cell[   28699] = 32'h96aae955;
    ram_cell[   28700] = 32'h1da598a4;
    ram_cell[   28701] = 32'hffff5e4b;
    ram_cell[   28702] = 32'h05b0a6d1;
    ram_cell[   28703] = 32'hc4b1af60;
    ram_cell[   28704] = 32'hb6b33649;
    ram_cell[   28705] = 32'h0434b345;
    ram_cell[   28706] = 32'hac49a974;
    ram_cell[   28707] = 32'h87bc9c8d;
    ram_cell[   28708] = 32'h0a7d9176;
    ram_cell[   28709] = 32'hfb097175;
    ram_cell[   28710] = 32'h1447e169;
    ram_cell[   28711] = 32'h8eaf3e94;
    ram_cell[   28712] = 32'ha05ff7b7;
    ram_cell[   28713] = 32'h5cfbc47b;
    ram_cell[   28714] = 32'h15c5b56c;
    ram_cell[   28715] = 32'h3c4b2a19;
    ram_cell[   28716] = 32'hbeca61b4;
    ram_cell[   28717] = 32'hc0169fce;
    ram_cell[   28718] = 32'ha2277286;
    ram_cell[   28719] = 32'h3fa189a2;
    ram_cell[   28720] = 32'h11519961;
    ram_cell[   28721] = 32'h0d15555c;
    ram_cell[   28722] = 32'h67846454;
    ram_cell[   28723] = 32'hebfbe4e5;
    ram_cell[   28724] = 32'hea300498;
    ram_cell[   28725] = 32'hab3937c6;
    ram_cell[   28726] = 32'h16a43572;
    ram_cell[   28727] = 32'h59308e78;
    ram_cell[   28728] = 32'he9da02c4;
    ram_cell[   28729] = 32'h1eeb588b;
    ram_cell[   28730] = 32'h12aca436;
    ram_cell[   28731] = 32'h0f3177a8;
    ram_cell[   28732] = 32'hd7b248c7;
    ram_cell[   28733] = 32'h5b1eb3a1;
    ram_cell[   28734] = 32'h2ecace58;
    ram_cell[   28735] = 32'h0927b908;
    ram_cell[   28736] = 32'h9dcaaa15;
    ram_cell[   28737] = 32'h0a6a7a93;
    ram_cell[   28738] = 32'h2fdb0585;
    ram_cell[   28739] = 32'h138afebf;
    ram_cell[   28740] = 32'h2f04b45c;
    ram_cell[   28741] = 32'h7b49abe8;
    ram_cell[   28742] = 32'h6a87956a;
    ram_cell[   28743] = 32'hb53a3578;
    ram_cell[   28744] = 32'ha6c1d88c;
    ram_cell[   28745] = 32'h129189ec;
    ram_cell[   28746] = 32'he356cc7b;
    ram_cell[   28747] = 32'ha1a00268;
    ram_cell[   28748] = 32'h86aa98c9;
    ram_cell[   28749] = 32'h5e17164b;
    ram_cell[   28750] = 32'h154b6c45;
    ram_cell[   28751] = 32'h6d90e91a;
    ram_cell[   28752] = 32'h51ffecec;
    ram_cell[   28753] = 32'h01f6e320;
    ram_cell[   28754] = 32'h27067b7e;
    ram_cell[   28755] = 32'hbf5111d9;
    ram_cell[   28756] = 32'h60a6339f;
    ram_cell[   28757] = 32'h17f9b4ff;
    ram_cell[   28758] = 32'hdf6884c3;
    ram_cell[   28759] = 32'hca7a98e4;
    ram_cell[   28760] = 32'h49e75219;
    ram_cell[   28761] = 32'hc9e61225;
    ram_cell[   28762] = 32'h456a3521;
    ram_cell[   28763] = 32'h140e05ef;
    ram_cell[   28764] = 32'h795f9994;
    ram_cell[   28765] = 32'h610cdbca;
    ram_cell[   28766] = 32'h08d4676f;
    ram_cell[   28767] = 32'h73f46dfa;
    ram_cell[   28768] = 32'h0c7bdea6;
    ram_cell[   28769] = 32'hbb4774f1;
    ram_cell[   28770] = 32'h44b1613e;
    ram_cell[   28771] = 32'h0efa08f8;
    ram_cell[   28772] = 32'h7de2606c;
    ram_cell[   28773] = 32'h75ce221f;
    ram_cell[   28774] = 32'h018d14d0;
    ram_cell[   28775] = 32'hfddd8bf2;
    ram_cell[   28776] = 32'ha45dedd3;
    ram_cell[   28777] = 32'hb85ca3f8;
    ram_cell[   28778] = 32'h8572d715;
    ram_cell[   28779] = 32'h2ee76e6c;
    ram_cell[   28780] = 32'h707f5879;
    ram_cell[   28781] = 32'hc0e9988c;
    ram_cell[   28782] = 32'h8df8e18f;
    ram_cell[   28783] = 32'h9f2681f8;
    ram_cell[   28784] = 32'h782cab41;
    ram_cell[   28785] = 32'hd3694a0a;
    ram_cell[   28786] = 32'h218fecd9;
    ram_cell[   28787] = 32'hf681c4fa;
    ram_cell[   28788] = 32'h48b759c2;
    ram_cell[   28789] = 32'hfd3f1562;
    ram_cell[   28790] = 32'hf73967f5;
    ram_cell[   28791] = 32'h00723c4f;
    ram_cell[   28792] = 32'h2bc9d9f4;
    ram_cell[   28793] = 32'hb66a49e6;
    ram_cell[   28794] = 32'h8adb583a;
    ram_cell[   28795] = 32'hf017fc3b;
    ram_cell[   28796] = 32'h2a6930ba;
    ram_cell[   28797] = 32'h7791afa1;
    ram_cell[   28798] = 32'h64d5449e;
    ram_cell[   28799] = 32'h9bb5d582;
    ram_cell[   28800] = 32'h0a23fdb3;
    ram_cell[   28801] = 32'hf86a0130;
    ram_cell[   28802] = 32'h0604d950;
    ram_cell[   28803] = 32'h05c0e944;
    ram_cell[   28804] = 32'hfe14867f;
    ram_cell[   28805] = 32'h9813e04e;
    ram_cell[   28806] = 32'h55e7bd77;
    ram_cell[   28807] = 32'h6c55dbb5;
    ram_cell[   28808] = 32'hd4743b49;
    ram_cell[   28809] = 32'hcabad50b;
    ram_cell[   28810] = 32'hc018fd3f;
    ram_cell[   28811] = 32'h322fb587;
    ram_cell[   28812] = 32'h6f14e2e1;
    ram_cell[   28813] = 32'hf717c521;
    ram_cell[   28814] = 32'h93e2af9d;
    ram_cell[   28815] = 32'he13927a0;
    ram_cell[   28816] = 32'h36c159c6;
    ram_cell[   28817] = 32'h0b9097f5;
    ram_cell[   28818] = 32'h2cb8ba2e;
    ram_cell[   28819] = 32'h8b39a5f6;
    ram_cell[   28820] = 32'ha8336c2a;
    ram_cell[   28821] = 32'h983dedd0;
    ram_cell[   28822] = 32'hc171253c;
    ram_cell[   28823] = 32'h26ad2350;
    ram_cell[   28824] = 32'h9eebad49;
    ram_cell[   28825] = 32'h6ec5fad7;
    ram_cell[   28826] = 32'hae58f642;
    ram_cell[   28827] = 32'h58fad765;
    ram_cell[   28828] = 32'hdd4f42af;
    ram_cell[   28829] = 32'hc855f9ad;
    ram_cell[   28830] = 32'h036742d4;
    ram_cell[   28831] = 32'hda50c0dc;
    ram_cell[   28832] = 32'hc9fd3f2a;
    ram_cell[   28833] = 32'h797bed77;
    ram_cell[   28834] = 32'h46e47716;
    ram_cell[   28835] = 32'h50f9469b;
    ram_cell[   28836] = 32'hdf29b631;
    ram_cell[   28837] = 32'ha244d767;
    ram_cell[   28838] = 32'h36b7496e;
    ram_cell[   28839] = 32'h1d834edc;
    ram_cell[   28840] = 32'h25a1758f;
    ram_cell[   28841] = 32'ha94b4628;
    ram_cell[   28842] = 32'hb5382479;
    ram_cell[   28843] = 32'h3bb406fa;
    ram_cell[   28844] = 32'ha03d80c7;
    ram_cell[   28845] = 32'h171a2e4d;
    ram_cell[   28846] = 32'haccd79ad;
    ram_cell[   28847] = 32'hb2c6a8e4;
    ram_cell[   28848] = 32'he42c777c;
    ram_cell[   28849] = 32'h798b4655;
    ram_cell[   28850] = 32'h915d9407;
    ram_cell[   28851] = 32'h1275f3c5;
    ram_cell[   28852] = 32'h93ce7463;
    ram_cell[   28853] = 32'hb5512245;
    ram_cell[   28854] = 32'ha95bd245;
    ram_cell[   28855] = 32'h6b353c79;
    ram_cell[   28856] = 32'h56c1a948;
    ram_cell[   28857] = 32'h62ab8220;
    ram_cell[   28858] = 32'hbfbcb5ae;
    ram_cell[   28859] = 32'h5a353282;
    ram_cell[   28860] = 32'ha5a3fe96;
    ram_cell[   28861] = 32'h76329af3;
    ram_cell[   28862] = 32'h7ee6c409;
    ram_cell[   28863] = 32'h9d193f55;
    ram_cell[   28864] = 32'hf4521bae;
    ram_cell[   28865] = 32'h0477e974;
    ram_cell[   28866] = 32'hee0657a3;
    ram_cell[   28867] = 32'hfa8a4cef;
    ram_cell[   28868] = 32'h0c2b8cdf;
    ram_cell[   28869] = 32'h1c7ca621;
    ram_cell[   28870] = 32'h73ce4627;
    ram_cell[   28871] = 32'h177435e6;
    ram_cell[   28872] = 32'h037fd6d6;
    ram_cell[   28873] = 32'hffd67cd5;
    ram_cell[   28874] = 32'h5f6b1282;
    ram_cell[   28875] = 32'h69e52067;
    ram_cell[   28876] = 32'h58aa5219;
    ram_cell[   28877] = 32'hc30c69b4;
    ram_cell[   28878] = 32'he79f998b;
    ram_cell[   28879] = 32'h5558a484;
    ram_cell[   28880] = 32'h10ad27f2;
    ram_cell[   28881] = 32'h8052beb7;
    ram_cell[   28882] = 32'h9bdd2162;
    ram_cell[   28883] = 32'h44c78a83;
    ram_cell[   28884] = 32'he3ebf6ee;
    ram_cell[   28885] = 32'h88aec18f;
    ram_cell[   28886] = 32'h4d11ed59;
    ram_cell[   28887] = 32'h4f4e42ca;
    ram_cell[   28888] = 32'h44e3202e;
    ram_cell[   28889] = 32'h44ad06ea;
    ram_cell[   28890] = 32'h49370283;
    ram_cell[   28891] = 32'h8cf203b7;
    ram_cell[   28892] = 32'h1f7d85bc;
    ram_cell[   28893] = 32'hfad629c6;
    ram_cell[   28894] = 32'h1b4a51b1;
    ram_cell[   28895] = 32'h5023fee5;
    ram_cell[   28896] = 32'he6b45fd6;
    ram_cell[   28897] = 32'ha30b9ae7;
    ram_cell[   28898] = 32'h4e4bcaa2;
    ram_cell[   28899] = 32'h8526ae91;
    ram_cell[   28900] = 32'h5a6a5370;
    ram_cell[   28901] = 32'h70ee1d91;
    ram_cell[   28902] = 32'h70c2ef55;
    ram_cell[   28903] = 32'hb1a33891;
    ram_cell[   28904] = 32'h986e1bd5;
    ram_cell[   28905] = 32'hb24d78c8;
    ram_cell[   28906] = 32'hacfd63cd;
    ram_cell[   28907] = 32'h62b0bc80;
    ram_cell[   28908] = 32'h8252f336;
    ram_cell[   28909] = 32'ha7c6f5cf;
    ram_cell[   28910] = 32'hc90fa815;
    ram_cell[   28911] = 32'hc9f08964;
    ram_cell[   28912] = 32'h6f5097b8;
    ram_cell[   28913] = 32'hec26496f;
    ram_cell[   28914] = 32'h693e7f2a;
    ram_cell[   28915] = 32'h7f47717d;
    ram_cell[   28916] = 32'hfbc371fd;
    ram_cell[   28917] = 32'h9d9a63eb;
    ram_cell[   28918] = 32'hfacad477;
    ram_cell[   28919] = 32'hcd171e66;
    ram_cell[   28920] = 32'h53f7de4d;
    ram_cell[   28921] = 32'hd251e999;
    ram_cell[   28922] = 32'hf0c98e1e;
    ram_cell[   28923] = 32'h4d3e78f8;
    ram_cell[   28924] = 32'ha8f53e53;
    ram_cell[   28925] = 32'h35d60ba5;
    ram_cell[   28926] = 32'he72264fb;
    ram_cell[   28927] = 32'h75a89500;
    ram_cell[   28928] = 32'h24305917;
    ram_cell[   28929] = 32'h84f800c6;
    ram_cell[   28930] = 32'hd2f34209;
    ram_cell[   28931] = 32'hd365cd8f;
    ram_cell[   28932] = 32'he77e6f12;
    ram_cell[   28933] = 32'hd4b633b1;
    ram_cell[   28934] = 32'h8f7c5579;
    ram_cell[   28935] = 32'hb59a9163;
    ram_cell[   28936] = 32'h8473af4e;
    ram_cell[   28937] = 32'h3a984c12;
    ram_cell[   28938] = 32'h35c77f56;
    ram_cell[   28939] = 32'h003479b2;
    ram_cell[   28940] = 32'h0046a86d;
    ram_cell[   28941] = 32'h9c6ce246;
    ram_cell[   28942] = 32'h45d3d6d8;
    ram_cell[   28943] = 32'had994cad;
    ram_cell[   28944] = 32'h179948ca;
    ram_cell[   28945] = 32'he14e85e2;
    ram_cell[   28946] = 32'h977762b4;
    ram_cell[   28947] = 32'hb16dc828;
    ram_cell[   28948] = 32'h8cdf0191;
    ram_cell[   28949] = 32'hacec4ca0;
    ram_cell[   28950] = 32'h0bee6881;
    ram_cell[   28951] = 32'h8e66fb82;
    ram_cell[   28952] = 32'h0e751b01;
    ram_cell[   28953] = 32'hf8a2c1f0;
    ram_cell[   28954] = 32'h78ee0cd7;
    ram_cell[   28955] = 32'h672fa513;
    ram_cell[   28956] = 32'hd9c3e92a;
    ram_cell[   28957] = 32'ha092bf8f;
    ram_cell[   28958] = 32'h26fc69e6;
    ram_cell[   28959] = 32'he7199948;
    ram_cell[   28960] = 32'hb31fac09;
    ram_cell[   28961] = 32'ha7d9a1ad;
    ram_cell[   28962] = 32'h9b1fed3d;
    ram_cell[   28963] = 32'hd27b8a85;
    ram_cell[   28964] = 32'h7010beb2;
    ram_cell[   28965] = 32'h73153711;
    ram_cell[   28966] = 32'hf126d918;
    ram_cell[   28967] = 32'h23214911;
    ram_cell[   28968] = 32'hf8e4ed39;
    ram_cell[   28969] = 32'h9dab7949;
    ram_cell[   28970] = 32'h7fcb152e;
    ram_cell[   28971] = 32'h00a71755;
    ram_cell[   28972] = 32'h7c6bea94;
    ram_cell[   28973] = 32'hae28580a;
    ram_cell[   28974] = 32'hca387dc9;
    ram_cell[   28975] = 32'h4930f70d;
    ram_cell[   28976] = 32'h7a5ad26c;
    ram_cell[   28977] = 32'hc78a1787;
    ram_cell[   28978] = 32'h976d5e88;
    ram_cell[   28979] = 32'hb0b1cd7b;
    ram_cell[   28980] = 32'h078f7acf;
    ram_cell[   28981] = 32'h4db225cc;
    ram_cell[   28982] = 32'h87a04cb5;
    ram_cell[   28983] = 32'h40516df6;
    ram_cell[   28984] = 32'h0f946936;
    ram_cell[   28985] = 32'h6d513a40;
    ram_cell[   28986] = 32'hfcec0bd9;
    ram_cell[   28987] = 32'h7d844487;
    ram_cell[   28988] = 32'hb16cb1dc;
    ram_cell[   28989] = 32'hf2cdab65;
    ram_cell[   28990] = 32'hce2ecb42;
    ram_cell[   28991] = 32'hb32a6d49;
    ram_cell[   28992] = 32'h7cd49359;
    ram_cell[   28993] = 32'h7f5ff42e;
    ram_cell[   28994] = 32'h75b53f35;
    ram_cell[   28995] = 32'h845cd2db;
    ram_cell[   28996] = 32'h012ffb4b;
    ram_cell[   28997] = 32'hb0ea2913;
    ram_cell[   28998] = 32'h7d8f18ad;
    ram_cell[   28999] = 32'habcfc3cc;
    ram_cell[   29000] = 32'h8646eea9;
    ram_cell[   29001] = 32'h991e879c;
    ram_cell[   29002] = 32'he6d76e7f;
    ram_cell[   29003] = 32'hd6ff458a;
    ram_cell[   29004] = 32'hfb09325e;
    ram_cell[   29005] = 32'h1517ead0;
    ram_cell[   29006] = 32'h4a244efd;
    ram_cell[   29007] = 32'hbe977f39;
    ram_cell[   29008] = 32'hb579a0de;
    ram_cell[   29009] = 32'h9c3751ef;
    ram_cell[   29010] = 32'h50654a5c;
    ram_cell[   29011] = 32'hb4721c70;
    ram_cell[   29012] = 32'had699715;
    ram_cell[   29013] = 32'hdef05ed7;
    ram_cell[   29014] = 32'hb337dfe5;
    ram_cell[   29015] = 32'h248ad3d7;
    ram_cell[   29016] = 32'h3e0f5ae6;
    ram_cell[   29017] = 32'habc2346a;
    ram_cell[   29018] = 32'hc70ca950;
    ram_cell[   29019] = 32'h0ff38e01;
    ram_cell[   29020] = 32'h5b91450d;
    ram_cell[   29021] = 32'h8b06961c;
    ram_cell[   29022] = 32'hecc2b85c;
    ram_cell[   29023] = 32'h7ddaf295;
    ram_cell[   29024] = 32'h1daa6d56;
    ram_cell[   29025] = 32'had2fca05;
    ram_cell[   29026] = 32'hcb24e593;
    ram_cell[   29027] = 32'h4922ea83;
    ram_cell[   29028] = 32'h32142b00;
    ram_cell[   29029] = 32'h6357cdd1;
    ram_cell[   29030] = 32'hfef7f5bf;
    ram_cell[   29031] = 32'h11939e91;
    ram_cell[   29032] = 32'h70d94af3;
    ram_cell[   29033] = 32'h2bc9dd45;
    ram_cell[   29034] = 32'h4e18f52e;
    ram_cell[   29035] = 32'hdcdb3707;
    ram_cell[   29036] = 32'h118d971d;
    ram_cell[   29037] = 32'h828ebd51;
    ram_cell[   29038] = 32'h3d0953f0;
    ram_cell[   29039] = 32'haf8f7afa;
    ram_cell[   29040] = 32'hd5ba934a;
    ram_cell[   29041] = 32'h90ccdb5a;
    ram_cell[   29042] = 32'h739e2520;
    ram_cell[   29043] = 32'he72d1fab;
    ram_cell[   29044] = 32'he1c45a63;
    ram_cell[   29045] = 32'hd5dc6fb3;
    ram_cell[   29046] = 32'h62ccf5b0;
    ram_cell[   29047] = 32'h15e11cbc;
    ram_cell[   29048] = 32'hdb43ead9;
    ram_cell[   29049] = 32'h4c7f5a37;
    ram_cell[   29050] = 32'h2241a04c;
    ram_cell[   29051] = 32'h5dbe852f;
    ram_cell[   29052] = 32'hdc461e57;
    ram_cell[   29053] = 32'hc2ecc15c;
    ram_cell[   29054] = 32'he96eda27;
    ram_cell[   29055] = 32'h3be12ae9;
    ram_cell[   29056] = 32'h5c4ea3b2;
    ram_cell[   29057] = 32'h2c8b702a;
    ram_cell[   29058] = 32'h1878186f;
    ram_cell[   29059] = 32'h88d526ac;
    ram_cell[   29060] = 32'hafcd755d;
    ram_cell[   29061] = 32'h0e386303;
    ram_cell[   29062] = 32'h43923461;
    ram_cell[   29063] = 32'h679e448b;
    ram_cell[   29064] = 32'hceada805;
    ram_cell[   29065] = 32'ha604bd26;
    ram_cell[   29066] = 32'h0a917f87;
    ram_cell[   29067] = 32'h2b116b8a;
    ram_cell[   29068] = 32'h128c1457;
    ram_cell[   29069] = 32'h276b6254;
    ram_cell[   29070] = 32'h4f49ce97;
    ram_cell[   29071] = 32'he5b5fff8;
    ram_cell[   29072] = 32'hdaa2b33e;
    ram_cell[   29073] = 32'hf8b41271;
    ram_cell[   29074] = 32'h2242bcb1;
    ram_cell[   29075] = 32'hbd33077f;
    ram_cell[   29076] = 32'h0b2bf08c;
    ram_cell[   29077] = 32'hd2925ffb;
    ram_cell[   29078] = 32'hf35ea4cd;
    ram_cell[   29079] = 32'h2a9b3ce7;
    ram_cell[   29080] = 32'hd27211dc;
    ram_cell[   29081] = 32'hde7d628f;
    ram_cell[   29082] = 32'h916f75e0;
    ram_cell[   29083] = 32'he7a3badd;
    ram_cell[   29084] = 32'h7dc1c463;
    ram_cell[   29085] = 32'h371f01f3;
    ram_cell[   29086] = 32'h4584c03e;
    ram_cell[   29087] = 32'h1512d291;
    ram_cell[   29088] = 32'h380ccc73;
    ram_cell[   29089] = 32'hfb4aa08b;
    ram_cell[   29090] = 32'hbab415db;
    ram_cell[   29091] = 32'h9bb03bd9;
    ram_cell[   29092] = 32'he21c6165;
    ram_cell[   29093] = 32'h6250e9ad;
    ram_cell[   29094] = 32'hc17c81b6;
    ram_cell[   29095] = 32'h658043e2;
    ram_cell[   29096] = 32'hef69d0b7;
    ram_cell[   29097] = 32'h4aa3b098;
    ram_cell[   29098] = 32'h177cde4f;
    ram_cell[   29099] = 32'hbc62689a;
    ram_cell[   29100] = 32'ha04946b8;
    ram_cell[   29101] = 32'h1f673d28;
    ram_cell[   29102] = 32'h9767425b;
    ram_cell[   29103] = 32'hb2cd068c;
    ram_cell[   29104] = 32'h5c917bd3;
    ram_cell[   29105] = 32'haf6c8d62;
    ram_cell[   29106] = 32'hf180b945;
    ram_cell[   29107] = 32'h3fc6a3b7;
    ram_cell[   29108] = 32'hb5074763;
    ram_cell[   29109] = 32'hcee4c6fc;
    ram_cell[   29110] = 32'h0db2f742;
    ram_cell[   29111] = 32'h6fab4b07;
    ram_cell[   29112] = 32'hc88ead30;
    ram_cell[   29113] = 32'h9c76cc08;
    ram_cell[   29114] = 32'h573568fc;
    ram_cell[   29115] = 32'h20fe34c4;
    ram_cell[   29116] = 32'h8739f05f;
    ram_cell[   29117] = 32'hac061632;
    ram_cell[   29118] = 32'hd10b374d;
    ram_cell[   29119] = 32'hea255cb6;
    ram_cell[   29120] = 32'h7014084d;
    ram_cell[   29121] = 32'h23b8dcfa;
    ram_cell[   29122] = 32'hb2ba1940;
    ram_cell[   29123] = 32'h65507d35;
    ram_cell[   29124] = 32'h72a32419;
    ram_cell[   29125] = 32'h7474b148;
    ram_cell[   29126] = 32'hf215381a;
    ram_cell[   29127] = 32'he29e47dd;
    ram_cell[   29128] = 32'h1730ff53;
    ram_cell[   29129] = 32'h8f16a9c4;
    ram_cell[   29130] = 32'h7f8f2fd6;
    ram_cell[   29131] = 32'h60cdea7b;
    ram_cell[   29132] = 32'h681b51c8;
    ram_cell[   29133] = 32'h0d263053;
    ram_cell[   29134] = 32'h8b024600;
    ram_cell[   29135] = 32'h3ded74f5;
    ram_cell[   29136] = 32'h1f55dae5;
    ram_cell[   29137] = 32'h52e772a2;
    ram_cell[   29138] = 32'h55383e29;
    ram_cell[   29139] = 32'h92e96238;
    ram_cell[   29140] = 32'hf97754d4;
    ram_cell[   29141] = 32'h809e4940;
    ram_cell[   29142] = 32'h50b35d9b;
    ram_cell[   29143] = 32'h0cb2dca7;
    ram_cell[   29144] = 32'h8700af28;
    ram_cell[   29145] = 32'h2ca4d8b8;
    ram_cell[   29146] = 32'h7fb3f2a4;
    ram_cell[   29147] = 32'h2e14fd4b;
    ram_cell[   29148] = 32'h1d8f9f78;
    ram_cell[   29149] = 32'hd596b10a;
    ram_cell[   29150] = 32'hf47e3ad6;
    ram_cell[   29151] = 32'hf1d554bf;
    ram_cell[   29152] = 32'hc85a2a5a;
    ram_cell[   29153] = 32'ha9ca37ec;
    ram_cell[   29154] = 32'ha09aacdb;
    ram_cell[   29155] = 32'h94bddad2;
    ram_cell[   29156] = 32'hb0a87990;
    ram_cell[   29157] = 32'h8feb8798;
    ram_cell[   29158] = 32'hc2907d7b;
    ram_cell[   29159] = 32'hfc8fce49;
    ram_cell[   29160] = 32'he8a87b50;
    ram_cell[   29161] = 32'hbac2700d;
    ram_cell[   29162] = 32'h578e9388;
    ram_cell[   29163] = 32'h7bf57e23;
    ram_cell[   29164] = 32'hd57b6858;
    ram_cell[   29165] = 32'h8692e7c4;
    ram_cell[   29166] = 32'hb6eefbad;
    ram_cell[   29167] = 32'hf45e6e17;
    ram_cell[   29168] = 32'hac4c9e92;
    ram_cell[   29169] = 32'hd4e92fb3;
    ram_cell[   29170] = 32'h73c6f576;
    ram_cell[   29171] = 32'hd8a0966a;
    ram_cell[   29172] = 32'hd45ce574;
    ram_cell[   29173] = 32'h6871a648;
    ram_cell[   29174] = 32'hac11c9b2;
    ram_cell[   29175] = 32'h9b632ba6;
    ram_cell[   29176] = 32'hcb71e10b;
    ram_cell[   29177] = 32'he6f48bc4;
    ram_cell[   29178] = 32'hb251ab00;
    ram_cell[   29179] = 32'h053186e9;
    ram_cell[   29180] = 32'h5599449d;
    ram_cell[   29181] = 32'hf17169fe;
    ram_cell[   29182] = 32'h2164d8ff;
    ram_cell[   29183] = 32'h76f60ace;
    ram_cell[   29184] = 32'hb5fd1f6e;
    ram_cell[   29185] = 32'hf79ed6f3;
    ram_cell[   29186] = 32'h50e957be;
    ram_cell[   29187] = 32'hc82b589b;
    ram_cell[   29188] = 32'h648d6475;
    ram_cell[   29189] = 32'hf45f6b42;
    ram_cell[   29190] = 32'ha3c2de54;
    ram_cell[   29191] = 32'h3c024452;
    ram_cell[   29192] = 32'h725dc66a;
    ram_cell[   29193] = 32'h6fb24c4e;
    ram_cell[   29194] = 32'h3b9e06aa;
    ram_cell[   29195] = 32'h459704a8;
    ram_cell[   29196] = 32'he5d86b95;
    ram_cell[   29197] = 32'h2deb076c;
    ram_cell[   29198] = 32'h0d4f469a;
    ram_cell[   29199] = 32'h69990ad3;
    ram_cell[   29200] = 32'h5e944c7b;
    ram_cell[   29201] = 32'h072a94da;
    ram_cell[   29202] = 32'h1b9c5219;
    ram_cell[   29203] = 32'hbbbfb404;
    ram_cell[   29204] = 32'ha148a04a;
    ram_cell[   29205] = 32'h66b3428b;
    ram_cell[   29206] = 32'h85cf64a9;
    ram_cell[   29207] = 32'h1fa76ce6;
    ram_cell[   29208] = 32'h02a91234;
    ram_cell[   29209] = 32'hca3f29de;
    ram_cell[   29210] = 32'h33e8f613;
    ram_cell[   29211] = 32'hc6f26673;
    ram_cell[   29212] = 32'hce48f844;
    ram_cell[   29213] = 32'h74490eab;
    ram_cell[   29214] = 32'hdc382ebf;
    ram_cell[   29215] = 32'hd9acfff3;
    ram_cell[   29216] = 32'hd418a84c;
    ram_cell[   29217] = 32'hebfcb66d;
    ram_cell[   29218] = 32'h20ced4f2;
    ram_cell[   29219] = 32'hae616697;
    ram_cell[   29220] = 32'h276be9f9;
    ram_cell[   29221] = 32'hd57c727d;
    ram_cell[   29222] = 32'h284a8587;
    ram_cell[   29223] = 32'hf8934ce5;
    ram_cell[   29224] = 32'hb0943e90;
    ram_cell[   29225] = 32'h0762d5b5;
    ram_cell[   29226] = 32'h661d6b67;
    ram_cell[   29227] = 32'h87370ea1;
    ram_cell[   29228] = 32'h8a1759d1;
    ram_cell[   29229] = 32'h7bb5f09e;
    ram_cell[   29230] = 32'h9a4df294;
    ram_cell[   29231] = 32'he6fdcaac;
    ram_cell[   29232] = 32'h4373a800;
    ram_cell[   29233] = 32'heb38e57e;
    ram_cell[   29234] = 32'h379bd939;
    ram_cell[   29235] = 32'h10e85683;
    ram_cell[   29236] = 32'h3015fc4a;
    ram_cell[   29237] = 32'h42cf5c5f;
    ram_cell[   29238] = 32'h74db5545;
    ram_cell[   29239] = 32'h3a53219a;
    ram_cell[   29240] = 32'hc3467082;
    ram_cell[   29241] = 32'hfd047028;
    ram_cell[   29242] = 32'haf6129c7;
    ram_cell[   29243] = 32'h496d235c;
    ram_cell[   29244] = 32'h627f8f7d;
    ram_cell[   29245] = 32'h6bcbf84e;
    ram_cell[   29246] = 32'h43edcf17;
    ram_cell[   29247] = 32'hbf6c43e7;
    ram_cell[   29248] = 32'hbe79319e;
    ram_cell[   29249] = 32'h814e8042;
    ram_cell[   29250] = 32'h99c1b46a;
    ram_cell[   29251] = 32'h19d59c20;
    ram_cell[   29252] = 32'h782d5b00;
    ram_cell[   29253] = 32'h30360295;
    ram_cell[   29254] = 32'h607b8dbb;
    ram_cell[   29255] = 32'h66c4c5b4;
    ram_cell[   29256] = 32'h597f5751;
    ram_cell[   29257] = 32'h7d745292;
    ram_cell[   29258] = 32'hf3d71248;
    ram_cell[   29259] = 32'h5e942bc1;
    ram_cell[   29260] = 32'h2f117e4a;
    ram_cell[   29261] = 32'haf4d1038;
    ram_cell[   29262] = 32'h23a0d084;
    ram_cell[   29263] = 32'h247b77ad;
    ram_cell[   29264] = 32'h3a1b0691;
    ram_cell[   29265] = 32'h3c5d3226;
    ram_cell[   29266] = 32'h96ea6ea0;
    ram_cell[   29267] = 32'h87ecb6f6;
    ram_cell[   29268] = 32'hd7008bdb;
    ram_cell[   29269] = 32'h57ac93d6;
    ram_cell[   29270] = 32'he81aacc0;
    ram_cell[   29271] = 32'h44be5f85;
    ram_cell[   29272] = 32'h444ce385;
    ram_cell[   29273] = 32'h24855543;
    ram_cell[   29274] = 32'h9504ded1;
    ram_cell[   29275] = 32'h44770e4d;
    ram_cell[   29276] = 32'h02212e1b;
    ram_cell[   29277] = 32'h6cb13ed5;
    ram_cell[   29278] = 32'hd701ee96;
    ram_cell[   29279] = 32'hf97c332f;
    ram_cell[   29280] = 32'h64f06373;
    ram_cell[   29281] = 32'h11f51bd1;
    ram_cell[   29282] = 32'h5115e0c9;
    ram_cell[   29283] = 32'h7c52978e;
    ram_cell[   29284] = 32'haaaf32b7;
    ram_cell[   29285] = 32'h41f2404b;
    ram_cell[   29286] = 32'h08406ce2;
    ram_cell[   29287] = 32'h8056da7f;
    ram_cell[   29288] = 32'h4f73cf5b;
    ram_cell[   29289] = 32'hb77d3c6c;
    ram_cell[   29290] = 32'h25ec8fd7;
    ram_cell[   29291] = 32'hc62c7fd6;
    ram_cell[   29292] = 32'hab6abf98;
    ram_cell[   29293] = 32'ha83426bd;
    ram_cell[   29294] = 32'hd2a8edee;
    ram_cell[   29295] = 32'h70b1dc14;
    ram_cell[   29296] = 32'ha2c258e8;
    ram_cell[   29297] = 32'h2c76d8ec;
    ram_cell[   29298] = 32'h4e451175;
    ram_cell[   29299] = 32'hc4ceb3ee;
    ram_cell[   29300] = 32'h49d4c57a;
    ram_cell[   29301] = 32'h84a45afa;
    ram_cell[   29302] = 32'h1baaf0ec;
    ram_cell[   29303] = 32'h949f4776;
    ram_cell[   29304] = 32'h052243f2;
    ram_cell[   29305] = 32'ha5919b89;
    ram_cell[   29306] = 32'h7b6c6ae3;
    ram_cell[   29307] = 32'h9a0e9219;
    ram_cell[   29308] = 32'he6fcd8c0;
    ram_cell[   29309] = 32'hfccf4f9b;
    ram_cell[   29310] = 32'hbf9608f1;
    ram_cell[   29311] = 32'h75bfa085;
    ram_cell[   29312] = 32'he009212d;
    ram_cell[   29313] = 32'h59e63d32;
    ram_cell[   29314] = 32'hf3ee73df;
    ram_cell[   29315] = 32'h13433fbc;
    ram_cell[   29316] = 32'h89ae1297;
    ram_cell[   29317] = 32'h43e69265;
    ram_cell[   29318] = 32'h2d77ba71;
    ram_cell[   29319] = 32'h4211092e;
    ram_cell[   29320] = 32'h22ad81ff;
    ram_cell[   29321] = 32'h1a8df2ca;
    ram_cell[   29322] = 32'h25056322;
    ram_cell[   29323] = 32'h5fdad594;
    ram_cell[   29324] = 32'h61c91828;
    ram_cell[   29325] = 32'ha9ba4c59;
    ram_cell[   29326] = 32'h6c43228d;
    ram_cell[   29327] = 32'h006ded90;
    ram_cell[   29328] = 32'hb34df47e;
    ram_cell[   29329] = 32'h49b71ca2;
    ram_cell[   29330] = 32'hf77c25e0;
    ram_cell[   29331] = 32'hbff359c6;
    ram_cell[   29332] = 32'hc6fa2057;
    ram_cell[   29333] = 32'hce5a8f3f;
    ram_cell[   29334] = 32'h73632214;
    ram_cell[   29335] = 32'h197d667e;
    ram_cell[   29336] = 32'h244a24ab;
    ram_cell[   29337] = 32'h62ca980b;
    ram_cell[   29338] = 32'h3475b93a;
    ram_cell[   29339] = 32'h5b1779b1;
    ram_cell[   29340] = 32'h4b70192c;
    ram_cell[   29341] = 32'h5075e321;
    ram_cell[   29342] = 32'h8c459aca;
    ram_cell[   29343] = 32'h4437aa4a;
    ram_cell[   29344] = 32'hfd9811c5;
    ram_cell[   29345] = 32'hba13deba;
    ram_cell[   29346] = 32'h36199e48;
    ram_cell[   29347] = 32'h97424b2c;
    ram_cell[   29348] = 32'h8ee239cd;
    ram_cell[   29349] = 32'hcd514b29;
    ram_cell[   29350] = 32'h2fefcf21;
    ram_cell[   29351] = 32'h70ac885c;
    ram_cell[   29352] = 32'hd0167891;
    ram_cell[   29353] = 32'h87bbce12;
    ram_cell[   29354] = 32'hdb289a17;
    ram_cell[   29355] = 32'h1fee04ef;
    ram_cell[   29356] = 32'hc19b1140;
    ram_cell[   29357] = 32'hb50fe7d1;
    ram_cell[   29358] = 32'h614d58d8;
    ram_cell[   29359] = 32'h25a84962;
    ram_cell[   29360] = 32'h6ad9df10;
    ram_cell[   29361] = 32'h44b41317;
    ram_cell[   29362] = 32'h9b1c00b4;
    ram_cell[   29363] = 32'h60873502;
    ram_cell[   29364] = 32'ha03f55bc;
    ram_cell[   29365] = 32'h32dc55f3;
    ram_cell[   29366] = 32'h16443713;
    ram_cell[   29367] = 32'h1ecbdddc;
    ram_cell[   29368] = 32'h7909ea1e;
    ram_cell[   29369] = 32'ha2a9b78b;
    ram_cell[   29370] = 32'hc20dace9;
    ram_cell[   29371] = 32'hd5a04deb;
    ram_cell[   29372] = 32'h82cabacc;
    ram_cell[   29373] = 32'hf469a4d5;
    ram_cell[   29374] = 32'he043268d;
    ram_cell[   29375] = 32'h19466bcc;
    ram_cell[   29376] = 32'hf1a90240;
    ram_cell[   29377] = 32'hfc5246db;
    ram_cell[   29378] = 32'hfea2a633;
    ram_cell[   29379] = 32'h3aa59151;
    ram_cell[   29380] = 32'h963060c7;
    ram_cell[   29381] = 32'h530ada22;
    ram_cell[   29382] = 32'h64a6db07;
    ram_cell[   29383] = 32'h6a37c91c;
    ram_cell[   29384] = 32'h4a919473;
    ram_cell[   29385] = 32'he26d4b32;
    ram_cell[   29386] = 32'h4e95ed56;
    ram_cell[   29387] = 32'h7ec82463;
    ram_cell[   29388] = 32'h16057058;
    ram_cell[   29389] = 32'h0de940a9;
    ram_cell[   29390] = 32'h3a6ff23f;
    ram_cell[   29391] = 32'hbecb0db0;
    ram_cell[   29392] = 32'h8a2159ed;
    ram_cell[   29393] = 32'haba7f77b;
    ram_cell[   29394] = 32'h5adfcb78;
    ram_cell[   29395] = 32'h10776f22;
    ram_cell[   29396] = 32'h875c53f0;
    ram_cell[   29397] = 32'h2a708bca;
    ram_cell[   29398] = 32'he78d9f26;
    ram_cell[   29399] = 32'h60e9986e;
    ram_cell[   29400] = 32'ha5af53ab;
    ram_cell[   29401] = 32'h420bd280;
    ram_cell[   29402] = 32'h912532a4;
    ram_cell[   29403] = 32'ha4ee35c4;
    ram_cell[   29404] = 32'h54340474;
    ram_cell[   29405] = 32'he30e8d73;
    ram_cell[   29406] = 32'hb93fedeb;
    ram_cell[   29407] = 32'hb10d7fb4;
    ram_cell[   29408] = 32'h2725b149;
    ram_cell[   29409] = 32'hbeadbf39;
    ram_cell[   29410] = 32'hf81169d8;
    ram_cell[   29411] = 32'h8ea40e46;
    ram_cell[   29412] = 32'h3662b51c;
    ram_cell[   29413] = 32'ha3451e3b;
    ram_cell[   29414] = 32'h687e8895;
    ram_cell[   29415] = 32'hcf2ea9e2;
    ram_cell[   29416] = 32'h3b3556cc;
    ram_cell[   29417] = 32'h9dfd47d4;
    ram_cell[   29418] = 32'hce10066d;
    ram_cell[   29419] = 32'hc22ab7bf;
    ram_cell[   29420] = 32'h41ea9c52;
    ram_cell[   29421] = 32'h6f366a84;
    ram_cell[   29422] = 32'h95c856be;
    ram_cell[   29423] = 32'h922c1fb3;
    ram_cell[   29424] = 32'hc07ea2af;
    ram_cell[   29425] = 32'h75fb92d9;
    ram_cell[   29426] = 32'ha3e02c16;
    ram_cell[   29427] = 32'h7d7af167;
    ram_cell[   29428] = 32'hc27f73d0;
    ram_cell[   29429] = 32'h2dceb9fa;
    ram_cell[   29430] = 32'h67846149;
    ram_cell[   29431] = 32'h7bccf601;
    ram_cell[   29432] = 32'h0232eb75;
    ram_cell[   29433] = 32'h7406f7ae;
    ram_cell[   29434] = 32'h7b7eb8f7;
    ram_cell[   29435] = 32'h24c4234d;
    ram_cell[   29436] = 32'hbc2a9809;
    ram_cell[   29437] = 32'hadb0dc28;
    ram_cell[   29438] = 32'h7dee26a4;
    ram_cell[   29439] = 32'hfb473988;
    ram_cell[   29440] = 32'h2aac40e5;
    ram_cell[   29441] = 32'hccc36445;
    ram_cell[   29442] = 32'ha07afaa2;
    ram_cell[   29443] = 32'hd3a102ef;
    ram_cell[   29444] = 32'h8ae9cb4d;
    ram_cell[   29445] = 32'h96039992;
    ram_cell[   29446] = 32'h2dbd0e5a;
    ram_cell[   29447] = 32'hf9938ae3;
    ram_cell[   29448] = 32'hfaeb9f7e;
    ram_cell[   29449] = 32'hd77076f5;
    ram_cell[   29450] = 32'h8816af4e;
    ram_cell[   29451] = 32'h43576c5d;
    ram_cell[   29452] = 32'h2344ad61;
    ram_cell[   29453] = 32'h1840b945;
    ram_cell[   29454] = 32'h5342f664;
    ram_cell[   29455] = 32'hba2fcbf4;
    ram_cell[   29456] = 32'h3ab44322;
    ram_cell[   29457] = 32'hda7c1c55;
    ram_cell[   29458] = 32'h370b8d3e;
    ram_cell[   29459] = 32'hba5822bb;
    ram_cell[   29460] = 32'h9995683b;
    ram_cell[   29461] = 32'hc5e0c99b;
    ram_cell[   29462] = 32'h0a74ba88;
    ram_cell[   29463] = 32'h52022a17;
    ram_cell[   29464] = 32'haa5e1c83;
    ram_cell[   29465] = 32'hbb3bf77a;
    ram_cell[   29466] = 32'h89f5d99e;
    ram_cell[   29467] = 32'h48aee713;
    ram_cell[   29468] = 32'h23c56524;
    ram_cell[   29469] = 32'hbd2ccf40;
    ram_cell[   29470] = 32'h92c6a6c5;
    ram_cell[   29471] = 32'h1a5475e7;
    ram_cell[   29472] = 32'h5d216ba3;
    ram_cell[   29473] = 32'hb208619f;
    ram_cell[   29474] = 32'haf0716d0;
    ram_cell[   29475] = 32'hf70b1960;
    ram_cell[   29476] = 32'h051e2b90;
    ram_cell[   29477] = 32'hf4c0e4be;
    ram_cell[   29478] = 32'ha948e37c;
    ram_cell[   29479] = 32'h81c6cf6a;
    ram_cell[   29480] = 32'hc59f7930;
    ram_cell[   29481] = 32'hf80f9e91;
    ram_cell[   29482] = 32'h85ebfbce;
    ram_cell[   29483] = 32'h63175304;
    ram_cell[   29484] = 32'h614577c1;
    ram_cell[   29485] = 32'h749b34ac;
    ram_cell[   29486] = 32'hb1594ffc;
    ram_cell[   29487] = 32'hb1b1eb05;
    ram_cell[   29488] = 32'h14fb5d79;
    ram_cell[   29489] = 32'h431ff0b2;
    ram_cell[   29490] = 32'h9d4561b6;
    ram_cell[   29491] = 32'h82dbf463;
    ram_cell[   29492] = 32'hf0f2da45;
    ram_cell[   29493] = 32'h8927806a;
    ram_cell[   29494] = 32'hc3f74f78;
    ram_cell[   29495] = 32'h6a96ffbf;
    ram_cell[   29496] = 32'h743d3e1c;
    ram_cell[   29497] = 32'h15f3514b;
    ram_cell[   29498] = 32'h7d7e7917;
    ram_cell[   29499] = 32'hc83413c8;
    ram_cell[   29500] = 32'h7ab99eb3;
    ram_cell[   29501] = 32'h06886642;
    ram_cell[   29502] = 32'h09549028;
    ram_cell[   29503] = 32'h870d829c;
    ram_cell[   29504] = 32'hbc0e0b46;
    ram_cell[   29505] = 32'haa6c2aec;
    ram_cell[   29506] = 32'h68538cf4;
    ram_cell[   29507] = 32'h3e13fe8c;
    ram_cell[   29508] = 32'h40814b99;
    ram_cell[   29509] = 32'h889fe071;
    ram_cell[   29510] = 32'h53bab755;
    ram_cell[   29511] = 32'hab6c26b0;
    ram_cell[   29512] = 32'h9ead1aa0;
    ram_cell[   29513] = 32'h49958a88;
    ram_cell[   29514] = 32'hd483e39c;
    ram_cell[   29515] = 32'h40b35e19;
    ram_cell[   29516] = 32'h08eaabbf;
    ram_cell[   29517] = 32'he1a08485;
    ram_cell[   29518] = 32'h9af12b25;
    ram_cell[   29519] = 32'ha3de235e;
    ram_cell[   29520] = 32'hd4f52889;
    ram_cell[   29521] = 32'hb847681b;
    ram_cell[   29522] = 32'h172f9db8;
    ram_cell[   29523] = 32'h8565a495;
    ram_cell[   29524] = 32'h31ea4a72;
    ram_cell[   29525] = 32'h814c653a;
    ram_cell[   29526] = 32'h2faf90b8;
    ram_cell[   29527] = 32'hc8cf1d54;
    ram_cell[   29528] = 32'h3938b048;
    ram_cell[   29529] = 32'ha3507781;
    ram_cell[   29530] = 32'h1e95d978;
    ram_cell[   29531] = 32'hbdb1326f;
    ram_cell[   29532] = 32'h21646b02;
    ram_cell[   29533] = 32'h1c02db0f;
    ram_cell[   29534] = 32'h25af68dc;
    ram_cell[   29535] = 32'h2900510c;
    ram_cell[   29536] = 32'hab4ab6ed;
    ram_cell[   29537] = 32'hb8b0a34a;
    ram_cell[   29538] = 32'h4b112966;
    ram_cell[   29539] = 32'ha4beef4a;
    ram_cell[   29540] = 32'h741e33d9;
    ram_cell[   29541] = 32'he080ed4e;
    ram_cell[   29542] = 32'h66a35aa9;
    ram_cell[   29543] = 32'h3c1f53ff;
    ram_cell[   29544] = 32'h2a25b7d3;
    ram_cell[   29545] = 32'ha914bc3a;
    ram_cell[   29546] = 32'h177af7e6;
    ram_cell[   29547] = 32'h902cf8dd;
    ram_cell[   29548] = 32'hf79f3eb1;
    ram_cell[   29549] = 32'h81e2904c;
    ram_cell[   29550] = 32'h89a43ac2;
    ram_cell[   29551] = 32'h70da04e4;
    ram_cell[   29552] = 32'h2d05201c;
    ram_cell[   29553] = 32'h0b865c2d;
    ram_cell[   29554] = 32'h9d384f6b;
    ram_cell[   29555] = 32'h7802d418;
    ram_cell[   29556] = 32'hba3d772b;
    ram_cell[   29557] = 32'h88127b3b;
    ram_cell[   29558] = 32'h1767dbe0;
    ram_cell[   29559] = 32'h39d5cca0;
    ram_cell[   29560] = 32'hb1e7e7a6;
    ram_cell[   29561] = 32'hfb9c343f;
    ram_cell[   29562] = 32'h868d312a;
    ram_cell[   29563] = 32'he04bac24;
    ram_cell[   29564] = 32'h58c33586;
    ram_cell[   29565] = 32'h04fde27a;
    ram_cell[   29566] = 32'hedf37e90;
    ram_cell[   29567] = 32'h915e6be9;
    ram_cell[   29568] = 32'h5c9910f3;
    ram_cell[   29569] = 32'h6cf10be8;
    ram_cell[   29570] = 32'h03c771dc;
    ram_cell[   29571] = 32'h11be114c;
    ram_cell[   29572] = 32'hae04566f;
    ram_cell[   29573] = 32'h0c2113c2;
    ram_cell[   29574] = 32'h52404d94;
    ram_cell[   29575] = 32'h83385b51;
    ram_cell[   29576] = 32'hce248ca7;
    ram_cell[   29577] = 32'h3fc14674;
    ram_cell[   29578] = 32'had4bec49;
    ram_cell[   29579] = 32'hf6421493;
    ram_cell[   29580] = 32'hd53871de;
    ram_cell[   29581] = 32'ha23c8021;
    ram_cell[   29582] = 32'h75ea1fa4;
    ram_cell[   29583] = 32'hec2aa4e9;
    ram_cell[   29584] = 32'h5a0e7900;
    ram_cell[   29585] = 32'hbd61acce;
    ram_cell[   29586] = 32'hd67b55ca;
    ram_cell[   29587] = 32'h6ccccfd8;
    ram_cell[   29588] = 32'hb3c9f599;
    ram_cell[   29589] = 32'hbce62893;
    ram_cell[   29590] = 32'hee5403e2;
    ram_cell[   29591] = 32'h5b1ec90d;
    ram_cell[   29592] = 32'h0c47d5e3;
    ram_cell[   29593] = 32'hf0d5781a;
    ram_cell[   29594] = 32'h3323408b;
    ram_cell[   29595] = 32'h39e2f6a2;
    ram_cell[   29596] = 32'h07926ab3;
    ram_cell[   29597] = 32'h4176e6b7;
    ram_cell[   29598] = 32'hcdf3fe20;
    ram_cell[   29599] = 32'h45158d46;
    ram_cell[   29600] = 32'ha32b6d94;
    ram_cell[   29601] = 32'h1744f1ff;
    ram_cell[   29602] = 32'h49552e52;
    ram_cell[   29603] = 32'h6825a920;
    ram_cell[   29604] = 32'hd7ea0e18;
    ram_cell[   29605] = 32'h47306a56;
    ram_cell[   29606] = 32'hba7e6df3;
    ram_cell[   29607] = 32'h29fed9d1;
    ram_cell[   29608] = 32'h5f6ef724;
    ram_cell[   29609] = 32'h231d46e1;
    ram_cell[   29610] = 32'h22d61825;
    ram_cell[   29611] = 32'hfa83cb74;
    ram_cell[   29612] = 32'h31efed0f;
    ram_cell[   29613] = 32'hacf528bb;
    ram_cell[   29614] = 32'h29428259;
    ram_cell[   29615] = 32'h7084a926;
    ram_cell[   29616] = 32'h8d70a29a;
    ram_cell[   29617] = 32'h6d82d177;
    ram_cell[   29618] = 32'hb617560c;
    ram_cell[   29619] = 32'hf1194b1c;
    ram_cell[   29620] = 32'h6205ab58;
    ram_cell[   29621] = 32'he662807b;
    ram_cell[   29622] = 32'h6a899bfe;
    ram_cell[   29623] = 32'h1a7fa046;
    ram_cell[   29624] = 32'h9fcf5fdb;
    ram_cell[   29625] = 32'haa48d8d2;
    ram_cell[   29626] = 32'h4de5a350;
    ram_cell[   29627] = 32'h4b33c6b3;
    ram_cell[   29628] = 32'h36c5f5c9;
    ram_cell[   29629] = 32'ha8802aeb;
    ram_cell[   29630] = 32'hd9d883a5;
    ram_cell[   29631] = 32'h3892e213;
    ram_cell[   29632] = 32'h2ecf4e65;
    ram_cell[   29633] = 32'h07a66b85;
    ram_cell[   29634] = 32'h575b4c41;
    ram_cell[   29635] = 32'h14b8a6b9;
    ram_cell[   29636] = 32'hb3bbfc7d;
    ram_cell[   29637] = 32'heb33e5f2;
    ram_cell[   29638] = 32'h54348f84;
    ram_cell[   29639] = 32'h6573e043;
    ram_cell[   29640] = 32'h46651289;
    ram_cell[   29641] = 32'h726ff0fc;
    ram_cell[   29642] = 32'h1a4c5aed;
    ram_cell[   29643] = 32'h38fed1a9;
    ram_cell[   29644] = 32'h1c51abbb;
    ram_cell[   29645] = 32'hb35afb01;
    ram_cell[   29646] = 32'hd3285c05;
    ram_cell[   29647] = 32'h96af9160;
    ram_cell[   29648] = 32'h2992a7f4;
    ram_cell[   29649] = 32'h512f6254;
    ram_cell[   29650] = 32'h2d03a84f;
    ram_cell[   29651] = 32'h0801c7d7;
    ram_cell[   29652] = 32'ha1d2e2cd;
    ram_cell[   29653] = 32'h9c6a51db;
    ram_cell[   29654] = 32'ha51d2a2b;
    ram_cell[   29655] = 32'h8de031cf;
    ram_cell[   29656] = 32'h3278bb10;
    ram_cell[   29657] = 32'hf1db0803;
    ram_cell[   29658] = 32'hd39b7e9a;
    ram_cell[   29659] = 32'h528e9cb9;
    ram_cell[   29660] = 32'h2f081154;
    ram_cell[   29661] = 32'h2c9576ae;
    ram_cell[   29662] = 32'h40f4975e;
    ram_cell[   29663] = 32'h25ff2095;
    ram_cell[   29664] = 32'h2734e612;
    ram_cell[   29665] = 32'hf50c19b9;
    ram_cell[   29666] = 32'h3125ebd2;
    ram_cell[   29667] = 32'h85477f65;
    ram_cell[   29668] = 32'h5f55bb9b;
    ram_cell[   29669] = 32'h5ec6b17c;
    ram_cell[   29670] = 32'hb2f3d878;
    ram_cell[   29671] = 32'h317d8b4b;
    ram_cell[   29672] = 32'h21861259;
    ram_cell[   29673] = 32'h8a8ab2e3;
    ram_cell[   29674] = 32'hc64082f0;
    ram_cell[   29675] = 32'h1f8f9a2e;
    ram_cell[   29676] = 32'h0904ae73;
    ram_cell[   29677] = 32'h7811e2f2;
    ram_cell[   29678] = 32'hc6159a43;
    ram_cell[   29679] = 32'h141445e4;
    ram_cell[   29680] = 32'h99440b17;
    ram_cell[   29681] = 32'hdf1737c8;
    ram_cell[   29682] = 32'h27cfb948;
    ram_cell[   29683] = 32'h409b6437;
    ram_cell[   29684] = 32'h80741504;
    ram_cell[   29685] = 32'h05246558;
    ram_cell[   29686] = 32'hde1208b7;
    ram_cell[   29687] = 32'h9122e1cd;
    ram_cell[   29688] = 32'hd87027d2;
    ram_cell[   29689] = 32'ha8dd05a3;
    ram_cell[   29690] = 32'h3697e7cc;
    ram_cell[   29691] = 32'h8901de91;
    ram_cell[   29692] = 32'haa9a83e7;
    ram_cell[   29693] = 32'h15f9ae29;
    ram_cell[   29694] = 32'hc5baf317;
    ram_cell[   29695] = 32'h1dc8e514;
    ram_cell[   29696] = 32'h9cf0c67e;
    ram_cell[   29697] = 32'h38ba0ce5;
    ram_cell[   29698] = 32'h5c27f049;
    ram_cell[   29699] = 32'hf3070abc;
    ram_cell[   29700] = 32'h0e1a8efd;
    ram_cell[   29701] = 32'h21833341;
    ram_cell[   29702] = 32'ha27fc80b;
    ram_cell[   29703] = 32'he54be920;
    ram_cell[   29704] = 32'h24706304;
    ram_cell[   29705] = 32'h9cdb5f2a;
    ram_cell[   29706] = 32'h2923a7f0;
    ram_cell[   29707] = 32'h381c3dc3;
    ram_cell[   29708] = 32'hd110527e;
    ram_cell[   29709] = 32'h4bf15302;
    ram_cell[   29710] = 32'hd474382b;
    ram_cell[   29711] = 32'ha47cb481;
    ram_cell[   29712] = 32'h44faec08;
    ram_cell[   29713] = 32'hc4514605;
    ram_cell[   29714] = 32'h7738d652;
    ram_cell[   29715] = 32'h4c3e9797;
    ram_cell[   29716] = 32'h8c3231fc;
    ram_cell[   29717] = 32'hb52b0cef;
    ram_cell[   29718] = 32'h12210441;
    ram_cell[   29719] = 32'h4556fab9;
    ram_cell[   29720] = 32'h013ac98d;
    ram_cell[   29721] = 32'haaea71c7;
    ram_cell[   29722] = 32'hfa1f02a7;
    ram_cell[   29723] = 32'he4c38e69;
    ram_cell[   29724] = 32'hec93aa38;
    ram_cell[   29725] = 32'hecd71fcc;
    ram_cell[   29726] = 32'h88c8c23d;
    ram_cell[   29727] = 32'h3e5709fc;
    ram_cell[   29728] = 32'h0a752d84;
    ram_cell[   29729] = 32'h31de0344;
    ram_cell[   29730] = 32'hacc41a5a;
    ram_cell[   29731] = 32'he98f2da5;
    ram_cell[   29732] = 32'h690ea05c;
    ram_cell[   29733] = 32'h07936ddf;
    ram_cell[   29734] = 32'hb7df96bd;
    ram_cell[   29735] = 32'hb33accf8;
    ram_cell[   29736] = 32'hf0284405;
    ram_cell[   29737] = 32'h9dec6e7d;
    ram_cell[   29738] = 32'hd2ef8baf;
    ram_cell[   29739] = 32'had99a9b2;
    ram_cell[   29740] = 32'h9e701acd;
    ram_cell[   29741] = 32'h4f73b51d;
    ram_cell[   29742] = 32'hb5e196a9;
    ram_cell[   29743] = 32'h17bfb30f;
    ram_cell[   29744] = 32'h627bb268;
    ram_cell[   29745] = 32'h441ad0b0;
    ram_cell[   29746] = 32'hefc018c1;
    ram_cell[   29747] = 32'h92a90269;
    ram_cell[   29748] = 32'hd78aa5eb;
    ram_cell[   29749] = 32'hff46a598;
    ram_cell[   29750] = 32'h2cb51704;
    ram_cell[   29751] = 32'h763918aa;
    ram_cell[   29752] = 32'h728a44b9;
    ram_cell[   29753] = 32'h99c0fc0c;
    ram_cell[   29754] = 32'hc97a6a6d;
    ram_cell[   29755] = 32'hdbe604b9;
    ram_cell[   29756] = 32'h52182c99;
    ram_cell[   29757] = 32'hde6e251f;
    ram_cell[   29758] = 32'hc5284029;
    ram_cell[   29759] = 32'hfc08d787;
    ram_cell[   29760] = 32'hb1c1caaa;
    ram_cell[   29761] = 32'hbc120bb1;
    ram_cell[   29762] = 32'hbfbfe0e5;
    ram_cell[   29763] = 32'h84acb7f7;
    ram_cell[   29764] = 32'h9fc424c0;
    ram_cell[   29765] = 32'h1930246c;
    ram_cell[   29766] = 32'h32431761;
    ram_cell[   29767] = 32'hb511bff6;
    ram_cell[   29768] = 32'hd93470d4;
    ram_cell[   29769] = 32'h3ca4c296;
    ram_cell[   29770] = 32'hea34bf3f;
    ram_cell[   29771] = 32'hf975c8ce;
    ram_cell[   29772] = 32'hce832e78;
    ram_cell[   29773] = 32'h601cbac8;
    ram_cell[   29774] = 32'h98a29461;
    ram_cell[   29775] = 32'heec955d6;
    ram_cell[   29776] = 32'h6ee45248;
    ram_cell[   29777] = 32'h28e6c9e3;
    ram_cell[   29778] = 32'h03f5c48e;
    ram_cell[   29779] = 32'ha9f56d80;
    ram_cell[   29780] = 32'h39699b51;
    ram_cell[   29781] = 32'heb24c8f3;
    ram_cell[   29782] = 32'h6acae9b2;
    ram_cell[   29783] = 32'hb93a43bb;
    ram_cell[   29784] = 32'h93b6e598;
    ram_cell[   29785] = 32'h54bf8cdd;
    ram_cell[   29786] = 32'h679927a8;
    ram_cell[   29787] = 32'h4c7dff50;
    ram_cell[   29788] = 32'h0cc6c8c9;
    ram_cell[   29789] = 32'h42422e27;
    ram_cell[   29790] = 32'h25a078e3;
    ram_cell[   29791] = 32'hc9a1cf5a;
    ram_cell[   29792] = 32'hb2fb705b;
    ram_cell[   29793] = 32'hefe8aec0;
    ram_cell[   29794] = 32'h0db6917b;
    ram_cell[   29795] = 32'h9f20fc9b;
    ram_cell[   29796] = 32'h21a7d432;
    ram_cell[   29797] = 32'ha4aa73da;
    ram_cell[   29798] = 32'h91fd8643;
    ram_cell[   29799] = 32'h9e28fb04;
    ram_cell[   29800] = 32'hbbd8553f;
    ram_cell[   29801] = 32'h04a2dfbe;
    ram_cell[   29802] = 32'h3554fcb1;
    ram_cell[   29803] = 32'hf23997b8;
    ram_cell[   29804] = 32'had735330;
    ram_cell[   29805] = 32'h767d713a;
    ram_cell[   29806] = 32'h03b67d02;
    ram_cell[   29807] = 32'hb39d2c1a;
    ram_cell[   29808] = 32'hfea1d658;
    ram_cell[   29809] = 32'h60f8826d;
    ram_cell[   29810] = 32'hb5872705;
    ram_cell[   29811] = 32'hb4453587;
    ram_cell[   29812] = 32'h9bec082c;
    ram_cell[   29813] = 32'hef7ae329;
    ram_cell[   29814] = 32'ha70c0a7c;
    ram_cell[   29815] = 32'h84c09dc1;
    ram_cell[   29816] = 32'hb39dd819;
    ram_cell[   29817] = 32'hc7435dbb;
    ram_cell[   29818] = 32'ha314778b;
    ram_cell[   29819] = 32'hf1452046;
    ram_cell[   29820] = 32'he80068d3;
    ram_cell[   29821] = 32'h01ed9c7b;
    ram_cell[   29822] = 32'ha9c9ae53;
    ram_cell[   29823] = 32'h783e20d9;
    ram_cell[   29824] = 32'h7259d6a1;
    ram_cell[   29825] = 32'h5e8dfbe3;
    ram_cell[   29826] = 32'h2ef14605;
    ram_cell[   29827] = 32'h0ef374ad;
    ram_cell[   29828] = 32'h462f0229;
    ram_cell[   29829] = 32'hec6e3b22;
    ram_cell[   29830] = 32'hdb901a2d;
    ram_cell[   29831] = 32'h62d02c15;
    ram_cell[   29832] = 32'hde3efe1a;
    ram_cell[   29833] = 32'h3787cd8d;
    ram_cell[   29834] = 32'hfe9bb2be;
    ram_cell[   29835] = 32'h6519c6a8;
    ram_cell[   29836] = 32'ha6cb54ff;
    ram_cell[   29837] = 32'h4ea1720f;
    ram_cell[   29838] = 32'h37b22e68;
    ram_cell[   29839] = 32'hff688409;
    ram_cell[   29840] = 32'hc2722726;
    ram_cell[   29841] = 32'h18292888;
    ram_cell[   29842] = 32'h95ace19c;
    ram_cell[   29843] = 32'h5de4787b;
    ram_cell[   29844] = 32'haed92768;
    ram_cell[   29845] = 32'h9b10d21e;
    ram_cell[   29846] = 32'hc11a6f78;
    ram_cell[   29847] = 32'h733ef7fd;
    ram_cell[   29848] = 32'h0bde548d;
    ram_cell[   29849] = 32'h8a1bf6d2;
    ram_cell[   29850] = 32'hcec7ba79;
    ram_cell[   29851] = 32'hcc1edc9d;
    ram_cell[   29852] = 32'haa3f6264;
    ram_cell[   29853] = 32'h8eebb8c4;
    ram_cell[   29854] = 32'hb3d48d64;
    ram_cell[   29855] = 32'h81ad2e33;
    ram_cell[   29856] = 32'h3c2be09b;
    ram_cell[   29857] = 32'h636da8b0;
    ram_cell[   29858] = 32'hc7ec44dd;
    ram_cell[   29859] = 32'h93d5a170;
    ram_cell[   29860] = 32'haeb8ff6c;
    ram_cell[   29861] = 32'hfd803ee3;
    ram_cell[   29862] = 32'h73eadb34;
    ram_cell[   29863] = 32'hc33b43c7;
    ram_cell[   29864] = 32'h0e5233dc;
    ram_cell[   29865] = 32'hc3a0b3cc;
    ram_cell[   29866] = 32'h9e7283b6;
    ram_cell[   29867] = 32'ha160a3b1;
    ram_cell[   29868] = 32'ha02f9ee5;
    ram_cell[   29869] = 32'h71980462;
    ram_cell[   29870] = 32'h8ac62f78;
    ram_cell[   29871] = 32'hccfa95a0;
    ram_cell[   29872] = 32'hb32d60c0;
    ram_cell[   29873] = 32'h1ab14a6c;
    ram_cell[   29874] = 32'h4919db58;
    ram_cell[   29875] = 32'h58328f40;
    ram_cell[   29876] = 32'hf67f5cbc;
    ram_cell[   29877] = 32'h29bf4281;
    ram_cell[   29878] = 32'h60db1516;
    ram_cell[   29879] = 32'h6cf8b716;
    ram_cell[   29880] = 32'he3e4f600;
    ram_cell[   29881] = 32'h6d0eed5a;
    ram_cell[   29882] = 32'h6961edec;
    ram_cell[   29883] = 32'h1fea79bf;
    ram_cell[   29884] = 32'ha2baea40;
    ram_cell[   29885] = 32'h6aeebefb;
    ram_cell[   29886] = 32'h3ac3827d;
    ram_cell[   29887] = 32'hc86ea784;
    ram_cell[   29888] = 32'ha383a1fa;
    ram_cell[   29889] = 32'h77ea40ce;
    ram_cell[   29890] = 32'h1278b6b6;
    ram_cell[   29891] = 32'h5b415085;
    ram_cell[   29892] = 32'h4179f8a2;
    ram_cell[   29893] = 32'h93f39248;
    ram_cell[   29894] = 32'h1147bc39;
    ram_cell[   29895] = 32'h39636471;
    ram_cell[   29896] = 32'h1af50fda;
    ram_cell[   29897] = 32'h612ed598;
    ram_cell[   29898] = 32'h71e8b668;
    ram_cell[   29899] = 32'hb04d8a55;
    ram_cell[   29900] = 32'h8a99d174;
    ram_cell[   29901] = 32'hb17bb4a6;
    ram_cell[   29902] = 32'haeed8d00;
    ram_cell[   29903] = 32'h7e8502b5;
    ram_cell[   29904] = 32'h88acd636;
    ram_cell[   29905] = 32'hc89870b0;
    ram_cell[   29906] = 32'h1bbd8fcb;
    ram_cell[   29907] = 32'h006ea0d6;
    ram_cell[   29908] = 32'hc406c854;
    ram_cell[   29909] = 32'hdd6e5495;
    ram_cell[   29910] = 32'h528c6e2d;
    ram_cell[   29911] = 32'h767e1881;
    ram_cell[   29912] = 32'h1adc3f10;
    ram_cell[   29913] = 32'he4266f00;
    ram_cell[   29914] = 32'h2be835bf;
    ram_cell[   29915] = 32'hb939e487;
    ram_cell[   29916] = 32'h047ce3fa;
    ram_cell[   29917] = 32'h75ade7fe;
    ram_cell[   29918] = 32'hec1d8896;
    ram_cell[   29919] = 32'ha48c387a;
    ram_cell[   29920] = 32'h206e094f;
    ram_cell[   29921] = 32'h56ffaa7b;
    ram_cell[   29922] = 32'ha52beb67;
    ram_cell[   29923] = 32'h9a2e74ce;
    ram_cell[   29924] = 32'h8496fa2f;
    ram_cell[   29925] = 32'hf7b2060c;
    ram_cell[   29926] = 32'he790af8b;
    ram_cell[   29927] = 32'h2fbac73f;
    ram_cell[   29928] = 32'h608fed48;
    ram_cell[   29929] = 32'h42ea1b9f;
    ram_cell[   29930] = 32'h4566d6e2;
    ram_cell[   29931] = 32'h816569e9;
    ram_cell[   29932] = 32'hd17094a0;
    ram_cell[   29933] = 32'hf312f4bc;
    ram_cell[   29934] = 32'h62128692;
    ram_cell[   29935] = 32'hc2c1946e;
    ram_cell[   29936] = 32'h4292416f;
    ram_cell[   29937] = 32'h026c0875;
    ram_cell[   29938] = 32'hd79d0d0f;
    ram_cell[   29939] = 32'hf7bdddcb;
    ram_cell[   29940] = 32'he469a929;
    ram_cell[   29941] = 32'h3efce0bd;
    ram_cell[   29942] = 32'h0024fdef;
    ram_cell[   29943] = 32'h99212155;
    ram_cell[   29944] = 32'hf35c26af;
    ram_cell[   29945] = 32'hebd787df;
    ram_cell[   29946] = 32'hb62af260;
    ram_cell[   29947] = 32'h5c984767;
    ram_cell[   29948] = 32'ha989d90d;
    ram_cell[   29949] = 32'h22aa3348;
    ram_cell[   29950] = 32'h4d7c2604;
    ram_cell[   29951] = 32'hb99b7a35;
    ram_cell[   29952] = 32'h823e17e2;
    ram_cell[   29953] = 32'h5a397006;
    ram_cell[   29954] = 32'h6d3b054c;
    ram_cell[   29955] = 32'h9e772bb4;
    ram_cell[   29956] = 32'hb81cd9d7;
    ram_cell[   29957] = 32'h12d2b7b0;
    ram_cell[   29958] = 32'h4cc4fedd;
    ram_cell[   29959] = 32'hd6d4eb6e;
    ram_cell[   29960] = 32'h0cd49700;
    ram_cell[   29961] = 32'h8511cfc9;
    ram_cell[   29962] = 32'hb310568e;
    ram_cell[   29963] = 32'hf0965c3a;
    ram_cell[   29964] = 32'hd3326751;
    ram_cell[   29965] = 32'h41de9cfc;
    ram_cell[   29966] = 32'h2cb92a01;
    ram_cell[   29967] = 32'h28a593c1;
    ram_cell[   29968] = 32'hb39b7f17;
    ram_cell[   29969] = 32'h184c326b;
    ram_cell[   29970] = 32'h3f055d8f;
    ram_cell[   29971] = 32'h77051bd7;
    ram_cell[   29972] = 32'h8aa15424;
    ram_cell[   29973] = 32'hbe00fac6;
    ram_cell[   29974] = 32'he02c75ce;
    ram_cell[   29975] = 32'h4f53d649;
    ram_cell[   29976] = 32'h0da3b493;
    ram_cell[   29977] = 32'h7f495387;
    ram_cell[   29978] = 32'hf4f32c54;
    ram_cell[   29979] = 32'h25586e07;
    ram_cell[   29980] = 32'hef13c80a;
    ram_cell[   29981] = 32'h7497432c;
    ram_cell[   29982] = 32'h4ea74eeb;
    ram_cell[   29983] = 32'hfd71e200;
    ram_cell[   29984] = 32'h54e8d45d;
    ram_cell[   29985] = 32'hdb1b40f6;
    ram_cell[   29986] = 32'h1af58701;
    ram_cell[   29987] = 32'he674f7fd;
    ram_cell[   29988] = 32'h433b9b46;
    ram_cell[   29989] = 32'h2993d856;
    ram_cell[   29990] = 32'h7b4bde19;
    ram_cell[   29991] = 32'h66a6e266;
    ram_cell[   29992] = 32'h58c1a762;
    ram_cell[   29993] = 32'h84aedaad;
    ram_cell[   29994] = 32'hd5b42c35;
    ram_cell[   29995] = 32'h8f8cd9d6;
    ram_cell[   29996] = 32'ha5e82d4d;
    ram_cell[   29997] = 32'he0601abc;
    ram_cell[   29998] = 32'hec3c1b59;
    ram_cell[   29999] = 32'h1a46cef3;
    ram_cell[   30000] = 32'h4dbf2baa;
    ram_cell[   30001] = 32'h145c4b2e;
    ram_cell[   30002] = 32'h94e1285f;
    ram_cell[   30003] = 32'h09d4f3a2;
    ram_cell[   30004] = 32'h1012eacd;
    ram_cell[   30005] = 32'heaa918df;
    ram_cell[   30006] = 32'h82fdad38;
    ram_cell[   30007] = 32'hbde4b4c8;
    ram_cell[   30008] = 32'h99c67ea4;
    ram_cell[   30009] = 32'h1f2c8b69;
    ram_cell[   30010] = 32'hcfe74da5;
    ram_cell[   30011] = 32'hd32b0c10;
    ram_cell[   30012] = 32'h33aeee2e;
    ram_cell[   30013] = 32'h354f5d0f;
    ram_cell[   30014] = 32'h072ed671;
    ram_cell[   30015] = 32'he1e8108b;
    ram_cell[   30016] = 32'h1d76fb71;
    ram_cell[   30017] = 32'h27ce7b6f;
    ram_cell[   30018] = 32'h8693efd2;
    ram_cell[   30019] = 32'he3eb35b7;
    ram_cell[   30020] = 32'h58a90099;
    ram_cell[   30021] = 32'h0c8857f2;
    ram_cell[   30022] = 32'h224983dc;
    ram_cell[   30023] = 32'h3a94ae16;
    ram_cell[   30024] = 32'h5e18d43a;
    ram_cell[   30025] = 32'h53bbe483;
    ram_cell[   30026] = 32'ha6b7bd7c;
    ram_cell[   30027] = 32'h8858b100;
    ram_cell[   30028] = 32'h2c751c10;
    ram_cell[   30029] = 32'h46750082;
    ram_cell[   30030] = 32'hb8006427;
    ram_cell[   30031] = 32'hfde4bf5c;
    ram_cell[   30032] = 32'h00aa5989;
    ram_cell[   30033] = 32'h9ab25203;
    ram_cell[   30034] = 32'hb523bd21;
    ram_cell[   30035] = 32'h6d31e4af;
    ram_cell[   30036] = 32'h7c1cde89;
    ram_cell[   30037] = 32'h6361c531;
    ram_cell[   30038] = 32'h552be8c0;
    ram_cell[   30039] = 32'h67d78737;
    ram_cell[   30040] = 32'h15ab0efa;
    ram_cell[   30041] = 32'h9c1dd42e;
    ram_cell[   30042] = 32'h5426ba7e;
    ram_cell[   30043] = 32'h4af17efe;
    ram_cell[   30044] = 32'h7dbdd7c4;
    ram_cell[   30045] = 32'h54a601f7;
    ram_cell[   30046] = 32'h295680c6;
    ram_cell[   30047] = 32'h44660fe0;
    ram_cell[   30048] = 32'heb4b8809;
    ram_cell[   30049] = 32'h22a85cd5;
    ram_cell[   30050] = 32'h5d3bd99a;
    ram_cell[   30051] = 32'h8f132140;
    ram_cell[   30052] = 32'h2c2b8cba;
    ram_cell[   30053] = 32'h6464fe56;
    ram_cell[   30054] = 32'h007d35ec;
    ram_cell[   30055] = 32'h8da5c0a4;
    ram_cell[   30056] = 32'h80df582b;
    ram_cell[   30057] = 32'h0d3a5c22;
    ram_cell[   30058] = 32'h0545d692;
    ram_cell[   30059] = 32'h8b33c9b7;
    ram_cell[   30060] = 32'h75f1a1e5;
    ram_cell[   30061] = 32'h1979ee9e;
    ram_cell[   30062] = 32'h2e8abe4b;
    ram_cell[   30063] = 32'h8436b3b1;
    ram_cell[   30064] = 32'h2a470756;
    ram_cell[   30065] = 32'hb87eefbc;
    ram_cell[   30066] = 32'h90f749d7;
    ram_cell[   30067] = 32'h18ca5eac;
    ram_cell[   30068] = 32'h36efc066;
    ram_cell[   30069] = 32'h9a690416;
    ram_cell[   30070] = 32'h976720a7;
    ram_cell[   30071] = 32'h62f36a98;
    ram_cell[   30072] = 32'hb1ad4dae;
    ram_cell[   30073] = 32'h0a3d1e3f;
    ram_cell[   30074] = 32'he4059980;
    ram_cell[   30075] = 32'hbc7a3e1d;
    ram_cell[   30076] = 32'hda3cff60;
    ram_cell[   30077] = 32'h5d58ee62;
    ram_cell[   30078] = 32'h3d33a065;
    ram_cell[   30079] = 32'hcfbec1a0;
    ram_cell[   30080] = 32'he6fc94b8;
    ram_cell[   30081] = 32'hf84f6e9e;
    ram_cell[   30082] = 32'hd4b699b7;
    ram_cell[   30083] = 32'h99863776;
    ram_cell[   30084] = 32'h0aba7f65;
    ram_cell[   30085] = 32'h5dcf858c;
    ram_cell[   30086] = 32'hf17f7e3f;
    ram_cell[   30087] = 32'h42a39289;
    ram_cell[   30088] = 32'h06294fc6;
    ram_cell[   30089] = 32'h526aa9d4;
    ram_cell[   30090] = 32'h31d4a20f;
    ram_cell[   30091] = 32'ha81e79c5;
    ram_cell[   30092] = 32'h3a45597b;
    ram_cell[   30093] = 32'h56a66660;
    ram_cell[   30094] = 32'h4a99a63e;
    ram_cell[   30095] = 32'h0252a0d4;
    ram_cell[   30096] = 32'h4be3b91d;
    ram_cell[   30097] = 32'h5f35771f;
    ram_cell[   30098] = 32'h872c5996;
    ram_cell[   30099] = 32'hd87bb54a;
    ram_cell[   30100] = 32'hdc88874b;
    ram_cell[   30101] = 32'hb35b7a8d;
    ram_cell[   30102] = 32'h0da41f7c;
    ram_cell[   30103] = 32'h36679198;
    ram_cell[   30104] = 32'h6f02a518;
    ram_cell[   30105] = 32'h3e2e97c4;
    ram_cell[   30106] = 32'h8229530d;
    ram_cell[   30107] = 32'hffe43cc3;
    ram_cell[   30108] = 32'h6ff390f6;
    ram_cell[   30109] = 32'ha9d3f0bf;
    ram_cell[   30110] = 32'h15b0c8fc;
    ram_cell[   30111] = 32'h40d4637e;
    ram_cell[   30112] = 32'ha57b4283;
    ram_cell[   30113] = 32'hc2b2c423;
    ram_cell[   30114] = 32'h32cc39cc;
    ram_cell[   30115] = 32'hb511ad4b;
    ram_cell[   30116] = 32'h057551ef;
    ram_cell[   30117] = 32'h26afde86;
    ram_cell[   30118] = 32'hca6dc807;
    ram_cell[   30119] = 32'hb1e0af69;
    ram_cell[   30120] = 32'h923d69c5;
    ram_cell[   30121] = 32'heb01b8a9;
    ram_cell[   30122] = 32'he80e599a;
    ram_cell[   30123] = 32'h28634d0f;
    ram_cell[   30124] = 32'hcf2ecb7c;
    ram_cell[   30125] = 32'h53c74f18;
    ram_cell[   30126] = 32'hf9f544a7;
    ram_cell[   30127] = 32'hb9d38d1a;
    ram_cell[   30128] = 32'hd078b105;
    ram_cell[   30129] = 32'h09c63f17;
    ram_cell[   30130] = 32'h6d572f83;
    ram_cell[   30131] = 32'h96549731;
    ram_cell[   30132] = 32'hc7c8728a;
    ram_cell[   30133] = 32'h3284ab15;
    ram_cell[   30134] = 32'hd2c8c265;
    ram_cell[   30135] = 32'h4233d113;
    ram_cell[   30136] = 32'h45e5f828;
    ram_cell[   30137] = 32'hdf022298;
    ram_cell[   30138] = 32'h86d66f65;
    ram_cell[   30139] = 32'h10d3802e;
    ram_cell[   30140] = 32'h5f39e1a9;
    ram_cell[   30141] = 32'h3c917fac;
    ram_cell[   30142] = 32'h95a4f19b;
    ram_cell[   30143] = 32'h00b67056;
    ram_cell[   30144] = 32'h4c7da32d;
    ram_cell[   30145] = 32'hee86ffb2;
    ram_cell[   30146] = 32'h95c12b0d;
    ram_cell[   30147] = 32'hb56997e7;
    ram_cell[   30148] = 32'h5fd22d00;
    ram_cell[   30149] = 32'hc9fa8b77;
    ram_cell[   30150] = 32'h01d71356;
    ram_cell[   30151] = 32'h267e3d4f;
    ram_cell[   30152] = 32'h667e2791;
    ram_cell[   30153] = 32'h0e42f9cd;
    ram_cell[   30154] = 32'h31604371;
    ram_cell[   30155] = 32'h8d6b5ddf;
    ram_cell[   30156] = 32'h008ffd83;
    ram_cell[   30157] = 32'hb66e665e;
    ram_cell[   30158] = 32'ha135eb3e;
    ram_cell[   30159] = 32'h73fd376b;
    ram_cell[   30160] = 32'h3940b630;
    ram_cell[   30161] = 32'h889e2bd2;
    ram_cell[   30162] = 32'he8010874;
    ram_cell[   30163] = 32'h68c23023;
    ram_cell[   30164] = 32'h96e88fa7;
    ram_cell[   30165] = 32'hfac47eb2;
    ram_cell[   30166] = 32'hf1cbbed6;
    ram_cell[   30167] = 32'h29c0acd4;
    ram_cell[   30168] = 32'h145efdb0;
    ram_cell[   30169] = 32'h06326f29;
    ram_cell[   30170] = 32'h36f4f8f0;
    ram_cell[   30171] = 32'h575b9f7f;
    ram_cell[   30172] = 32'hd0f88a60;
    ram_cell[   30173] = 32'he7fcf141;
    ram_cell[   30174] = 32'h9faeee54;
    ram_cell[   30175] = 32'h7cac9a08;
    ram_cell[   30176] = 32'h14a882d4;
    ram_cell[   30177] = 32'h2fe72ef9;
    ram_cell[   30178] = 32'h6e5c7fcf;
    ram_cell[   30179] = 32'h00a6c604;
    ram_cell[   30180] = 32'h8d967d6e;
    ram_cell[   30181] = 32'h62157206;
    ram_cell[   30182] = 32'h48eabf3a;
    ram_cell[   30183] = 32'h906f8bd9;
    ram_cell[   30184] = 32'hbeaa399b;
    ram_cell[   30185] = 32'hba01fc57;
    ram_cell[   30186] = 32'h106e5245;
    ram_cell[   30187] = 32'h85ca67e7;
    ram_cell[   30188] = 32'h3e2fe730;
    ram_cell[   30189] = 32'hff4f3a9e;
    ram_cell[   30190] = 32'h0dcf0032;
    ram_cell[   30191] = 32'he60247e6;
    ram_cell[   30192] = 32'h5b9c820f;
    ram_cell[   30193] = 32'hb4b1ca6a;
    ram_cell[   30194] = 32'h3c440d4f;
    ram_cell[   30195] = 32'h4112215c;
    ram_cell[   30196] = 32'h681379e8;
    ram_cell[   30197] = 32'hc70991c6;
    ram_cell[   30198] = 32'h1a4360e6;
    ram_cell[   30199] = 32'h3e2552e4;
    ram_cell[   30200] = 32'h2d70e404;
    ram_cell[   30201] = 32'h5335bd4f;
    ram_cell[   30202] = 32'h2506d64e;
    ram_cell[   30203] = 32'h4a123dd8;
    ram_cell[   30204] = 32'hb124c25d;
    ram_cell[   30205] = 32'h415fd187;
    ram_cell[   30206] = 32'h4858ecb1;
    ram_cell[   30207] = 32'habcca189;
    ram_cell[   30208] = 32'h1572cd98;
    ram_cell[   30209] = 32'haa9404e1;
    ram_cell[   30210] = 32'hb952efbd;
    ram_cell[   30211] = 32'hc43bf6c0;
    ram_cell[   30212] = 32'hdda59131;
    ram_cell[   30213] = 32'h9d60d599;
    ram_cell[   30214] = 32'hb917220d;
    ram_cell[   30215] = 32'h031c40f1;
    ram_cell[   30216] = 32'ha9206859;
    ram_cell[   30217] = 32'h6b801669;
    ram_cell[   30218] = 32'hb8553455;
    ram_cell[   30219] = 32'h27f7cef1;
    ram_cell[   30220] = 32'h5c0f09a1;
    ram_cell[   30221] = 32'h89d9814e;
    ram_cell[   30222] = 32'he8068649;
    ram_cell[   30223] = 32'he8a553ab;
    ram_cell[   30224] = 32'h7e769356;
    ram_cell[   30225] = 32'hd33d4945;
    ram_cell[   30226] = 32'h457154ea;
    ram_cell[   30227] = 32'h5168f3cf;
    ram_cell[   30228] = 32'h6acdd25e;
    ram_cell[   30229] = 32'h911ea35c;
    ram_cell[   30230] = 32'ha27a2ca8;
    ram_cell[   30231] = 32'h9bcdad7f;
    ram_cell[   30232] = 32'h69ce6286;
    ram_cell[   30233] = 32'h45f04e96;
    ram_cell[   30234] = 32'h0827ba14;
    ram_cell[   30235] = 32'h4a376d23;
    ram_cell[   30236] = 32'h113032ef;
    ram_cell[   30237] = 32'h0d84e11e;
    ram_cell[   30238] = 32'h59524602;
    ram_cell[   30239] = 32'h41058751;
    ram_cell[   30240] = 32'ha7fb1feb;
    ram_cell[   30241] = 32'he8fa7ae8;
    ram_cell[   30242] = 32'h57a33fdb;
    ram_cell[   30243] = 32'h4876d4d5;
    ram_cell[   30244] = 32'h943e530f;
    ram_cell[   30245] = 32'h7b4b8120;
    ram_cell[   30246] = 32'h88fc0ada;
    ram_cell[   30247] = 32'hccbc46a0;
    ram_cell[   30248] = 32'h857b4e44;
    ram_cell[   30249] = 32'h95a731b0;
    ram_cell[   30250] = 32'h12ebdf21;
    ram_cell[   30251] = 32'h821bff72;
    ram_cell[   30252] = 32'hfe2c72f1;
    ram_cell[   30253] = 32'h50e08fe5;
    ram_cell[   30254] = 32'ha719cb9a;
    ram_cell[   30255] = 32'h2da86895;
    ram_cell[   30256] = 32'h7ccf9e96;
    ram_cell[   30257] = 32'ha9b8a4b2;
    ram_cell[   30258] = 32'h9e3ff03a;
    ram_cell[   30259] = 32'h1d2bee60;
    ram_cell[   30260] = 32'h7cb7a089;
    ram_cell[   30261] = 32'hdedcfc24;
    ram_cell[   30262] = 32'h62b5cca0;
    ram_cell[   30263] = 32'h6b429b35;
    ram_cell[   30264] = 32'hb42df291;
    ram_cell[   30265] = 32'h4a28f7f3;
    ram_cell[   30266] = 32'h2280fba2;
    ram_cell[   30267] = 32'h094863ac;
    ram_cell[   30268] = 32'h8df6bfc7;
    ram_cell[   30269] = 32'h5686a1ce;
    ram_cell[   30270] = 32'h7657df6e;
    ram_cell[   30271] = 32'h397dccfc;
    ram_cell[   30272] = 32'h5eaf5fd1;
    ram_cell[   30273] = 32'h712bc7b5;
    ram_cell[   30274] = 32'h20e513a8;
    ram_cell[   30275] = 32'hd5d45480;
    ram_cell[   30276] = 32'hae1cf4d4;
    ram_cell[   30277] = 32'h8b1fe3e5;
    ram_cell[   30278] = 32'h96eca62e;
    ram_cell[   30279] = 32'he1f5e1d7;
    ram_cell[   30280] = 32'h1bf406d0;
    ram_cell[   30281] = 32'he19184fa;
    ram_cell[   30282] = 32'h4d307d3e;
    ram_cell[   30283] = 32'hd147a0b4;
    ram_cell[   30284] = 32'h776d2e95;
    ram_cell[   30285] = 32'hf98af6b9;
    ram_cell[   30286] = 32'hb00885c6;
    ram_cell[   30287] = 32'h9b59d2b6;
    ram_cell[   30288] = 32'h8c76f02d;
    ram_cell[   30289] = 32'h89bf8bd5;
    ram_cell[   30290] = 32'h46bc2975;
    ram_cell[   30291] = 32'h3bc2e21d;
    ram_cell[   30292] = 32'h0348a734;
    ram_cell[   30293] = 32'h92221a3f;
    ram_cell[   30294] = 32'h22fbc55f;
    ram_cell[   30295] = 32'h1d55e770;
    ram_cell[   30296] = 32'hf282e262;
    ram_cell[   30297] = 32'ha02b27b8;
    ram_cell[   30298] = 32'hb328bdba;
    ram_cell[   30299] = 32'h90c10a17;
    ram_cell[   30300] = 32'h366747a1;
    ram_cell[   30301] = 32'h8657f119;
    ram_cell[   30302] = 32'hf4c0b867;
    ram_cell[   30303] = 32'hf0401205;
    ram_cell[   30304] = 32'hf6c7ec72;
    ram_cell[   30305] = 32'h7079ae1c;
    ram_cell[   30306] = 32'h94078594;
    ram_cell[   30307] = 32'h18307ae2;
    ram_cell[   30308] = 32'h9029f954;
    ram_cell[   30309] = 32'h97fa00c1;
    ram_cell[   30310] = 32'h0c7fc2aa;
    ram_cell[   30311] = 32'h0a6b2ef7;
    ram_cell[   30312] = 32'ha59442d2;
    ram_cell[   30313] = 32'h8f81eba5;
    ram_cell[   30314] = 32'h8d4ebcfa;
    ram_cell[   30315] = 32'h98f2bed7;
    ram_cell[   30316] = 32'h0fde96f5;
    ram_cell[   30317] = 32'hb895af29;
    ram_cell[   30318] = 32'h4cc7b3b9;
    ram_cell[   30319] = 32'h05ae3e3b;
    ram_cell[   30320] = 32'h4cdc4869;
    ram_cell[   30321] = 32'h344be772;
    ram_cell[   30322] = 32'hd0b08255;
    ram_cell[   30323] = 32'h56596abc;
    ram_cell[   30324] = 32'he583ebaa;
    ram_cell[   30325] = 32'hd4fd72ae;
    ram_cell[   30326] = 32'h8cc97652;
    ram_cell[   30327] = 32'h72878671;
    ram_cell[   30328] = 32'h582d94e7;
    ram_cell[   30329] = 32'h3c8e5c3a;
    ram_cell[   30330] = 32'haba8b7b1;
    ram_cell[   30331] = 32'h455c6909;
    ram_cell[   30332] = 32'h2ee7076f;
    ram_cell[   30333] = 32'hf66c61a4;
    ram_cell[   30334] = 32'h82193ddf;
    ram_cell[   30335] = 32'hf62bf78a;
    ram_cell[   30336] = 32'h6e1cda92;
    ram_cell[   30337] = 32'hd64005d0;
    ram_cell[   30338] = 32'h14cebb75;
    ram_cell[   30339] = 32'he915dd5d;
    ram_cell[   30340] = 32'h6d3ae7dd;
    ram_cell[   30341] = 32'haeb194a8;
    ram_cell[   30342] = 32'hb3a1419f;
    ram_cell[   30343] = 32'h5366093e;
    ram_cell[   30344] = 32'hae7b483b;
    ram_cell[   30345] = 32'h90f6172f;
    ram_cell[   30346] = 32'h985c955f;
    ram_cell[   30347] = 32'h357a2a6e;
    ram_cell[   30348] = 32'hfe0e9bc5;
    ram_cell[   30349] = 32'h07a0511e;
    ram_cell[   30350] = 32'h0a7dd2c3;
    ram_cell[   30351] = 32'h672567f6;
    ram_cell[   30352] = 32'hfca9de50;
    ram_cell[   30353] = 32'h12e8ac10;
    ram_cell[   30354] = 32'h72b7b76e;
    ram_cell[   30355] = 32'h7cfdc3ef;
    ram_cell[   30356] = 32'hcabfd2c3;
    ram_cell[   30357] = 32'h63b775d5;
    ram_cell[   30358] = 32'h0c86605a;
    ram_cell[   30359] = 32'ha9a46a5e;
    ram_cell[   30360] = 32'h67df5460;
    ram_cell[   30361] = 32'h5df9aafb;
    ram_cell[   30362] = 32'h26fafcbf;
    ram_cell[   30363] = 32'h152f9d33;
    ram_cell[   30364] = 32'h70823142;
    ram_cell[   30365] = 32'h536429c1;
    ram_cell[   30366] = 32'hb74646ec;
    ram_cell[   30367] = 32'hff316124;
    ram_cell[   30368] = 32'hb6b19982;
    ram_cell[   30369] = 32'hb663c8f0;
    ram_cell[   30370] = 32'h2e16adad;
    ram_cell[   30371] = 32'h435eaa63;
    ram_cell[   30372] = 32'hf078763b;
    ram_cell[   30373] = 32'h09490011;
    ram_cell[   30374] = 32'h839de9e7;
    ram_cell[   30375] = 32'ha9a95456;
    ram_cell[   30376] = 32'hb623b0fb;
    ram_cell[   30377] = 32'h4f8c2e36;
    ram_cell[   30378] = 32'ha77f29e1;
    ram_cell[   30379] = 32'hecaf32ba;
    ram_cell[   30380] = 32'h3b6a18aa;
    ram_cell[   30381] = 32'haac60055;
    ram_cell[   30382] = 32'h5b9e3dd8;
    ram_cell[   30383] = 32'haf4ae3ec;
    ram_cell[   30384] = 32'h5c166161;
    ram_cell[   30385] = 32'h713d9ccb;
    ram_cell[   30386] = 32'h383f5215;
    ram_cell[   30387] = 32'h1094db1c;
    ram_cell[   30388] = 32'h5e3c6066;
    ram_cell[   30389] = 32'h28d50ab1;
    ram_cell[   30390] = 32'h2881d664;
    ram_cell[   30391] = 32'hc62208bd;
    ram_cell[   30392] = 32'h77d38ed8;
    ram_cell[   30393] = 32'h88f0dd51;
    ram_cell[   30394] = 32'ha7b321d9;
    ram_cell[   30395] = 32'h0dbb5a47;
    ram_cell[   30396] = 32'h0acb8c7b;
    ram_cell[   30397] = 32'hcddd39e4;
    ram_cell[   30398] = 32'h497f622a;
    ram_cell[   30399] = 32'h980d7787;
    ram_cell[   30400] = 32'h32181c1f;
    ram_cell[   30401] = 32'h424efe3e;
    ram_cell[   30402] = 32'hd8e8ee1d;
    ram_cell[   30403] = 32'hbac5c7bf;
    ram_cell[   30404] = 32'h01ba20cb;
    ram_cell[   30405] = 32'ha8cb784a;
    ram_cell[   30406] = 32'hffac109c;
    ram_cell[   30407] = 32'h8c13d3d6;
    ram_cell[   30408] = 32'hd34660c6;
    ram_cell[   30409] = 32'h6c5e994f;
    ram_cell[   30410] = 32'h01114dc7;
    ram_cell[   30411] = 32'hdd513114;
    ram_cell[   30412] = 32'hed9336a9;
    ram_cell[   30413] = 32'hf0d08a31;
    ram_cell[   30414] = 32'h24a9dd06;
    ram_cell[   30415] = 32'hf4dedc35;
    ram_cell[   30416] = 32'ha8e17375;
    ram_cell[   30417] = 32'h32c79221;
    ram_cell[   30418] = 32'h4b0f29d1;
    ram_cell[   30419] = 32'h372e7419;
    ram_cell[   30420] = 32'h67d20a99;
    ram_cell[   30421] = 32'h653f1ca9;
    ram_cell[   30422] = 32'h85f0366c;
    ram_cell[   30423] = 32'h3c00533f;
    ram_cell[   30424] = 32'h3f1d1129;
    ram_cell[   30425] = 32'h8ee36e8b;
    ram_cell[   30426] = 32'hc453a3cb;
    ram_cell[   30427] = 32'h57d49502;
    ram_cell[   30428] = 32'haab55c7c;
    ram_cell[   30429] = 32'h950fc6b0;
    ram_cell[   30430] = 32'h7fdcdc0c;
    ram_cell[   30431] = 32'hdde06a8c;
    ram_cell[   30432] = 32'h3d20f5ba;
    ram_cell[   30433] = 32'h99a1f0b9;
    ram_cell[   30434] = 32'hde3ac4f4;
    ram_cell[   30435] = 32'h47ca2f66;
    ram_cell[   30436] = 32'h2e595717;
    ram_cell[   30437] = 32'hbc2b0284;
    ram_cell[   30438] = 32'h6b292400;
    ram_cell[   30439] = 32'h847adc18;
    ram_cell[   30440] = 32'he3a48afd;
    ram_cell[   30441] = 32'hebcffe9e;
    ram_cell[   30442] = 32'h316cbf58;
    ram_cell[   30443] = 32'h6bb1d9af;
    ram_cell[   30444] = 32'hc6bfa9d3;
    ram_cell[   30445] = 32'heeaf9822;
    ram_cell[   30446] = 32'h89270a6d;
    ram_cell[   30447] = 32'h053623a0;
    ram_cell[   30448] = 32'h557491a7;
    ram_cell[   30449] = 32'h70dcb9b9;
    ram_cell[   30450] = 32'h55da6739;
    ram_cell[   30451] = 32'haccce14d;
    ram_cell[   30452] = 32'hd4a72c1d;
    ram_cell[   30453] = 32'h14912639;
    ram_cell[   30454] = 32'h6b77ffc2;
    ram_cell[   30455] = 32'h0792392b;
    ram_cell[   30456] = 32'hff78a491;
    ram_cell[   30457] = 32'he62d05b1;
    ram_cell[   30458] = 32'h2d04fbcf;
    ram_cell[   30459] = 32'h02ee75c4;
    ram_cell[   30460] = 32'h96cb69b9;
    ram_cell[   30461] = 32'h7aa383d9;
    ram_cell[   30462] = 32'hc81d506c;
    ram_cell[   30463] = 32'ha0a0a0ac;
    ram_cell[   30464] = 32'h017d95c5;
    ram_cell[   30465] = 32'he1eb639f;
    ram_cell[   30466] = 32'h54120dba;
    ram_cell[   30467] = 32'hc87f09c8;
    ram_cell[   30468] = 32'h7ec9da46;
    ram_cell[   30469] = 32'h404885dc;
    ram_cell[   30470] = 32'h87faa294;
    ram_cell[   30471] = 32'h59e37611;
    ram_cell[   30472] = 32'h37d85186;
    ram_cell[   30473] = 32'h1947c919;
    ram_cell[   30474] = 32'hc0d2cffa;
    ram_cell[   30475] = 32'h988cefa6;
    ram_cell[   30476] = 32'h905a5871;
    ram_cell[   30477] = 32'hfadd2565;
    ram_cell[   30478] = 32'h251a2eab;
    ram_cell[   30479] = 32'hd78db4d2;
    ram_cell[   30480] = 32'he4d12107;
    ram_cell[   30481] = 32'hfec10bc5;
    ram_cell[   30482] = 32'h5dd50b8e;
    ram_cell[   30483] = 32'haefd2249;
    ram_cell[   30484] = 32'h515352ce;
    ram_cell[   30485] = 32'hf182dc12;
    ram_cell[   30486] = 32'hc831d8f0;
    ram_cell[   30487] = 32'h3a7ac742;
    ram_cell[   30488] = 32'hc50d9d58;
    ram_cell[   30489] = 32'h022394e1;
    ram_cell[   30490] = 32'h83fce503;
    ram_cell[   30491] = 32'ha7fa1aa4;
    ram_cell[   30492] = 32'h6825652d;
    ram_cell[   30493] = 32'h0b7979b6;
    ram_cell[   30494] = 32'h4598a51f;
    ram_cell[   30495] = 32'h35178bcd;
    ram_cell[   30496] = 32'h00ae1e8e;
    ram_cell[   30497] = 32'h5eddaac3;
    ram_cell[   30498] = 32'h762a9ac8;
    ram_cell[   30499] = 32'h7931e318;
    ram_cell[   30500] = 32'h4c8c53fb;
    ram_cell[   30501] = 32'h3443077b;
    ram_cell[   30502] = 32'h4efbf47a;
    ram_cell[   30503] = 32'h5d134502;
    ram_cell[   30504] = 32'hf00be6d9;
    ram_cell[   30505] = 32'h1411c685;
    ram_cell[   30506] = 32'h52a703c9;
    ram_cell[   30507] = 32'h792b6f70;
    ram_cell[   30508] = 32'h074d0c02;
    ram_cell[   30509] = 32'h0933d792;
    ram_cell[   30510] = 32'h79cb803d;
    ram_cell[   30511] = 32'h380fb4d7;
    ram_cell[   30512] = 32'h184fb2c2;
    ram_cell[   30513] = 32'h3423e9df;
    ram_cell[   30514] = 32'h37869cd2;
    ram_cell[   30515] = 32'h3dd631f1;
    ram_cell[   30516] = 32'h7d00a629;
    ram_cell[   30517] = 32'hea92e133;
    ram_cell[   30518] = 32'h7f0cb3f0;
    ram_cell[   30519] = 32'h02437730;
    ram_cell[   30520] = 32'hbf8c646c;
    ram_cell[   30521] = 32'h83bff1f5;
    ram_cell[   30522] = 32'h124ef58b;
    ram_cell[   30523] = 32'h58edd1d9;
    ram_cell[   30524] = 32'h4f4be370;
    ram_cell[   30525] = 32'h5175f865;
    ram_cell[   30526] = 32'h40068f1d;
    ram_cell[   30527] = 32'h7054dd91;
    ram_cell[   30528] = 32'h2c8aa4b8;
    ram_cell[   30529] = 32'h664c109e;
    ram_cell[   30530] = 32'h22ea8d33;
    ram_cell[   30531] = 32'ha3521718;
    ram_cell[   30532] = 32'h8ed324c8;
    ram_cell[   30533] = 32'h46006f7f;
    ram_cell[   30534] = 32'ha36414eb;
    ram_cell[   30535] = 32'h25031153;
    ram_cell[   30536] = 32'h3a59ca06;
    ram_cell[   30537] = 32'h396e6ba7;
    ram_cell[   30538] = 32'h5e524578;
    ram_cell[   30539] = 32'h43860d37;
    ram_cell[   30540] = 32'h90ccdefa;
    ram_cell[   30541] = 32'h68029fb6;
    ram_cell[   30542] = 32'h28d80b54;
    ram_cell[   30543] = 32'h678667ea;
    ram_cell[   30544] = 32'hf9829146;
    ram_cell[   30545] = 32'h8b5cf870;
    ram_cell[   30546] = 32'hf49b4320;
    ram_cell[   30547] = 32'h604248e8;
    ram_cell[   30548] = 32'he9787067;
    ram_cell[   30549] = 32'h64879639;
    ram_cell[   30550] = 32'h291aefca;
    ram_cell[   30551] = 32'hd857022f;
    ram_cell[   30552] = 32'h025ce4a7;
    ram_cell[   30553] = 32'h164ef250;
    ram_cell[   30554] = 32'h66b8d485;
    ram_cell[   30555] = 32'hbe7fa559;
    ram_cell[   30556] = 32'h361473f6;
    ram_cell[   30557] = 32'h96d5e3eb;
    ram_cell[   30558] = 32'h7c137507;
    ram_cell[   30559] = 32'h286b8dc1;
    ram_cell[   30560] = 32'h59fa73b7;
    ram_cell[   30561] = 32'hd07a149b;
    ram_cell[   30562] = 32'h4ecd9025;
    ram_cell[   30563] = 32'h6d205ae1;
    ram_cell[   30564] = 32'hc69db967;
    ram_cell[   30565] = 32'h855b8830;
    ram_cell[   30566] = 32'h94c70f7d;
    ram_cell[   30567] = 32'h94ab7c77;
    ram_cell[   30568] = 32'h2672ee9c;
    ram_cell[   30569] = 32'hd7f8f721;
    ram_cell[   30570] = 32'h371bf7fe;
    ram_cell[   30571] = 32'h5b2cf565;
    ram_cell[   30572] = 32'heef1cc40;
    ram_cell[   30573] = 32'hd82b4c72;
    ram_cell[   30574] = 32'ha8ad1272;
    ram_cell[   30575] = 32'h4f883809;
    ram_cell[   30576] = 32'h7e7f235f;
    ram_cell[   30577] = 32'hfd8f46d0;
    ram_cell[   30578] = 32'he09a9365;
    ram_cell[   30579] = 32'hbdb36642;
    ram_cell[   30580] = 32'h5da74e2b;
    ram_cell[   30581] = 32'h8064562f;
    ram_cell[   30582] = 32'hdafb753b;
    ram_cell[   30583] = 32'he7ab780b;
    ram_cell[   30584] = 32'h73c966c5;
    ram_cell[   30585] = 32'hf5a75f6c;
    ram_cell[   30586] = 32'h00e0f394;
    ram_cell[   30587] = 32'hd2e4bd73;
    ram_cell[   30588] = 32'h53dab94f;
    ram_cell[   30589] = 32'he80e1f64;
    ram_cell[   30590] = 32'h8dfdca6a;
    ram_cell[   30591] = 32'h21971558;
    ram_cell[   30592] = 32'hacca7bce;
    ram_cell[   30593] = 32'h5cff6905;
    ram_cell[   30594] = 32'h889f3674;
    ram_cell[   30595] = 32'h0fa615f4;
    ram_cell[   30596] = 32'hc124b24c;
    ram_cell[   30597] = 32'hb4cf98c5;
    ram_cell[   30598] = 32'hffb92bf9;
    ram_cell[   30599] = 32'hf10e0d18;
    ram_cell[   30600] = 32'hc0597095;
    ram_cell[   30601] = 32'h6df07d38;
    ram_cell[   30602] = 32'h68b9288b;
    ram_cell[   30603] = 32'h1d9422b8;
    ram_cell[   30604] = 32'h87f01ad3;
    ram_cell[   30605] = 32'h40b8c9ff;
    ram_cell[   30606] = 32'hb2fd573f;
    ram_cell[   30607] = 32'h24045159;
    ram_cell[   30608] = 32'hb18a171c;
    ram_cell[   30609] = 32'h2b04beb3;
    ram_cell[   30610] = 32'he6282853;
    ram_cell[   30611] = 32'hd0dc62ce;
    ram_cell[   30612] = 32'h60892d77;
    ram_cell[   30613] = 32'hbd194ddd;
    ram_cell[   30614] = 32'h8dab77ea;
    ram_cell[   30615] = 32'h2f9a08ba;
    ram_cell[   30616] = 32'ha7dab661;
    ram_cell[   30617] = 32'h29e033fa;
    ram_cell[   30618] = 32'h5e96b5fd;
    ram_cell[   30619] = 32'hebe00414;
    ram_cell[   30620] = 32'h90a84302;
    ram_cell[   30621] = 32'hdd67e82d;
    ram_cell[   30622] = 32'h36078cb5;
    ram_cell[   30623] = 32'hbe64471c;
    ram_cell[   30624] = 32'h5b4d3d16;
    ram_cell[   30625] = 32'haad6c2e6;
    ram_cell[   30626] = 32'h8af1f649;
    ram_cell[   30627] = 32'hfe360cea;
    ram_cell[   30628] = 32'hd6580a3c;
    ram_cell[   30629] = 32'hf43df580;
    ram_cell[   30630] = 32'hd98f9a28;
    ram_cell[   30631] = 32'h88850a6e;
    ram_cell[   30632] = 32'haa803785;
    ram_cell[   30633] = 32'hd5b7457f;
    ram_cell[   30634] = 32'he4d3fca7;
    ram_cell[   30635] = 32'hd904ba62;
    ram_cell[   30636] = 32'h4d7cbfe9;
    ram_cell[   30637] = 32'h33c39bb6;
    ram_cell[   30638] = 32'h6ad1d6e6;
    ram_cell[   30639] = 32'h11d6738e;
    ram_cell[   30640] = 32'h6c4fd841;
    ram_cell[   30641] = 32'he19a2444;
    ram_cell[   30642] = 32'h91b6f1c1;
    ram_cell[   30643] = 32'hf9261494;
    ram_cell[   30644] = 32'h3c4f1409;
    ram_cell[   30645] = 32'hae742e4c;
    ram_cell[   30646] = 32'hcbcd8c1c;
    ram_cell[   30647] = 32'hf2cd6698;
    ram_cell[   30648] = 32'hbecef2cb;
    ram_cell[   30649] = 32'h1c59df9c;
    ram_cell[   30650] = 32'h5aa67c1b;
    ram_cell[   30651] = 32'h57214729;
    ram_cell[   30652] = 32'h412f2af2;
    ram_cell[   30653] = 32'h8a87e589;
    ram_cell[   30654] = 32'h36bfd227;
    ram_cell[   30655] = 32'h21f83970;
    ram_cell[   30656] = 32'h6676b01a;
    ram_cell[   30657] = 32'h4d433ec9;
    ram_cell[   30658] = 32'h9d47736a;
    ram_cell[   30659] = 32'hb3c685a6;
    ram_cell[   30660] = 32'h00ee1b3e;
    ram_cell[   30661] = 32'h18164313;
    ram_cell[   30662] = 32'h80c6720f;
    ram_cell[   30663] = 32'h9fd65f02;
    ram_cell[   30664] = 32'h4c70163f;
    ram_cell[   30665] = 32'hd5f98a1e;
    ram_cell[   30666] = 32'h3b7fd4a6;
    ram_cell[   30667] = 32'h90136de5;
    ram_cell[   30668] = 32'h2b858df7;
    ram_cell[   30669] = 32'h40de92bf;
    ram_cell[   30670] = 32'hbd4d57fa;
    ram_cell[   30671] = 32'h7efa2ac1;
    ram_cell[   30672] = 32'h9bacb9cf;
    ram_cell[   30673] = 32'he61396d0;
    ram_cell[   30674] = 32'h3642e7b6;
    ram_cell[   30675] = 32'h9243e194;
    ram_cell[   30676] = 32'h3ed75034;
    ram_cell[   30677] = 32'h708d47b1;
    ram_cell[   30678] = 32'hcc160411;
    ram_cell[   30679] = 32'hf9d9353c;
    ram_cell[   30680] = 32'ha14248d8;
    ram_cell[   30681] = 32'h147b8b75;
    ram_cell[   30682] = 32'h53b0f4b6;
    ram_cell[   30683] = 32'h2b9a98b4;
    ram_cell[   30684] = 32'h6c9ff907;
    ram_cell[   30685] = 32'h6fce2edb;
    ram_cell[   30686] = 32'h04dfe3d6;
    ram_cell[   30687] = 32'hdd5bc173;
    ram_cell[   30688] = 32'h63b3589c;
    ram_cell[   30689] = 32'h16483849;
    ram_cell[   30690] = 32'hb0d1bfff;
    ram_cell[   30691] = 32'he6bd1567;
    ram_cell[   30692] = 32'h2f4f6eac;
    ram_cell[   30693] = 32'h0844d0f2;
    ram_cell[   30694] = 32'hafb885d9;
    ram_cell[   30695] = 32'hc667bf55;
    ram_cell[   30696] = 32'h342d3ba9;
    ram_cell[   30697] = 32'hd47ad837;
    ram_cell[   30698] = 32'hcafd86a8;
    ram_cell[   30699] = 32'hcf20452b;
    ram_cell[   30700] = 32'he312a899;
    ram_cell[   30701] = 32'h32a670fe;
    ram_cell[   30702] = 32'h37ee9f6f;
    ram_cell[   30703] = 32'h3125af7e;
    ram_cell[   30704] = 32'hb7b0e942;
    ram_cell[   30705] = 32'ha5313aca;
    ram_cell[   30706] = 32'h23ad1152;
    ram_cell[   30707] = 32'hb8bdc18a;
    ram_cell[   30708] = 32'h843ff931;
    ram_cell[   30709] = 32'h6cb12ca2;
    ram_cell[   30710] = 32'h4acc8845;
    ram_cell[   30711] = 32'h93536538;
    ram_cell[   30712] = 32'h45943bbc;
    ram_cell[   30713] = 32'hf5ed8480;
    ram_cell[   30714] = 32'h1548fdd7;
    ram_cell[   30715] = 32'h242fc0d8;
    ram_cell[   30716] = 32'hec1fa883;
    ram_cell[   30717] = 32'h3374e95e;
    ram_cell[   30718] = 32'h419c14aa;
    ram_cell[   30719] = 32'h3f084464;
    ram_cell[   30720] = 32'h32887683;
    ram_cell[   30721] = 32'h4223ce11;
    ram_cell[   30722] = 32'h3cf6ecd3;
    ram_cell[   30723] = 32'h22e88279;
    ram_cell[   30724] = 32'h3e4d50d4;
    ram_cell[   30725] = 32'hb34202b0;
    ram_cell[   30726] = 32'h3e29ba70;
    ram_cell[   30727] = 32'h6878d891;
    ram_cell[   30728] = 32'he5252f39;
    ram_cell[   30729] = 32'hc7e66723;
    ram_cell[   30730] = 32'h156bfee7;
    ram_cell[   30731] = 32'h9267e5ea;
    ram_cell[   30732] = 32'h4be65ac0;
    ram_cell[   30733] = 32'h6bfd757d;
    ram_cell[   30734] = 32'hb4b676a7;
    ram_cell[   30735] = 32'hc9602f23;
    ram_cell[   30736] = 32'hb691db08;
    ram_cell[   30737] = 32'h92f4313e;
    ram_cell[   30738] = 32'h66fee719;
    ram_cell[   30739] = 32'hd6817224;
    ram_cell[   30740] = 32'h2b75f222;
    ram_cell[   30741] = 32'h0305c637;
    ram_cell[   30742] = 32'h8e1a9f3c;
    ram_cell[   30743] = 32'ha9fbc664;
    ram_cell[   30744] = 32'h8d17f38e;
    ram_cell[   30745] = 32'hb139024e;
    ram_cell[   30746] = 32'h82704de2;
    ram_cell[   30747] = 32'h8d30eafe;
    ram_cell[   30748] = 32'h1103588d;
    ram_cell[   30749] = 32'h93628db9;
    ram_cell[   30750] = 32'he77794b5;
    ram_cell[   30751] = 32'he2634874;
    ram_cell[   30752] = 32'hbaca490b;
    ram_cell[   30753] = 32'h4731967c;
    ram_cell[   30754] = 32'h1d8261ba;
    ram_cell[   30755] = 32'h40afe091;
    ram_cell[   30756] = 32'he59a3a5c;
    ram_cell[   30757] = 32'h42b572e6;
    ram_cell[   30758] = 32'h95c9e3cd;
    ram_cell[   30759] = 32'h692b911e;
    ram_cell[   30760] = 32'h5f221931;
    ram_cell[   30761] = 32'hfa54533a;
    ram_cell[   30762] = 32'h39bb12c5;
    ram_cell[   30763] = 32'hce1e3397;
    ram_cell[   30764] = 32'ha7c38f71;
    ram_cell[   30765] = 32'h3706bd34;
    ram_cell[   30766] = 32'h25c66e72;
    ram_cell[   30767] = 32'he302daee;
    ram_cell[   30768] = 32'h67c0d964;
    ram_cell[   30769] = 32'h3946f71a;
    ram_cell[   30770] = 32'h538e11d6;
    ram_cell[   30771] = 32'h0ab228bd;
    ram_cell[   30772] = 32'h88eaa728;
    ram_cell[   30773] = 32'h3256fc0d;
    ram_cell[   30774] = 32'ha49291f6;
    ram_cell[   30775] = 32'hb8ab1b54;
    ram_cell[   30776] = 32'h560fc8b2;
    ram_cell[   30777] = 32'ha9f1244b;
    ram_cell[   30778] = 32'h6659894b;
    ram_cell[   30779] = 32'h53742c53;
    ram_cell[   30780] = 32'hf957ac21;
    ram_cell[   30781] = 32'h46435c90;
    ram_cell[   30782] = 32'h1c12f35b;
    ram_cell[   30783] = 32'hf16e9656;
    ram_cell[   30784] = 32'hc362ee19;
    ram_cell[   30785] = 32'h615e04b1;
    ram_cell[   30786] = 32'hf48e2a11;
    ram_cell[   30787] = 32'hcaa5880d;
    ram_cell[   30788] = 32'h8a9a07ad;
    ram_cell[   30789] = 32'h6397867f;
    ram_cell[   30790] = 32'hf43726c6;
    ram_cell[   30791] = 32'h882c72cc;
    ram_cell[   30792] = 32'h2a1968f3;
    ram_cell[   30793] = 32'h005a6115;
    ram_cell[   30794] = 32'h0495f08d;
    ram_cell[   30795] = 32'h1827e7db;
    ram_cell[   30796] = 32'h61adc2ec;
    ram_cell[   30797] = 32'h3cc5221f;
    ram_cell[   30798] = 32'h9325588b;
    ram_cell[   30799] = 32'hea6e9086;
    ram_cell[   30800] = 32'h8e675b20;
    ram_cell[   30801] = 32'h605333a3;
    ram_cell[   30802] = 32'h865b35b6;
    ram_cell[   30803] = 32'h97c13ced;
    ram_cell[   30804] = 32'ha364b287;
    ram_cell[   30805] = 32'h88a477d8;
    ram_cell[   30806] = 32'h535483df;
    ram_cell[   30807] = 32'hc0df7cda;
    ram_cell[   30808] = 32'h80f0941d;
    ram_cell[   30809] = 32'h69d81d2a;
    ram_cell[   30810] = 32'hb610a692;
    ram_cell[   30811] = 32'hd0166e6f;
    ram_cell[   30812] = 32'h203855cf;
    ram_cell[   30813] = 32'h3abcfa75;
    ram_cell[   30814] = 32'h8bc3cb7a;
    ram_cell[   30815] = 32'h1c8fed5f;
    ram_cell[   30816] = 32'hf541efbb;
    ram_cell[   30817] = 32'h995ea461;
    ram_cell[   30818] = 32'h1140eb0a;
    ram_cell[   30819] = 32'h0df9baf0;
    ram_cell[   30820] = 32'h9213ae27;
    ram_cell[   30821] = 32'h8709af14;
    ram_cell[   30822] = 32'hf2cb8887;
    ram_cell[   30823] = 32'he76c047a;
    ram_cell[   30824] = 32'h9f4eb598;
    ram_cell[   30825] = 32'h2669ca34;
    ram_cell[   30826] = 32'h73fd784c;
    ram_cell[   30827] = 32'h4f9191d4;
    ram_cell[   30828] = 32'h07f7a41d;
    ram_cell[   30829] = 32'h2fb90d33;
    ram_cell[   30830] = 32'h62b3e95b;
    ram_cell[   30831] = 32'hb148cd26;
    ram_cell[   30832] = 32'he200d5a0;
    ram_cell[   30833] = 32'hf3ddce78;
    ram_cell[   30834] = 32'h5005ce2d;
    ram_cell[   30835] = 32'hc1b43428;
    ram_cell[   30836] = 32'hcc75b7b7;
    ram_cell[   30837] = 32'h8d1ddab6;
    ram_cell[   30838] = 32'h73e381e8;
    ram_cell[   30839] = 32'hb710a89b;
    ram_cell[   30840] = 32'h7acb8691;
    ram_cell[   30841] = 32'h243fc309;
    ram_cell[   30842] = 32'hd8e0e2ed;
    ram_cell[   30843] = 32'h1aecf34d;
    ram_cell[   30844] = 32'h09c0906c;
    ram_cell[   30845] = 32'h1b69b266;
    ram_cell[   30846] = 32'h54ba253a;
    ram_cell[   30847] = 32'h7275e0ae;
    ram_cell[   30848] = 32'haced635d;
    ram_cell[   30849] = 32'hcb5ca45b;
    ram_cell[   30850] = 32'h7af186a2;
    ram_cell[   30851] = 32'hd9cc83fe;
    ram_cell[   30852] = 32'he0bd202d;
    ram_cell[   30853] = 32'hdfdd5463;
    ram_cell[   30854] = 32'h8fc75a06;
    ram_cell[   30855] = 32'h20c98d58;
    ram_cell[   30856] = 32'hf190a511;
    ram_cell[   30857] = 32'h1ca7e70b;
    ram_cell[   30858] = 32'h1b5d32a8;
    ram_cell[   30859] = 32'hf1adab5f;
    ram_cell[   30860] = 32'h342b0b70;
    ram_cell[   30861] = 32'hedde1f7d;
    ram_cell[   30862] = 32'hc6e9f513;
    ram_cell[   30863] = 32'h39739523;
    ram_cell[   30864] = 32'h06d9afc1;
    ram_cell[   30865] = 32'h30335467;
    ram_cell[   30866] = 32'h984fbb06;
    ram_cell[   30867] = 32'h8262bc68;
    ram_cell[   30868] = 32'h3e577ddc;
    ram_cell[   30869] = 32'hb0f85f25;
    ram_cell[   30870] = 32'hd9aba3b9;
    ram_cell[   30871] = 32'h28f78b5a;
    ram_cell[   30872] = 32'hd88ae485;
    ram_cell[   30873] = 32'h4c7c3d54;
    ram_cell[   30874] = 32'he6cf7bcd;
    ram_cell[   30875] = 32'h0ccb9507;
    ram_cell[   30876] = 32'hcc652aab;
    ram_cell[   30877] = 32'hd8463731;
    ram_cell[   30878] = 32'he4341bd1;
    ram_cell[   30879] = 32'hf8153d67;
    ram_cell[   30880] = 32'h1958d056;
    ram_cell[   30881] = 32'h966e7876;
    ram_cell[   30882] = 32'h0bb360ff;
    ram_cell[   30883] = 32'he28bf3ee;
    ram_cell[   30884] = 32'h41218319;
    ram_cell[   30885] = 32'h3fcec9ab;
    ram_cell[   30886] = 32'hd129c1cf;
    ram_cell[   30887] = 32'hc09e5859;
    ram_cell[   30888] = 32'hbb30d0e5;
    ram_cell[   30889] = 32'h0959dab2;
    ram_cell[   30890] = 32'h784a4b04;
    ram_cell[   30891] = 32'h7de58b61;
    ram_cell[   30892] = 32'ha182f01b;
    ram_cell[   30893] = 32'h19957398;
    ram_cell[   30894] = 32'hec529f5e;
    ram_cell[   30895] = 32'h02d74502;
    ram_cell[   30896] = 32'h66eb86c2;
    ram_cell[   30897] = 32'h4699d5bd;
    ram_cell[   30898] = 32'h37a2552d;
    ram_cell[   30899] = 32'h633308a2;
    ram_cell[   30900] = 32'h3a2923d2;
    ram_cell[   30901] = 32'hbffe8dc3;
    ram_cell[   30902] = 32'hc81664f0;
    ram_cell[   30903] = 32'h7a8e8312;
    ram_cell[   30904] = 32'hc1a7e4d0;
    ram_cell[   30905] = 32'h2ba343eb;
    ram_cell[   30906] = 32'he820d745;
    ram_cell[   30907] = 32'hd19d37cd;
    ram_cell[   30908] = 32'h2a083900;
    ram_cell[   30909] = 32'h6addb3b4;
    ram_cell[   30910] = 32'h1a6616ab;
    ram_cell[   30911] = 32'h898f3b5a;
    ram_cell[   30912] = 32'h05ffcf31;
    ram_cell[   30913] = 32'hc6f3bce9;
    ram_cell[   30914] = 32'h770028cf;
    ram_cell[   30915] = 32'h1968ee34;
    ram_cell[   30916] = 32'h166196f1;
    ram_cell[   30917] = 32'h86308c21;
    ram_cell[   30918] = 32'h671e9ce9;
    ram_cell[   30919] = 32'hdaec98a9;
    ram_cell[   30920] = 32'h53d4d6e8;
    ram_cell[   30921] = 32'h41c11cd5;
    ram_cell[   30922] = 32'ha3404a16;
    ram_cell[   30923] = 32'haa9c0d54;
    ram_cell[   30924] = 32'hd0a859a2;
    ram_cell[   30925] = 32'h937b5687;
    ram_cell[   30926] = 32'h6d1516e3;
    ram_cell[   30927] = 32'h70762c42;
    ram_cell[   30928] = 32'h446b1e54;
    ram_cell[   30929] = 32'ha2a36576;
    ram_cell[   30930] = 32'h8fc07e58;
    ram_cell[   30931] = 32'hc6d5275b;
    ram_cell[   30932] = 32'h66e346dc;
    ram_cell[   30933] = 32'h2487e1d6;
    ram_cell[   30934] = 32'h86e21853;
    ram_cell[   30935] = 32'h8c02a83e;
    ram_cell[   30936] = 32'hf5f823cb;
    ram_cell[   30937] = 32'hed334376;
    ram_cell[   30938] = 32'h82ab1e18;
    ram_cell[   30939] = 32'hed190ea7;
    ram_cell[   30940] = 32'hee13be4b;
    ram_cell[   30941] = 32'hf17195df;
    ram_cell[   30942] = 32'h27a6f4dc;
    ram_cell[   30943] = 32'h1a1da0da;
    ram_cell[   30944] = 32'h7a749f4a;
    ram_cell[   30945] = 32'he577ff73;
    ram_cell[   30946] = 32'h99d707c6;
    ram_cell[   30947] = 32'h9ce5ea70;
    ram_cell[   30948] = 32'h71bfefaf;
    ram_cell[   30949] = 32'h5a3fcd04;
    ram_cell[   30950] = 32'h65e65e4b;
    ram_cell[   30951] = 32'h4807fa78;
    ram_cell[   30952] = 32'h37b268e5;
    ram_cell[   30953] = 32'h0f0459f5;
    ram_cell[   30954] = 32'hd15252d7;
    ram_cell[   30955] = 32'h9476b24b;
    ram_cell[   30956] = 32'h414f47b0;
    ram_cell[   30957] = 32'hfeee5329;
    ram_cell[   30958] = 32'h772a227c;
    ram_cell[   30959] = 32'hcf7c85d4;
    ram_cell[   30960] = 32'ha3422b65;
    ram_cell[   30961] = 32'h955f1fb2;
    ram_cell[   30962] = 32'h107c3635;
    ram_cell[   30963] = 32'hdd633638;
    ram_cell[   30964] = 32'h28fe69e1;
    ram_cell[   30965] = 32'h659b662f;
    ram_cell[   30966] = 32'haa65970b;
    ram_cell[   30967] = 32'h91c9d76b;
    ram_cell[   30968] = 32'hc9f9534e;
    ram_cell[   30969] = 32'h56936843;
    ram_cell[   30970] = 32'hb0b9feea;
    ram_cell[   30971] = 32'he6e2f9e4;
    ram_cell[   30972] = 32'h6037664f;
    ram_cell[   30973] = 32'h67cc55e7;
    ram_cell[   30974] = 32'h93019ceb;
    ram_cell[   30975] = 32'hd7699304;
    ram_cell[   30976] = 32'h6a15beb2;
    ram_cell[   30977] = 32'hce706d6b;
    ram_cell[   30978] = 32'h42818962;
    ram_cell[   30979] = 32'h6d19edc2;
    ram_cell[   30980] = 32'h653478b3;
    ram_cell[   30981] = 32'h176975cc;
    ram_cell[   30982] = 32'hf42c116c;
    ram_cell[   30983] = 32'he7b84245;
    ram_cell[   30984] = 32'hcd66b8fe;
    ram_cell[   30985] = 32'h4a5f52f3;
    ram_cell[   30986] = 32'h73aba28f;
    ram_cell[   30987] = 32'hf0e4396a;
    ram_cell[   30988] = 32'hfeba1286;
    ram_cell[   30989] = 32'h7be566dc;
    ram_cell[   30990] = 32'hc0ab087d;
    ram_cell[   30991] = 32'h0023b0a7;
    ram_cell[   30992] = 32'h36582f7f;
    ram_cell[   30993] = 32'h8c94ffda;
    ram_cell[   30994] = 32'h3d23f75f;
    ram_cell[   30995] = 32'h42bedc66;
    ram_cell[   30996] = 32'h3dd3d0a8;
    ram_cell[   30997] = 32'h4676abdf;
    ram_cell[   30998] = 32'h40470fc4;
    ram_cell[   30999] = 32'h78d8d8d0;
    ram_cell[   31000] = 32'h2464a2c7;
    ram_cell[   31001] = 32'h66d9b6d7;
    ram_cell[   31002] = 32'h82b064de;
    ram_cell[   31003] = 32'h1f70c43a;
    ram_cell[   31004] = 32'h5c257116;
    ram_cell[   31005] = 32'h8f71af61;
    ram_cell[   31006] = 32'hb732068d;
    ram_cell[   31007] = 32'h29dd613c;
    ram_cell[   31008] = 32'h3b5d249a;
    ram_cell[   31009] = 32'h550e30f6;
    ram_cell[   31010] = 32'habccc50b;
    ram_cell[   31011] = 32'h632784a9;
    ram_cell[   31012] = 32'h1f3e1dce;
    ram_cell[   31013] = 32'h338bbe57;
    ram_cell[   31014] = 32'hc6ab9762;
    ram_cell[   31015] = 32'h68b02934;
    ram_cell[   31016] = 32'h69a8cf17;
    ram_cell[   31017] = 32'h9ddaedb0;
    ram_cell[   31018] = 32'h36441b37;
    ram_cell[   31019] = 32'hb5e26985;
    ram_cell[   31020] = 32'hd72b0501;
    ram_cell[   31021] = 32'h3c643d9a;
    ram_cell[   31022] = 32'h960f7d20;
    ram_cell[   31023] = 32'h9432c454;
    ram_cell[   31024] = 32'hf6fd2185;
    ram_cell[   31025] = 32'h48a7a932;
    ram_cell[   31026] = 32'h70eba272;
    ram_cell[   31027] = 32'hbb1ec144;
    ram_cell[   31028] = 32'hb8b8509c;
    ram_cell[   31029] = 32'h38cbad12;
    ram_cell[   31030] = 32'hd9d69a09;
    ram_cell[   31031] = 32'h42a0d90e;
    ram_cell[   31032] = 32'h53c6e550;
    ram_cell[   31033] = 32'h1f86745e;
    ram_cell[   31034] = 32'h8085e1eb;
    ram_cell[   31035] = 32'h4be430c8;
    ram_cell[   31036] = 32'h8bce6584;
    ram_cell[   31037] = 32'hb033af8b;
    ram_cell[   31038] = 32'h084512a4;
    ram_cell[   31039] = 32'ha284870d;
    ram_cell[   31040] = 32'hf9d70780;
    ram_cell[   31041] = 32'he3106d5f;
    ram_cell[   31042] = 32'h1b21cd8a;
    ram_cell[   31043] = 32'h7ee87373;
    ram_cell[   31044] = 32'h7de00d09;
    ram_cell[   31045] = 32'hb0a7db68;
    ram_cell[   31046] = 32'h757cb36d;
    ram_cell[   31047] = 32'h9fe296d7;
    ram_cell[   31048] = 32'h2f75b243;
    ram_cell[   31049] = 32'h2a4ab0c6;
    ram_cell[   31050] = 32'hba6bf4c3;
    ram_cell[   31051] = 32'h1697f5d7;
    ram_cell[   31052] = 32'hdabd4376;
    ram_cell[   31053] = 32'hf4a8c06e;
    ram_cell[   31054] = 32'h3f283f12;
    ram_cell[   31055] = 32'hfa36165d;
    ram_cell[   31056] = 32'h5eb0bbe3;
    ram_cell[   31057] = 32'he7379f1a;
    ram_cell[   31058] = 32'h0aab5c93;
    ram_cell[   31059] = 32'hf178c942;
    ram_cell[   31060] = 32'hd8e6fd85;
    ram_cell[   31061] = 32'hb2324de9;
    ram_cell[   31062] = 32'h25ed1afe;
    ram_cell[   31063] = 32'h86ca951f;
    ram_cell[   31064] = 32'hdaddeae5;
    ram_cell[   31065] = 32'hac04adc2;
    ram_cell[   31066] = 32'h17d97159;
    ram_cell[   31067] = 32'h800835a4;
    ram_cell[   31068] = 32'hc5a2cc05;
    ram_cell[   31069] = 32'h59e126e4;
    ram_cell[   31070] = 32'h3f1221f3;
    ram_cell[   31071] = 32'hf3528451;
    ram_cell[   31072] = 32'h50e7a274;
    ram_cell[   31073] = 32'h7bfbdccf;
    ram_cell[   31074] = 32'h00701736;
    ram_cell[   31075] = 32'h33c04dfc;
    ram_cell[   31076] = 32'h5c827f85;
    ram_cell[   31077] = 32'hb60dbc7c;
    ram_cell[   31078] = 32'h6ba842d3;
    ram_cell[   31079] = 32'h9e7af4c6;
    ram_cell[   31080] = 32'h258c75df;
    ram_cell[   31081] = 32'h1bbcadea;
    ram_cell[   31082] = 32'h6bbf7516;
    ram_cell[   31083] = 32'h1810c8a0;
    ram_cell[   31084] = 32'h2ff34954;
    ram_cell[   31085] = 32'h0b20334d;
    ram_cell[   31086] = 32'h02480d8f;
    ram_cell[   31087] = 32'he27c3316;
    ram_cell[   31088] = 32'h8838e996;
    ram_cell[   31089] = 32'he169295c;
    ram_cell[   31090] = 32'h58250c1c;
    ram_cell[   31091] = 32'hec1ffde0;
    ram_cell[   31092] = 32'hf4d8aec6;
    ram_cell[   31093] = 32'hb131ae61;
    ram_cell[   31094] = 32'h90d4d40a;
    ram_cell[   31095] = 32'h8efc17d6;
    ram_cell[   31096] = 32'h4422afd5;
    ram_cell[   31097] = 32'h0de337c6;
    ram_cell[   31098] = 32'hb774e752;
    ram_cell[   31099] = 32'hba8efcc2;
    ram_cell[   31100] = 32'h07ddba67;
    ram_cell[   31101] = 32'h795ca0bc;
    ram_cell[   31102] = 32'h472c501a;
    ram_cell[   31103] = 32'h4421db93;
    ram_cell[   31104] = 32'h4678b360;
    ram_cell[   31105] = 32'hf0e392cd;
    ram_cell[   31106] = 32'hc73b8f42;
    ram_cell[   31107] = 32'h07d9d9e1;
    ram_cell[   31108] = 32'ha48e7d07;
    ram_cell[   31109] = 32'h4d47c617;
    ram_cell[   31110] = 32'h0d1ed325;
    ram_cell[   31111] = 32'hbbac9f62;
    ram_cell[   31112] = 32'ha20d7a1b;
    ram_cell[   31113] = 32'h87948a27;
    ram_cell[   31114] = 32'hce723307;
    ram_cell[   31115] = 32'hb8bf327f;
    ram_cell[   31116] = 32'heeceaa0f;
    ram_cell[   31117] = 32'hc6476bc0;
    ram_cell[   31118] = 32'h9ece6a00;
    ram_cell[   31119] = 32'h18459723;
    ram_cell[   31120] = 32'h242036d7;
    ram_cell[   31121] = 32'h035c5c34;
    ram_cell[   31122] = 32'h3fff01e6;
    ram_cell[   31123] = 32'h7e5e96f4;
    ram_cell[   31124] = 32'h2f4b1ec4;
    ram_cell[   31125] = 32'h3bd08361;
    ram_cell[   31126] = 32'hf9764be3;
    ram_cell[   31127] = 32'h3ae091f2;
    ram_cell[   31128] = 32'hb30134e3;
    ram_cell[   31129] = 32'ha1d6f2de;
    ram_cell[   31130] = 32'hc919006b;
    ram_cell[   31131] = 32'h40697eae;
    ram_cell[   31132] = 32'h7037d496;
    ram_cell[   31133] = 32'he77da7c3;
    ram_cell[   31134] = 32'h7990a6fc;
    ram_cell[   31135] = 32'h9147a321;
    ram_cell[   31136] = 32'h094c0d0f;
    ram_cell[   31137] = 32'ha98b164c;
    ram_cell[   31138] = 32'h7274e951;
    ram_cell[   31139] = 32'h3d873a2f;
    ram_cell[   31140] = 32'hafcd6e96;
    ram_cell[   31141] = 32'h06f97495;
    ram_cell[   31142] = 32'hbcbd2d11;
    ram_cell[   31143] = 32'hbc160886;
    ram_cell[   31144] = 32'h9cf1797f;
    ram_cell[   31145] = 32'h6c73b44e;
    ram_cell[   31146] = 32'hbad33898;
    ram_cell[   31147] = 32'ha1c4bfae;
    ram_cell[   31148] = 32'hde085e68;
    ram_cell[   31149] = 32'hd8764875;
    ram_cell[   31150] = 32'h5b06e3ef;
    ram_cell[   31151] = 32'h8dd976e3;
    ram_cell[   31152] = 32'h61a247a6;
    ram_cell[   31153] = 32'ha5ec3ffd;
    ram_cell[   31154] = 32'hd078a380;
    ram_cell[   31155] = 32'hc338e010;
    ram_cell[   31156] = 32'h9f6ef3a3;
    ram_cell[   31157] = 32'h0a3ce0d1;
    ram_cell[   31158] = 32'h56deccbf;
    ram_cell[   31159] = 32'h55b7fd15;
    ram_cell[   31160] = 32'hac34ec86;
    ram_cell[   31161] = 32'h8084293b;
    ram_cell[   31162] = 32'h7e5b0950;
    ram_cell[   31163] = 32'h8774e37f;
    ram_cell[   31164] = 32'h1c4c3bd3;
    ram_cell[   31165] = 32'he7962b05;
    ram_cell[   31166] = 32'h64a768e5;
    ram_cell[   31167] = 32'h20477e96;
    ram_cell[   31168] = 32'h9d8e6f00;
    ram_cell[   31169] = 32'h7a6ee338;
    ram_cell[   31170] = 32'h497f5282;
    ram_cell[   31171] = 32'h667642e2;
    ram_cell[   31172] = 32'h1182219a;
    ram_cell[   31173] = 32'hfdb43daf;
    ram_cell[   31174] = 32'hb86840e4;
    ram_cell[   31175] = 32'h034080a0;
    ram_cell[   31176] = 32'h98412708;
    ram_cell[   31177] = 32'h0b50b274;
    ram_cell[   31178] = 32'h196065f5;
    ram_cell[   31179] = 32'h85eaa3e8;
    ram_cell[   31180] = 32'h428e927c;
    ram_cell[   31181] = 32'hcb99e3c4;
    ram_cell[   31182] = 32'h50c7dd39;
    ram_cell[   31183] = 32'h39cd4f40;
    ram_cell[   31184] = 32'h84fefb88;
    ram_cell[   31185] = 32'h511f7659;
    ram_cell[   31186] = 32'h06c7a1a3;
    ram_cell[   31187] = 32'h1261f6ac;
    ram_cell[   31188] = 32'hfeb4f502;
    ram_cell[   31189] = 32'h9927689a;
    ram_cell[   31190] = 32'h54aa5024;
    ram_cell[   31191] = 32'h90d5b27d;
    ram_cell[   31192] = 32'h9d2d323d;
    ram_cell[   31193] = 32'h0349d10f;
    ram_cell[   31194] = 32'h3c3e348e;
    ram_cell[   31195] = 32'hcc5830b4;
    ram_cell[   31196] = 32'h9a2b495d;
    ram_cell[   31197] = 32'hb532e3bb;
    ram_cell[   31198] = 32'h23ba1040;
    ram_cell[   31199] = 32'h0ba7a8cd;
    ram_cell[   31200] = 32'h90016428;
    ram_cell[   31201] = 32'h11fcbf7d;
    ram_cell[   31202] = 32'hdfa273ef;
    ram_cell[   31203] = 32'hc2eb75a2;
    ram_cell[   31204] = 32'hfe412877;
    ram_cell[   31205] = 32'h3989d278;
    ram_cell[   31206] = 32'h4ac37463;
    ram_cell[   31207] = 32'h75002967;
    ram_cell[   31208] = 32'h4c1d0bdb;
    ram_cell[   31209] = 32'h8058d734;
    ram_cell[   31210] = 32'h13277540;
    ram_cell[   31211] = 32'h1483e20d;
    ram_cell[   31212] = 32'ha6c9e7d3;
    ram_cell[   31213] = 32'h682feeab;
    ram_cell[   31214] = 32'ha944eb04;
    ram_cell[   31215] = 32'h7354e5f4;
    ram_cell[   31216] = 32'h8831342d;
    ram_cell[   31217] = 32'h787a7bee;
    ram_cell[   31218] = 32'hf62b1e1d;
    ram_cell[   31219] = 32'h4bc8a76c;
    ram_cell[   31220] = 32'h51b533e9;
    ram_cell[   31221] = 32'he480d85d;
    ram_cell[   31222] = 32'h7729aa62;
    ram_cell[   31223] = 32'hc54fcc5b;
    ram_cell[   31224] = 32'ha7d15404;
    ram_cell[   31225] = 32'h0ee171e5;
    ram_cell[   31226] = 32'ha34c1142;
    ram_cell[   31227] = 32'h6005c85d;
    ram_cell[   31228] = 32'h0ca12edb;
    ram_cell[   31229] = 32'h7cff1712;
    ram_cell[   31230] = 32'hbfbd82bd;
    ram_cell[   31231] = 32'hbc907ea9;
    ram_cell[   31232] = 32'h08714cd9;
    ram_cell[   31233] = 32'h9618f8c5;
    ram_cell[   31234] = 32'h54065832;
    ram_cell[   31235] = 32'h7c3cb282;
    ram_cell[   31236] = 32'h3aed7d3a;
    ram_cell[   31237] = 32'h107542ba;
    ram_cell[   31238] = 32'h9efbf9a0;
    ram_cell[   31239] = 32'h933b2212;
    ram_cell[   31240] = 32'hb4a7bcf7;
    ram_cell[   31241] = 32'h62cb92b3;
    ram_cell[   31242] = 32'hc503685d;
    ram_cell[   31243] = 32'h060cfc76;
    ram_cell[   31244] = 32'hb8a70550;
    ram_cell[   31245] = 32'ha31b49ec;
    ram_cell[   31246] = 32'h5225acd0;
    ram_cell[   31247] = 32'h80ce11b0;
    ram_cell[   31248] = 32'haaf4ddfc;
    ram_cell[   31249] = 32'hd0e44882;
    ram_cell[   31250] = 32'h46ac063b;
    ram_cell[   31251] = 32'h021dc52c;
    ram_cell[   31252] = 32'h2a53671d;
    ram_cell[   31253] = 32'h24674893;
    ram_cell[   31254] = 32'hb45a8e13;
    ram_cell[   31255] = 32'h4d8ab48a;
    ram_cell[   31256] = 32'h59250acd;
    ram_cell[   31257] = 32'h705d77b3;
    ram_cell[   31258] = 32'h334976e5;
    ram_cell[   31259] = 32'haae477ca;
    ram_cell[   31260] = 32'h32e7f1e7;
    ram_cell[   31261] = 32'h7a6d04da;
    ram_cell[   31262] = 32'hf5df3ca4;
    ram_cell[   31263] = 32'h903cc933;
    ram_cell[   31264] = 32'h96035a09;
    ram_cell[   31265] = 32'h370d2fef;
    ram_cell[   31266] = 32'hb8501829;
    ram_cell[   31267] = 32'hd979c4d7;
    ram_cell[   31268] = 32'h0437efa2;
    ram_cell[   31269] = 32'hf7efb231;
    ram_cell[   31270] = 32'h4a29349c;
    ram_cell[   31271] = 32'hb517d705;
    ram_cell[   31272] = 32'ha39aa6a7;
    ram_cell[   31273] = 32'h071de54c;
    ram_cell[   31274] = 32'h49063693;
    ram_cell[   31275] = 32'hd6dbe099;
    ram_cell[   31276] = 32'hdba13a32;
    ram_cell[   31277] = 32'h110b36ef;
    ram_cell[   31278] = 32'h4c2da3f9;
    ram_cell[   31279] = 32'h715cd9c3;
    ram_cell[   31280] = 32'h229819ec;
    ram_cell[   31281] = 32'hf5a78071;
    ram_cell[   31282] = 32'h74e7e20a;
    ram_cell[   31283] = 32'h0e975100;
    ram_cell[   31284] = 32'he4dc59c8;
    ram_cell[   31285] = 32'hea03b38a;
    ram_cell[   31286] = 32'h5bfbd0ca;
    ram_cell[   31287] = 32'hdf4974ef;
    ram_cell[   31288] = 32'h5c1a2a3a;
    ram_cell[   31289] = 32'h33617135;
    ram_cell[   31290] = 32'h7aecfeb6;
    ram_cell[   31291] = 32'h72b2f362;
    ram_cell[   31292] = 32'h6fc9e3b3;
    ram_cell[   31293] = 32'hfb15beac;
    ram_cell[   31294] = 32'h86c038f3;
    ram_cell[   31295] = 32'h51661045;
    ram_cell[   31296] = 32'hd98d4884;
    ram_cell[   31297] = 32'h2cb475d7;
    ram_cell[   31298] = 32'h59e063cb;
    ram_cell[   31299] = 32'h58877fbb;
    ram_cell[   31300] = 32'hda111531;
    ram_cell[   31301] = 32'h2db4f663;
    ram_cell[   31302] = 32'h5bbe501c;
    ram_cell[   31303] = 32'he114675e;
    ram_cell[   31304] = 32'hbf588977;
    ram_cell[   31305] = 32'h4cefbabe;
    ram_cell[   31306] = 32'h18b6993d;
    ram_cell[   31307] = 32'h3bd821ac;
    ram_cell[   31308] = 32'h849925c0;
    ram_cell[   31309] = 32'h170225ec;
    ram_cell[   31310] = 32'h3332e2e3;
    ram_cell[   31311] = 32'h7ce1abd3;
    ram_cell[   31312] = 32'hf53066ec;
    ram_cell[   31313] = 32'h93e440ba;
    ram_cell[   31314] = 32'hb3e4a637;
    ram_cell[   31315] = 32'h8842ad1a;
    ram_cell[   31316] = 32'h601feced;
    ram_cell[   31317] = 32'haf9ec01b;
    ram_cell[   31318] = 32'hdc1c7eca;
    ram_cell[   31319] = 32'h15a91337;
    ram_cell[   31320] = 32'hd5fcd04e;
    ram_cell[   31321] = 32'hd08c3e5e;
    ram_cell[   31322] = 32'hb6dda93d;
    ram_cell[   31323] = 32'h663a6172;
    ram_cell[   31324] = 32'hf7a347b3;
    ram_cell[   31325] = 32'hf31fac29;
    ram_cell[   31326] = 32'h9f02bf5f;
    ram_cell[   31327] = 32'h72a32cdc;
    ram_cell[   31328] = 32'hd0a30de0;
    ram_cell[   31329] = 32'h648ae730;
    ram_cell[   31330] = 32'h6174b049;
    ram_cell[   31331] = 32'h55d13d2a;
    ram_cell[   31332] = 32'h917c4a53;
    ram_cell[   31333] = 32'h30f9c018;
    ram_cell[   31334] = 32'h107d8c82;
    ram_cell[   31335] = 32'h6bb7e0e0;
    ram_cell[   31336] = 32'h33f7b7ca;
    ram_cell[   31337] = 32'he6b1780e;
    ram_cell[   31338] = 32'h0fb99b7b;
    ram_cell[   31339] = 32'hbf59c88a;
    ram_cell[   31340] = 32'he24b3e1f;
    ram_cell[   31341] = 32'h257a05a2;
    ram_cell[   31342] = 32'h95479ce4;
    ram_cell[   31343] = 32'h787df387;
    ram_cell[   31344] = 32'h792238c1;
    ram_cell[   31345] = 32'h5fca58dd;
    ram_cell[   31346] = 32'h08976a6d;
    ram_cell[   31347] = 32'h956285b0;
    ram_cell[   31348] = 32'h61d33008;
    ram_cell[   31349] = 32'h3cc4f928;
    ram_cell[   31350] = 32'hd14c14c8;
    ram_cell[   31351] = 32'h3506ba7c;
    ram_cell[   31352] = 32'h1ef47d5e;
    ram_cell[   31353] = 32'h04e4032c;
    ram_cell[   31354] = 32'hd79982e6;
    ram_cell[   31355] = 32'hf37d4a54;
    ram_cell[   31356] = 32'ha9cf9988;
    ram_cell[   31357] = 32'hef18c6a8;
    ram_cell[   31358] = 32'h56742c78;
    ram_cell[   31359] = 32'h6a01b32e;
    ram_cell[   31360] = 32'h70ed7b13;
    ram_cell[   31361] = 32'hde9d629c;
    ram_cell[   31362] = 32'h77a94c80;
    ram_cell[   31363] = 32'h023a2f6c;
    ram_cell[   31364] = 32'h02985091;
    ram_cell[   31365] = 32'h0e0e8f1d;
    ram_cell[   31366] = 32'hc03836f3;
    ram_cell[   31367] = 32'h92b7ba09;
    ram_cell[   31368] = 32'h8b0de160;
    ram_cell[   31369] = 32'haa857565;
    ram_cell[   31370] = 32'h011bc52f;
    ram_cell[   31371] = 32'he21d17ed;
    ram_cell[   31372] = 32'ha247ad8b;
    ram_cell[   31373] = 32'h97650b70;
    ram_cell[   31374] = 32'hfb2ea40a;
    ram_cell[   31375] = 32'hbd72e046;
    ram_cell[   31376] = 32'h7975994d;
    ram_cell[   31377] = 32'h85a256a0;
    ram_cell[   31378] = 32'ha5e60ec1;
    ram_cell[   31379] = 32'h5e1ee535;
    ram_cell[   31380] = 32'h72ebce38;
    ram_cell[   31381] = 32'ha4507aae;
    ram_cell[   31382] = 32'h272991b2;
    ram_cell[   31383] = 32'h7483ee28;
    ram_cell[   31384] = 32'hdd974232;
    ram_cell[   31385] = 32'h6a51f2c8;
    ram_cell[   31386] = 32'he0da2e4e;
    ram_cell[   31387] = 32'h1cca48d5;
    ram_cell[   31388] = 32'h1ed33fed;
    ram_cell[   31389] = 32'ha6bd6a28;
    ram_cell[   31390] = 32'hb7b9a0f0;
    ram_cell[   31391] = 32'h09cb54f0;
    ram_cell[   31392] = 32'h6e597b98;
    ram_cell[   31393] = 32'ha37e1dff;
    ram_cell[   31394] = 32'hf9018913;
    ram_cell[   31395] = 32'h4862a1d3;
    ram_cell[   31396] = 32'hb4fd568f;
    ram_cell[   31397] = 32'hcced3e13;
    ram_cell[   31398] = 32'hd3c68ffa;
    ram_cell[   31399] = 32'h358902c2;
    ram_cell[   31400] = 32'h23db34e1;
    ram_cell[   31401] = 32'h8cb7e9d7;
    ram_cell[   31402] = 32'h75f804e5;
    ram_cell[   31403] = 32'hb8135e78;
    ram_cell[   31404] = 32'h9bf38547;
    ram_cell[   31405] = 32'haa49b88f;
    ram_cell[   31406] = 32'h23d45ac3;
    ram_cell[   31407] = 32'h6998ba5c;
    ram_cell[   31408] = 32'hbd45707c;
    ram_cell[   31409] = 32'h9a39ede1;
    ram_cell[   31410] = 32'h57bdf71d;
    ram_cell[   31411] = 32'hec4586b0;
    ram_cell[   31412] = 32'h3fb759dd;
    ram_cell[   31413] = 32'hc50229cd;
    ram_cell[   31414] = 32'he24483fc;
    ram_cell[   31415] = 32'h4905ff7a;
    ram_cell[   31416] = 32'h816f3442;
    ram_cell[   31417] = 32'hc6c9a00a;
    ram_cell[   31418] = 32'hf50a903a;
    ram_cell[   31419] = 32'h43f51845;
    ram_cell[   31420] = 32'h465d5a5a;
    ram_cell[   31421] = 32'h6887b4fc;
    ram_cell[   31422] = 32'he2f335d9;
    ram_cell[   31423] = 32'h7466f8cc;
    ram_cell[   31424] = 32'hb63ba1ca;
    ram_cell[   31425] = 32'h24538a81;
    ram_cell[   31426] = 32'h5c022229;
    ram_cell[   31427] = 32'hb1d92fe6;
    ram_cell[   31428] = 32'hce6ec129;
    ram_cell[   31429] = 32'hd4dac7fd;
    ram_cell[   31430] = 32'h3e2b5781;
    ram_cell[   31431] = 32'h803cd24a;
    ram_cell[   31432] = 32'h5cce1f50;
    ram_cell[   31433] = 32'h7e419fc5;
    ram_cell[   31434] = 32'h1180fd5a;
    ram_cell[   31435] = 32'h4112f8e0;
    ram_cell[   31436] = 32'hc0df7e0c;
    ram_cell[   31437] = 32'h08a12511;
    ram_cell[   31438] = 32'h2903480c;
    ram_cell[   31439] = 32'had659a05;
    ram_cell[   31440] = 32'h47f0582a;
    ram_cell[   31441] = 32'hfd518e19;
    ram_cell[   31442] = 32'h15e3f994;
    ram_cell[   31443] = 32'heec73184;
    ram_cell[   31444] = 32'h2f03b7a6;
    ram_cell[   31445] = 32'hdbe6a8f2;
    ram_cell[   31446] = 32'hcb941d99;
    ram_cell[   31447] = 32'h189fc347;
    ram_cell[   31448] = 32'h6a376e5b;
    ram_cell[   31449] = 32'h49405088;
    ram_cell[   31450] = 32'h16d2f6b9;
    ram_cell[   31451] = 32'h0089165a;
    ram_cell[   31452] = 32'h9c218dcc;
    ram_cell[   31453] = 32'h2053c79d;
    ram_cell[   31454] = 32'h323a7c1f;
    ram_cell[   31455] = 32'h962bc97b;
    ram_cell[   31456] = 32'h5ab50767;
    ram_cell[   31457] = 32'hcfd72b78;
    ram_cell[   31458] = 32'h6f8ed290;
    ram_cell[   31459] = 32'h29d4186b;
    ram_cell[   31460] = 32'h8a3d6f1f;
    ram_cell[   31461] = 32'hb8dffd99;
    ram_cell[   31462] = 32'hab0252d9;
    ram_cell[   31463] = 32'hd4ba211e;
    ram_cell[   31464] = 32'h6bcf8cbc;
    ram_cell[   31465] = 32'heee18a3d;
    ram_cell[   31466] = 32'he8331ff5;
    ram_cell[   31467] = 32'h030fd75d;
    ram_cell[   31468] = 32'he55802dc;
    ram_cell[   31469] = 32'h70fffe9b;
    ram_cell[   31470] = 32'h1ab98c44;
    ram_cell[   31471] = 32'h88f59eb1;
    ram_cell[   31472] = 32'h7d7be07f;
    ram_cell[   31473] = 32'h87a31b3a;
    ram_cell[   31474] = 32'h06362445;
    ram_cell[   31475] = 32'h9e3f09f4;
    ram_cell[   31476] = 32'hfb5b37d2;
    ram_cell[   31477] = 32'h0220000c;
    ram_cell[   31478] = 32'h719441fc;
    ram_cell[   31479] = 32'hfaee7da6;
    ram_cell[   31480] = 32'h9e5e10a9;
    ram_cell[   31481] = 32'h31c3e653;
    ram_cell[   31482] = 32'he7e503b5;
    ram_cell[   31483] = 32'hba48281d;
    ram_cell[   31484] = 32'he792ee96;
    ram_cell[   31485] = 32'hfaafa734;
    ram_cell[   31486] = 32'h5df9632f;
    ram_cell[   31487] = 32'h86d6cdf2;
    ram_cell[   31488] = 32'hdb5dc49c;
    ram_cell[   31489] = 32'h5467f5c2;
    ram_cell[   31490] = 32'hc21c3208;
    ram_cell[   31491] = 32'he08381f4;
    ram_cell[   31492] = 32'hc15bc8f3;
    ram_cell[   31493] = 32'h0b7198f9;
    ram_cell[   31494] = 32'h63a6df2b;
    ram_cell[   31495] = 32'hd7431fb9;
    ram_cell[   31496] = 32'hc921d0e9;
    ram_cell[   31497] = 32'h27b142d3;
    ram_cell[   31498] = 32'hdb032f82;
    ram_cell[   31499] = 32'hb032ae66;
    ram_cell[   31500] = 32'h699547eb;
    ram_cell[   31501] = 32'h96b56816;
    ram_cell[   31502] = 32'ha6d78af5;
    ram_cell[   31503] = 32'h8aef75c8;
    ram_cell[   31504] = 32'h3e841a5e;
    ram_cell[   31505] = 32'he8c2a64d;
    ram_cell[   31506] = 32'h77a56a4c;
    ram_cell[   31507] = 32'habb0eab6;
    ram_cell[   31508] = 32'hb1c03015;
    ram_cell[   31509] = 32'hf3c6e519;
    ram_cell[   31510] = 32'h7283324e;
    ram_cell[   31511] = 32'hd2b519be;
    ram_cell[   31512] = 32'h7e69f962;
    ram_cell[   31513] = 32'h86b9794d;
    ram_cell[   31514] = 32'h2a23136a;
    ram_cell[   31515] = 32'h06b11442;
    ram_cell[   31516] = 32'h94ed5ba5;
    ram_cell[   31517] = 32'h34ff2f3c;
    ram_cell[   31518] = 32'h4ceed4ff;
    ram_cell[   31519] = 32'h60fa910c;
    ram_cell[   31520] = 32'hfd2e66f1;
    ram_cell[   31521] = 32'hbbaa4c26;
    ram_cell[   31522] = 32'h1bcb5a87;
    ram_cell[   31523] = 32'h6b0eb28c;
    ram_cell[   31524] = 32'h667c0c49;
    ram_cell[   31525] = 32'h260b3f11;
    ram_cell[   31526] = 32'hd6faf233;
    ram_cell[   31527] = 32'he122ead8;
    ram_cell[   31528] = 32'hc402eab6;
    ram_cell[   31529] = 32'heb8b7442;
    ram_cell[   31530] = 32'h88ea5959;
    ram_cell[   31531] = 32'hb186fc29;
    ram_cell[   31532] = 32'hd8dd9956;
    ram_cell[   31533] = 32'ha2886b69;
    ram_cell[   31534] = 32'hf99f262c;
    ram_cell[   31535] = 32'h438cfb2b;
    ram_cell[   31536] = 32'h79fd962c;
    ram_cell[   31537] = 32'h431a8c7a;
    ram_cell[   31538] = 32'hda8a5d3b;
    ram_cell[   31539] = 32'ha16c729a;
    ram_cell[   31540] = 32'h36012c6e;
    ram_cell[   31541] = 32'h48bf9641;
    ram_cell[   31542] = 32'h70dbb732;
    ram_cell[   31543] = 32'he44f157b;
    ram_cell[   31544] = 32'h7a586ff3;
    ram_cell[   31545] = 32'h28ac2233;
    ram_cell[   31546] = 32'h91c3df32;
    ram_cell[   31547] = 32'h566292e7;
    ram_cell[   31548] = 32'h2d061ac8;
    ram_cell[   31549] = 32'hc0580da9;
    ram_cell[   31550] = 32'h45be2965;
    ram_cell[   31551] = 32'h06f3a8e6;
    ram_cell[   31552] = 32'h11e2ad8d;
    ram_cell[   31553] = 32'hc00c8a63;
    ram_cell[   31554] = 32'h073d41c9;
    ram_cell[   31555] = 32'h519ea48b;
    ram_cell[   31556] = 32'hd8a92cab;
    ram_cell[   31557] = 32'h649a3b0f;
    ram_cell[   31558] = 32'h477308a6;
    ram_cell[   31559] = 32'h6e5a7188;
    ram_cell[   31560] = 32'hfc23a072;
    ram_cell[   31561] = 32'hfb827c12;
    ram_cell[   31562] = 32'hd8b9abf6;
    ram_cell[   31563] = 32'h2c9bc9ec;
    ram_cell[   31564] = 32'h82bf8605;
    ram_cell[   31565] = 32'hea100cbd;
    ram_cell[   31566] = 32'h8e25993f;
    ram_cell[   31567] = 32'h97a3a88a;
    ram_cell[   31568] = 32'h702c4fed;
    ram_cell[   31569] = 32'hb4fd253b;
    ram_cell[   31570] = 32'h3c91063b;
    ram_cell[   31571] = 32'h58d23f65;
    ram_cell[   31572] = 32'h5387b8b8;
    ram_cell[   31573] = 32'h3d46e014;
    ram_cell[   31574] = 32'he12992cf;
    ram_cell[   31575] = 32'hdc97226d;
    ram_cell[   31576] = 32'h1776cf7e;
    ram_cell[   31577] = 32'h2d598e24;
    ram_cell[   31578] = 32'hbedf6602;
    ram_cell[   31579] = 32'h88ffcd54;
    ram_cell[   31580] = 32'h8409011f;
    ram_cell[   31581] = 32'h0a4ad2e6;
    ram_cell[   31582] = 32'h98a7bc86;
    ram_cell[   31583] = 32'ha7129af4;
    ram_cell[   31584] = 32'h3600d8d6;
    ram_cell[   31585] = 32'h26b62494;
    ram_cell[   31586] = 32'hbe3d8d4b;
    ram_cell[   31587] = 32'h500ecb02;
    ram_cell[   31588] = 32'hd40fc277;
    ram_cell[   31589] = 32'h72e6b18f;
    ram_cell[   31590] = 32'h0bff4d68;
    ram_cell[   31591] = 32'h3f39fae4;
    ram_cell[   31592] = 32'he2aaa79e;
    ram_cell[   31593] = 32'h2b1043b6;
    ram_cell[   31594] = 32'h08ea0a46;
    ram_cell[   31595] = 32'h013050e4;
    ram_cell[   31596] = 32'h11307af7;
    ram_cell[   31597] = 32'hab97c1cd;
    ram_cell[   31598] = 32'h58462c32;
    ram_cell[   31599] = 32'h0315ad3e;
    ram_cell[   31600] = 32'h42bf658c;
    ram_cell[   31601] = 32'h4ca3690b;
    ram_cell[   31602] = 32'h25b87d41;
    ram_cell[   31603] = 32'h0d0073b5;
    ram_cell[   31604] = 32'hdf1403e8;
    ram_cell[   31605] = 32'hb7283b36;
    ram_cell[   31606] = 32'hc6fb519a;
    ram_cell[   31607] = 32'h56fb44c4;
    ram_cell[   31608] = 32'h5ef793ab;
    ram_cell[   31609] = 32'h58b158f3;
    ram_cell[   31610] = 32'h537cf590;
    ram_cell[   31611] = 32'h53c4fb6a;
    ram_cell[   31612] = 32'h5f052eab;
    ram_cell[   31613] = 32'h693e48a1;
    ram_cell[   31614] = 32'he9a9a84c;
    ram_cell[   31615] = 32'h280a3901;
    ram_cell[   31616] = 32'hc847b6ec;
    ram_cell[   31617] = 32'ha1af752d;
    ram_cell[   31618] = 32'h33af55dc;
    ram_cell[   31619] = 32'h501d5a97;
    ram_cell[   31620] = 32'h2e0ba49e;
    ram_cell[   31621] = 32'hc8015e15;
    ram_cell[   31622] = 32'h4dfcf5bc;
    ram_cell[   31623] = 32'h427c1cd1;
    ram_cell[   31624] = 32'h463a6782;
    ram_cell[   31625] = 32'h19714f02;
    ram_cell[   31626] = 32'hf7796bf0;
    ram_cell[   31627] = 32'h2446ca7c;
    ram_cell[   31628] = 32'h2b797eb0;
    ram_cell[   31629] = 32'h7bc91a33;
    ram_cell[   31630] = 32'hef6c45ee;
    ram_cell[   31631] = 32'h8fbeb1f2;
    ram_cell[   31632] = 32'h30962f3a;
    ram_cell[   31633] = 32'hd885165c;
    ram_cell[   31634] = 32'hfe8c4d61;
    ram_cell[   31635] = 32'h1b55005e;
    ram_cell[   31636] = 32'h95b38ad2;
    ram_cell[   31637] = 32'h6e403713;
    ram_cell[   31638] = 32'h1fc4ae52;
    ram_cell[   31639] = 32'hfb78751e;
    ram_cell[   31640] = 32'h44d65632;
    ram_cell[   31641] = 32'h5fe25622;
    ram_cell[   31642] = 32'h738890ce;
    ram_cell[   31643] = 32'h8ee52ef0;
    ram_cell[   31644] = 32'hf7ce6383;
    ram_cell[   31645] = 32'h45d31fd0;
    ram_cell[   31646] = 32'hd742449f;
    ram_cell[   31647] = 32'h5c42021a;
    ram_cell[   31648] = 32'h5d3876ad;
    ram_cell[   31649] = 32'h573bb88e;
    ram_cell[   31650] = 32'h6fee15d7;
    ram_cell[   31651] = 32'h94750d03;
    ram_cell[   31652] = 32'h9de7dbe1;
    ram_cell[   31653] = 32'h30fa0466;
    ram_cell[   31654] = 32'hf61e5aa9;
    ram_cell[   31655] = 32'h2f97bdcf;
    ram_cell[   31656] = 32'hff94f1fe;
    ram_cell[   31657] = 32'haff4cb90;
    ram_cell[   31658] = 32'h354c5e73;
    ram_cell[   31659] = 32'h4e6f1cfd;
    ram_cell[   31660] = 32'hf46614eb;
    ram_cell[   31661] = 32'h3822c875;
    ram_cell[   31662] = 32'ha7220412;
    ram_cell[   31663] = 32'h5628252f;
    ram_cell[   31664] = 32'heec73ce5;
    ram_cell[   31665] = 32'h08ca47ba;
    ram_cell[   31666] = 32'h918cce40;
    ram_cell[   31667] = 32'h62e8b162;
    ram_cell[   31668] = 32'h57aa6806;
    ram_cell[   31669] = 32'h092e3c9c;
    ram_cell[   31670] = 32'h582ea5db;
    ram_cell[   31671] = 32'h7cc2284d;
    ram_cell[   31672] = 32'h45c40cd7;
    ram_cell[   31673] = 32'h385e1e7f;
    ram_cell[   31674] = 32'hd4e13cb8;
    ram_cell[   31675] = 32'h7c22a175;
    ram_cell[   31676] = 32'hd001f8fb;
    ram_cell[   31677] = 32'h36b0cedd;
    ram_cell[   31678] = 32'h29c84220;
    ram_cell[   31679] = 32'hd73b9d79;
    ram_cell[   31680] = 32'h355e57f2;
    ram_cell[   31681] = 32'h945b6f9a;
    ram_cell[   31682] = 32'h322e98b8;
    ram_cell[   31683] = 32'h6a3e8a9a;
    ram_cell[   31684] = 32'hcc9d40cc;
    ram_cell[   31685] = 32'hdbeed780;
    ram_cell[   31686] = 32'ha26f1ef6;
    ram_cell[   31687] = 32'hd859e4c7;
    ram_cell[   31688] = 32'hedf54441;
    ram_cell[   31689] = 32'h1ddee921;
    ram_cell[   31690] = 32'hd09c9c41;
    ram_cell[   31691] = 32'h1a1f785e;
    ram_cell[   31692] = 32'hd7bd52a6;
    ram_cell[   31693] = 32'h03019925;
    ram_cell[   31694] = 32'h26925b7f;
    ram_cell[   31695] = 32'h566f7f4b;
    ram_cell[   31696] = 32'hf08336ec;
    ram_cell[   31697] = 32'h1a86aea1;
    ram_cell[   31698] = 32'hc017a0a0;
    ram_cell[   31699] = 32'h3339c57e;
    ram_cell[   31700] = 32'hb8d695e2;
    ram_cell[   31701] = 32'h277df0cd;
    ram_cell[   31702] = 32'h05432221;
    ram_cell[   31703] = 32'h1e472345;
    ram_cell[   31704] = 32'hf176c90e;
    ram_cell[   31705] = 32'h358f5de8;
    ram_cell[   31706] = 32'h47eae7a5;
    ram_cell[   31707] = 32'hb19c00ba;
    ram_cell[   31708] = 32'h76f71fbb;
    ram_cell[   31709] = 32'h57a35a0c;
    ram_cell[   31710] = 32'h5697dbfd;
    ram_cell[   31711] = 32'haa5b0800;
    ram_cell[   31712] = 32'h48a6764a;
    ram_cell[   31713] = 32'h5ff1d093;
    ram_cell[   31714] = 32'h99063300;
    ram_cell[   31715] = 32'h6003d7a7;
    ram_cell[   31716] = 32'h42c8cf99;
    ram_cell[   31717] = 32'h2e74edd8;
    ram_cell[   31718] = 32'h153283f3;
    ram_cell[   31719] = 32'hd997348e;
    ram_cell[   31720] = 32'h23e52bdc;
    ram_cell[   31721] = 32'he13d4ffa;
    ram_cell[   31722] = 32'hdedceff0;
    ram_cell[   31723] = 32'hbfd3fa1e;
    ram_cell[   31724] = 32'h5aaaeac9;
    ram_cell[   31725] = 32'h46415fed;
    ram_cell[   31726] = 32'hf09dc1d1;
    ram_cell[   31727] = 32'hab519ffa;
    ram_cell[   31728] = 32'ha21b6d79;
    ram_cell[   31729] = 32'h3ab3392c;
    ram_cell[   31730] = 32'hbb7d343f;
    ram_cell[   31731] = 32'he72d3825;
    ram_cell[   31732] = 32'hc1fdfbc2;
    ram_cell[   31733] = 32'h40be665d;
    ram_cell[   31734] = 32'h264de162;
    ram_cell[   31735] = 32'h4c4caf1b;
    ram_cell[   31736] = 32'h42c7f421;
    ram_cell[   31737] = 32'hd8c6b1fc;
    ram_cell[   31738] = 32'h80dca18e;
    ram_cell[   31739] = 32'ha313d2ac;
    ram_cell[   31740] = 32'h75c163c4;
    ram_cell[   31741] = 32'ha5842ee3;
    ram_cell[   31742] = 32'h1db1fbbb;
    ram_cell[   31743] = 32'hd0510482;
    ram_cell[   31744] = 32'h81d06247;
    ram_cell[   31745] = 32'h8e1f5815;
    ram_cell[   31746] = 32'h30c04c28;
    ram_cell[   31747] = 32'hb023eecb;
    ram_cell[   31748] = 32'hd10ad628;
    ram_cell[   31749] = 32'h4b9580e7;
    ram_cell[   31750] = 32'haa5386c7;
    ram_cell[   31751] = 32'hea0669ba;
    ram_cell[   31752] = 32'hf03ea8a6;
    ram_cell[   31753] = 32'h8995b325;
    ram_cell[   31754] = 32'h9ef160a0;
    ram_cell[   31755] = 32'h03a90b2d;
    ram_cell[   31756] = 32'h5184b05b;
    ram_cell[   31757] = 32'h971d361a;
    ram_cell[   31758] = 32'hf981b6ff;
    ram_cell[   31759] = 32'hdc0425aa;
    ram_cell[   31760] = 32'h69589cbd;
    ram_cell[   31761] = 32'h14035b84;
    ram_cell[   31762] = 32'hb43f8a5d;
    ram_cell[   31763] = 32'hf22403b2;
    ram_cell[   31764] = 32'ha5632e77;
    ram_cell[   31765] = 32'h559074a5;
    ram_cell[   31766] = 32'h3fef41c0;
    ram_cell[   31767] = 32'h8500865c;
    ram_cell[   31768] = 32'h9d0f66d1;
    ram_cell[   31769] = 32'h558f9a7a;
    ram_cell[   31770] = 32'h3f4e0111;
    ram_cell[   31771] = 32'h7a3f8aa3;
    ram_cell[   31772] = 32'h65bf893f;
    ram_cell[   31773] = 32'hf4121638;
    ram_cell[   31774] = 32'haa92cedf;
    ram_cell[   31775] = 32'h7f95d458;
    ram_cell[   31776] = 32'h3219f027;
    ram_cell[   31777] = 32'h20693cde;
    ram_cell[   31778] = 32'hf4ca6703;
    ram_cell[   31779] = 32'hb2c6526e;
    ram_cell[   31780] = 32'h8e149b4d;
    ram_cell[   31781] = 32'h9a6d5c5e;
    ram_cell[   31782] = 32'h6617c323;
    ram_cell[   31783] = 32'hf05c198f;
    ram_cell[   31784] = 32'h1c56967a;
    ram_cell[   31785] = 32'h918cdca9;
    ram_cell[   31786] = 32'he6becb00;
    ram_cell[   31787] = 32'hb76e9da6;
    ram_cell[   31788] = 32'hce9683c4;
    ram_cell[   31789] = 32'h7a5c469b;
    ram_cell[   31790] = 32'h8d4b991c;
    ram_cell[   31791] = 32'h5ee808b3;
    ram_cell[   31792] = 32'hc0ae3d7a;
    ram_cell[   31793] = 32'hd96ce424;
    ram_cell[   31794] = 32'hc25f3509;
    ram_cell[   31795] = 32'hd2e164ef;
    ram_cell[   31796] = 32'h3d5f6c2a;
    ram_cell[   31797] = 32'h1cb5d962;
    ram_cell[   31798] = 32'h87445f27;
    ram_cell[   31799] = 32'h37f28def;
    ram_cell[   31800] = 32'hecca1ee8;
    ram_cell[   31801] = 32'hcf597837;
    ram_cell[   31802] = 32'h1277f61e;
    ram_cell[   31803] = 32'h17ada489;
    ram_cell[   31804] = 32'h866e1658;
    ram_cell[   31805] = 32'h117f775b;
    ram_cell[   31806] = 32'h0fb60eed;
    ram_cell[   31807] = 32'hd3a5f712;
    ram_cell[   31808] = 32'hafd1f8ac;
    ram_cell[   31809] = 32'h7ab0397f;
    ram_cell[   31810] = 32'h266df834;
    ram_cell[   31811] = 32'h39db8ad7;
    ram_cell[   31812] = 32'h28b9a8ab;
    ram_cell[   31813] = 32'h3473808a;
    ram_cell[   31814] = 32'h8885e3a3;
    ram_cell[   31815] = 32'hb364dfe1;
    ram_cell[   31816] = 32'h0c0b171a;
    ram_cell[   31817] = 32'h717e0032;
    ram_cell[   31818] = 32'h9180f9fe;
    ram_cell[   31819] = 32'h6d8106f1;
    ram_cell[   31820] = 32'h9b94fb6b;
    ram_cell[   31821] = 32'h121c8040;
    ram_cell[   31822] = 32'h52ca7c16;
    ram_cell[   31823] = 32'h31750005;
    ram_cell[   31824] = 32'h11979b99;
    ram_cell[   31825] = 32'hc9f8a53a;
    ram_cell[   31826] = 32'h35b783e3;
    ram_cell[   31827] = 32'h3ebf1240;
    ram_cell[   31828] = 32'h63fb86cc;
    ram_cell[   31829] = 32'ha54002c1;
    ram_cell[   31830] = 32'hfeea78e9;
    ram_cell[   31831] = 32'h73e0dd3c;
    ram_cell[   31832] = 32'ha6025b5f;
    ram_cell[   31833] = 32'h735018c6;
    ram_cell[   31834] = 32'h7f17daa3;
    ram_cell[   31835] = 32'h0290c610;
    ram_cell[   31836] = 32'h33ec346a;
    ram_cell[   31837] = 32'h77286125;
    ram_cell[   31838] = 32'he19d018a;
    ram_cell[   31839] = 32'h2a115e93;
    ram_cell[   31840] = 32'h135eed76;
    ram_cell[   31841] = 32'h779e63ab;
    ram_cell[   31842] = 32'h7f428b21;
    ram_cell[   31843] = 32'hb3248550;
    ram_cell[   31844] = 32'h2dbed4ee;
    ram_cell[   31845] = 32'h3fed6789;
    ram_cell[   31846] = 32'h7085023e;
    ram_cell[   31847] = 32'h9005b24f;
    ram_cell[   31848] = 32'h1c9e6811;
    ram_cell[   31849] = 32'hb463bccd;
    ram_cell[   31850] = 32'h426a2fd8;
    ram_cell[   31851] = 32'h8c5f7793;
    ram_cell[   31852] = 32'h21b0110b;
    ram_cell[   31853] = 32'h13ac0b15;
    ram_cell[   31854] = 32'h46061c7c;
    ram_cell[   31855] = 32'h534ec5f6;
    ram_cell[   31856] = 32'hb24fcba7;
    ram_cell[   31857] = 32'h1bdda6d9;
    ram_cell[   31858] = 32'h3c4a5ce6;
    ram_cell[   31859] = 32'h9c600171;
    ram_cell[   31860] = 32'h3e239ef8;
    ram_cell[   31861] = 32'h75b6cea1;
    ram_cell[   31862] = 32'h5154eaf1;
    ram_cell[   31863] = 32'h368da7f4;
    ram_cell[   31864] = 32'h89139563;
    ram_cell[   31865] = 32'h01eee4c5;
    ram_cell[   31866] = 32'h459c3d1f;
    ram_cell[   31867] = 32'h9b24969c;
    ram_cell[   31868] = 32'h44452313;
    ram_cell[   31869] = 32'h06141be7;
    ram_cell[   31870] = 32'h3df6570c;
    ram_cell[   31871] = 32'h3cfc69dd;
    ram_cell[   31872] = 32'hf926e1bc;
    ram_cell[   31873] = 32'h0764a4b4;
    ram_cell[   31874] = 32'h3fab1c0d;
    ram_cell[   31875] = 32'h2acf6d63;
    ram_cell[   31876] = 32'h2fa0f2a8;
    ram_cell[   31877] = 32'hd406e754;
    ram_cell[   31878] = 32'he17b65f9;
    ram_cell[   31879] = 32'h4b1b17a5;
    ram_cell[   31880] = 32'h3c0f5df2;
    ram_cell[   31881] = 32'h29937127;
    ram_cell[   31882] = 32'h578e92de;
    ram_cell[   31883] = 32'hef61d703;
    ram_cell[   31884] = 32'hed79be38;
    ram_cell[   31885] = 32'h7c7605e7;
    ram_cell[   31886] = 32'h1b6b33de;
    ram_cell[   31887] = 32'h7c784d9c;
    ram_cell[   31888] = 32'hc36d86cd;
    ram_cell[   31889] = 32'h94d13984;
    ram_cell[   31890] = 32'h20189d43;
    ram_cell[   31891] = 32'h512c2f63;
    ram_cell[   31892] = 32'hd76c5931;
    ram_cell[   31893] = 32'h6c24f072;
    ram_cell[   31894] = 32'h21bf191e;
    ram_cell[   31895] = 32'hd2f2f517;
    ram_cell[   31896] = 32'h984728f0;
    ram_cell[   31897] = 32'h63794b93;
    ram_cell[   31898] = 32'h12651721;
    ram_cell[   31899] = 32'h4656ff02;
    ram_cell[   31900] = 32'hdf54fe3b;
    ram_cell[   31901] = 32'h83795ba5;
    ram_cell[   31902] = 32'hf7964980;
    ram_cell[   31903] = 32'h53f9a0c1;
    ram_cell[   31904] = 32'h28512af7;
    ram_cell[   31905] = 32'h5268dcf7;
    ram_cell[   31906] = 32'ha87ae8c1;
    ram_cell[   31907] = 32'h68802230;
    ram_cell[   31908] = 32'h70720f1e;
    ram_cell[   31909] = 32'he2657038;
    ram_cell[   31910] = 32'hedcfe77d;
    ram_cell[   31911] = 32'h9587ed94;
    ram_cell[   31912] = 32'haaeae126;
    ram_cell[   31913] = 32'hab12b293;
    ram_cell[   31914] = 32'h7618fc2f;
    ram_cell[   31915] = 32'h85a34647;
    ram_cell[   31916] = 32'h6a23f525;
    ram_cell[   31917] = 32'h1ebd104d;
    ram_cell[   31918] = 32'h0b0dad19;
    ram_cell[   31919] = 32'ha481478c;
    ram_cell[   31920] = 32'h6e77e0c2;
    ram_cell[   31921] = 32'h821ff361;
    ram_cell[   31922] = 32'h7e743a5b;
    ram_cell[   31923] = 32'hee9e011f;
    ram_cell[   31924] = 32'hbe06fa62;
    ram_cell[   31925] = 32'h5a632f7e;
    ram_cell[   31926] = 32'h33285de9;
    ram_cell[   31927] = 32'h4e98f359;
    ram_cell[   31928] = 32'he6fed29a;
    ram_cell[   31929] = 32'h40df02f2;
    ram_cell[   31930] = 32'ha5e0c555;
    ram_cell[   31931] = 32'h382b9d3f;
    ram_cell[   31932] = 32'ha407b6c5;
    ram_cell[   31933] = 32'h84daa42b;
    ram_cell[   31934] = 32'h618eb253;
    ram_cell[   31935] = 32'hcf620a5d;
    ram_cell[   31936] = 32'h081db95e;
    ram_cell[   31937] = 32'h7ce84b09;
    ram_cell[   31938] = 32'h465baaf4;
    ram_cell[   31939] = 32'hc9653ab7;
    ram_cell[   31940] = 32'hb51dc52d;
    ram_cell[   31941] = 32'h26463b87;
    ram_cell[   31942] = 32'h05540206;
    ram_cell[   31943] = 32'hcf33c34f;
    ram_cell[   31944] = 32'h7b262775;
    ram_cell[   31945] = 32'h946ed602;
    ram_cell[   31946] = 32'h38c34f58;
    ram_cell[   31947] = 32'h49b936b0;
    ram_cell[   31948] = 32'hcb10297a;
    ram_cell[   31949] = 32'ha6a5dccc;
    ram_cell[   31950] = 32'h96778c04;
    ram_cell[   31951] = 32'h2c849999;
    ram_cell[   31952] = 32'h6c666052;
    ram_cell[   31953] = 32'h505485f5;
    ram_cell[   31954] = 32'h95d491c7;
    ram_cell[   31955] = 32'h0a4187df;
    ram_cell[   31956] = 32'hec1cc438;
    ram_cell[   31957] = 32'hd20d7f89;
    ram_cell[   31958] = 32'h02f92d1e;
    ram_cell[   31959] = 32'h60c24624;
    ram_cell[   31960] = 32'h8abdd789;
    ram_cell[   31961] = 32'hb60aa914;
    ram_cell[   31962] = 32'h37a8133a;
    ram_cell[   31963] = 32'h8c61c679;
    ram_cell[   31964] = 32'he60796ec;
    ram_cell[   31965] = 32'h927cac7c;
    ram_cell[   31966] = 32'he3347904;
    ram_cell[   31967] = 32'h70808a3e;
    ram_cell[   31968] = 32'h4ffbc991;
    ram_cell[   31969] = 32'he2894d5f;
    ram_cell[   31970] = 32'h3904448a;
    ram_cell[   31971] = 32'h210c5b52;
    ram_cell[   31972] = 32'he34a286d;
    ram_cell[   31973] = 32'h8e0117c9;
    ram_cell[   31974] = 32'h2cb596c6;
    ram_cell[   31975] = 32'hbc5b6e25;
    ram_cell[   31976] = 32'h25b2d88f;
    ram_cell[   31977] = 32'hf5e985cf;
    ram_cell[   31978] = 32'he87a0403;
    ram_cell[   31979] = 32'h94bc44ea;
    ram_cell[   31980] = 32'hcebb7813;
    ram_cell[   31981] = 32'h80f69de5;
    ram_cell[   31982] = 32'hecb35f58;
    ram_cell[   31983] = 32'hc6fbe373;
    ram_cell[   31984] = 32'h2bc7e647;
    ram_cell[   31985] = 32'h35995d3a;
    ram_cell[   31986] = 32'h3ab04c17;
    ram_cell[   31987] = 32'h34b5c8fa;
    ram_cell[   31988] = 32'h4977f5fc;
    ram_cell[   31989] = 32'h81184194;
    ram_cell[   31990] = 32'h03448f00;
    ram_cell[   31991] = 32'h51d9013b;
    ram_cell[   31992] = 32'h5dac60c3;
    ram_cell[   31993] = 32'h6e8bb259;
    ram_cell[   31994] = 32'hf6d7a940;
    ram_cell[   31995] = 32'ha940b0d1;
    ram_cell[   31996] = 32'ha00a0a64;
    ram_cell[   31997] = 32'h33eeb0bf;
    ram_cell[   31998] = 32'hb1962124;
    ram_cell[   31999] = 32'h90752edb;
    ram_cell[   32000] = 32'h695b4bf5;
    ram_cell[   32001] = 32'h99092a1d;
    ram_cell[   32002] = 32'h8ca8b4bd;
    ram_cell[   32003] = 32'h7414aa9c;
    ram_cell[   32004] = 32'hfb188b09;
    ram_cell[   32005] = 32'h6c1115b2;
    ram_cell[   32006] = 32'h7fd248dd;
    ram_cell[   32007] = 32'h18334e52;
    ram_cell[   32008] = 32'h2c8086f2;
    ram_cell[   32009] = 32'h10c32228;
    ram_cell[   32010] = 32'hb57d8fb0;
    ram_cell[   32011] = 32'h3a46955f;
    ram_cell[   32012] = 32'ha7e4582d;
    ram_cell[   32013] = 32'h8d354a03;
    ram_cell[   32014] = 32'h9d88a5a4;
    ram_cell[   32015] = 32'h7bc3c949;
    ram_cell[   32016] = 32'h9b3cb0b6;
    ram_cell[   32017] = 32'hb0ef458b;
    ram_cell[   32018] = 32'hd15c31f8;
    ram_cell[   32019] = 32'ha8b8a313;
    ram_cell[   32020] = 32'hc6bcc1f1;
    ram_cell[   32021] = 32'h0c979b57;
    ram_cell[   32022] = 32'hf64c2032;
    ram_cell[   32023] = 32'heaafc326;
    ram_cell[   32024] = 32'hb1d2e3fe;
    ram_cell[   32025] = 32'ha485f960;
    ram_cell[   32026] = 32'he3b82f62;
    ram_cell[   32027] = 32'hb3a580cb;
    ram_cell[   32028] = 32'hb0e5a4c5;
    ram_cell[   32029] = 32'hf23dbadb;
    ram_cell[   32030] = 32'h6e862fd1;
    ram_cell[   32031] = 32'h5c69260e;
    ram_cell[   32032] = 32'hc82eb5c4;
    ram_cell[   32033] = 32'h9e2d58f0;
    ram_cell[   32034] = 32'hc45721c1;
    ram_cell[   32035] = 32'ha5ff8045;
    ram_cell[   32036] = 32'hf8cd5150;
    ram_cell[   32037] = 32'hbef10858;
    ram_cell[   32038] = 32'h01d4d640;
    ram_cell[   32039] = 32'hf5ecf71d;
    ram_cell[   32040] = 32'hd476082f;
    ram_cell[   32041] = 32'h5b4faafd;
    ram_cell[   32042] = 32'h127e8df2;
    ram_cell[   32043] = 32'h0ba5c37f;
    ram_cell[   32044] = 32'h0217fe34;
    ram_cell[   32045] = 32'hc6672784;
    ram_cell[   32046] = 32'h8b0c3b19;
    ram_cell[   32047] = 32'hb716a0c6;
    ram_cell[   32048] = 32'hd3252e8e;
    ram_cell[   32049] = 32'hab3642a3;
    ram_cell[   32050] = 32'hfc8f4f3c;
    ram_cell[   32051] = 32'hd204a800;
    ram_cell[   32052] = 32'h2c332648;
    ram_cell[   32053] = 32'hca201687;
    ram_cell[   32054] = 32'h6e61a6a5;
    ram_cell[   32055] = 32'h7cb05682;
    ram_cell[   32056] = 32'h5db22a6a;
    ram_cell[   32057] = 32'h7973feb4;
    ram_cell[   32058] = 32'hd101c6bc;
    ram_cell[   32059] = 32'hb96937db;
    ram_cell[   32060] = 32'hfa37c92c;
    ram_cell[   32061] = 32'h5a27086b;
    ram_cell[   32062] = 32'h48377ae4;
    ram_cell[   32063] = 32'h1571efb8;
    ram_cell[   32064] = 32'hbf0acb0a;
    ram_cell[   32065] = 32'h9eac2c2a;
    ram_cell[   32066] = 32'h9a739d32;
    ram_cell[   32067] = 32'ha31ab6b3;
    ram_cell[   32068] = 32'h0f8f9158;
    ram_cell[   32069] = 32'hbc8e9481;
    ram_cell[   32070] = 32'hf75cbe2b;
    ram_cell[   32071] = 32'h549006e4;
    ram_cell[   32072] = 32'hc4d5bdbd;
    ram_cell[   32073] = 32'ha33c5ca2;
    ram_cell[   32074] = 32'h4cfc3e5c;
    ram_cell[   32075] = 32'h9c91d1f7;
    ram_cell[   32076] = 32'h5ebd11fd;
    ram_cell[   32077] = 32'he8cd4755;
    ram_cell[   32078] = 32'h893e5190;
    ram_cell[   32079] = 32'h1d9b3f7a;
    ram_cell[   32080] = 32'hd947ce47;
    ram_cell[   32081] = 32'hcca0bc73;
    ram_cell[   32082] = 32'hb1dfefc3;
    ram_cell[   32083] = 32'h38e17fc8;
    ram_cell[   32084] = 32'h0cd45ab5;
    ram_cell[   32085] = 32'hd07ece3b;
    ram_cell[   32086] = 32'h2a2a1cd4;
    ram_cell[   32087] = 32'h357ed804;
    ram_cell[   32088] = 32'hc6843d52;
    ram_cell[   32089] = 32'h4db55ef9;
    ram_cell[   32090] = 32'hb6f44128;
    ram_cell[   32091] = 32'hf3bdf4fd;
    ram_cell[   32092] = 32'h470ee4fa;
    ram_cell[   32093] = 32'h4fb86064;
    ram_cell[   32094] = 32'h37f6c8cd;
    ram_cell[   32095] = 32'h6a477743;
    ram_cell[   32096] = 32'h63f76f2e;
    ram_cell[   32097] = 32'hfbf6d90e;
    ram_cell[   32098] = 32'h1ba73731;
    ram_cell[   32099] = 32'h83d54483;
    ram_cell[   32100] = 32'h57566c8f;
    ram_cell[   32101] = 32'h6c38a160;
    ram_cell[   32102] = 32'h67b48c8e;
    ram_cell[   32103] = 32'hc6ef167f;
    ram_cell[   32104] = 32'h45a6ccb5;
    ram_cell[   32105] = 32'h25600557;
    ram_cell[   32106] = 32'h111cd378;
    ram_cell[   32107] = 32'h95b2c23a;
    ram_cell[   32108] = 32'hbec388ba;
    ram_cell[   32109] = 32'ha2b9ab36;
    ram_cell[   32110] = 32'h7cd52a83;
    ram_cell[   32111] = 32'hfdbf3ca2;
    ram_cell[   32112] = 32'h9a2d013a;
    ram_cell[   32113] = 32'h8c83c762;
    ram_cell[   32114] = 32'h782579d3;
    ram_cell[   32115] = 32'hbc67ecb7;
    ram_cell[   32116] = 32'h566123ee;
    ram_cell[   32117] = 32'hbd9a1ee4;
    ram_cell[   32118] = 32'ha55b839c;
    ram_cell[   32119] = 32'h6a5966a3;
    ram_cell[   32120] = 32'h36542364;
    ram_cell[   32121] = 32'h70beadab;
    ram_cell[   32122] = 32'h656dffbb;
    ram_cell[   32123] = 32'hb481f0a2;
    ram_cell[   32124] = 32'hca7c0b50;
    ram_cell[   32125] = 32'h1d9f1291;
    ram_cell[   32126] = 32'hf5749b8c;
    ram_cell[   32127] = 32'h2c8dc943;
    ram_cell[   32128] = 32'h9a965f17;
    ram_cell[   32129] = 32'h80fc267c;
    ram_cell[   32130] = 32'h9bfdf032;
    ram_cell[   32131] = 32'hf501a89b;
    ram_cell[   32132] = 32'h6c122f45;
    ram_cell[   32133] = 32'h5493b537;
    ram_cell[   32134] = 32'hda663206;
    ram_cell[   32135] = 32'h87cfd54e;
    ram_cell[   32136] = 32'h3d48d055;
    ram_cell[   32137] = 32'h51075f70;
    ram_cell[   32138] = 32'h04ebb496;
    ram_cell[   32139] = 32'ha81c7d32;
    ram_cell[   32140] = 32'hbb87f463;
    ram_cell[   32141] = 32'h9657b518;
    ram_cell[   32142] = 32'h3eccd134;
    ram_cell[   32143] = 32'h80e16679;
    ram_cell[   32144] = 32'h46ad4542;
    ram_cell[   32145] = 32'h7d575c3b;
    ram_cell[   32146] = 32'hafc1322a;
    ram_cell[   32147] = 32'h8e5aa6a7;
    ram_cell[   32148] = 32'h05c076da;
    ram_cell[   32149] = 32'h7ef8b3e6;
    ram_cell[   32150] = 32'hc963e6cf;
    ram_cell[   32151] = 32'hc5b64ac9;
    ram_cell[   32152] = 32'ha7ac8beb;
    ram_cell[   32153] = 32'hb8dc7c5d;
    ram_cell[   32154] = 32'h6925f11a;
    ram_cell[   32155] = 32'h67597d42;
    ram_cell[   32156] = 32'h596cf20a;
    ram_cell[   32157] = 32'h324977f5;
    ram_cell[   32158] = 32'h2348f945;
    ram_cell[   32159] = 32'hc3edd5e2;
    ram_cell[   32160] = 32'h95627035;
    ram_cell[   32161] = 32'he4397728;
    ram_cell[   32162] = 32'hc90255b9;
    ram_cell[   32163] = 32'h7c99edf9;
    ram_cell[   32164] = 32'h7d931394;
    ram_cell[   32165] = 32'h78db3f90;
    ram_cell[   32166] = 32'h63fba8d8;
    ram_cell[   32167] = 32'hf204efb8;
    ram_cell[   32168] = 32'hf520d8ed;
    ram_cell[   32169] = 32'ha7ff3d7d;
    ram_cell[   32170] = 32'h3292e2bb;
    ram_cell[   32171] = 32'h3069ad56;
    ram_cell[   32172] = 32'he633eb06;
    ram_cell[   32173] = 32'hf6ffc6c4;
    ram_cell[   32174] = 32'hd27d4c7b;
    ram_cell[   32175] = 32'ha5436419;
    ram_cell[   32176] = 32'hc6520751;
    ram_cell[   32177] = 32'h11b965ac;
    ram_cell[   32178] = 32'h54522a59;
    ram_cell[   32179] = 32'h2fd3f04e;
    ram_cell[   32180] = 32'h8e911c3a;
    ram_cell[   32181] = 32'hdfc7420e;
    ram_cell[   32182] = 32'hd5129934;
    ram_cell[   32183] = 32'h6787dc43;
    ram_cell[   32184] = 32'h449e0a4d;
    ram_cell[   32185] = 32'hd46b85f4;
    ram_cell[   32186] = 32'hd7ab1276;
    ram_cell[   32187] = 32'hdaa7ec7a;
    ram_cell[   32188] = 32'h84be94ec;
    ram_cell[   32189] = 32'hf6b89ad9;
    ram_cell[   32190] = 32'hbec0fdab;
    ram_cell[   32191] = 32'h442c651a;
    ram_cell[   32192] = 32'h5ed60355;
    ram_cell[   32193] = 32'h7c9a8a4a;
    ram_cell[   32194] = 32'h9db1baa2;
    ram_cell[   32195] = 32'hfd0d4e65;
    ram_cell[   32196] = 32'hf0f70abc;
    ram_cell[   32197] = 32'h4a5ad813;
    ram_cell[   32198] = 32'h4709d356;
    ram_cell[   32199] = 32'h315ec3aa;
    ram_cell[   32200] = 32'h5aa25277;
    ram_cell[   32201] = 32'h1553a5f5;
    ram_cell[   32202] = 32'h8048ec91;
    ram_cell[   32203] = 32'h33ec74c4;
    ram_cell[   32204] = 32'hb8d27807;
    ram_cell[   32205] = 32'h948b08c8;
    ram_cell[   32206] = 32'hcbedc9d5;
    ram_cell[   32207] = 32'h0fd02e54;
    ram_cell[   32208] = 32'hd3957ed0;
    ram_cell[   32209] = 32'h5d1a4a3a;
    ram_cell[   32210] = 32'hc8a3e660;
    ram_cell[   32211] = 32'h89af4029;
    ram_cell[   32212] = 32'hddebfc91;
    ram_cell[   32213] = 32'had64c7a5;
    ram_cell[   32214] = 32'hac371ee6;
    ram_cell[   32215] = 32'h5810fb51;
    ram_cell[   32216] = 32'h816e9598;
    ram_cell[   32217] = 32'hca920b3b;
    ram_cell[   32218] = 32'h4a93e08c;
    ram_cell[   32219] = 32'h780f0de5;
    ram_cell[   32220] = 32'h5cf4026d;
    ram_cell[   32221] = 32'ha9aed288;
    ram_cell[   32222] = 32'hd90efbf1;
    ram_cell[   32223] = 32'h3151e01a;
    ram_cell[   32224] = 32'hd15bae56;
    ram_cell[   32225] = 32'hecebeb02;
    ram_cell[   32226] = 32'h99c0e3db;
    ram_cell[   32227] = 32'h487cdca8;
    ram_cell[   32228] = 32'h5dabc0fa;
    ram_cell[   32229] = 32'h48490a42;
    ram_cell[   32230] = 32'habd676b7;
    ram_cell[   32231] = 32'h2b0d1bb6;
    ram_cell[   32232] = 32'h5d3b5222;
    ram_cell[   32233] = 32'hfb62d406;
    ram_cell[   32234] = 32'h745ca825;
    ram_cell[   32235] = 32'h6935a5d8;
    ram_cell[   32236] = 32'h2e79e935;
    ram_cell[   32237] = 32'h6c2edb84;
    ram_cell[   32238] = 32'h9b95a398;
    ram_cell[   32239] = 32'h1174b411;
    ram_cell[   32240] = 32'h70c5d4b2;
    ram_cell[   32241] = 32'hbfb97c14;
    ram_cell[   32242] = 32'h37769f7d;
    ram_cell[   32243] = 32'h09f4f77d;
    ram_cell[   32244] = 32'he8fae4e9;
    ram_cell[   32245] = 32'h6a4ee0cb;
    ram_cell[   32246] = 32'h72db9782;
    ram_cell[   32247] = 32'hb93b21ec;
    ram_cell[   32248] = 32'hc2ce8ce6;
    ram_cell[   32249] = 32'h8de0e683;
    ram_cell[   32250] = 32'h0e43597f;
    ram_cell[   32251] = 32'hb7e8560c;
    ram_cell[   32252] = 32'h1ece5883;
    ram_cell[   32253] = 32'h0ef8675c;
    ram_cell[   32254] = 32'he299014f;
    ram_cell[   32255] = 32'hb23d0037;
    ram_cell[   32256] = 32'h83df4240;
    ram_cell[   32257] = 32'h5aeab3fd;
    ram_cell[   32258] = 32'hb0d76298;
    ram_cell[   32259] = 32'h571c0edd;
    ram_cell[   32260] = 32'h34711c51;
    ram_cell[   32261] = 32'hcd83d847;
    ram_cell[   32262] = 32'h46e1964f;
    ram_cell[   32263] = 32'h9788b401;
    ram_cell[   32264] = 32'h5575d7d2;
    ram_cell[   32265] = 32'h1183ecb5;
    ram_cell[   32266] = 32'h14c8abd6;
    ram_cell[   32267] = 32'h8c33519a;
    ram_cell[   32268] = 32'hf6c13f82;
    ram_cell[   32269] = 32'h9d004d1a;
    ram_cell[   32270] = 32'h36281b8c;
    ram_cell[   32271] = 32'h73583baa;
    ram_cell[   32272] = 32'h62539400;
    ram_cell[   32273] = 32'hecd87d0e;
    ram_cell[   32274] = 32'h9504dca5;
    ram_cell[   32275] = 32'h5ec1fd36;
    ram_cell[   32276] = 32'he27e5159;
    ram_cell[   32277] = 32'h0f6c96a8;
    ram_cell[   32278] = 32'h4feffe9e;
    ram_cell[   32279] = 32'h709bc8eb;
    ram_cell[   32280] = 32'h62391eb1;
    ram_cell[   32281] = 32'hc3ad247d;
    ram_cell[   32282] = 32'h93079ad5;
    ram_cell[   32283] = 32'h693896b0;
    ram_cell[   32284] = 32'hf886e35a;
    ram_cell[   32285] = 32'h5f8dccdc;
    ram_cell[   32286] = 32'hc25a0ee2;
    ram_cell[   32287] = 32'h7d7ffdeb;
    ram_cell[   32288] = 32'h08703d18;
    ram_cell[   32289] = 32'h73b2e104;
    ram_cell[   32290] = 32'h7873988f;
    ram_cell[   32291] = 32'ha81926c2;
    ram_cell[   32292] = 32'h17f1e5da;
    ram_cell[   32293] = 32'h1e12f095;
    ram_cell[   32294] = 32'hcf10aab9;
    ram_cell[   32295] = 32'h80668803;
    ram_cell[   32296] = 32'h0867f84d;
    ram_cell[   32297] = 32'h2404771e;
    ram_cell[   32298] = 32'h459ff3f3;
    ram_cell[   32299] = 32'h1b253e17;
    ram_cell[   32300] = 32'hd62ac762;
    ram_cell[   32301] = 32'hbdc2f4cc;
    ram_cell[   32302] = 32'h48505365;
    ram_cell[   32303] = 32'h0d797ce4;
    ram_cell[   32304] = 32'he3bb0739;
    ram_cell[   32305] = 32'h0f83c732;
    ram_cell[   32306] = 32'hf6e821f0;
    ram_cell[   32307] = 32'hb9c90972;
    ram_cell[   32308] = 32'h3eed0d93;
    ram_cell[   32309] = 32'he5a4a4da;
    ram_cell[   32310] = 32'h1ece871b;
    ram_cell[   32311] = 32'he242282a;
    ram_cell[   32312] = 32'h64bdb66c;
    ram_cell[   32313] = 32'h2e0f6cd0;
    ram_cell[   32314] = 32'h54bf567a;
    ram_cell[   32315] = 32'hcaa0d1fe;
    ram_cell[   32316] = 32'hf2137f39;
    ram_cell[   32317] = 32'h8f19e016;
    ram_cell[   32318] = 32'h47522844;
    ram_cell[   32319] = 32'hb8784a91;
    ram_cell[   32320] = 32'hbbad08c4;
    ram_cell[   32321] = 32'h37cca59d;
    ram_cell[   32322] = 32'hf8661eb9;
    ram_cell[   32323] = 32'he7f2a888;
    ram_cell[   32324] = 32'h4ccac4e1;
    ram_cell[   32325] = 32'h54e3b540;
    ram_cell[   32326] = 32'hbba9ead4;
    ram_cell[   32327] = 32'hef4bf8ae;
    ram_cell[   32328] = 32'h291e05f2;
    ram_cell[   32329] = 32'hd1ba06d0;
    ram_cell[   32330] = 32'h8f70a967;
    ram_cell[   32331] = 32'h08f5e546;
    ram_cell[   32332] = 32'h3b4a50ca;
    ram_cell[   32333] = 32'hf35a8d2f;
    ram_cell[   32334] = 32'h08b2e6e1;
    ram_cell[   32335] = 32'h9c2c26d9;
    ram_cell[   32336] = 32'hb4b5e0d0;
    ram_cell[   32337] = 32'h2bbc2304;
    ram_cell[   32338] = 32'h37f5819f;
    ram_cell[   32339] = 32'h99e33ce8;
    ram_cell[   32340] = 32'hdb7fda45;
    ram_cell[   32341] = 32'hcf24b759;
    ram_cell[   32342] = 32'hfb1ca8a1;
    ram_cell[   32343] = 32'h197130e0;
    ram_cell[   32344] = 32'h9189a452;
    ram_cell[   32345] = 32'h6db5bf59;
    ram_cell[   32346] = 32'h56af8976;
    ram_cell[   32347] = 32'h1e80cb82;
    ram_cell[   32348] = 32'h19d0081d;
    ram_cell[   32349] = 32'h33b2f4b2;
    ram_cell[   32350] = 32'hb94edd74;
    ram_cell[   32351] = 32'hbf1bacf4;
    ram_cell[   32352] = 32'h28330819;
    ram_cell[   32353] = 32'hd67f5f7f;
    ram_cell[   32354] = 32'hb355bcd0;
    ram_cell[   32355] = 32'hdca9a65f;
    ram_cell[   32356] = 32'h3be76f78;
    ram_cell[   32357] = 32'hbcf93f7a;
    ram_cell[   32358] = 32'hc51e48be;
    ram_cell[   32359] = 32'hb0a661ba;
    ram_cell[   32360] = 32'h023b8467;
    ram_cell[   32361] = 32'hf3f6101d;
    ram_cell[   32362] = 32'h8fab76b4;
    ram_cell[   32363] = 32'h821c885a;
    ram_cell[   32364] = 32'h2f8d9c8d;
    ram_cell[   32365] = 32'h9bf97414;
    ram_cell[   32366] = 32'h6855f775;
    ram_cell[   32367] = 32'h826eef09;
    ram_cell[   32368] = 32'hd6517205;
    ram_cell[   32369] = 32'h02ffd4d6;
    ram_cell[   32370] = 32'h921ed5b6;
    ram_cell[   32371] = 32'hf25085ba;
    ram_cell[   32372] = 32'hb4348e67;
    ram_cell[   32373] = 32'hec9f6bbf;
    ram_cell[   32374] = 32'h4204aa31;
    ram_cell[   32375] = 32'h830e3c4b;
    ram_cell[   32376] = 32'h60faddba;
    ram_cell[   32377] = 32'he1660c9d;
    ram_cell[   32378] = 32'hb3bef642;
    ram_cell[   32379] = 32'h65402ab1;
    ram_cell[   32380] = 32'h0a120e10;
    ram_cell[   32381] = 32'h8f31201b;
    ram_cell[   32382] = 32'h333865c5;
    ram_cell[   32383] = 32'h652c375b;
    ram_cell[   32384] = 32'hf56d48f3;
    ram_cell[   32385] = 32'h62d94294;
    ram_cell[   32386] = 32'hc3bf0253;
    ram_cell[   32387] = 32'h89ca3632;
    ram_cell[   32388] = 32'h721ad9d4;
    ram_cell[   32389] = 32'h914c002c;
    ram_cell[   32390] = 32'h27582e81;
    ram_cell[   32391] = 32'hee738145;
    ram_cell[   32392] = 32'hdd0b750c;
    ram_cell[   32393] = 32'h17ef9588;
    ram_cell[   32394] = 32'h352007f9;
    ram_cell[   32395] = 32'h07b0fe33;
    ram_cell[   32396] = 32'h01ddbc70;
    ram_cell[   32397] = 32'hdf8d093b;
    ram_cell[   32398] = 32'hb44b6b58;
    ram_cell[   32399] = 32'hec6a246e;
    ram_cell[   32400] = 32'h819950b7;
    ram_cell[   32401] = 32'he25fb28b;
    ram_cell[   32402] = 32'hfb23f8bd;
    ram_cell[   32403] = 32'h96d61a0c;
    ram_cell[   32404] = 32'hc8f2946f;
    ram_cell[   32405] = 32'h88cdd1b9;
    ram_cell[   32406] = 32'h880f7b88;
    ram_cell[   32407] = 32'h3322e4cf;
    ram_cell[   32408] = 32'h8bb1dcd8;
    ram_cell[   32409] = 32'h1912595c;
    ram_cell[   32410] = 32'h0077cdec;
    ram_cell[   32411] = 32'h24ef04b3;
    ram_cell[   32412] = 32'h65870a51;
    ram_cell[   32413] = 32'hdc8080d3;
    ram_cell[   32414] = 32'hed7473c7;
    ram_cell[   32415] = 32'h4c871aa8;
    ram_cell[   32416] = 32'hfd25d5f0;
    ram_cell[   32417] = 32'h4380706a;
    ram_cell[   32418] = 32'h5833d580;
    ram_cell[   32419] = 32'h76b1a0f0;
    ram_cell[   32420] = 32'hc36eac66;
    ram_cell[   32421] = 32'h0bbbbc07;
    ram_cell[   32422] = 32'h1bb3f9d8;
    ram_cell[   32423] = 32'h533dfc87;
    ram_cell[   32424] = 32'h58ae540d;
    ram_cell[   32425] = 32'hea375e06;
    ram_cell[   32426] = 32'he84933f1;
    ram_cell[   32427] = 32'hbbb56dc0;
    ram_cell[   32428] = 32'h5aa2858b;
    ram_cell[   32429] = 32'hf58dbc8e;
    ram_cell[   32430] = 32'hf26d2848;
    ram_cell[   32431] = 32'h7b2a08e7;
    ram_cell[   32432] = 32'h68e042a4;
    ram_cell[   32433] = 32'h5f3bea10;
    ram_cell[   32434] = 32'h3333b1e6;
    ram_cell[   32435] = 32'h64bb8a35;
    ram_cell[   32436] = 32'hdabd1522;
    ram_cell[   32437] = 32'hedf998fd;
    ram_cell[   32438] = 32'hfe1e08ae;
    ram_cell[   32439] = 32'he8bd814f;
    ram_cell[   32440] = 32'h98f15d16;
    ram_cell[   32441] = 32'h0973fe7a;
    ram_cell[   32442] = 32'h4229343b;
    ram_cell[   32443] = 32'hbd1569fa;
    ram_cell[   32444] = 32'h17789f27;
    ram_cell[   32445] = 32'haeeb70e4;
    ram_cell[   32446] = 32'h89ed91a8;
    ram_cell[   32447] = 32'hac73b089;
    ram_cell[   32448] = 32'h3765968b;
    ram_cell[   32449] = 32'hd301e228;
    ram_cell[   32450] = 32'h96e18423;
    ram_cell[   32451] = 32'h64edaa0e;
    ram_cell[   32452] = 32'hbdb30941;
    ram_cell[   32453] = 32'h2689b3d3;
    ram_cell[   32454] = 32'h1ed18c7e;
    ram_cell[   32455] = 32'hb2ba1aa5;
    ram_cell[   32456] = 32'hdf950525;
    ram_cell[   32457] = 32'h9db0e479;
    ram_cell[   32458] = 32'h0eabc14f;
    ram_cell[   32459] = 32'h7e43800a;
    ram_cell[   32460] = 32'h8ac4a809;
    ram_cell[   32461] = 32'hb15bbd38;
    ram_cell[   32462] = 32'hefd33d58;
    ram_cell[   32463] = 32'h366195a7;
    ram_cell[   32464] = 32'h740842f2;
    ram_cell[   32465] = 32'hc5322abb;
    ram_cell[   32466] = 32'h6a736c3c;
    ram_cell[   32467] = 32'h76700c9f;
    ram_cell[   32468] = 32'haa475158;
    ram_cell[   32469] = 32'h45e775f5;
    ram_cell[   32470] = 32'h992e8426;
    ram_cell[   32471] = 32'h1208d314;
    ram_cell[   32472] = 32'h36c8b0d2;
    ram_cell[   32473] = 32'h9cc38c97;
    ram_cell[   32474] = 32'h760163dd;
    ram_cell[   32475] = 32'hfc8371b4;
    ram_cell[   32476] = 32'he515fe69;
    ram_cell[   32477] = 32'h2ca31dcd;
    ram_cell[   32478] = 32'hef0bdc0a;
    ram_cell[   32479] = 32'he6591d9c;
    ram_cell[   32480] = 32'h6d4656dd;
    ram_cell[   32481] = 32'hf9f682c6;
    ram_cell[   32482] = 32'h2421b028;
    ram_cell[   32483] = 32'h08b76622;
    ram_cell[   32484] = 32'h22d78f06;
    ram_cell[   32485] = 32'h50242888;
    ram_cell[   32486] = 32'hbf99899f;
    ram_cell[   32487] = 32'h0d727c33;
    ram_cell[   32488] = 32'hefd742da;
    ram_cell[   32489] = 32'hc81c028a;
    ram_cell[   32490] = 32'h4d1aee45;
    ram_cell[   32491] = 32'he3c3523e;
    ram_cell[   32492] = 32'h864450ed;
    ram_cell[   32493] = 32'h119b0df3;
    ram_cell[   32494] = 32'h5fe9d03a;
    ram_cell[   32495] = 32'hf34a0a05;
    ram_cell[   32496] = 32'he99cc385;
    ram_cell[   32497] = 32'h0613fb07;
    ram_cell[   32498] = 32'h010826ed;
    ram_cell[   32499] = 32'h6c382820;
    ram_cell[   32500] = 32'hcb876e7c;
    ram_cell[   32501] = 32'h186334be;
    ram_cell[   32502] = 32'h2da01c4d;
    ram_cell[   32503] = 32'h9fa586bf;
    ram_cell[   32504] = 32'hc4003f60;
    ram_cell[   32505] = 32'ha858a86a;
    ram_cell[   32506] = 32'h846dac46;
    ram_cell[   32507] = 32'h09fd0816;
    ram_cell[   32508] = 32'hc1e87dc4;
    ram_cell[   32509] = 32'h75fc8a62;
    ram_cell[   32510] = 32'he4b878fc;
    ram_cell[   32511] = 32'h0f2602e7;
    ram_cell[   32512] = 32'hfe0b93b1;
    ram_cell[   32513] = 32'h8d8adf31;
    ram_cell[   32514] = 32'h1a6c9655;
    ram_cell[   32515] = 32'h3917cf2e;
    ram_cell[   32516] = 32'he4829c29;
    ram_cell[   32517] = 32'h68110826;
    ram_cell[   32518] = 32'hc4ffcb26;
    ram_cell[   32519] = 32'h5e6a8640;
    ram_cell[   32520] = 32'hfbc54305;
    ram_cell[   32521] = 32'hae8f952f;
    ram_cell[   32522] = 32'hb2ec86e1;
    ram_cell[   32523] = 32'hb2ae668a;
    ram_cell[   32524] = 32'hfa7ff8a5;
    ram_cell[   32525] = 32'h92c68d4a;
    ram_cell[   32526] = 32'h12a89e5e;
    ram_cell[   32527] = 32'h46a5adb6;
    ram_cell[   32528] = 32'he48be78e;
    ram_cell[   32529] = 32'hccfbbd91;
    ram_cell[   32530] = 32'ha2234d43;
    ram_cell[   32531] = 32'h4cb8009e;
    ram_cell[   32532] = 32'hac523a89;
    ram_cell[   32533] = 32'h43e2dbbd;
    ram_cell[   32534] = 32'he1b89428;
    ram_cell[   32535] = 32'hecf76a37;
    ram_cell[   32536] = 32'h7c67e347;
    ram_cell[   32537] = 32'ha509ecc1;
    ram_cell[   32538] = 32'h1e1ddffb;
    ram_cell[   32539] = 32'h0c268ec2;
    ram_cell[   32540] = 32'h4145ed4b;
    ram_cell[   32541] = 32'h5451b47a;
    ram_cell[   32542] = 32'h95c0e3fa;
    ram_cell[   32543] = 32'h099cb684;
    ram_cell[   32544] = 32'hd97f2e5d;
    ram_cell[   32545] = 32'hc940570d;
    ram_cell[   32546] = 32'heacf0f06;
    ram_cell[   32547] = 32'h7dd07d65;
    ram_cell[   32548] = 32'h6ad6d0ec;
    ram_cell[   32549] = 32'h6c0d8817;
    ram_cell[   32550] = 32'h7c074541;
    ram_cell[   32551] = 32'had98c9ec;
    ram_cell[   32552] = 32'h7226f445;
    ram_cell[   32553] = 32'h254b7679;
    ram_cell[   32554] = 32'h3c701375;
    ram_cell[   32555] = 32'heffa7a72;
    ram_cell[   32556] = 32'he5f28e83;
    ram_cell[   32557] = 32'h6430c9e7;
    ram_cell[   32558] = 32'h933189bd;
    ram_cell[   32559] = 32'h3e937d54;
    ram_cell[   32560] = 32'he7319c90;
    ram_cell[   32561] = 32'hd4eaa0b6;
    ram_cell[   32562] = 32'h5f8e1b97;
    ram_cell[   32563] = 32'h04a212d0;
    ram_cell[   32564] = 32'h441aca76;
    ram_cell[   32565] = 32'hb1feb8ca;
    ram_cell[   32566] = 32'h3f59b561;
    ram_cell[   32567] = 32'h400177b4;
    ram_cell[   32568] = 32'h2ebecedd;
    ram_cell[   32569] = 32'h81516eb8;
    ram_cell[   32570] = 32'hb7e97513;
    ram_cell[   32571] = 32'h5285731d;
    ram_cell[   32572] = 32'h48c0394b;
    ram_cell[   32573] = 32'h5652c003;
    ram_cell[   32574] = 32'he229b0b4;
    ram_cell[   32575] = 32'hcf5017a9;
    ram_cell[   32576] = 32'haab07006;
    ram_cell[   32577] = 32'hc2e82865;
    ram_cell[   32578] = 32'h9f1ce575;
    ram_cell[   32579] = 32'hbf77b1ac;
    ram_cell[   32580] = 32'h679afb92;
    ram_cell[   32581] = 32'h9508a9c6;
    ram_cell[   32582] = 32'hacb6c2c3;
    ram_cell[   32583] = 32'h8964e96f;
    ram_cell[   32584] = 32'h26cd7aeb;
    ram_cell[   32585] = 32'h9823cb7d;
    ram_cell[   32586] = 32'h1433141b;
    ram_cell[   32587] = 32'h71d236d9;
    ram_cell[   32588] = 32'h344195e7;
    ram_cell[   32589] = 32'h4f0dff92;
    ram_cell[   32590] = 32'h575b9cb6;
    ram_cell[   32591] = 32'hbd72b92b;
    ram_cell[   32592] = 32'h603005f4;
    ram_cell[   32593] = 32'h1ede98bf;
    ram_cell[   32594] = 32'h1bfe13d2;
    ram_cell[   32595] = 32'hd812b8c6;
    ram_cell[   32596] = 32'hd0df8ab7;
    ram_cell[   32597] = 32'h636a1851;
    ram_cell[   32598] = 32'h5c0a9498;
    ram_cell[   32599] = 32'h725b6691;
    ram_cell[   32600] = 32'h62dbb62a;
    ram_cell[   32601] = 32'h63d28a19;
    ram_cell[   32602] = 32'h5d1ef516;
    ram_cell[   32603] = 32'h901a1e31;
    ram_cell[   32604] = 32'hd2479d24;
    ram_cell[   32605] = 32'h3b531a20;
    ram_cell[   32606] = 32'h86e344f3;
    ram_cell[   32607] = 32'h5805c8c4;
    ram_cell[   32608] = 32'h71617d99;
    ram_cell[   32609] = 32'h17b668df;
    ram_cell[   32610] = 32'h145ff32c;
    ram_cell[   32611] = 32'h9e15bb98;
    ram_cell[   32612] = 32'hf1d9788f;
    ram_cell[   32613] = 32'hece47dd8;
    ram_cell[   32614] = 32'h51eb9ea2;
    ram_cell[   32615] = 32'h66980a78;
    ram_cell[   32616] = 32'h48caa218;
    ram_cell[   32617] = 32'h28a8cbd1;
    ram_cell[   32618] = 32'hbba895b3;
    ram_cell[   32619] = 32'h6de15348;
    ram_cell[   32620] = 32'h43b65a6c;
    ram_cell[   32621] = 32'hcbcadaa9;
    ram_cell[   32622] = 32'h913909ad;
    ram_cell[   32623] = 32'h92b0f3d9;
    ram_cell[   32624] = 32'h3510a6e0;
    ram_cell[   32625] = 32'hc6012232;
    ram_cell[   32626] = 32'h61a60c76;
    ram_cell[   32627] = 32'h2a09c660;
    ram_cell[   32628] = 32'h2ad21743;
    ram_cell[   32629] = 32'heb5d6842;
    ram_cell[   32630] = 32'h563e946e;
    ram_cell[   32631] = 32'h28401b10;
    ram_cell[   32632] = 32'hcded2135;
    ram_cell[   32633] = 32'h90a1ae9e;
    ram_cell[   32634] = 32'h7465ad2d;
    ram_cell[   32635] = 32'h2624165b;
    ram_cell[   32636] = 32'hea5d0812;
    ram_cell[   32637] = 32'ha996d99c;
    ram_cell[   32638] = 32'h119a5e6f;
    ram_cell[   32639] = 32'h6ab24b0f;
    ram_cell[   32640] = 32'hed090d16;
    ram_cell[   32641] = 32'hb06e4d30;
    ram_cell[   32642] = 32'h3438b341;
    ram_cell[   32643] = 32'h8eccf68a;
    ram_cell[   32644] = 32'haa30a705;
    ram_cell[   32645] = 32'hc9d3a247;
    ram_cell[   32646] = 32'he2653e71;
    ram_cell[   32647] = 32'h6f0418eb;
    ram_cell[   32648] = 32'hf573b16d;
    ram_cell[   32649] = 32'hec092d3c;
    ram_cell[   32650] = 32'hf387a766;
    ram_cell[   32651] = 32'h7205d61c;
    ram_cell[   32652] = 32'hf6f821e6;
    ram_cell[   32653] = 32'hcb9e495e;
    ram_cell[   32654] = 32'hf414d571;
    ram_cell[   32655] = 32'h24324fef;
    ram_cell[   32656] = 32'h451200f0;
    ram_cell[   32657] = 32'h2251167a;
    ram_cell[   32658] = 32'hbe8eb749;
    ram_cell[   32659] = 32'hff09c218;
    ram_cell[   32660] = 32'h368f6471;
    ram_cell[   32661] = 32'h8ed3f313;
    ram_cell[   32662] = 32'hbcbef52f;
    ram_cell[   32663] = 32'h71e1236b;
    ram_cell[   32664] = 32'h899a08cd;
    ram_cell[   32665] = 32'h10ac9573;
    ram_cell[   32666] = 32'h718e2174;
    ram_cell[   32667] = 32'h91720d74;
    ram_cell[   32668] = 32'h93a5462f;
    ram_cell[   32669] = 32'he14a7e6e;
    ram_cell[   32670] = 32'he4a399de;
    ram_cell[   32671] = 32'ha9d27428;
    ram_cell[   32672] = 32'h97c058ba;
    ram_cell[   32673] = 32'hdb8d2bc2;
    ram_cell[   32674] = 32'h4f823856;
    ram_cell[   32675] = 32'hf73c2dac;
    ram_cell[   32676] = 32'hc64f57ca;
    ram_cell[   32677] = 32'hd8005fbc;
    ram_cell[   32678] = 32'h52dc4707;
    ram_cell[   32679] = 32'hf1d24759;
    ram_cell[   32680] = 32'h1012c5a8;
    ram_cell[   32681] = 32'h3df0ccdd;
    ram_cell[   32682] = 32'h542853e7;
    ram_cell[   32683] = 32'h29419622;
    ram_cell[   32684] = 32'h109be840;
    ram_cell[   32685] = 32'h18f43053;
    ram_cell[   32686] = 32'he8de4e2a;
    ram_cell[   32687] = 32'h616dd71b;
    ram_cell[   32688] = 32'h25b2f263;
    ram_cell[   32689] = 32'hc225c866;
    ram_cell[   32690] = 32'hdbea9cbe;
    ram_cell[   32691] = 32'h6318a257;
    ram_cell[   32692] = 32'he69c54cd;
    ram_cell[   32693] = 32'h014aaeaf;
    ram_cell[   32694] = 32'h6fdcf479;
    ram_cell[   32695] = 32'h8555ebc7;
    ram_cell[   32696] = 32'h8fed0cea;
    ram_cell[   32697] = 32'hb5890aee;
    ram_cell[   32698] = 32'ha9adc236;
    ram_cell[   32699] = 32'h8bb2e79a;
    ram_cell[   32700] = 32'h92c14d46;
    ram_cell[   32701] = 32'h16398f7f;
    ram_cell[   32702] = 32'hd25690cf;
    ram_cell[   32703] = 32'h29c074fd;
    ram_cell[   32704] = 32'h1fbc0f84;
    ram_cell[   32705] = 32'haa67c345;
    ram_cell[   32706] = 32'hf104303c;
    ram_cell[   32707] = 32'h548cdfb0;
    ram_cell[   32708] = 32'hdb56bb61;
    ram_cell[   32709] = 32'hd5f859b1;
    ram_cell[   32710] = 32'h40c7b57d;
    ram_cell[   32711] = 32'h805abdec;
    ram_cell[   32712] = 32'hf2827a5d;
    ram_cell[   32713] = 32'h140c6000;
    ram_cell[   32714] = 32'h85baf2f8;
    ram_cell[   32715] = 32'hefa31423;
    ram_cell[   32716] = 32'he9894bdd;
    ram_cell[   32717] = 32'h01248be4;
    ram_cell[   32718] = 32'h2cc28469;
    ram_cell[   32719] = 32'hbe0f564a;
    ram_cell[   32720] = 32'hb9b5399d;
    ram_cell[   32721] = 32'hff8218b0;
    ram_cell[   32722] = 32'h76b151c3;
    ram_cell[   32723] = 32'hde6f413f;
    ram_cell[   32724] = 32'hd6bb1097;
    ram_cell[   32725] = 32'h61cf0d32;
    ram_cell[   32726] = 32'h45b72194;
    ram_cell[   32727] = 32'h958e089d;
    ram_cell[   32728] = 32'hfa50c6bd;
    ram_cell[   32729] = 32'h12c61e0c;
    ram_cell[   32730] = 32'h9690de9f;
    ram_cell[   32731] = 32'h22ee20d8;
    ram_cell[   32732] = 32'h5928f1e9;
    ram_cell[   32733] = 32'h411976ed;
    ram_cell[   32734] = 32'hc6bb65ca;
    ram_cell[   32735] = 32'hb8b682e1;
    ram_cell[   32736] = 32'h9709ebf2;
    ram_cell[   32737] = 32'hd3223eb1;
    ram_cell[   32738] = 32'h2a9ed127;
    ram_cell[   32739] = 32'h10cbcbba;
    ram_cell[   32740] = 32'h11bdbab4;
    ram_cell[   32741] = 32'h9e8175ad;
    ram_cell[   32742] = 32'h6657dc62;
    ram_cell[   32743] = 32'h8e6c3ff8;
    ram_cell[   32744] = 32'h3e45a2a1;
    ram_cell[   32745] = 32'hd91a268c;
    ram_cell[   32746] = 32'hc06cd281;
    ram_cell[   32747] = 32'hcd952ef0;
    ram_cell[   32748] = 32'h0d0e18e0;
    ram_cell[   32749] = 32'h306f0c66;
    ram_cell[   32750] = 32'h223d1281;
    ram_cell[   32751] = 32'he1063fdd;
    ram_cell[   32752] = 32'h71a3946d;
    ram_cell[   32753] = 32'hbc24ab2c;
    ram_cell[   32754] = 32'h1f5713c6;
    ram_cell[   32755] = 32'hf0e3ea8d;
    ram_cell[   32756] = 32'h2e4a9252;
    ram_cell[   32757] = 32'hf4912ece;
    ram_cell[   32758] = 32'h99a8c1ee;
    ram_cell[   32759] = 32'hb0348461;
    ram_cell[   32760] = 32'he6f5bd3c;
    ram_cell[   32761] = 32'h21b3bc87;
    ram_cell[   32762] = 32'h7c428e26;
    ram_cell[   32763] = 32'ha02c3048;
    ram_cell[   32764] = 32'h0b2e8034;
    ram_cell[   32765] = 32'hc43fe62f;
    ram_cell[   32766] = 32'h3722b0ea;
    ram_cell[   32767] = 32'h9fe5ba9b;
    // src matrix B
    ram_cell[   32768] = 32'h8f0c74c9;
    ram_cell[   32769] = 32'hc8c8e370;
    ram_cell[   32770] = 32'h014b08fd;
    ram_cell[   32771] = 32'h3f92e0f9;
    ram_cell[   32772] = 32'h43e011f1;
    ram_cell[   32773] = 32'h60191023;
    ram_cell[   32774] = 32'h61e9bd65;
    ram_cell[   32775] = 32'hf122e293;
    ram_cell[   32776] = 32'h8ebdecc7;
    ram_cell[   32777] = 32'h77b65f68;
    ram_cell[   32778] = 32'h7bc688d0;
    ram_cell[   32779] = 32'h905f4447;
    ram_cell[   32780] = 32'hbab42b32;
    ram_cell[   32781] = 32'h5f0b905f;
    ram_cell[   32782] = 32'hfa43ce8b;
    ram_cell[   32783] = 32'hc4474fd0;
    ram_cell[   32784] = 32'hef83b2d0;
    ram_cell[   32785] = 32'h5966eb8d;
    ram_cell[   32786] = 32'h82945585;
    ram_cell[   32787] = 32'hda104384;
    ram_cell[   32788] = 32'h2e4c3679;
    ram_cell[   32789] = 32'h37df0806;
    ram_cell[   32790] = 32'h877ef048;
    ram_cell[   32791] = 32'h9dcbcbf1;
    ram_cell[   32792] = 32'h26dddd08;
    ram_cell[   32793] = 32'h6f1a5086;
    ram_cell[   32794] = 32'h57aa3680;
    ram_cell[   32795] = 32'hfca7d3e6;
    ram_cell[   32796] = 32'h547972a3;
    ram_cell[   32797] = 32'h5f657b24;
    ram_cell[   32798] = 32'hea4e7ca6;
    ram_cell[   32799] = 32'h5a03443a;
    ram_cell[   32800] = 32'h7f26c0fa;
    ram_cell[   32801] = 32'h614864bd;
    ram_cell[   32802] = 32'hf8f0fe88;
    ram_cell[   32803] = 32'h00be0606;
    ram_cell[   32804] = 32'h5dbe8c4d;
    ram_cell[   32805] = 32'h1336ec29;
    ram_cell[   32806] = 32'h20103af0;
    ram_cell[   32807] = 32'h15ad8e06;
    ram_cell[   32808] = 32'h8fb770d4;
    ram_cell[   32809] = 32'h1f42fd97;
    ram_cell[   32810] = 32'h6a24495e;
    ram_cell[   32811] = 32'h618e6846;
    ram_cell[   32812] = 32'hf33600e5;
    ram_cell[   32813] = 32'h19e880bf;
    ram_cell[   32814] = 32'h47ffa0af;
    ram_cell[   32815] = 32'h29a07618;
    ram_cell[   32816] = 32'hfda57bcf;
    ram_cell[   32817] = 32'hdd51fed9;
    ram_cell[   32818] = 32'h9e81b076;
    ram_cell[   32819] = 32'h01376844;
    ram_cell[   32820] = 32'h6f98ff5a;
    ram_cell[   32821] = 32'h1d8f091f;
    ram_cell[   32822] = 32'h6ee89d7a;
    ram_cell[   32823] = 32'h84d4e9f7;
    ram_cell[   32824] = 32'h7a5f5164;
    ram_cell[   32825] = 32'hf763c651;
    ram_cell[   32826] = 32'hb585cec4;
    ram_cell[   32827] = 32'h4c8385d3;
    ram_cell[   32828] = 32'h5951360b;
    ram_cell[   32829] = 32'h793e83e1;
    ram_cell[   32830] = 32'h0dd5e2cd;
    ram_cell[   32831] = 32'h729a2caa;
    ram_cell[   32832] = 32'hbc715983;
    ram_cell[   32833] = 32'h0f2ded96;
    ram_cell[   32834] = 32'hc91fd060;
    ram_cell[   32835] = 32'h66da5502;
    ram_cell[   32836] = 32'hf11898fb;
    ram_cell[   32837] = 32'hae93b3bb;
    ram_cell[   32838] = 32'h052b62b7;
    ram_cell[   32839] = 32'h6d995b28;
    ram_cell[   32840] = 32'hdd017f6d;
    ram_cell[   32841] = 32'h5cfbc185;
    ram_cell[   32842] = 32'haad4bc49;
    ram_cell[   32843] = 32'hf5e9f89d;
    ram_cell[   32844] = 32'h03cacd2d;
    ram_cell[   32845] = 32'h9fe976a8;
    ram_cell[   32846] = 32'hd803f81a;
    ram_cell[   32847] = 32'h41e1ff6b;
    ram_cell[   32848] = 32'hf6dd2257;
    ram_cell[   32849] = 32'hbc8d1947;
    ram_cell[   32850] = 32'h4862b91a;
    ram_cell[   32851] = 32'h4886d471;
    ram_cell[   32852] = 32'h02463292;
    ram_cell[   32853] = 32'hc75470b8;
    ram_cell[   32854] = 32'hcff40652;
    ram_cell[   32855] = 32'h7e53da2a;
    ram_cell[   32856] = 32'h193524fb;
    ram_cell[   32857] = 32'h29cf171a;
    ram_cell[   32858] = 32'hbb122e82;
    ram_cell[   32859] = 32'hd26b3e0a;
    ram_cell[   32860] = 32'h26ec3b4f;
    ram_cell[   32861] = 32'h27102857;
    ram_cell[   32862] = 32'h215cc166;
    ram_cell[   32863] = 32'he12d89a1;
    ram_cell[   32864] = 32'h257b3f36;
    ram_cell[   32865] = 32'h1bee6580;
    ram_cell[   32866] = 32'h4a1a8f69;
    ram_cell[   32867] = 32'hdf94267c;
    ram_cell[   32868] = 32'hd78f2c4a;
    ram_cell[   32869] = 32'ha7e583ea;
    ram_cell[   32870] = 32'h084abdcc;
    ram_cell[   32871] = 32'h624f1e9a;
    ram_cell[   32872] = 32'hce5988e7;
    ram_cell[   32873] = 32'h65ed1ae5;
    ram_cell[   32874] = 32'h4144825a;
    ram_cell[   32875] = 32'hcd2097e6;
    ram_cell[   32876] = 32'heda0b487;
    ram_cell[   32877] = 32'h8c7537bd;
    ram_cell[   32878] = 32'h37855da1;
    ram_cell[   32879] = 32'haaa5214e;
    ram_cell[   32880] = 32'h4b5591a0;
    ram_cell[   32881] = 32'h52e41224;
    ram_cell[   32882] = 32'h902a7b93;
    ram_cell[   32883] = 32'h82bff0bf;
    ram_cell[   32884] = 32'h85589f2e;
    ram_cell[   32885] = 32'h2241bea5;
    ram_cell[   32886] = 32'hdbf4ca8d;
    ram_cell[   32887] = 32'h2b474a20;
    ram_cell[   32888] = 32'he3c06fb9;
    ram_cell[   32889] = 32'h58b43f61;
    ram_cell[   32890] = 32'hde5b0e26;
    ram_cell[   32891] = 32'hdf4852fc;
    ram_cell[   32892] = 32'hc88c548b;
    ram_cell[   32893] = 32'h45340543;
    ram_cell[   32894] = 32'h7e233744;
    ram_cell[   32895] = 32'h953f8c12;
    ram_cell[   32896] = 32'h4be69369;
    ram_cell[   32897] = 32'h51880402;
    ram_cell[   32898] = 32'h885679b7;
    ram_cell[   32899] = 32'h81bd993b;
    ram_cell[   32900] = 32'hd0e6b6cb;
    ram_cell[   32901] = 32'he9f463b9;
    ram_cell[   32902] = 32'ha2aec0d2;
    ram_cell[   32903] = 32'h1e1bb59d;
    ram_cell[   32904] = 32'h0a74fb49;
    ram_cell[   32905] = 32'hb1adc550;
    ram_cell[   32906] = 32'ha8eb5de1;
    ram_cell[   32907] = 32'hd2d1320c;
    ram_cell[   32908] = 32'h5f4d29dc;
    ram_cell[   32909] = 32'h5ba008d0;
    ram_cell[   32910] = 32'h5d11d711;
    ram_cell[   32911] = 32'hf7f914b7;
    ram_cell[   32912] = 32'h3cc51cb3;
    ram_cell[   32913] = 32'h63faf095;
    ram_cell[   32914] = 32'h59a9f265;
    ram_cell[   32915] = 32'h0e147fd9;
    ram_cell[   32916] = 32'hb112eba9;
    ram_cell[   32917] = 32'hee295a6b;
    ram_cell[   32918] = 32'hf8da3408;
    ram_cell[   32919] = 32'h8449462c;
    ram_cell[   32920] = 32'h9c9fff4e;
    ram_cell[   32921] = 32'hcaf62e57;
    ram_cell[   32922] = 32'hf1d4f715;
    ram_cell[   32923] = 32'h25d346de;
    ram_cell[   32924] = 32'h692ed40e;
    ram_cell[   32925] = 32'h5360e6cd;
    ram_cell[   32926] = 32'h8ce0bc90;
    ram_cell[   32927] = 32'hbbc60c9e;
    ram_cell[   32928] = 32'hde836885;
    ram_cell[   32929] = 32'h4c7612f2;
    ram_cell[   32930] = 32'h3e0b934c;
    ram_cell[   32931] = 32'hd034d71a;
    ram_cell[   32932] = 32'h2a6d2ffe;
    ram_cell[   32933] = 32'hbcc16902;
    ram_cell[   32934] = 32'h08daa066;
    ram_cell[   32935] = 32'hae6f7b1a;
    ram_cell[   32936] = 32'hea56d1eb;
    ram_cell[   32937] = 32'h9c314437;
    ram_cell[   32938] = 32'h3a2ad4dd;
    ram_cell[   32939] = 32'h7597e563;
    ram_cell[   32940] = 32'h78e7674c;
    ram_cell[   32941] = 32'h5f4e218d;
    ram_cell[   32942] = 32'h3963048e;
    ram_cell[   32943] = 32'hc804d8a5;
    ram_cell[   32944] = 32'h81945a2b;
    ram_cell[   32945] = 32'h9cdb72b8;
    ram_cell[   32946] = 32'hc583b168;
    ram_cell[   32947] = 32'h05d96b4a;
    ram_cell[   32948] = 32'h724fb601;
    ram_cell[   32949] = 32'ha269efd2;
    ram_cell[   32950] = 32'h68b705bf;
    ram_cell[   32951] = 32'h966e180e;
    ram_cell[   32952] = 32'h4781babf;
    ram_cell[   32953] = 32'h9755959a;
    ram_cell[   32954] = 32'h8d9ba4a4;
    ram_cell[   32955] = 32'h46412d31;
    ram_cell[   32956] = 32'h026fd0df;
    ram_cell[   32957] = 32'ha5678421;
    ram_cell[   32958] = 32'h572d2557;
    ram_cell[   32959] = 32'h4b7ea094;
    ram_cell[   32960] = 32'h4bc53c41;
    ram_cell[   32961] = 32'h15d20671;
    ram_cell[   32962] = 32'h7bb0c381;
    ram_cell[   32963] = 32'ha76af328;
    ram_cell[   32964] = 32'h6ef66734;
    ram_cell[   32965] = 32'h3cb431d2;
    ram_cell[   32966] = 32'h004d2428;
    ram_cell[   32967] = 32'hdf34c148;
    ram_cell[   32968] = 32'he6264b1f;
    ram_cell[   32969] = 32'h5a66ed0d;
    ram_cell[   32970] = 32'hfcb52a95;
    ram_cell[   32971] = 32'hea6a46d7;
    ram_cell[   32972] = 32'hd561d59a;
    ram_cell[   32973] = 32'h6e8f8001;
    ram_cell[   32974] = 32'hb719bba1;
    ram_cell[   32975] = 32'h90672253;
    ram_cell[   32976] = 32'h2bd332fd;
    ram_cell[   32977] = 32'hc2e7282c;
    ram_cell[   32978] = 32'hc4654d32;
    ram_cell[   32979] = 32'h30213e34;
    ram_cell[   32980] = 32'hcf429b36;
    ram_cell[   32981] = 32'h1202eb7a;
    ram_cell[   32982] = 32'hb304502b;
    ram_cell[   32983] = 32'hc31cc4ae;
    ram_cell[   32984] = 32'h23c09cf3;
    ram_cell[   32985] = 32'ha99c76c1;
    ram_cell[   32986] = 32'hbc2a2948;
    ram_cell[   32987] = 32'hc5d04d97;
    ram_cell[   32988] = 32'hf451c43b;
    ram_cell[   32989] = 32'h27be00b5;
    ram_cell[   32990] = 32'had9b81a2;
    ram_cell[   32991] = 32'h295baf85;
    ram_cell[   32992] = 32'hb8bc12b9;
    ram_cell[   32993] = 32'hcfd073c2;
    ram_cell[   32994] = 32'hc69f4fdd;
    ram_cell[   32995] = 32'h3113870c;
    ram_cell[   32996] = 32'h4ff0e944;
    ram_cell[   32997] = 32'h320cc23c;
    ram_cell[   32998] = 32'h5cf0ecf9;
    ram_cell[   32999] = 32'hd8b5f588;
    ram_cell[   33000] = 32'h2e2588e4;
    ram_cell[   33001] = 32'h6fef6a58;
    ram_cell[   33002] = 32'h75222773;
    ram_cell[   33003] = 32'h61d7fc5a;
    ram_cell[   33004] = 32'hf93d3824;
    ram_cell[   33005] = 32'h6ce4225a;
    ram_cell[   33006] = 32'hd7079c2c;
    ram_cell[   33007] = 32'h78a122f3;
    ram_cell[   33008] = 32'h609e8797;
    ram_cell[   33009] = 32'h627080af;
    ram_cell[   33010] = 32'h913a116d;
    ram_cell[   33011] = 32'h4301b1e6;
    ram_cell[   33012] = 32'haa5d5694;
    ram_cell[   33013] = 32'h4f35f406;
    ram_cell[   33014] = 32'hbbca9d53;
    ram_cell[   33015] = 32'h7f95fb01;
    ram_cell[   33016] = 32'hd54f7072;
    ram_cell[   33017] = 32'h8c634a76;
    ram_cell[   33018] = 32'h852fdc79;
    ram_cell[   33019] = 32'h9e95379f;
    ram_cell[   33020] = 32'h4cd62124;
    ram_cell[   33021] = 32'h7db3158d;
    ram_cell[   33022] = 32'hb9154ccd;
    ram_cell[   33023] = 32'heec50343;
    ram_cell[   33024] = 32'h3beb2dfc;
    ram_cell[   33025] = 32'hfd58aa04;
    ram_cell[   33026] = 32'hee703a5a;
    ram_cell[   33027] = 32'h77249019;
    ram_cell[   33028] = 32'hcad7dd60;
    ram_cell[   33029] = 32'h3b49d66a;
    ram_cell[   33030] = 32'hdb185e4e;
    ram_cell[   33031] = 32'he5d87791;
    ram_cell[   33032] = 32'hd46baeca;
    ram_cell[   33033] = 32'hca1505e5;
    ram_cell[   33034] = 32'he27de08e;
    ram_cell[   33035] = 32'he26a1c57;
    ram_cell[   33036] = 32'h33505cf9;
    ram_cell[   33037] = 32'h81d211eb;
    ram_cell[   33038] = 32'hf9cce781;
    ram_cell[   33039] = 32'h844f63a2;
    ram_cell[   33040] = 32'he18a0e31;
    ram_cell[   33041] = 32'h8b861807;
    ram_cell[   33042] = 32'h4112bfbf;
    ram_cell[   33043] = 32'h54025de2;
    ram_cell[   33044] = 32'h906adb33;
    ram_cell[   33045] = 32'h51f41cfa;
    ram_cell[   33046] = 32'hfb7c8488;
    ram_cell[   33047] = 32'h0c25192b;
    ram_cell[   33048] = 32'h995b8a6c;
    ram_cell[   33049] = 32'hb0c391e5;
    ram_cell[   33050] = 32'h8e02ce83;
    ram_cell[   33051] = 32'h2cece7aa;
    ram_cell[   33052] = 32'h0e4d27b2;
    ram_cell[   33053] = 32'hee697257;
    ram_cell[   33054] = 32'ha4f1c903;
    ram_cell[   33055] = 32'h615c9767;
    ram_cell[   33056] = 32'hff8ffb85;
    ram_cell[   33057] = 32'hb6eb5abc;
    ram_cell[   33058] = 32'hee27fb2c;
    ram_cell[   33059] = 32'h270824a1;
    ram_cell[   33060] = 32'ha733e8a7;
    ram_cell[   33061] = 32'h145a212d;
    ram_cell[   33062] = 32'h71bf687e;
    ram_cell[   33063] = 32'h194c1fa7;
    ram_cell[   33064] = 32'h0b6ba9cf;
    ram_cell[   33065] = 32'h060c5260;
    ram_cell[   33066] = 32'h8b6bf72b;
    ram_cell[   33067] = 32'hd9776102;
    ram_cell[   33068] = 32'h722637ca;
    ram_cell[   33069] = 32'h6d08c85b;
    ram_cell[   33070] = 32'h8277ef1c;
    ram_cell[   33071] = 32'hdc3824d2;
    ram_cell[   33072] = 32'h5dae2863;
    ram_cell[   33073] = 32'he664f443;
    ram_cell[   33074] = 32'h7b1f7d73;
    ram_cell[   33075] = 32'h7d148d49;
    ram_cell[   33076] = 32'h6a4a662a;
    ram_cell[   33077] = 32'hf3c1522c;
    ram_cell[   33078] = 32'h4922c248;
    ram_cell[   33079] = 32'hbd12668f;
    ram_cell[   33080] = 32'h56ff657b;
    ram_cell[   33081] = 32'hc83c3684;
    ram_cell[   33082] = 32'hcc564805;
    ram_cell[   33083] = 32'h1e17d22b;
    ram_cell[   33084] = 32'hc861a8b8;
    ram_cell[   33085] = 32'hdd2b5227;
    ram_cell[   33086] = 32'h80bd410e;
    ram_cell[   33087] = 32'h68778ce8;
    ram_cell[   33088] = 32'h28dfc6ef;
    ram_cell[   33089] = 32'h2632d8ab;
    ram_cell[   33090] = 32'h2d1cb3dc;
    ram_cell[   33091] = 32'h4b6cfc39;
    ram_cell[   33092] = 32'h598a53ee;
    ram_cell[   33093] = 32'hd88fa161;
    ram_cell[   33094] = 32'hd34dc35e;
    ram_cell[   33095] = 32'hd19b884d;
    ram_cell[   33096] = 32'h27574104;
    ram_cell[   33097] = 32'h09e5bf29;
    ram_cell[   33098] = 32'h9eeb1083;
    ram_cell[   33099] = 32'hac268144;
    ram_cell[   33100] = 32'h270a4a58;
    ram_cell[   33101] = 32'hfbc81ade;
    ram_cell[   33102] = 32'h557904fb;
    ram_cell[   33103] = 32'he9169011;
    ram_cell[   33104] = 32'h7eee3dc1;
    ram_cell[   33105] = 32'h68ce3727;
    ram_cell[   33106] = 32'h77179711;
    ram_cell[   33107] = 32'he8e7cc34;
    ram_cell[   33108] = 32'hbf1cd508;
    ram_cell[   33109] = 32'h066cbc80;
    ram_cell[   33110] = 32'h23f1af0c;
    ram_cell[   33111] = 32'h5c3b12c9;
    ram_cell[   33112] = 32'hfd53002e;
    ram_cell[   33113] = 32'had5c1561;
    ram_cell[   33114] = 32'h842b8151;
    ram_cell[   33115] = 32'h6914e5f3;
    ram_cell[   33116] = 32'hf8f84611;
    ram_cell[   33117] = 32'h0994e1ea;
    ram_cell[   33118] = 32'h36e0e005;
    ram_cell[   33119] = 32'h7f4cd43b;
    ram_cell[   33120] = 32'h153ffa13;
    ram_cell[   33121] = 32'ha3d5ff03;
    ram_cell[   33122] = 32'h2fed5d94;
    ram_cell[   33123] = 32'he3bcd55f;
    ram_cell[   33124] = 32'h116a986b;
    ram_cell[   33125] = 32'he9eb22f4;
    ram_cell[   33126] = 32'h5e1e1ca2;
    ram_cell[   33127] = 32'ha90dee6c;
    ram_cell[   33128] = 32'hb8a51f15;
    ram_cell[   33129] = 32'h20f2714a;
    ram_cell[   33130] = 32'h16a62612;
    ram_cell[   33131] = 32'he0fb0f4c;
    ram_cell[   33132] = 32'h706a4404;
    ram_cell[   33133] = 32'hf8689223;
    ram_cell[   33134] = 32'h45b2d0c8;
    ram_cell[   33135] = 32'h4dd989dd;
    ram_cell[   33136] = 32'hc742b2a5;
    ram_cell[   33137] = 32'h2504792c;
    ram_cell[   33138] = 32'h123def3e;
    ram_cell[   33139] = 32'haf397a69;
    ram_cell[   33140] = 32'h5b91c5e9;
    ram_cell[   33141] = 32'he6c017a2;
    ram_cell[   33142] = 32'h46fdb148;
    ram_cell[   33143] = 32'h3eddeac7;
    ram_cell[   33144] = 32'h319e138e;
    ram_cell[   33145] = 32'hd2613ae3;
    ram_cell[   33146] = 32'he2f25d0f;
    ram_cell[   33147] = 32'hacf2d71d;
    ram_cell[   33148] = 32'h271bdba2;
    ram_cell[   33149] = 32'h7498d0ba;
    ram_cell[   33150] = 32'h8613446b;
    ram_cell[   33151] = 32'h7b938b36;
    ram_cell[   33152] = 32'h52b2757d;
    ram_cell[   33153] = 32'h2d21706a;
    ram_cell[   33154] = 32'h8aaf9040;
    ram_cell[   33155] = 32'hde043c58;
    ram_cell[   33156] = 32'h01821a0f;
    ram_cell[   33157] = 32'h3368a8f8;
    ram_cell[   33158] = 32'h3a9d2a23;
    ram_cell[   33159] = 32'h5a8a89d2;
    ram_cell[   33160] = 32'heaee99f4;
    ram_cell[   33161] = 32'h7032a460;
    ram_cell[   33162] = 32'hba16e204;
    ram_cell[   33163] = 32'h3d159074;
    ram_cell[   33164] = 32'h4385a19f;
    ram_cell[   33165] = 32'h33830b40;
    ram_cell[   33166] = 32'h02977519;
    ram_cell[   33167] = 32'hae02b1c9;
    ram_cell[   33168] = 32'h41996cdc;
    ram_cell[   33169] = 32'h1ceefb1c;
    ram_cell[   33170] = 32'h68633699;
    ram_cell[   33171] = 32'h2407b229;
    ram_cell[   33172] = 32'h715ee2e0;
    ram_cell[   33173] = 32'h900beea5;
    ram_cell[   33174] = 32'h767ec051;
    ram_cell[   33175] = 32'hed64a18c;
    ram_cell[   33176] = 32'hdf8582a5;
    ram_cell[   33177] = 32'hb298c198;
    ram_cell[   33178] = 32'hbe982f21;
    ram_cell[   33179] = 32'h6d8b76f7;
    ram_cell[   33180] = 32'h04552792;
    ram_cell[   33181] = 32'h67dc16f6;
    ram_cell[   33182] = 32'h06fa51cf;
    ram_cell[   33183] = 32'h6d57ad4b;
    ram_cell[   33184] = 32'h276e6fad;
    ram_cell[   33185] = 32'hb6c9df25;
    ram_cell[   33186] = 32'hb3c650a9;
    ram_cell[   33187] = 32'h8f4319fc;
    ram_cell[   33188] = 32'h8d164fe0;
    ram_cell[   33189] = 32'h64482388;
    ram_cell[   33190] = 32'h8d9498ad;
    ram_cell[   33191] = 32'h3ba7c694;
    ram_cell[   33192] = 32'h56f19242;
    ram_cell[   33193] = 32'hdcf369b5;
    ram_cell[   33194] = 32'hf6998a11;
    ram_cell[   33195] = 32'hf4d9708c;
    ram_cell[   33196] = 32'h38582f22;
    ram_cell[   33197] = 32'hf5621066;
    ram_cell[   33198] = 32'h086e120c;
    ram_cell[   33199] = 32'haccb66c5;
    ram_cell[   33200] = 32'hb4b8bf69;
    ram_cell[   33201] = 32'h1297dca4;
    ram_cell[   33202] = 32'h3e1bd859;
    ram_cell[   33203] = 32'h2bb0307b;
    ram_cell[   33204] = 32'h590be8ed;
    ram_cell[   33205] = 32'h8590aeb7;
    ram_cell[   33206] = 32'h604d8519;
    ram_cell[   33207] = 32'haf173a22;
    ram_cell[   33208] = 32'h7857ed31;
    ram_cell[   33209] = 32'h697cbf2e;
    ram_cell[   33210] = 32'he5b540cb;
    ram_cell[   33211] = 32'h22888bcc;
    ram_cell[   33212] = 32'hb9681239;
    ram_cell[   33213] = 32'h26e7a5c2;
    ram_cell[   33214] = 32'hdadcef1b;
    ram_cell[   33215] = 32'h932b50bb;
    ram_cell[   33216] = 32'he1fb471a;
    ram_cell[   33217] = 32'hf61667aa;
    ram_cell[   33218] = 32'h22e120e0;
    ram_cell[   33219] = 32'h33b25707;
    ram_cell[   33220] = 32'hdbfadafe;
    ram_cell[   33221] = 32'h0ce6fa42;
    ram_cell[   33222] = 32'he2c565b1;
    ram_cell[   33223] = 32'ha3e1f217;
    ram_cell[   33224] = 32'h7730a6cb;
    ram_cell[   33225] = 32'h57fd7c7f;
    ram_cell[   33226] = 32'hdf7ab71e;
    ram_cell[   33227] = 32'h8fc5a7ca;
    ram_cell[   33228] = 32'hb377f53b;
    ram_cell[   33229] = 32'hbe7d3e7d;
    ram_cell[   33230] = 32'he580a277;
    ram_cell[   33231] = 32'hd0cc0776;
    ram_cell[   33232] = 32'hc3d700b9;
    ram_cell[   33233] = 32'h19a11cd2;
    ram_cell[   33234] = 32'ha4f3fbf5;
    ram_cell[   33235] = 32'ha16343c7;
    ram_cell[   33236] = 32'h02f61a17;
    ram_cell[   33237] = 32'h233e9bcd;
    ram_cell[   33238] = 32'h1de8d5ae;
    ram_cell[   33239] = 32'h6ec7298c;
    ram_cell[   33240] = 32'h703b7ff4;
    ram_cell[   33241] = 32'h6ae6f037;
    ram_cell[   33242] = 32'h6df7ab27;
    ram_cell[   33243] = 32'h3526fef6;
    ram_cell[   33244] = 32'hbf960386;
    ram_cell[   33245] = 32'h8e504dfa;
    ram_cell[   33246] = 32'he46d507c;
    ram_cell[   33247] = 32'h37115bc8;
    ram_cell[   33248] = 32'haadcfdac;
    ram_cell[   33249] = 32'h4af6351e;
    ram_cell[   33250] = 32'h45c82ec4;
    ram_cell[   33251] = 32'h4d3e92a9;
    ram_cell[   33252] = 32'h9f0b1f82;
    ram_cell[   33253] = 32'hc478ae9c;
    ram_cell[   33254] = 32'hc1d77bfa;
    ram_cell[   33255] = 32'hf196cf9e;
    ram_cell[   33256] = 32'h6ce9b31f;
    ram_cell[   33257] = 32'h3bb301c2;
    ram_cell[   33258] = 32'hf1cdc883;
    ram_cell[   33259] = 32'hb272a7ee;
    ram_cell[   33260] = 32'h7864adc8;
    ram_cell[   33261] = 32'h81a33c4e;
    ram_cell[   33262] = 32'h7af546fb;
    ram_cell[   33263] = 32'h3d4ad52f;
    ram_cell[   33264] = 32'hef3b177c;
    ram_cell[   33265] = 32'h5cd14cd8;
    ram_cell[   33266] = 32'h4d6c98a9;
    ram_cell[   33267] = 32'h9f19f494;
    ram_cell[   33268] = 32'h8e02569f;
    ram_cell[   33269] = 32'h30a36d86;
    ram_cell[   33270] = 32'h97be7d29;
    ram_cell[   33271] = 32'ha1e3c51f;
    ram_cell[   33272] = 32'hd877827c;
    ram_cell[   33273] = 32'h625402b9;
    ram_cell[   33274] = 32'h1791d1cf;
    ram_cell[   33275] = 32'h9a872f70;
    ram_cell[   33276] = 32'h5a6d4560;
    ram_cell[   33277] = 32'h1f687713;
    ram_cell[   33278] = 32'hd460285d;
    ram_cell[   33279] = 32'hfd37fe7c;
    ram_cell[   33280] = 32'h9d664914;
    ram_cell[   33281] = 32'h98ee7d0a;
    ram_cell[   33282] = 32'hb7b368ff;
    ram_cell[   33283] = 32'hd10719e6;
    ram_cell[   33284] = 32'h88dd4b64;
    ram_cell[   33285] = 32'hfaba88cb;
    ram_cell[   33286] = 32'h36166a63;
    ram_cell[   33287] = 32'h6bd4b827;
    ram_cell[   33288] = 32'hdf53845f;
    ram_cell[   33289] = 32'hbd167c7b;
    ram_cell[   33290] = 32'h47b153e6;
    ram_cell[   33291] = 32'h23f05a38;
    ram_cell[   33292] = 32'hdd95d517;
    ram_cell[   33293] = 32'he4a16dc0;
    ram_cell[   33294] = 32'hef20c1ea;
    ram_cell[   33295] = 32'hb50635dd;
    ram_cell[   33296] = 32'haa1b0963;
    ram_cell[   33297] = 32'h13cbecda;
    ram_cell[   33298] = 32'hd2e3a725;
    ram_cell[   33299] = 32'h3baf044e;
    ram_cell[   33300] = 32'h2fdaa144;
    ram_cell[   33301] = 32'h0278b713;
    ram_cell[   33302] = 32'h4f41777e;
    ram_cell[   33303] = 32'hc023bf4d;
    ram_cell[   33304] = 32'h1684f6ba;
    ram_cell[   33305] = 32'h0171a18d;
    ram_cell[   33306] = 32'h143a5de2;
    ram_cell[   33307] = 32'hc679bc4a;
    ram_cell[   33308] = 32'h3fb65878;
    ram_cell[   33309] = 32'h19a5000c;
    ram_cell[   33310] = 32'hf5a89c42;
    ram_cell[   33311] = 32'h327fd786;
    ram_cell[   33312] = 32'hf12f5a55;
    ram_cell[   33313] = 32'hdb4f6891;
    ram_cell[   33314] = 32'h297965a9;
    ram_cell[   33315] = 32'h266d02d1;
    ram_cell[   33316] = 32'hdb650d5a;
    ram_cell[   33317] = 32'h7aee0a99;
    ram_cell[   33318] = 32'h4887a674;
    ram_cell[   33319] = 32'hefae8891;
    ram_cell[   33320] = 32'h3c46b656;
    ram_cell[   33321] = 32'hdfe337e4;
    ram_cell[   33322] = 32'hbff78bc8;
    ram_cell[   33323] = 32'h9fb8cb49;
    ram_cell[   33324] = 32'hc53d6b3e;
    ram_cell[   33325] = 32'hec91dc96;
    ram_cell[   33326] = 32'h7ffb0ef8;
    ram_cell[   33327] = 32'h71d3b32b;
    ram_cell[   33328] = 32'hba574f5e;
    ram_cell[   33329] = 32'h3f85a2b7;
    ram_cell[   33330] = 32'hcb15d0d6;
    ram_cell[   33331] = 32'hb81a5cba;
    ram_cell[   33332] = 32'h1acb2880;
    ram_cell[   33333] = 32'h92652d21;
    ram_cell[   33334] = 32'h14f35c81;
    ram_cell[   33335] = 32'hf0f0ed8d;
    ram_cell[   33336] = 32'h93b24d4c;
    ram_cell[   33337] = 32'h7235acb9;
    ram_cell[   33338] = 32'h50849a21;
    ram_cell[   33339] = 32'h3da6d471;
    ram_cell[   33340] = 32'h8cdcbeff;
    ram_cell[   33341] = 32'hb331a34c;
    ram_cell[   33342] = 32'h06555325;
    ram_cell[   33343] = 32'h2e5bdd08;
    ram_cell[   33344] = 32'hcd2eb8e6;
    ram_cell[   33345] = 32'hf5d9d44c;
    ram_cell[   33346] = 32'h858814fc;
    ram_cell[   33347] = 32'hb5bebd5a;
    ram_cell[   33348] = 32'hf64c7a08;
    ram_cell[   33349] = 32'h768eb9f4;
    ram_cell[   33350] = 32'h22cb6604;
    ram_cell[   33351] = 32'h7b57e52c;
    ram_cell[   33352] = 32'h736fe7cf;
    ram_cell[   33353] = 32'hb94d34cf;
    ram_cell[   33354] = 32'h8dd60712;
    ram_cell[   33355] = 32'hda9c4ea7;
    ram_cell[   33356] = 32'hca4de6c8;
    ram_cell[   33357] = 32'h0ebe1638;
    ram_cell[   33358] = 32'hfbf835a9;
    ram_cell[   33359] = 32'h2cd9d39a;
    ram_cell[   33360] = 32'h9828dbeb;
    ram_cell[   33361] = 32'h7f4dd487;
    ram_cell[   33362] = 32'h58a6a969;
    ram_cell[   33363] = 32'hd3c149a0;
    ram_cell[   33364] = 32'hb8684c90;
    ram_cell[   33365] = 32'hb503258b;
    ram_cell[   33366] = 32'heb1c2be0;
    ram_cell[   33367] = 32'h54c16400;
    ram_cell[   33368] = 32'hf51e2c51;
    ram_cell[   33369] = 32'h9ebcadea;
    ram_cell[   33370] = 32'h50bd3202;
    ram_cell[   33371] = 32'hee9e86a4;
    ram_cell[   33372] = 32'h445a82ca;
    ram_cell[   33373] = 32'hcae9feda;
    ram_cell[   33374] = 32'hcfb7cb4e;
    ram_cell[   33375] = 32'hfdd3f508;
    ram_cell[   33376] = 32'he5879b43;
    ram_cell[   33377] = 32'h50bb1f5c;
    ram_cell[   33378] = 32'h0da19f72;
    ram_cell[   33379] = 32'h93542bf2;
    ram_cell[   33380] = 32'h921f2b2f;
    ram_cell[   33381] = 32'h178a0284;
    ram_cell[   33382] = 32'h815a6ca7;
    ram_cell[   33383] = 32'h2a598fd2;
    ram_cell[   33384] = 32'h7f85d904;
    ram_cell[   33385] = 32'hc3d39080;
    ram_cell[   33386] = 32'h187a6aa9;
    ram_cell[   33387] = 32'hfe9535d6;
    ram_cell[   33388] = 32'h3d90f8aa;
    ram_cell[   33389] = 32'h8caa17b0;
    ram_cell[   33390] = 32'h058ee9db;
    ram_cell[   33391] = 32'hb16d585c;
    ram_cell[   33392] = 32'h1aae97ef;
    ram_cell[   33393] = 32'hcbb0278a;
    ram_cell[   33394] = 32'h02c3c1ac;
    ram_cell[   33395] = 32'h07bf1509;
    ram_cell[   33396] = 32'hd9a6ee69;
    ram_cell[   33397] = 32'h7e1e87f9;
    ram_cell[   33398] = 32'h837cd467;
    ram_cell[   33399] = 32'hcf543f66;
    ram_cell[   33400] = 32'hf96dca22;
    ram_cell[   33401] = 32'h62878456;
    ram_cell[   33402] = 32'h0c0461d4;
    ram_cell[   33403] = 32'he932906c;
    ram_cell[   33404] = 32'h13fcebd9;
    ram_cell[   33405] = 32'h39b4cd5c;
    ram_cell[   33406] = 32'h308092de;
    ram_cell[   33407] = 32'hd6b69e2a;
    ram_cell[   33408] = 32'hdef61a1c;
    ram_cell[   33409] = 32'h58e6d6af;
    ram_cell[   33410] = 32'hb0f91c0d;
    ram_cell[   33411] = 32'h498eb82d;
    ram_cell[   33412] = 32'ha2db4748;
    ram_cell[   33413] = 32'hce5bc75f;
    ram_cell[   33414] = 32'h90146cf2;
    ram_cell[   33415] = 32'heae5b759;
    ram_cell[   33416] = 32'h55c00de8;
    ram_cell[   33417] = 32'h80a8cc46;
    ram_cell[   33418] = 32'h0a070e50;
    ram_cell[   33419] = 32'hbcb51891;
    ram_cell[   33420] = 32'hb7d7f212;
    ram_cell[   33421] = 32'h3d48cf77;
    ram_cell[   33422] = 32'ha23df2d9;
    ram_cell[   33423] = 32'hc81bf3f3;
    ram_cell[   33424] = 32'he27c887a;
    ram_cell[   33425] = 32'hde335b7c;
    ram_cell[   33426] = 32'h31d68895;
    ram_cell[   33427] = 32'h1631424f;
    ram_cell[   33428] = 32'h0d399b8d;
    ram_cell[   33429] = 32'hda33f05b;
    ram_cell[   33430] = 32'hb7b61855;
    ram_cell[   33431] = 32'h76b54f2d;
    ram_cell[   33432] = 32'h4e566a9b;
    ram_cell[   33433] = 32'hb1795bd3;
    ram_cell[   33434] = 32'hd6c3d0a9;
    ram_cell[   33435] = 32'h40181572;
    ram_cell[   33436] = 32'h5a9da634;
    ram_cell[   33437] = 32'h0dd66632;
    ram_cell[   33438] = 32'h363922b9;
    ram_cell[   33439] = 32'h2b69fb19;
    ram_cell[   33440] = 32'haecfb68c;
    ram_cell[   33441] = 32'h8ee4bd18;
    ram_cell[   33442] = 32'hc9a8dcf1;
    ram_cell[   33443] = 32'h27881025;
    ram_cell[   33444] = 32'h31632b85;
    ram_cell[   33445] = 32'hcbc381d5;
    ram_cell[   33446] = 32'h6a36c310;
    ram_cell[   33447] = 32'hb012fa1c;
    ram_cell[   33448] = 32'hdafb2874;
    ram_cell[   33449] = 32'h6b475fab;
    ram_cell[   33450] = 32'h893d221a;
    ram_cell[   33451] = 32'h6de25978;
    ram_cell[   33452] = 32'h4c4120b4;
    ram_cell[   33453] = 32'h0058f796;
    ram_cell[   33454] = 32'haff42118;
    ram_cell[   33455] = 32'he11c9a1d;
    ram_cell[   33456] = 32'he2e7f8b0;
    ram_cell[   33457] = 32'hfae18472;
    ram_cell[   33458] = 32'he6d1ddc4;
    ram_cell[   33459] = 32'h7fff6e61;
    ram_cell[   33460] = 32'h2447f583;
    ram_cell[   33461] = 32'h45651b6a;
    ram_cell[   33462] = 32'hd1c42d93;
    ram_cell[   33463] = 32'hef4a33ab;
    ram_cell[   33464] = 32'h0e404254;
    ram_cell[   33465] = 32'h3087a494;
    ram_cell[   33466] = 32'h01c10cdd;
    ram_cell[   33467] = 32'h656ac4df;
    ram_cell[   33468] = 32'ha3a424cd;
    ram_cell[   33469] = 32'h4ca8fdcd;
    ram_cell[   33470] = 32'h7eb206e9;
    ram_cell[   33471] = 32'h917bc0f4;
    ram_cell[   33472] = 32'hfcdebd6e;
    ram_cell[   33473] = 32'hbfd7fba1;
    ram_cell[   33474] = 32'h25671d27;
    ram_cell[   33475] = 32'h2e570269;
    ram_cell[   33476] = 32'h6e7a27c3;
    ram_cell[   33477] = 32'h8e705d99;
    ram_cell[   33478] = 32'h35da8f6f;
    ram_cell[   33479] = 32'h5c5d8ca2;
    ram_cell[   33480] = 32'hd7949503;
    ram_cell[   33481] = 32'he44b75c6;
    ram_cell[   33482] = 32'hee4fdc60;
    ram_cell[   33483] = 32'h7d02995f;
    ram_cell[   33484] = 32'h28d4761d;
    ram_cell[   33485] = 32'h867e5159;
    ram_cell[   33486] = 32'h79a05656;
    ram_cell[   33487] = 32'hccfe81e6;
    ram_cell[   33488] = 32'hce21e516;
    ram_cell[   33489] = 32'h702a1617;
    ram_cell[   33490] = 32'h0191acb1;
    ram_cell[   33491] = 32'h36af52da;
    ram_cell[   33492] = 32'h340768f9;
    ram_cell[   33493] = 32'h71c75b9a;
    ram_cell[   33494] = 32'he23e7f45;
    ram_cell[   33495] = 32'hb800ae80;
    ram_cell[   33496] = 32'h72ad706c;
    ram_cell[   33497] = 32'h5672d0c9;
    ram_cell[   33498] = 32'ha6d902b0;
    ram_cell[   33499] = 32'hf11a9a14;
    ram_cell[   33500] = 32'h0b5f9066;
    ram_cell[   33501] = 32'ha5ce4e40;
    ram_cell[   33502] = 32'h8ff23e44;
    ram_cell[   33503] = 32'hb237b83b;
    ram_cell[   33504] = 32'hfaabca2e;
    ram_cell[   33505] = 32'h51ff1268;
    ram_cell[   33506] = 32'h65453c87;
    ram_cell[   33507] = 32'h69024ea9;
    ram_cell[   33508] = 32'hf134a611;
    ram_cell[   33509] = 32'h75ba0b7c;
    ram_cell[   33510] = 32'hd955e44d;
    ram_cell[   33511] = 32'h946e8f98;
    ram_cell[   33512] = 32'h3ae17905;
    ram_cell[   33513] = 32'hccf680c4;
    ram_cell[   33514] = 32'h31f0a101;
    ram_cell[   33515] = 32'h850459e9;
    ram_cell[   33516] = 32'h15b1184d;
    ram_cell[   33517] = 32'h233a5333;
    ram_cell[   33518] = 32'hda97ded6;
    ram_cell[   33519] = 32'h1c332d65;
    ram_cell[   33520] = 32'hfeb8dc41;
    ram_cell[   33521] = 32'hcb3f211e;
    ram_cell[   33522] = 32'h0f8713e4;
    ram_cell[   33523] = 32'h7ced3f99;
    ram_cell[   33524] = 32'h1d03eecf;
    ram_cell[   33525] = 32'h54670136;
    ram_cell[   33526] = 32'h6449ce00;
    ram_cell[   33527] = 32'h95357b64;
    ram_cell[   33528] = 32'h954291fb;
    ram_cell[   33529] = 32'h5d8cc440;
    ram_cell[   33530] = 32'hf4233322;
    ram_cell[   33531] = 32'h287e29fa;
    ram_cell[   33532] = 32'h3d8f06b8;
    ram_cell[   33533] = 32'h771cadf8;
    ram_cell[   33534] = 32'h2ae0a711;
    ram_cell[   33535] = 32'h1ce86b19;
    ram_cell[   33536] = 32'hb14517ff;
    ram_cell[   33537] = 32'hacc67262;
    ram_cell[   33538] = 32'h90766968;
    ram_cell[   33539] = 32'he44397df;
    ram_cell[   33540] = 32'hc2cf6630;
    ram_cell[   33541] = 32'h9b5802cf;
    ram_cell[   33542] = 32'hae932b66;
    ram_cell[   33543] = 32'h0312dacc;
    ram_cell[   33544] = 32'h0af68494;
    ram_cell[   33545] = 32'hc53a9665;
    ram_cell[   33546] = 32'h52054d29;
    ram_cell[   33547] = 32'h2e2b8715;
    ram_cell[   33548] = 32'hb617930e;
    ram_cell[   33549] = 32'hc2950835;
    ram_cell[   33550] = 32'h97cf6e82;
    ram_cell[   33551] = 32'h290a80d1;
    ram_cell[   33552] = 32'h3868591d;
    ram_cell[   33553] = 32'hbb58fca5;
    ram_cell[   33554] = 32'h3bf60357;
    ram_cell[   33555] = 32'hb9b27bee;
    ram_cell[   33556] = 32'h4c85e9b2;
    ram_cell[   33557] = 32'ha542e11e;
    ram_cell[   33558] = 32'h4c2e01ff;
    ram_cell[   33559] = 32'h89ad50a9;
    ram_cell[   33560] = 32'h74fdabe8;
    ram_cell[   33561] = 32'hfbbe537e;
    ram_cell[   33562] = 32'hfcfa87fa;
    ram_cell[   33563] = 32'h3767c044;
    ram_cell[   33564] = 32'h13ec1813;
    ram_cell[   33565] = 32'ha5cf6a53;
    ram_cell[   33566] = 32'h9ef7c833;
    ram_cell[   33567] = 32'h5ae9a307;
    ram_cell[   33568] = 32'hbf68ed6a;
    ram_cell[   33569] = 32'h74894eab;
    ram_cell[   33570] = 32'h92f62bd2;
    ram_cell[   33571] = 32'he0cbfe63;
    ram_cell[   33572] = 32'he9fc962f;
    ram_cell[   33573] = 32'h91402795;
    ram_cell[   33574] = 32'hc2d55ec6;
    ram_cell[   33575] = 32'h6c6faedf;
    ram_cell[   33576] = 32'hd55f850b;
    ram_cell[   33577] = 32'h4d73ee09;
    ram_cell[   33578] = 32'h2b8ddf89;
    ram_cell[   33579] = 32'hc618ae79;
    ram_cell[   33580] = 32'h285f8377;
    ram_cell[   33581] = 32'h15fec8a9;
    ram_cell[   33582] = 32'h023cbcfb;
    ram_cell[   33583] = 32'h5f65a11a;
    ram_cell[   33584] = 32'hbbc76a20;
    ram_cell[   33585] = 32'hf5904f89;
    ram_cell[   33586] = 32'h48f2f695;
    ram_cell[   33587] = 32'ha0b6e061;
    ram_cell[   33588] = 32'hf9a20c54;
    ram_cell[   33589] = 32'h17dcbc90;
    ram_cell[   33590] = 32'he1b887ed;
    ram_cell[   33591] = 32'h12ce2fc3;
    ram_cell[   33592] = 32'hb90a8b7c;
    ram_cell[   33593] = 32'h8e3eb14c;
    ram_cell[   33594] = 32'h87736d11;
    ram_cell[   33595] = 32'hfa1d2968;
    ram_cell[   33596] = 32'h78643d84;
    ram_cell[   33597] = 32'h60a41572;
    ram_cell[   33598] = 32'hf6b78e86;
    ram_cell[   33599] = 32'h239ed45b;
    ram_cell[   33600] = 32'hc6353131;
    ram_cell[   33601] = 32'hc172fdac;
    ram_cell[   33602] = 32'hd21ce66e;
    ram_cell[   33603] = 32'hbcba7ef9;
    ram_cell[   33604] = 32'h0cf4c5c6;
    ram_cell[   33605] = 32'h322e4c00;
    ram_cell[   33606] = 32'h4a65003c;
    ram_cell[   33607] = 32'hd5f920e3;
    ram_cell[   33608] = 32'h745e1b15;
    ram_cell[   33609] = 32'h3c513b58;
    ram_cell[   33610] = 32'h9f8b12f5;
    ram_cell[   33611] = 32'hf4b468e5;
    ram_cell[   33612] = 32'h64dee14f;
    ram_cell[   33613] = 32'h87f04b25;
    ram_cell[   33614] = 32'hd06c9bef;
    ram_cell[   33615] = 32'hd208873d;
    ram_cell[   33616] = 32'h2dfd3ae2;
    ram_cell[   33617] = 32'h57e62daa;
    ram_cell[   33618] = 32'hcc680f0f;
    ram_cell[   33619] = 32'hbbdebb4a;
    ram_cell[   33620] = 32'h553525d2;
    ram_cell[   33621] = 32'h210c1e4e;
    ram_cell[   33622] = 32'h04a60826;
    ram_cell[   33623] = 32'h9d251ec6;
    ram_cell[   33624] = 32'h4b8002d7;
    ram_cell[   33625] = 32'h838edc9f;
    ram_cell[   33626] = 32'h4ea580cd;
    ram_cell[   33627] = 32'h7fc6650c;
    ram_cell[   33628] = 32'hcc6053ec;
    ram_cell[   33629] = 32'h72b19059;
    ram_cell[   33630] = 32'h0e0eb004;
    ram_cell[   33631] = 32'h98320f76;
    ram_cell[   33632] = 32'h2caa3580;
    ram_cell[   33633] = 32'hc189d253;
    ram_cell[   33634] = 32'h083c0d44;
    ram_cell[   33635] = 32'h98d5c159;
    ram_cell[   33636] = 32'hfcfcc946;
    ram_cell[   33637] = 32'h6bcf2f8a;
    ram_cell[   33638] = 32'h8e1f6dab;
    ram_cell[   33639] = 32'hf048fedc;
    ram_cell[   33640] = 32'h51ad8189;
    ram_cell[   33641] = 32'he85e48e7;
    ram_cell[   33642] = 32'h334b8950;
    ram_cell[   33643] = 32'hda77a617;
    ram_cell[   33644] = 32'hdc5bd9eb;
    ram_cell[   33645] = 32'h2a221530;
    ram_cell[   33646] = 32'h882e0111;
    ram_cell[   33647] = 32'hd59aa8f8;
    ram_cell[   33648] = 32'h6d45b2c0;
    ram_cell[   33649] = 32'hee4597de;
    ram_cell[   33650] = 32'h8e737a64;
    ram_cell[   33651] = 32'hb97392f6;
    ram_cell[   33652] = 32'hfff49386;
    ram_cell[   33653] = 32'ha67d0ffd;
    ram_cell[   33654] = 32'h41e95d2a;
    ram_cell[   33655] = 32'h1077033c;
    ram_cell[   33656] = 32'hebdee191;
    ram_cell[   33657] = 32'h7449c397;
    ram_cell[   33658] = 32'ha46a8375;
    ram_cell[   33659] = 32'h8920a34c;
    ram_cell[   33660] = 32'h2221573b;
    ram_cell[   33661] = 32'h159ddc65;
    ram_cell[   33662] = 32'h4d9fc1b8;
    ram_cell[   33663] = 32'h2da8e512;
    ram_cell[   33664] = 32'h0058fab1;
    ram_cell[   33665] = 32'h37e2bf59;
    ram_cell[   33666] = 32'h5bf83f4d;
    ram_cell[   33667] = 32'hc2c7a2a9;
    ram_cell[   33668] = 32'hedfab5c8;
    ram_cell[   33669] = 32'hda45e3e3;
    ram_cell[   33670] = 32'hd5cc6f43;
    ram_cell[   33671] = 32'h85c7677d;
    ram_cell[   33672] = 32'h77ed787c;
    ram_cell[   33673] = 32'h4ca284bc;
    ram_cell[   33674] = 32'h15737cf8;
    ram_cell[   33675] = 32'h36c7b237;
    ram_cell[   33676] = 32'h598b945b;
    ram_cell[   33677] = 32'h58361e4b;
    ram_cell[   33678] = 32'h437978e5;
    ram_cell[   33679] = 32'h564df28f;
    ram_cell[   33680] = 32'h1c9db7fc;
    ram_cell[   33681] = 32'h0aad6af2;
    ram_cell[   33682] = 32'hceaf290b;
    ram_cell[   33683] = 32'h81913b8a;
    ram_cell[   33684] = 32'had450c79;
    ram_cell[   33685] = 32'hb7a150fe;
    ram_cell[   33686] = 32'h92221c9e;
    ram_cell[   33687] = 32'h1b1a1622;
    ram_cell[   33688] = 32'hebcfe8e5;
    ram_cell[   33689] = 32'hb9973576;
    ram_cell[   33690] = 32'h4678b385;
    ram_cell[   33691] = 32'h7d3d2e18;
    ram_cell[   33692] = 32'h23640ae3;
    ram_cell[   33693] = 32'h81d168e3;
    ram_cell[   33694] = 32'h13fd07d4;
    ram_cell[   33695] = 32'hb7342fc3;
    ram_cell[   33696] = 32'h9fba95f9;
    ram_cell[   33697] = 32'h20f0a88e;
    ram_cell[   33698] = 32'hc64d91bf;
    ram_cell[   33699] = 32'h07b00e0b;
    ram_cell[   33700] = 32'hca491c73;
    ram_cell[   33701] = 32'h78be934a;
    ram_cell[   33702] = 32'hdc8de5f3;
    ram_cell[   33703] = 32'h39f459f8;
    ram_cell[   33704] = 32'h4e7d6e5e;
    ram_cell[   33705] = 32'h7607af3a;
    ram_cell[   33706] = 32'hcd7a89c7;
    ram_cell[   33707] = 32'h3847fa81;
    ram_cell[   33708] = 32'h43c4f0e3;
    ram_cell[   33709] = 32'hdd061d0c;
    ram_cell[   33710] = 32'h76d5dd87;
    ram_cell[   33711] = 32'he47c84d5;
    ram_cell[   33712] = 32'h223e5a22;
    ram_cell[   33713] = 32'hf2dd42fe;
    ram_cell[   33714] = 32'h31579209;
    ram_cell[   33715] = 32'h02f41232;
    ram_cell[   33716] = 32'hb90c348c;
    ram_cell[   33717] = 32'hc7cce12d;
    ram_cell[   33718] = 32'hf058096d;
    ram_cell[   33719] = 32'hc49f9913;
    ram_cell[   33720] = 32'hac885559;
    ram_cell[   33721] = 32'hd1df2aad;
    ram_cell[   33722] = 32'hb84e81f1;
    ram_cell[   33723] = 32'h382ec88d;
    ram_cell[   33724] = 32'h2cea04f9;
    ram_cell[   33725] = 32'h37b0cf8e;
    ram_cell[   33726] = 32'hf27caf53;
    ram_cell[   33727] = 32'h12d17c64;
    ram_cell[   33728] = 32'h7f95983f;
    ram_cell[   33729] = 32'hf28fb629;
    ram_cell[   33730] = 32'he868ef9b;
    ram_cell[   33731] = 32'h6af9a9d0;
    ram_cell[   33732] = 32'h6afe1a51;
    ram_cell[   33733] = 32'h4a9017dc;
    ram_cell[   33734] = 32'h349fca8d;
    ram_cell[   33735] = 32'h6be80817;
    ram_cell[   33736] = 32'hbe2491b7;
    ram_cell[   33737] = 32'heb9d0988;
    ram_cell[   33738] = 32'hada8f913;
    ram_cell[   33739] = 32'h791bea42;
    ram_cell[   33740] = 32'h946864f6;
    ram_cell[   33741] = 32'h6895290c;
    ram_cell[   33742] = 32'hdfe42673;
    ram_cell[   33743] = 32'h037808b2;
    ram_cell[   33744] = 32'h4a26f073;
    ram_cell[   33745] = 32'hdf313978;
    ram_cell[   33746] = 32'h29360ac7;
    ram_cell[   33747] = 32'h1f29ae99;
    ram_cell[   33748] = 32'h1f38694b;
    ram_cell[   33749] = 32'h2343349d;
    ram_cell[   33750] = 32'h31ee5172;
    ram_cell[   33751] = 32'h7e9a3102;
    ram_cell[   33752] = 32'h265dabec;
    ram_cell[   33753] = 32'hf5691939;
    ram_cell[   33754] = 32'h9497f228;
    ram_cell[   33755] = 32'h375af209;
    ram_cell[   33756] = 32'h4712dadf;
    ram_cell[   33757] = 32'h5dab48f2;
    ram_cell[   33758] = 32'h5000fe04;
    ram_cell[   33759] = 32'hd21dd069;
    ram_cell[   33760] = 32'h4686a17a;
    ram_cell[   33761] = 32'h6cd4c4ef;
    ram_cell[   33762] = 32'hfc31e88c;
    ram_cell[   33763] = 32'h973ec04c;
    ram_cell[   33764] = 32'hdd2abfc9;
    ram_cell[   33765] = 32'h5df2d70a;
    ram_cell[   33766] = 32'h6246efaf;
    ram_cell[   33767] = 32'h6a918996;
    ram_cell[   33768] = 32'h09cc24c8;
    ram_cell[   33769] = 32'h2e9da8cd;
    ram_cell[   33770] = 32'h1de83eb5;
    ram_cell[   33771] = 32'hafb146d5;
    ram_cell[   33772] = 32'hb22bd386;
    ram_cell[   33773] = 32'h4eb9726d;
    ram_cell[   33774] = 32'hd38df6a8;
    ram_cell[   33775] = 32'h66562278;
    ram_cell[   33776] = 32'h547209b2;
    ram_cell[   33777] = 32'h4ba31995;
    ram_cell[   33778] = 32'h472d47fc;
    ram_cell[   33779] = 32'h2c14c387;
    ram_cell[   33780] = 32'ha749f5a3;
    ram_cell[   33781] = 32'h737dd4c2;
    ram_cell[   33782] = 32'h2f9710bb;
    ram_cell[   33783] = 32'heef8a04a;
    ram_cell[   33784] = 32'h6064d47e;
    ram_cell[   33785] = 32'hb0d86d4a;
    ram_cell[   33786] = 32'h9a885654;
    ram_cell[   33787] = 32'h0e985f2e;
    ram_cell[   33788] = 32'h805b9301;
    ram_cell[   33789] = 32'h7fb4d76c;
    ram_cell[   33790] = 32'h04b14145;
    ram_cell[   33791] = 32'h37cd7b3e;
    ram_cell[   33792] = 32'h39a3c1e0;
    ram_cell[   33793] = 32'h5e4de20b;
    ram_cell[   33794] = 32'hbd19ce78;
    ram_cell[   33795] = 32'h6d8adfb2;
    ram_cell[   33796] = 32'h79f4a00d;
    ram_cell[   33797] = 32'h3362fc32;
    ram_cell[   33798] = 32'h0594793f;
    ram_cell[   33799] = 32'h9325f2ac;
    ram_cell[   33800] = 32'hb8092687;
    ram_cell[   33801] = 32'hf71e5525;
    ram_cell[   33802] = 32'hc436d00e;
    ram_cell[   33803] = 32'h7d624caf;
    ram_cell[   33804] = 32'h232b2fcb;
    ram_cell[   33805] = 32'h4fe7962e;
    ram_cell[   33806] = 32'he40e0fe5;
    ram_cell[   33807] = 32'hf8bb43c0;
    ram_cell[   33808] = 32'h2520ea64;
    ram_cell[   33809] = 32'h95393469;
    ram_cell[   33810] = 32'h0022e067;
    ram_cell[   33811] = 32'h38c5e921;
    ram_cell[   33812] = 32'h7a926c2a;
    ram_cell[   33813] = 32'hb91cceb7;
    ram_cell[   33814] = 32'h23bb028d;
    ram_cell[   33815] = 32'hbce4ade2;
    ram_cell[   33816] = 32'heb5842c7;
    ram_cell[   33817] = 32'h42585246;
    ram_cell[   33818] = 32'h09c26764;
    ram_cell[   33819] = 32'h3c59c6f7;
    ram_cell[   33820] = 32'h540993e9;
    ram_cell[   33821] = 32'h402551a8;
    ram_cell[   33822] = 32'h2884d5e5;
    ram_cell[   33823] = 32'h793acf3b;
    ram_cell[   33824] = 32'h2e2909cc;
    ram_cell[   33825] = 32'h919fe56b;
    ram_cell[   33826] = 32'hf7356fec;
    ram_cell[   33827] = 32'h60f054fa;
    ram_cell[   33828] = 32'h9f6543da;
    ram_cell[   33829] = 32'h83d1268c;
    ram_cell[   33830] = 32'h0a7adab5;
    ram_cell[   33831] = 32'hf815f198;
    ram_cell[   33832] = 32'h717b62c7;
    ram_cell[   33833] = 32'h50a104e7;
    ram_cell[   33834] = 32'h342dc11d;
    ram_cell[   33835] = 32'h23c0698f;
    ram_cell[   33836] = 32'h6e33effc;
    ram_cell[   33837] = 32'he3969f9a;
    ram_cell[   33838] = 32'h1af5facf;
    ram_cell[   33839] = 32'hfbcbfe85;
    ram_cell[   33840] = 32'hba736743;
    ram_cell[   33841] = 32'hacdcf8b2;
    ram_cell[   33842] = 32'hc1022e97;
    ram_cell[   33843] = 32'hba9d2f15;
    ram_cell[   33844] = 32'hd6760250;
    ram_cell[   33845] = 32'hc1810be9;
    ram_cell[   33846] = 32'hc735f005;
    ram_cell[   33847] = 32'hf0250f03;
    ram_cell[   33848] = 32'hfdf31428;
    ram_cell[   33849] = 32'h2503deb4;
    ram_cell[   33850] = 32'ha38257bd;
    ram_cell[   33851] = 32'ha4c84a00;
    ram_cell[   33852] = 32'h92285c61;
    ram_cell[   33853] = 32'hdb69e20b;
    ram_cell[   33854] = 32'h5479fa6e;
    ram_cell[   33855] = 32'hb7d14243;
    ram_cell[   33856] = 32'h8fe02243;
    ram_cell[   33857] = 32'hb24d8ed5;
    ram_cell[   33858] = 32'h57627e94;
    ram_cell[   33859] = 32'h88df39c3;
    ram_cell[   33860] = 32'h8a246f4b;
    ram_cell[   33861] = 32'hfe48bde2;
    ram_cell[   33862] = 32'hdadf98f8;
    ram_cell[   33863] = 32'h3b45cd34;
    ram_cell[   33864] = 32'h747fa7eb;
    ram_cell[   33865] = 32'h333b0be7;
    ram_cell[   33866] = 32'h7e5c16f1;
    ram_cell[   33867] = 32'h8202f205;
    ram_cell[   33868] = 32'hddb54d35;
    ram_cell[   33869] = 32'h64b34167;
    ram_cell[   33870] = 32'h9926894f;
    ram_cell[   33871] = 32'h670db3c1;
    ram_cell[   33872] = 32'hfbbbb6f6;
    ram_cell[   33873] = 32'hf1941518;
    ram_cell[   33874] = 32'hec6250f9;
    ram_cell[   33875] = 32'hd9a87b24;
    ram_cell[   33876] = 32'h17c5aaac;
    ram_cell[   33877] = 32'h7891655c;
    ram_cell[   33878] = 32'hd8609e75;
    ram_cell[   33879] = 32'h1de78c0b;
    ram_cell[   33880] = 32'h291cd461;
    ram_cell[   33881] = 32'h56e5ccd0;
    ram_cell[   33882] = 32'hd26d1c57;
    ram_cell[   33883] = 32'h25937e0e;
    ram_cell[   33884] = 32'hd38b7374;
    ram_cell[   33885] = 32'h70f3af28;
    ram_cell[   33886] = 32'h7d91d3ef;
    ram_cell[   33887] = 32'he6e3deab;
    ram_cell[   33888] = 32'hb5b1459c;
    ram_cell[   33889] = 32'h2158c0e0;
    ram_cell[   33890] = 32'h42278115;
    ram_cell[   33891] = 32'habd0c233;
    ram_cell[   33892] = 32'h6de7ad4e;
    ram_cell[   33893] = 32'hc9930110;
    ram_cell[   33894] = 32'h04fb97aa;
    ram_cell[   33895] = 32'h0be11a1e;
    ram_cell[   33896] = 32'h20aca84f;
    ram_cell[   33897] = 32'h5f0045d9;
    ram_cell[   33898] = 32'hc7d57cb4;
    ram_cell[   33899] = 32'h4635c705;
    ram_cell[   33900] = 32'h46dfc49a;
    ram_cell[   33901] = 32'h1a93b74a;
    ram_cell[   33902] = 32'hb9b7882c;
    ram_cell[   33903] = 32'h42a3279f;
    ram_cell[   33904] = 32'h48089fed;
    ram_cell[   33905] = 32'hf1af1809;
    ram_cell[   33906] = 32'h7dfdc82b;
    ram_cell[   33907] = 32'he52c1bd4;
    ram_cell[   33908] = 32'hf097029d;
    ram_cell[   33909] = 32'ha1293142;
    ram_cell[   33910] = 32'h3a24b2b7;
    ram_cell[   33911] = 32'h3336452c;
    ram_cell[   33912] = 32'hddc27ed7;
    ram_cell[   33913] = 32'h1aa4cddd;
    ram_cell[   33914] = 32'h1d6d45ed;
    ram_cell[   33915] = 32'h1bdd6f9c;
    ram_cell[   33916] = 32'h7d5e2e54;
    ram_cell[   33917] = 32'h7d6d1b7e;
    ram_cell[   33918] = 32'h6afe1906;
    ram_cell[   33919] = 32'h3c9053e3;
    ram_cell[   33920] = 32'hc75d8221;
    ram_cell[   33921] = 32'h863ddf08;
    ram_cell[   33922] = 32'h879ef4b5;
    ram_cell[   33923] = 32'hac0e25ba;
    ram_cell[   33924] = 32'h3a565a42;
    ram_cell[   33925] = 32'h5867abd2;
    ram_cell[   33926] = 32'h77d4be11;
    ram_cell[   33927] = 32'hdc0e08b4;
    ram_cell[   33928] = 32'hc9577879;
    ram_cell[   33929] = 32'h9161ec6e;
    ram_cell[   33930] = 32'haf4a7b09;
    ram_cell[   33931] = 32'h3e571137;
    ram_cell[   33932] = 32'hb868bfee;
    ram_cell[   33933] = 32'h9488bb15;
    ram_cell[   33934] = 32'hfd580659;
    ram_cell[   33935] = 32'ha0b2892f;
    ram_cell[   33936] = 32'h28d43910;
    ram_cell[   33937] = 32'h31c9573d;
    ram_cell[   33938] = 32'h449f650a;
    ram_cell[   33939] = 32'h38e43f83;
    ram_cell[   33940] = 32'h3948f6e0;
    ram_cell[   33941] = 32'hfcd7d0c8;
    ram_cell[   33942] = 32'h547b30d7;
    ram_cell[   33943] = 32'hd4ebe7a9;
    ram_cell[   33944] = 32'he225073b;
    ram_cell[   33945] = 32'hc687062b;
    ram_cell[   33946] = 32'h6f298aa9;
    ram_cell[   33947] = 32'h64efd29d;
    ram_cell[   33948] = 32'h80e23907;
    ram_cell[   33949] = 32'hd1693e7d;
    ram_cell[   33950] = 32'h8f9504a3;
    ram_cell[   33951] = 32'h10514e16;
    ram_cell[   33952] = 32'h4e2d1500;
    ram_cell[   33953] = 32'hb72f6a21;
    ram_cell[   33954] = 32'hf2191bcd;
    ram_cell[   33955] = 32'h515e5c61;
    ram_cell[   33956] = 32'hcc4f8b71;
    ram_cell[   33957] = 32'hed470a4d;
    ram_cell[   33958] = 32'h8bb6b8ab;
    ram_cell[   33959] = 32'h580c8baa;
    ram_cell[   33960] = 32'h120ee541;
    ram_cell[   33961] = 32'hd1c417bc;
    ram_cell[   33962] = 32'he20a684a;
    ram_cell[   33963] = 32'hd18ed657;
    ram_cell[   33964] = 32'hcf510850;
    ram_cell[   33965] = 32'h8d20372a;
    ram_cell[   33966] = 32'hfa36d542;
    ram_cell[   33967] = 32'he197b80c;
    ram_cell[   33968] = 32'h0b0f0930;
    ram_cell[   33969] = 32'h841c0ba2;
    ram_cell[   33970] = 32'hb1c73598;
    ram_cell[   33971] = 32'h20c3af2c;
    ram_cell[   33972] = 32'hf0e592ba;
    ram_cell[   33973] = 32'h67fbeb72;
    ram_cell[   33974] = 32'ha07aacac;
    ram_cell[   33975] = 32'h9c510c54;
    ram_cell[   33976] = 32'h74d3d2f0;
    ram_cell[   33977] = 32'h79d8d6ec;
    ram_cell[   33978] = 32'h68eaa5e2;
    ram_cell[   33979] = 32'h28501093;
    ram_cell[   33980] = 32'h66daa0ef;
    ram_cell[   33981] = 32'h149cf52d;
    ram_cell[   33982] = 32'ha831d9ff;
    ram_cell[   33983] = 32'h3a302c47;
    ram_cell[   33984] = 32'h1f069a15;
    ram_cell[   33985] = 32'hb0780635;
    ram_cell[   33986] = 32'h0ce222c2;
    ram_cell[   33987] = 32'ha194dbdb;
    ram_cell[   33988] = 32'h2a76308a;
    ram_cell[   33989] = 32'h43aae5c4;
    ram_cell[   33990] = 32'h5047db6f;
    ram_cell[   33991] = 32'hb2181971;
    ram_cell[   33992] = 32'h694f1d96;
    ram_cell[   33993] = 32'h48ef4bd0;
    ram_cell[   33994] = 32'h6b59868e;
    ram_cell[   33995] = 32'h828f2c2c;
    ram_cell[   33996] = 32'h1e90875d;
    ram_cell[   33997] = 32'h679f2d29;
    ram_cell[   33998] = 32'h148a7579;
    ram_cell[   33999] = 32'h7c85108d;
    ram_cell[   34000] = 32'hcdc1c2bb;
    ram_cell[   34001] = 32'h4c9c4f78;
    ram_cell[   34002] = 32'h0f212c73;
    ram_cell[   34003] = 32'h165572d2;
    ram_cell[   34004] = 32'h0037e661;
    ram_cell[   34005] = 32'h15ea31b7;
    ram_cell[   34006] = 32'hb26f0cf8;
    ram_cell[   34007] = 32'hbe9420e6;
    ram_cell[   34008] = 32'h0b3ff98c;
    ram_cell[   34009] = 32'h71d1df69;
    ram_cell[   34010] = 32'hb92dafc2;
    ram_cell[   34011] = 32'h9902b83d;
    ram_cell[   34012] = 32'h8aa912fa;
    ram_cell[   34013] = 32'h1da5a8dc;
    ram_cell[   34014] = 32'hf0710c00;
    ram_cell[   34015] = 32'h32947aec;
    ram_cell[   34016] = 32'h217b0665;
    ram_cell[   34017] = 32'heb0e7ed4;
    ram_cell[   34018] = 32'h6b3e103e;
    ram_cell[   34019] = 32'hddedeb9f;
    ram_cell[   34020] = 32'h51b7d02b;
    ram_cell[   34021] = 32'h02e56bc0;
    ram_cell[   34022] = 32'hcbe7f53f;
    ram_cell[   34023] = 32'hd69173fd;
    ram_cell[   34024] = 32'h0dcfcdc0;
    ram_cell[   34025] = 32'he0d7f64d;
    ram_cell[   34026] = 32'h43e794c1;
    ram_cell[   34027] = 32'h5ed478b5;
    ram_cell[   34028] = 32'h4215c633;
    ram_cell[   34029] = 32'hd9651a3e;
    ram_cell[   34030] = 32'h8836ef4d;
    ram_cell[   34031] = 32'h27c53dc7;
    ram_cell[   34032] = 32'h0b4c378d;
    ram_cell[   34033] = 32'h25064683;
    ram_cell[   34034] = 32'ha66e9e3a;
    ram_cell[   34035] = 32'hd5a467fd;
    ram_cell[   34036] = 32'h3da4c2ed;
    ram_cell[   34037] = 32'ha423e86f;
    ram_cell[   34038] = 32'h9387a984;
    ram_cell[   34039] = 32'he0143a1f;
    ram_cell[   34040] = 32'h69f96f66;
    ram_cell[   34041] = 32'h16c5dee4;
    ram_cell[   34042] = 32'hff46da1b;
    ram_cell[   34043] = 32'h3bc96e77;
    ram_cell[   34044] = 32'hb55e9174;
    ram_cell[   34045] = 32'h43cfdfe4;
    ram_cell[   34046] = 32'h4b13cd36;
    ram_cell[   34047] = 32'h18ec5be7;
    ram_cell[   34048] = 32'hdda5f4c5;
    ram_cell[   34049] = 32'hce4c2f08;
    ram_cell[   34050] = 32'hcd36de61;
    ram_cell[   34051] = 32'h345b91c4;
    ram_cell[   34052] = 32'hb5dd6fe9;
    ram_cell[   34053] = 32'hfde61b6d;
    ram_cell[   34054] = 32'h400e1199;
    ram_cell[   34055] = 32'h05a75f93;
    ram_cell[   34056] = 32'h41723702;
    ram_cell[   34057] = 32'hb3d24027;
    ram_cell[   34058] = 32'h5bb096d0;
    ram_cell[   34059] = 32'hb4c46eb9;
    ram_cell[   34060] = 32'hf0a79ab9;
    ram_cell[   34061] = 32'had37b8ca;
    ram_cell[   34062] = 32'h86c6df6a;
    ram_cell[   34063] = 32'h05e7a7b1;
    ram_cell[   34064] = 32'h55e90ac5;
    ram_cell[   34065] = 32'hddcc5ed7;
    ram_cell[   34066] = 32'hc2906e35;
    ram_cell[   34067] = 32'h59054cc7;
    ram_cell[   34068] = 32'h2f6cdbc4;
    ram_cell[   34069] = 32'hafd9808f;
    ram_cell[   34070] = 32'h17acb6fd;
    ram_cell[   34071] = 32'he33e1274;
    ram_cell[   34072] = 32'h8b60e0aa;
    ram_cell[   34073] = 32'h76343a1b;
    ram_cell[   34074] = 32'h8e6e1e8e;
    ram_cell[   34075] = 32'h7621c61b;
    ram_cell[   34076] = 32'h8467f4d9;
    ram_cell[   34077] = 32'haf8fb8ea;
    ram_cell[   34078] = 32'h473050ab;
    ram_cell[   34079] = 32'h04fa4a2a;
    ram_cell[   34080] = 32'hba4e1819;
    ram_cell[   34081] = 32'h1523378f;
    ram_cell[   34082] = 32'ha0f68bc9;
    ram_cell[   34083] = 32'hb06f0457;
    ram_cell[   34084] = 32'ha74f01c1;
    ram_cell[   34085] = 32'h2d7506c2;
    ram_cell[   34086] = 32'h3dc3e186;
    ram_cell[   34087] = 32'h13f3e0bb;
    ram_cell[   34088] = 32'hba7b69a8;
    ram_cell[   34089] = 32'he3075807;
    ram_cell[   34090] = 32'h173603bf;
    ram_cell[   34091] = 32'h8f16f83d;
    ram_cell[   34092] = 32'h7d9b056c;
    ram_cell[   34093] = 32'hcd54699c;
    ram_cell[   34094] = 32'h4de8d538;
    ram_cell[   34095] = 32'h8f81351e;
    ram_cell[   34096] = 32'h38e3c496;
    ram_cell[   34097] = 32'h6f4f230a;
    ram_cell[   34098] = 32'h7ac8e015;
    ram_cell[   34099] = 32'hdfe4d2a1;
    ram_cell[   34100] = 32'hfdeeeed7;
    ram_cell[   34101] = 32'he39857a0;
    ram_cell[   34102] = 32'h2f743cc9;
    ram_cell[   34103] = 32'hf4c68f9b;
    ram_cell[   34104] = 32'h6fd4a687;
    ram_cell[   34105] = 32'h838f0de3;
    ram_cell[   34106] = 32'hbdc1c842;
    ram_cell[   34107] = 32'hf16d7d7f;
    ram_cell[   34108] = 32'ha7ada1ba;
    ram_cell[   34109] = 32'h9659ebd8;
    ram_cell[   34110] = 32'hdb5d28df;
    ram_cell[   34111] = 32'hd17ecfa3;
    ram_cell[   34112] = 32'hfebc8b3b;
    ram_cell[   34113] = 32'he2c41767;
    ram_cell[   34114] = 32'h048703eb;
    ram_cell[   34115] = 32'h52892bef;
    ram_cell[   34116] = 32'haa18b1f5;
    ram_cell[   34117] = 32'h6260b3e0;
    ram_cell[   34118] = 32'h6594ffcc;
    ram_cell[   34119] = 32'h4af1f18b;
    ram_cell[   34120] = 32'h084bb486;
    ram_cell[   34121] = 32'h8ad75ea3;
    ram_cell[   34122] = 32'hda92ad7d;
    ram_cell[   34123] = 32'haadffef3;
    ram_cell[   34124] = 32'h292818d9;
    ram_cell[   34125] = 32'h70f79768;
    ram_cell[   34126] = 32'h1b31f8e2;
    ram_cell[   34127] = 32'h2c2e9db9;
    ram_cell[   34128] = 32'h8c42b9dd;
    ram_cell[   34129] = 32'hdb247c36;
    ram_cell[   34130] = 32'hed92f0ed;
    ram_cell[   34131] = 32'h6a4150cd;
    ram_cell[   34132] = 32'hdeb785ea;
    ram_cell[   34133] = 32'h75cbc670;
    ram_cell[   34134] = 32'h737efe24;
    ram_cell[   34135] = 32'hdf3f1696;
    ram_cell[   34136] = 32'hd0940c10;
    ram_cell[   34137] = 32'h4d86c766;
    ram_cell[   34138] = 32'h831d59bb;
    ram_cell[   34139] = 32'hf11ae733;
    ram_cell[   34140] = 32'hdba23621;
    ram_cell[   34141] = 32'hef3f11ce;
    ram_cell[   34142] = 32'h8b21a8e9;
    ram_cell[   34143] = 32'h2e8b1b95;
    ram_cell[   34144] = 32'h8ce54809;
    ram_cell[   34145] = 32'h056cd8a5;
    ram_cell[   34146] = 32'h4f1ab79d;
    ram_cell[   34147] = 32'h2d72cbd0;
    ram_cell[   34148] = 32'hb299e0c7;
    ram_cell[   34149] = 32'h9ce37385;
    ram_cell[   34150] = 32'hd849f3fb;
    ram_cell[   34151] = 32'h7780ec10;
    ram_cell[   34152] = 32'h6172953e;
    ram_cell[   34153] = 32'ha0beb310;
    ram_cell[   34154] = 32'h2561fc87;
    ram_cell[   34155] = 32'h25b47483;
    ram_cell[   34156] = 32'hc0bd3c75;
    ram_cell[   34157] = 32'h19f7b480;
    ram_cell[   34158] = 32'h1ea83746;
    ram_cell[   34159] = 32'ha02d775f;
    ram_cell[   34160] = 32'hc57a641a;
    ram_cell[   34161] = 32'h4f07c134;
    ram_cell[   34162] = 32'h94054615;
    ram_cell[   34163] = 32'hed0c5446;
    ram_cell[   34164] = 32'h15ccb680;
    ram_cell[   34165] = 32'h0bde1653;
    ram_cell[   34166] = 32'h9bb77a39;
    ram_cell[   34167] = 32'hd3fa7439;
    ram_cell[   34168] = 32'h1e098cda;
    ram_cell[   34169] = 32'h0333cde2;
    ram_cell[   34170] = 32'haffb0777;
    ram_cell[   34171] = 32'h414586f7;
    ram_cell[   34172] = 32'h16ed2ddd;
    ram_cell[   34173] = 32'h8886cb97;
    ram_cell[   34174] = 32'h18b107d5;
    ram_cell[   34175] = 32'he6bb3bbd;
    ram_cell[   34176] = 32'h3de0db2d;
    ram_cell[   34177] = 32'h144e0f0e;
    ram_cell[   34178] = 32'hccdf9c01;
    ram_cell[   34179] = 32'hf6e14f03;
    ram_cell[   34180] = 32'h2e2b8210;
    ram_cell[   34181] = 32'h8ed92832;
    ram_cell[   34182] = 32'h66b39a67;
    ram_cell[   34183] = 32'hb1e1246e;
    ram_cell[   34184] = 32'hcf8a9e9b;
    ram_cell[   34185] = 32'hb8652c94;
    ram_cell[   34186] = 32'h5d8e6807;
    ram_cell[   34187] = 32'h50c8418e;
    ram_cell[   34188] = 32'h93d9040b;
    ram_cell[   34189] = 32'h79f26c49;
    ram_cell[   34190] = 32'he42f1caf;
    ram_cell[   34191] = 32'h2780f945;
    ram_cell[   34192] = 32'h0421366e;
    ram_cell[   34193] = 32'hfc83e212;
    ram_cell[   34194] = 32'hc29506f7;
    ram_cell[   34195] = 32'h717157e1;
    ram_cell[   34196] = 32'h405e66c7;
    ram_cell[   34197] = 32'hc35f77aa;
    ram_cell[   34198] = 32'hcb35edd3;
    ram_cell[   34199] = 32'h33266a35;
    ram_cell[   34200] = 32'he7652147;
    ram_cell[   34201] = 32'h0efde0d2;
    ram_cell[   34202] = 32'h88425853;
    ram_cell[   34203] = 32'hf8729145;
    ram_cell[   34204] = 32'hcd715ca1;
    ram_cell[   34205] = 32'h14200c72;
    ram_cell[   34206] = 32'hc3e1dd1b;
    ram_cell[   34207] = 32'hfe1ea758;
    ram_cell[   34208] = 32'h9d34c154;
    ram_cell[   34209] = 32'h4d2ccdf2;
    ram_cell[   34210] = 32'h959eccee;
    ram_cell[   34211] = 32'h5ac0cabf;
    ram_cell[   34212] = 32'hb689fa7c;
    ram_cell[   34213] = 32'h89b0daeb;
    ram_cell[   34214] = 32'h06582a7f;
    ram_cell[   34215] = 32'hfa3d3b15;
    ram_cell[   34216] = 32'h442a3a4e;
    ram_cell[   34217] = 32'h2a74cbeb;
    ram_cell[   34218] = 32'hf97b4fb9;
    ram_cell[   34219] = 32'h6bd034e3;
    ram_cell[   34220] = 32'h855915f9;
    ram_cell[   34221] = 32'hddb07287;
    ram_cell[   34222] = 32'hb1b1a300;
    ram_cell[   34223] = 32'h9d1613e4;
    ram_cell[   34224] = 32'h69caee7d;
    ram_cell[   34225] = 32'he2da0253;
    ram_cell[   34226] = 32'hc741aeba;
    ram_cell[   34227] = 32'h4fa8b9b2;
    ram_cell[   34228] = 32'h96144783;
    ram_cell[   34229] = 32'h2caaa045;
    ram_cell[   34230] = 32'h85e4d5b5;
    ram_cell[   34231] = 32'hf2ceab00;
    ram_cell[   34232] = 32'h9b1549ed;
    ram_cell[   34233] = 32'haea9b304;
    ram_cell[   34234] = 32'h4907bbd4;
    ram_cell[   34235] = 32'h99ec0648;
    ram_cell[   34236] = 32'hb8d31e49;
    ram_cell[   34237] = 32'h488eba39;
    ram_cell[   34238] = 32'h739aa019;
    ram_cell[   34239] = 32'hf042d5e6;
    ram_cell[   34240] = 32'h478b3366;
    ram_cell[   34241] = 32'h3a05c1c5;
    ram_cell[   34242] = 32'h4a3bf396;
    ram_cell[   34243] = 32'h8e5f4c9d;
    ram_cell[   34244] = 32'h6cbb1fc2;
    ram_cell[   34245] = 32'hf9e7aed4;
    ram_cell[   34246] = 32'h91dd07c6;
    ram_cell[   34247] = 32'h1556794d;
    ram_cell[   34248] = 32'h37c04a41;
    ram_cell[   34249] = 32'h27925e6f;
    ram_cell[   34250] = 32'hfd7c75e9;
    ram_cell[   34251] = 32'hbbe46600;
    ram_cell[   34252] = 32'hcf943f22;
    ram_cell[   34253] = 32'h8239081b;
    ram_cell[   34254] = 32'ha5f8f238;
    ram_cell[   34255] = 32'h8ec967ae;
    ram_cell[   34256] = 32'h9ca72d83;
    ram_cell[   34257] = 32'h763f2f76;
    ram_cell[   34258] = 32'hb99ee5a3;
    ram_cell[   34259] = 32'h63001518;
    ram_cell[   34260] = 32'hfb128253;
    ram_cell[   34261] = 32'hf15944c3;
    ram_cell[   34262] = 32'hca6d9767;
    ram_cell[   34263] = 32'h49d12b50;
    ram_cell[   34264] = 32'h03b20309;
    ram_cell[   34265] = 32'h06b5c676;
    ram_cell[   34266] = 32'h0b9718b0;
    ram_cell[   34267] = 32'hd49b9052;
    ram_cell[   34268] = 32'h589596ea;
    ram_cell[   34269] = 32'hbc4a3a57;
    ram_cell[   34270] = 32'hebd27484;
    ram_cell[   34271] = 32'h8b79356c;
    ram_cell[   34272] = 32'hbe394cc0;
    ram_cell[   34273] = 32'h0c25c6a4;
    ram_cell[   34274] = 32'h87237cd3;
    ram_cell[   34275] = 32'h90624eab;
    ram_cell[   34276] = 32'h861050eb;
    ram_cell[   34277] = 32'h66d456c8;
    ram_cell[   34278] = 32'h6991bda8;
    ram_cell[   34279] = 32'hb334d568;
    ram_cell[   34280] = 32'hb0a0d41e;
    ram_cell[   34281] = 32'h210ffa98;
    ram_cell[   34282] = 32'h0ac6c7fd;
    ram_cell[   34283] = 32'hb168c326;
    ram_cell[   34284] = 32'h0b685cbf;
    ram_cell[   34285] = 32'h95bd7e49;
    ram_cell[   34286] = 32'h919b4d8b;
    ram_cell[   34287] = 32'hb67e85ed;
    ram_cell[   34288] = 32'hf37b06bf;
    ram_cell[   34289] = 32'h0d2990fd;
    ram_cell[   34290] = 32'h042809ea;
    ram_cell[   34291] = 32'hd7774530;
    ram_cell[   34292] = 32'hf2bb5d03;
    ram_cell[   34293] = 32'hdeaff997;
    ram_cell[   34294] = 32'h65fd4a50;
    ram_cell[   34295] = 32'h5f34004b;
    ram_cell[   34296] = 32'he95f8c99;
    ram_cell[   34297] = 32'he7bf9b1f;
    ram_cell[   34298] = 32'h0c2393cd;
    ram_cell[   34299] = 32'h4e79347b;
    ram_cell[   34300] = 32'h7a6aea50;
    ram_cell[   34301] = 32'h44d6aa6f;
    ram_cell[   34302] = 32'h3b5a4316;
    ram_cell[   34303] = 32'hec9525bc;
    ram_cell[   34304] = 32'h1fe543e0;
    ram_cell[   34305] = 32'he3e210ae;
    ram_cell[   34306] = 32'hc4f1aa32;
    ram_cell[   34307] = 32'h835bbf3a;
    ram_cell[   34308] = 32'h803e0702;
    ram_cell[   34309] = 32'h20dd235f;
    ram_cell[   34310] = 32'ha2554667;
    ram_cell[   34311] = 32'hc9929b34;
    ram_cell[   34312] = 32'h693637cd;
    ram_cell[   34313] = 32'h1d743644;
    ram_cell[   34314] = 32'h8e1ae530;
    ram_cell[   34315] = 32'hb4e66624;
    ram_cell[   34316] = 32'hb25132f5;
    ram_cell[   34317] = 32'hced03a54;
    ram_cell[   34318] = 32'h68b9967e;
    ram_cell[   34319] = 32'hff1a960e;
    ram_cell[   34320] = 32'h0eaff423;
    ram_cell[   34321] = 32'h354515cb;
    ram_cell[   34322] = 32'h477fdfbb;
    ram_cell[   34323] = 32'h44b41f7e;
    ram_cell[   34324] = 32'hd1bd7477;
    ram_cell[   34325] = 32'h4a959791;
    ram_cell[   34326] = 32'h1aa64bda;
    ram_cell[   34327] = 32'ha1522cca;
    ram_cell[   34328] = 32'hade5702c;
    ram_cell[   34329] = 32'h0ddab793;
    ram_cell[   34330] = 32'h897acb7c;
    ram_cell[   34331] = 32'he86da23e;
    ram_cell[   34332] = 32'h329d8a67;
    ram_cell[   34333] = 32'hd88f1fae;
    ram_cell[   34334] = 32'hbbe469cb;
    ram_cell[   34335] = 32'h7f8a2fa4;
    ram_cell[   34336] = 32'h24e48238;
    ram_cell[   34337] = 32'h5f036a46;
    ram_cell[   34338] = 32'hc727cc1e;
    ram_cell[   34339] = 32'h8e230f26;
    ram_cell[   34340] = 32'h89c29819;
    ram_cell[   34341] = 32'hab2682f9;
    ram_cell[   34342] = 32'h4b6ff956;
    ram_cell[   34343] = 32'h1854a7bd;
    ram_cell[   34344] = 32'h2a8e8f49;
    ram_cell[   34345] = 32'h11f06110;
    ram_cell[   34346] = 32'hfb349a38;
    ram_cell[   34347] = 32'hf14b0cc6;
    ram_cell[   34348] = 32'h602294db;
    ram_cell[   34349] = 32'hfe3ebb0d;
    ram_cell[   34350] = 32'h5b45a895;
    ram_cell[   34351] = 32'h8c683c7b;
    ram_cell[   34352] = 32'hbb3d03a0;
    ram_cell[   34353] = 32'ha7f295c4;
    ram_cell[   34354] = 32'h1296eafd;
    ram_cell[   34355] = 32'hf3e8d454;
    ram_cell[   34356] = 32'h869fdae3;
    ram_cell[   34357] = 32'hb2eb5fde;
    ram_cell[   34358] = 32'hcf32237b;
    ram_cell[   34359] = 32'hc646f0b1;
    ram_cell[   34360] = 32'h9fffcb3e;
    ram_cell[   34361] = 32'h25836682;
    ram_cell[   34362] = 32'ha85e83a6;
    ram_cell[   34363] = 32'h7c037ffe;
    ram_cell[   34364] = 32'h355ae20c;
    ram_cell[   34365] = 32'h9f7a8c6c;
    ram_cell[   34366] = 32'h8269d01f;
    ram_cell[   34367] = 32'h0531d7a0;
    ram_cell[   34368] = 32'hbabd27bd;
    ram_cell[   34369] = 32'hafe55ae6;
    ram_cell[   34370] = 32'hc40e1b6c;
    ram_cell[   34371] = 32'h5c3b0c8b;
    ram_cell[   34372] = 32'hb172d96c;
    ram_cell[   34373] = 32'h1473e1b2;
    ram_cell[   34374] = 32'h7a827597;
    ram_cell[   34375] = 32'hefb3f6bc;
    ram_cell[   34376] = 32'h381ba755;
    ram_cell[   34377] = 32'h0d8955a5;
    ram_cell[   34378] = 32'ha625f771;
    ram_cell[   34379] = 32'h2f6f5d66;
    ram_cell[   34380] = 32'hddd0c945;
    ram_cell[   34381] = 32'h55b81425;
    ram_cell[   34382] = 32'he4fe4cb1;
    ram_cell[   34383] = 32'h39eb1ded;
    ram_cell[   34384] = 32'h61c2ad83;
    ram_cell[   34385] = 32'hac158707;
    ram_cell[   34386] = 32'hce015c29;
    ram_cell[   34387] = 32'h2cd16509;
    ram_cell[   34388] = 32'hdb8bc3ad;
    ram_cell[   34389] = 32'h9a6fcf11;
    ram_cell[   34390] = 32'h556e3db3;
    ram_cell[   34391] = 32'h9295d10c;
    ram_cell[   34392] = 32'hb1121c02;
    ram_cell[   34393] = 32'h970906cb;
    ram_cell[   34394] = 32'hc85b4b7e;
    ram_cell[   34395] = 32'h14e06aad;
    ram_cell[   34396] = 32'h41abe416;
    ram_cell[   34397] = 32'h87185c12;
    ram_cell[   34398] = 32'h9a9d4086;
    ram_cell[   34399] = 32'h41174a30;
    ram_cell[   34400] = 32'h20d6c0e5;
    ram_cell[   34401] = 32'hb338d3f3;
    ram_cell[   34402] = 32'h23f13249;
    ram_cell[   34403] = 32'h00962f72;
    ram_cell[   34404] = 32'h164f2e99;
    ram_cell[   34405] = 32'ha97004a1;
    ram_cell[   34406] = 32'h7b2d67c0;
    ram_cell[   34407] = 32'h0f0c6817;
    ram_cell[   34408] = 32'h49163570;
    ram_cell[   34409] = 32'hbc154e09;
    ram_cell[   34410] = 32'h9af8e430;
    ram_cell[   34411] = 32'h891ddeb6;
    ram_cell[   34412] = 32'hb02a92b8;
    ram_cell[   34413] = 32'h7a347e4c;
    ram_cell[   34414] = 32'h0e92be94;
    ram_cell[   34415] = 32'h4d364ba4;
    ram_cell[   34416] = 32'h533314d2;
    ram_cell[   34417] = 32'h4fc03366;
    ram_cell[   34418] = 32'h32826789;
    ram_cell[   34419] = 32'h66efaf65;
    ram_cell[   34420] = 32'h86394750;
    ram_cell[   34421] = 32'hda8a32b0;
    ram_cell[   34422] = 32'h84ab9de8;
    ram_cell[   34423] = 32'h2ca1aecf;
    ram_cell[   34424] = 32'h6cc17b98;
    ram_cell[   34425] = 32'hf99263ec;
    ram_cell[   34426] = 32'h62708260;
    ram_cell[   34427] = 32'h098da670;
    ram_cell[   34428] = 32'h3e05d901;
    ram_cell[   34429] = 32'h0d1646e3;
    ram_cell[   34430] = 32'h9de0f514;
    ram_cell[   34431] = 32'h83aa9c92;
    ram_cell[   34432] = 32'heff3ea8d;
    ram_cell[   34433] = 32'h621ba73a;
    ram_cell[   34434] = 32'h7eb0162b;
    ram_cell[   34435] = 32'haf28ef15;
    ram_cell[   34436] = 32'h92414cb1;
    ram_cell[   34437] = 32'h2e9e0cdd;
    ram_cell[   34438] = 32'ha1b3065a;
    ram_cell[   34439] = 32'h4ea270af;
    ram_cell[   34440] = 32'h0826f4b2;
    ram_cell[   34441] = 32'h2c348eea;
    ram_cell[   34442] = 32'hcd268d15;
    ram_cell[   34443] = 32'h17de7b1f;
    ram_cell[   34444] = 32'ha8c52e7d;
    ram_cell[   34445] = 32'h9b32512f;
    ram_cell[   34446] = 32'hc8dd9248;
    ram_cell[   34447] = 32'h52c36ee6;
    ram_cell[   34448] = 32'he2691fc3;
    ram_cell[   34449] = 32'h2c096b6b;
    ram_cell[   34450] = 32'h00f4b14f;
    ram_cell[   34451] = 32'h53a2a80b;
    ram_cell[   34452] = 32'h388400b8;
    ram_cell[   34453] = 32'h2991e09e;
    ram_cell[   34454] = 32'hd0975746;
    ram_cell[   34455] = 32'h88e66060;
    ram_cell[   34456] = 32'hb45510e3;
    ram_cell[   34457] = 32'hcfe7a43c;
    ram_cell[   34458] = 32'h371dda9e;
    ram_cell[   34459] = 32'hc933d70e;
    ram_cell[   34460] = 32'h058a4908;
    ram_cell[   34461] = 32'h59a3e2c6;
    ram_cell[   34462] = 32'h40560002;
    ram_cell[   34463] = 32'hbb49f753;
    ram_cell[   34464] = 32'h37f93756;
    ram_cell[   34465] = 32'h9e5f090a;
    ram_cell[   34466] = 32'h15befc33;
    ram_cell[   34467] = 32'h30ff1cc3;
    ram_cell[   34468] = 32'he9789f55;
    ram_cell[   34469] = 32'hef213b35;
    ram_cell[   34470] = 32'ha1861d8c;
    ram_cell[   34471] = 32'h10004bb6;
    ram_cell[   34472] = 32'h4f7c3419;
    ram_cell[   34473] = 32'h417be782;
    ram_cell[   34474] = 32'hd7c134ac;
    ram_cell[   34475] = 32'h21086e23;
    ram_cell[   34476] = 32'h4d20b6f9;
    ram_cell[   34477] = 32'hcc2ce857;
    ram_cell[   34478] = 32'h6f38f851;
    ram_cell[   34479] = 32'h98a5a889;
    ram_cell[   34480] = 32'h98d47f93;
    ram_cell[   34481] = 32'h73fd1413;
    ram_cell[   34482] = 32'h067cceef;
    ram_cell[   34483] = 32'h613645f4;
    ram_cell[   34484] = 32'hf6816e64;
    ram_cell[   34485] = 32'h7d9e2b8a;
    ram_cell[   34486] = 32'h2d8a2f32;
    ram_cell[   34487] = 32'hb356e1c5;
    ram_cell[   34488] = 32'h225807dc;
    ram_cell[   34489] = 32'h8cb96f9c;
    ram_cell[   34490] = 32'h96b73e11;
    ram_cell[   34491] = 32'hb6de7e37;
    ram_cell[   34492] = 32'hff5383d1;
    ram_cell[   34493] = 32'h2c520444;
    ram_cell[   34494] = 32'heb7f79b6;
    ram_cell[   34495] = 32'hd6dc3769;
    ram_cell[   34496] = 32'h2205fe9c;
    ram_cell[   34497] = 32'h14f7818c;
    ram_cell[   34498] = 32'hce34742d;
    ram_cell[   34499] = 32'hce80e9b6;
    ram_cell[   34500] = 32'h4690bb89;
    ram_cell[   34501] = 32'h621f7d0b;
    ram_cell[   34502] = 32'hc6e27136;
    ram_cell[   34503] = 32'heaa38158;
    ram_cell[   34504] = 32'hcbcd839a;
    ram_cell[   34505] = 32'h2620dec0;
    ram_cell[   34506] = 32'ha0e20147;
    ram_cell[   34507] = 32'hc98f3d0e;
    ram_cell[   34508] = 32'h8b58bc75;
    ram_cell[   34509] = 32'hefa64bfa;
    ram_cell[   34510] = 32'h41ca4745;
    ram_cell[   34511] = 32'h566af639;
    ram_cell[   34512] = 32'ha5221257;
    ram_cell[   34513] = 32'hf4474ba0;
    ram_cell[   34514] = 32'h1dcb8eca;
    ram_cell[   34515] = 32'h0d0ea70f;
    ram_cell[   34516] = 32'hf421fe98;
    ram_cell[   34517] = 32'h9a6a2bc9;
    ram_cell[   34518] = 32'hfd242899;
    ram_cell[   34519] = 32'hbe0a5219;
    ram_cell[   34520] = 32'h85a38161;
    ram_cell[   34521] = 32'hee965082;
    ram_cell[   34522] = 32'h225ff75f;
    ram_cell[   34523] = 32'h5792bc7d;
    ram_cell[   34524] = 32'h197450fe;
    ram_cell[   34525] = 32'h4ade2c90;
    ram_cell[   34526] = 32'ha2ba5d8d;
    ram_cell[   34527] = 32'hc19b2f7e;
    ram_cell[   34528] = 32'h841b4c8f;
    ram_cell[   34529] = 32'h6c27e5c2;
    ram_cell[   34530] = 32'hcd352f4d;
    ram_cell[   34531] = 32'h92787a56;
    ram_cell[   34532] = 32'h4fda1b98;
    ram_cell[   34533] = 32'h6619a926;
    ram_cell[   34534] = 32'h2a4357fa;
    ram_cell[   34535] = 32'h4c6cd81d;
    ram_cell[   34536] = 32'he39b656d;
    ram_cell[   34537] = 32'h1d07a2c8;
    ram_cell[   34538] = 32'h03072e42;
    ram_cell[   34539] = 32'hf06eb77b;
    ram_cell[   34540] = 32'hc45d81c6;
    ram_cell[   34541] = 32'hf51dfe27;
    ram_cell[   34542] = 32'hc4993219;
    ram_cell[   34543] = 32'h446635f1;
    ram_cell[   34544] = 32'h580cc89b;
    ram_cell[   34545] = 32'h2a26845c;
    ram_cell[   34546] = 32'h79112e2c;
    ram_cell[   34547] = 32'hc1d9da09;
    ram_cell[   34548] = 32'hf63fa92f;
    ram_cell[   34549] = 32'hbf307421;
    ram_cell[   34550] = 32'h97d83991;
    ram_cell[   34551] = 32'he0920a48;
    ram_cell[   34552] = 32'h978b6a3e;
    ram_cell[   34553] = 32'h55e44677;
    ram_cell[   34554] = 32'had071475;
    ram_cell[   34555] = 32'ha82853a1;
    ram_cell[   34556] = 32'h1ead35cb;
    ram_cell[   34557] = 32'h39889ac1;
    ram_cell[   34558] = 32'hcbf0129e;
    ram_cell[   34559] = 32'h6fe16b47;
    ram_cell[   34560] = 32'hed4f2eeb;
    ram_cell[   34561] = 32'hfb4faf6c;
    ram_cell[   34562] = 32'hf3765b7d;
    ram_cell[   34563] = 32'hd6b1bf8f;
    ram_cell[   34564] = 32'hcb8b0f3e;
    ram_cell[   34565] = 32'hcf1145a0;
    ram_cell[   34566] = 32'h7f595558;
    ram_cell[   34567] = 32'h9780bc75;
    ram_cell[   34568] = 32'h848e043e;
    ram_cell[   34569] = 32'h9ff1f368;
    ram_cell[   34570] = 32'ha10f4772;
    ram_cell[   34571] = 32'h02d0bd54;
    ram_cell[   34572] = 32'h66dd8c85;
    ram_cell[   34573] = 32'hda2b3c36;
    ram_cell[   34574] = 32'h0faa62e1;
    ram_cell[   34575] = 32'hbe7fc7d0;
    ram_cell[   34576] = 32'hca7bd6b8;
    ram_cell[   34577] = 32'h61be81f0;
    ram_cell[   34578] = 32'h1f999788;
    ram_cell[   34579] = 32'ha16c3db9;
    ram_cell[   34580] = 32'h1c57d6da;
    ram_cell[   34581] = 32'h84401dd3;
    ram_cell[   34582] = 32'h3f205cb6;
    ram_cell[   34583] = 32'hfcf897ea;
    ram_cell[   34584] = 32'h7552d518;
    ram_cell[   34585] = 32'h425d49e0;
    ram_cell[   34586] = 32'h456254b8;
    ram_cell[   34587] = 32'h1339087e;
    ram_cell[   34588] = 32'h8b1adfe0;
    ram_cell[   34589] = 32'h43503fe4;
    ram_cell[   34590] = 32'h915f68e2;
    ram_cell[   34591] = 32'h2b0fa1cc;
    ram_cell[   34592] = 32'h77e5b91d;
    ram_cell[   34593] = 32'h23717bc9;
    ram_cell[   34594] = 32'h971b3877;
    ram_cell[   34595] = 32'h9a58c9c6;
    ram_cell[   34596] = 32'hf878e047;
    ram_cell[   34597] = 32'h6557322a;
    ram_cell[   34598] = 32'ha554c5bb;
    ram_cell[   34599] = 32'h66690ce6;
    ram_cell[   34600] = 32'h83a9011c;
    ram_cell[   34601] = 32'h6b3963e0;
    ram_cell[   34602] = 32'h141ad440;
    ram_cell[   34603] = 32'hf7b72275;
    ram_cell[   34604] = 32'h5ad4c668;
    ram_cell[   34605] = 32'h11fd8412;
    ram_cell[   34606] = 32'hb8c0d4cd;
    ram_cell[   34607] = 32'hc40e811a;
    ram_cell[   34608] = 32'h9d9b95cb;
    ram_cell[   34609] = 32'h3bbc9c2d;
    ram_cell[   34610] = 32'hc7caead3;
    ram_cell[   34611] = 32'h298c6790;
    ram_cell[   34612] = 32'h2bf48876;
    ram_cell[   34613] = 32'h433c5134;
    ram_cell[   34614] = 32'h7c325405;
    ram_cell[   34615] = 32'h6a5b6396;
    ram_cell[   34616] = 32'h19b61e04;
    ram_cell[   34617] = 32'h6310ea4e;
    ram_cell[   34618] = 32'h80028dbb;
    ram_cell[   34619] = 32'h8a3e0f27;
    ram_cell[   34620] = 32'hccff1933;
    ram_cell[   34621] = 32'ha0ab0243;
    ram_cell[   34622] = 32'hea8f3d13;
    ram_cell[   34623] = 32'h9e53fb06;
    ram_cell[   34624] = 32'h898baab0;
    ram_cell[   34625] = 32'hf9bd3f3a;
    ram_cell[   34626] = 32'hda380490;
    ram_cell[   34627] = 32'he3d24f8a;
    ram_cell[   34628] = 32'hf6b62392;
    ram_cell[   34629] = 32'h6b62164e;
    ram_cell[   34630] = 32'h584da46a;
    ram_cell[   34631] = 32'h2f1710cd;
    ram_cell[   34632] = 32'h345b48e9;
    ram_cell[   34633] = 32'hc80a0a13;
    ram_cell[   34634] = 32'h43861815;
    ram_cell[   34635] = 32'h7fc602b7;
    ram_cell[   34636] = 32'h540b4ade;
    ram_cell[   34637] = 32'haaa12bbf;
    ram_cell[   34638] = 32'h322568b2;
    ram_cell[   34639] = 32'h23d94091;
    ram_cell[   34640] = 32'hdff85ecf;
    ram_cell[   34641] = 32'ha3d56ca0;
    ram_cell[   34642] = 32'h7e7199ab;
    ram_cell[   34643] = 32'habb176cd;
    ram_cell[   34644] = 32'hf8cc8fe9;
    ram_cell[   34645] = 32'h3daec266;
    ram_cell[   34646] = 32'h5b28bdd4;
    ram_cell[   34647] = 32'hc4613258;
    ram_cell[   34648] = 32'hccecf418;
    ram_cell[   34649] = 32'h36c59aa1;
    ram_cell[   34650] = 32'h6f1af949;
    ram_cell[   34651] = 32'hb74d8634;
    ram_cell[   34652] = 32'h0e67c5d5;
    ram_cell[   34653] = 32'hb6b3f6b9;
    ram_cell[   34654] = 32'h83186def;
    ram_cell[   34655] = 32'h5c2f5a9f;
    ram_cell[   34656] = 32'hc4552a9b;
    ram_cell[   34657] = 32'h65f67431;
    ram_cell[   34658] = 32'haf5ca8e8;
    ram_cell[   34659] = 32'hb9a3d917;
    ram_cell[   34660] = 32'h8af7164b;
    ram_cell[   34661] = 32'h36d2a2f5;
    ram_cell[   34662] = 32'h5111efea;
    ram_cell[   34663] = 32'hb2d4c87b;
    ram_cell[   34664] = 32'h8a1f4610;
    ram_cell[   34665] = 32'h4fc5a2a1;
    ram_cell[   34666] = 32'h565981f1;
    ram_cell[   34667] = 32'h725c955a;
    ram_cell[   34668] = 32'h321db4e5;
    ram_cell[   34669] = 32'h23a3cb88;
    ram_cell[   34670] = 32'h9735bcdd;
    ram_cell[   34671] = 32'h30926528;
    ram_cell[   34672] = 32'h5bcd8559;
    ram_cell[   34673] = 32'h4f525d28;
    ram_cell[   34674] = 32'ha9ef4c16;
    ram_cell[   34675] = 32'hb00d6380;
    ram_cell[   34676] = 32'h6cf867f3;
    ram_cell[   34677] = 32'h302f0150;
    ram_cell[   34678] = 32'hb455b6b8;
    ram_cell[   34679] = 32'h1d5ab843;
    ram_cell[   34680] = 32'hd081c008;
    ram_cell[   34681] = 32'h799ae516;
    ram_cell[   34682] = 32'h9ee0ec27;
    ram_cell[   34683] = 32'h175618cd;
    ram_cell[   34684] = 32'he608b6e3;
    ram_cell[   34685] = 32'h15d16c42;
    ram_cell[   34686] = 32'hae26902e;
    ram_cell[   34687] = 32'h67371d7b;
    ram_cell[   34688] = 32'h03562583;
    ram_cell[   34689] = 32'h15b75772;
    ram_cell[   34690] = 32'hc6a9d5a0;
    ram_cell[   34691] = 32'hf6a8675c;
    ram_cell[   34692] = 32'h71d6c28c;
    ram_cell[   34693] = 32'hc56cb315;
    ram_cell[   34694] = 32'hda1c3857;
    ram_cell[   34695] = 32'h4cc87caf;
    ram_cell[   34696] = 32'h68fccd61;
    ram_cell[   34697] = 32'h39fdc614;
    ram_cell[   34698] = 32'h96684f39;
    ram_cell[   34699] = 32'hb90626db;
    ram_cell[   34700] = 32'he2ed5cba;
    ram_cell[   34701] = 32'hc5cde91e;
    ram_cell[   34702] = 32'h2646474a;
    ram_cell[   34703] = 32'h147daa44;
    ram_cell[   34704] = 32'hb62243a6;
    ram_cell[   34705] = 32'hb6351501;
    ram_cell[   34706] = 32'h388ca772;
    ram_cell[   34707] = 32'h36bb2af2;
    ram_cell[   34708] = 32'he78f7ba5;
    ram_cell[   34709] = 32'h6c2dbc46;
    ram_cell[   34710] = 32'hf1a54809;
    ram_cell[   34711] = 32'hba2d7e2b;
    ram_cell[   34712] = 32'hed30f3f0;
    ram_cell[   34713] = 32'h99b75b81;
    ram_cell[   34714] = 32'he6c26ba8;
    ram_cell[   34715] = 32'h02ec006b;
    ram_cell[   34716] = 32'h5efe98f2;
    ram_cell[   34717] = 32'h50e5c162;
    ram_cell[   34718] = 32'h43b6b394;
    ram_cell[   34719] = 32'h43a99fb6;
    ram_cell[   34720] = 32'h2eb47d5b;
    ram_cell[   34721] = 32'h0c1f28ee;
    ram_cell[   34722] = 32'h36b3ac2d;
    ram_cell[   34723] = 32'he3528059;
    ram_cell[   34724] = 32'ha099de5c;
    ram_cell[   34725] = 32'hbd6438b4;
    ram_cell[   34726] = 32'ha96ffffc;
    ram_cell[   34727] = 32'hf2713908;
    ram_cell[   34728] = 32'h723e62d1;
    ram_cell[   34729] = 32'h4c475c10;
    ram_cell[   34730] = 32'h556edc1e;
    ram_cell[   34731] = 32'hf4f41036;
    ram_cell[   34732] = 32'hc2c33af6;
    ram_cell[   34733] = 32'h9a654a77;
    ram_cell[   34734] = 32'h4edea3e0;
    ram_cell[   34735] = 32'h218dd1d2;
    ram_cell[   34736] = 32'h2085325b;
    ram_cell[   34737] = 32'h9d6772b3;
    ram_cell[   34738] = 32'hb1920585;
    ram_cell[   34739] = 32'ha0daa341;
    ram_cell[   34740] = 32'h43510168;
    ram_cell[   34741] = 32'h7059676e;
    ram_cell[   34742] = 32'h730f1a59;
    ram_cell[   34743] = 32'h2c72a592;
    ram_cell[   34744] = 32'h8b3e76d9;
    ram_cell[   34745] = 32'hffed8d68;
    ram_cell[   34746] = 32'h22c40b08;
    ram_cell[   34747] = 32'hc604b0a7;
    ram_cell[   34748] = 32'ha2e9c2be;
    ram_cell[   34749] = 32'h42d35c4c;
    ram_cell[   34750] = 32'hfe7a5e9a;
    ram_cell[   34751] = 32'h6d877a25;
    ram_cell[   34752] = 32'h7103215f;
    ram_cell[   34753] = 32'hdfb5854e;
    ram_cell[   34754] = 32'h8039beed;
    ram_cell[   34755] = 32'hc100aadd;
    ram_cell[   34756] = 32'hae850684;
    ram_cell[   34757] = 32'hc81f1e22;
    ram_cell[   34758] = 32'h01324c0c;
    ram_cell[   34759] = 32'hf79de52f;
    ram_cell[   34760] = 32'h98f010a2;
    ram_cell[   34761] = 32'hadd6cbc7;
    ram_cell[   34762] = 32'hea8de36b;
    ram_cell[   34763] = 32'hfe3fc967;
    ram_cell[   34764] = 32'hab708e1e;
    ram_cell[   34765] = 32'hac0ad3e5;
    ram_cell[   34766] = 32'h76e4c661;
    ram_cell[   34767] = 32'h03a8ddb2;
    ram_cell[   34768] = 32'h3a036046;
    ram_cell[   34769] = 32'h05af9d9e;
    ram_cell[   34770] = 32'hb035aca4;
    ram_cell[   34771] = 32'h593cb2fe;
    ram_cell[   34772] = 32'h976592ec;
    ram_cell[   34773] = 32'h0b1ada74;
    ram_cell[   34774] = 32'h3240543b;
    ram_cell[   34775] = 32'h93847aa5;
    ram_cell[   34776] = 32'h03f12971;
    ram_cell[   34777] = 32'h21a7b224;
    ram_cell[   34778] = 32'hd6daef6e;
    ram_cell[   34779] = 32'hc72dd424;
    ram_cell[   34780] = 32'h9a880d8e;
    ram_cell[   34781] = 32'h2eea35c1;
    ram_cell[   34782] = 32'h284e54f0;
    ram_cell[   34783] = 32'he7501f87;
    ram_cell[   34784] = 32'hda731fed;
    ram_cell[   34785] = 32'hd2a5d47a;
    ram_cell[   34786] = 32'he97c0210;
    ram_cell[   34787] = 32'h14825988;
    ram_cell[   34788] = 32'hb9c48b70;
    ram_cell[   34789] = 32'hd2c8ced1;
    ram_cell[   34790] = 32'haae6111d;
    ram_cell[   34791] = 32'hec3ad40b;
    ram_cell[   34792] = 32'h2b2e2063;
    ram_cell[   34793] = 32'hc5a779d9;
    ram_cell[   34794] = 32'h998ac361;
    ram_cell[   34795] = 32'hc66a7783;
    ram_cell[   34796] = 32'h839f25fe;
    ram_cell[   34797] = 32'hc4905995;
    ram_cell[   34798] = 32'hfd14f92e;
    ram_cell[   34799] = 32'h2d29ab64;
    ram_cell[   34800] = 32'hd112271c;
    ram_cell[   34801] = 32'hbd206890;
    ram_cell[   34802] = 32'h16f8488d;
    ram_cell[   34803] = 32'h2b8794f1;
    ram_cell[   34804] = 32'h6d0e9d1b;
    ram_cell[   34805] = 32'h53aff7c3;
    ram_cell[   34806] = 32'h0c50df3c;
    ram_cell[   34807] = 32'h42ec4911;
    ram_cell[   34808] = 32'hebcc4f51;
    ram_cell[   34809] = 32'h3a2e32a5;
    ram_cell[   34810] = 32'h20734cf9;
    ram_cell[   34811] = 32'h11cadefd;
    ram_cell[   34812] = 32'h50dfe963;
    ram_cell[   34813] = 32'h8c674444;
    ram_cell[   34814] = 32'hc5fd18d6;
    ram_cell[   34815] = 32'h6f64d9ce;
    ram_cell[   34816] = 32'h88687bc7;
    ram_cell[   34817] = 32'h4a2b5985;
    ram_cell[   34818] = 32'hb2c639b9;
    ram_cell[   34819] = 32'h2d3911b8;
    ram_cell[   34820] = 32'h76924f11;
    ram_cell[   34821] = 32'h2c5f2099;
    ram_cell[   34822] = 32'h4e1bf9df;
    ram_cell[   34823] = 32'hf08e2f37;
    ram_cell[   34824] = 32'h771b6d69;
    ram_cell[   34825] = 32'h3e5a711c;
    ram_cell[   34826] = 32'hc83c784c;
    ram_cell[   34827] = 32'hc396839e;
    ram_cell[   34828] = 32'h46a276d6;
    ram_cell[   34829] = 32'hb76bbc7b;
    ram_cell[   34830] = 32'hd426a245;
    ram_cell[   34831] = 32'h6c7615ab;
    ram_cell[   34832] = 32'h6cd94eb4;
    ram_cell[   34833] = 32'h81b6ea21;
    ram_cell[   34834] = 32'h2fd5f795;
    ram_cell[   34835] = 32'h19f50eee;
    ram_cell[   34836] = 32'hc83b098e;
    ram_cell[   34837] = 32'hf85dccb6;
    ram_cell[   34838] = 32'h980c83ab;
    ram_cell[   34839] = 32'h0f3ddf71;
    ram_cell[   34840] = 32'hf6f51ca9;
    ram_cell[   34841] = 32'hb761690b;
    ram_cell[   34842] = 32'hf1574544;
    ram_cell[   34843] = 32'h9c43aa33;
    ram_cell[   34844] = 32'h5f8effd2;
    ram_cell[   34845] = 32'h707fd40a;
    ram_cell[   34846] = 32'h45eb0596;
    ram_cell[   34847] = 32'h688e5fd0;
    ram_cell[   34848] = 32'h8cfc2435;
    ram_cell[   34849] = 32'h7fb8b921;
    ram_cell[   34850] = 32'h6cded6ea;
    ram_cell[   34851] = 32'h5f6e05ad;
    ram_cell[   34852] = 32'h79939714;
    ram_cell[   34853] = 32'h37442788;
    ram_cell[   34854] = 32'hdcdb0676;
    ram_cell[   34855] = 32'h1c11a618;
    ram_cell[   34856] = 32'h568b80b9;
    ram_cell[   34857] = 32'hb5175ca7;
    ram_cell[   34858] = 32'h11b13c09;
    ram_cell[   34859] = 32'haff0407a;
    ram_cell[   34860] = 32'h747360dd;
    ram_cell[   34861] = 32'h54265d30;
    ram_cell[   34862] = 32'hfa053d11;
    ram_cell[   34863] = 32'h08dc03bc;
    ram_cell[   34864] = 32'hab782a42;
    ram_cell[   34865] = 32'h8ed7e89f;
    ram_cell[   34866] = 32'h59765426;
    ram_cell[   34867] = 32'h4422a918;
    ram_cell[   34868] = 32'h81be347b;
    ram_cell[   34869] = 32'h42f600d9;
    ram_cell[   34870] = 32'hc609cbf7;
    ram_cell[   34871] = 32'hba664b49;
    ram_cell[   34872] = 32'h622c3a39;
    ram_cell[   34873] = 32'h8e4a014b;
    ram_cell[   34874] = 32'hde08643e;
    ram_cell[   34875] = 32'h5527abd7;
    ram_cell[   34876] = 32'h312b3b4d;
    ram_cell[   34877] = 32'h8382dd26;
    ram_cell[   34878] = 32'h89d38136;
    ram_cell[   34879] = 32'h0de7bfc7;
    ram_cell[   34880] = 32'h91e319be;
    ram_cell[   34881] = 32'h8a14c05a;
    ram_cell[   34882] = 32'h9d823125;
    ram_cell[   34883] = 32'h1be0b44e;
    ram_cell[   34884] = 32'h4b9f10df;
    ram_cell[   34885] = 32'h4921a837;
    ram_cell[   34886] = 32'hb72efa80;
    ram_cell[   34887] = 32'h3b87056c;
    ram_cell[   34888] = 32'ha92f7f88;
    ram_cell[   34889] = 32'hb3e22130;
    ram_cell[   34890] = 32'hb6877fd8;
    ram_cell[   34891] = 32'hcfd63e7d;
    ram_cell[   34892] = 32'h4cdcddf5;
    ram_cell[   34893] = 32'he814cf5e;
    ram_cell[   34894] = 32'h1ea1bf75;
    ram_cell[   34895] = 32'h59c2d89a;
    ram_cell[   34896] = 32'h254389e6;
    ram_cell[   34897] = 32'h05425077;
    ram_cell[   34898] = 32'h2dd14b34;
    ram_cell[   34899] = 32'h3d370db2;
    ram_cell[   34900] = 32'h14902b30;
    ram_cell[   34901] = 32'h6086b50b;
    ram_cell[   34902] = 32'h078f7c45;
    ram_cell[   34903] = 32'h64d26293;
    ram_cell[   34904] = 32'hf0acae6d;
    ram_cell[   34905] = 32'h89f41fc8;
    ram_cell[   34906] = 32'hcad29fcd;
    ram_cell[   34907] = 32'hd678bccf;
    ram_cell[   34908] = 32'hdbed5291;
    ram_cell[   34909] = 32'h7474ea0a;
    ram_cell[   34910] = 32'hf3ea38f5;
    ram_cell[   34911] = 32'h602bd437;
    ram_cell[   34912] = 32'hc7e8ebde;
    ram_cell[   34913] = 32'h93187552;
    ram_cell[   34914] = 32'had7a5d60;
    ram_cell[   34915] = 32'h96904d87;
    ram_cell[   34916] = 32'h9c17fdc3;
    ram_cell[   34917] = 32'h6a14c957;
    ram_cell[   34918] = 32'hc6ab2d06;
    ram_cell[   34919] = 32'h41847613;
    ram_cell[   34920] = 32'h24c461e1;
    ram_cell[   34921] = 32'hc187c153;
    ram_cell[   34922] = 32'hbef80915;
    ram_cell[   34923] = 32'h3d2215b2;
    ram_cell[   34924] = 32'h57d91ea2;
    ram_cell[   34925] = 32'hed6d3696;
    ram_cell[   34926] = 32'hdf91bb40;
    ram_cell[   34927] = 32'h71ecc08c;
    ram_cell[   34928] = 32'h1111d56e;
    ram_cell[   34929] = 32'h10a614d2;
    ram_cell[   34930] = 32'hddf5cd9e;
    ram_cell[   34931] = 32'h0aa61dce;
    ram_cell[   34932] = 32'h991b2779;
    ram_cell[   34933] = 32'h357b436f;
    ram_cell[   34934] = 32'h6a67d7f3;
    ram_cell[   34935] = 32'h2da62b5f;
    ram_cell[   34936] = 32'h3fc55598;
    ram_cell[   34937] = 32'h5dcc3ef3;
    ram_cell[   34938] = 32'ha87fa776;
    ram_cell[   34939] = 32'h20641d9e;
    ram_cell[   34940] = 32'hd76418cc;
    ram_cell[   34941] = 32'hd6aa14d5;
    ram_cell[   34942] = 32'h013698bd;
    ram_cell[   34943] = 32'hb9fc96d1;
    ram_cell[   34944] = 32'h7d7c21c9;
    ram_cell[   34945] = 32'ha6c89268;
    ram_cell[   34946] = 32'hd0b2d337;
    ram_cell[   34947] = 32'he33841b7;
    ram_cell[   34948] = 32'h9a4d887f;
    ram_cell[   34949] = 32'h82bb3827;
    ram_cell[   34950] = 32'h84d5b45e;
    ram_cell[   34951] = 32'h670ef34a;
    ram_cell[   34952] = 32'h82f04ac7;
    ram_cell[   34953] = 32'hd00d7ca1;
    ram_cell[   34954] = 32'h634c9455;
    ram_cell[   34955] = 32'h8184cca1;
    ram_cell[   34956] = 32'h039be3f1;
    ram_cell[   34957] = 32'hee7c2b59;
    ram_cell[   34958] = 32'h55e13f69;
    ram_cell[   34959] = 32'h7de8e97f;
    ram_cell[   34960] = 32'h0b264f5d;
    ram_cell[   34961] = 32'h6b1fc403;
    ram_cell[   34962] = 32'h759ac697;
    ram_cell[   34963] = 32'h3467ab6e;
    ram_cell[   34964] = 32'hb3e24b5b;
    ram_cell[   34965] = 32'h67e52204;
    ram_cell[   34966] = 32'h9d849458;
    ram_cell[   34967] = 32'h0633f1fb;
    ram_cell[   34968] = 32'h737918c7;
    ram_cell[   34969] = 32'hbd801a94;
    ram_cell[   34970] = 32'h6ef7db4b;
    ram_cell[   34971] = 32'h81817d73;
    ram_cell[   34972] = 32'hea3a6977;
    ram_cell[   34973] = 32'h39ab5ff0;
    ram_cell[   34974] = 32'hcf0b241d;
    ram_cell[   34975] = 32'h4ef9c005;
    ram_cell[   34976] = 32'h0dd8e985;
    ram_cell[   34977] = 32'hd6ae96db;
    ram_cell[   34978] = 32'hc1ffe9af;
    ram_cell[   34979] = 32'h31283d49;
    ram_cell[   34980] = 32'hb596a554;
    ram_cell[   34981] = 32'hdf4593da;
    ram_cell[   34982] = 32'heeb898d3;
    ram_cell[   34983] = 32'hafc8afad;
    ram_cell[   34984] = 32'hac70d3b6;
    ram_cell[   34985] = 32'h5bf0e909;
    ram_cell[   34986] = 32'h7b4414a3;
    ram_cell[   34987] = 32'ha66f7f93;
    ram_cell[   34988] = 32'h2caa64ab;
    ram_cell[   34989] = 32'hf5a32240;
    ram_cell[   34990] = 32'h09696288;
    ram_cell[   34991] = 32'h5e7880ca;
    ram_cell[   34992] = 32'h9059cb78;
    ram_cell[   34993] = 32'hb4ce8967;
    ram_cell[   34994] = 32'h48a4be1a;
    ram_cell[   34995] = 32'hced7d11b;
    ram_cell[   34996] = 32'h4d10d33a;
    ram_cell[   34997] = 32'hae29675c;
    ram_cell[   34998] = 32'hdd18196f;
    ram_cell[   34999] = 32'h0c52d2ea;
    ram_cell[   35000] = 32'h5cd14d7e;
    ram_cell[   35001] = 32'h7d8fa88c;
    ram_cell[   35002] = 32'h203460b6;
    ram_cell[   35003] = 32'h6c537733;
    ram_cell[   35004] = 32'he3a5b9cf;
    ram_cell[   35005] = 32'hdd686727;
    ram_cell[   35006] = 32'h741617a7;
    ram_cell[   35007] = 32'hfa603711;
    ram_cell[   35008] = 32'h7d6cafd8;
    ram_cell[   35009] = 32'h2813ea01;
    ram_cell[   35010] = 32'h2878913d;
    ram_cell[   35011] = 32'ha64cca12;
    ram_cell[   35012] = 32'h53929c84;
    ram_cell[   35013] = 32'h2da7bd29;
    ram_cell[   35014] = 32'hfb46807c;
    ram_cell[   35015] = 32'h1172bed6;
    ram_cell[   35016] = 32'hae1278b7;
    ram_cell[   35017] = 32'h06d0a251;
    ram_cell[   35018] = 32'h54c6c21c;
    ram_cell[   35019] = 32'h7182ea60;
    ram_cell[   35020] = 32'h9f2c27d9;
    ram_cell[   35021] = 32'h3b0985c8;
    ram_cell[   35022] = 32'h409c1e28;
    ram_cell[   35023] = 32'h6d70ada1;
    ram_cell[   35024] = 32'h7280a43c;
    ram_cell[   35025] = 32'h266a0e14;
    ram_cell[   35026] = 32'h9d9e267f;
    ram_cell[   35027] = 32'h78919e12;
    ram_cell[   35028] = 32'h26e0c68e;
    ram_cell[   35029] = 32'hed0bcee9;
    ram_cell[   35030] = 32'h9ebdd087;
    ram_cell[   35031] = 32'h95846034;
    ram_cell[   35032] = 32'he6ee8f23;
    ram_cell[   35033] = 32'h77ddb75d;
    ram_cell[   35034] = 32'h17df4448;
    ram_cell[   35035] = 32'hf6cf979c;
    ram_cell[   35036] = 32'h193a7d51;
    ram_cell[   35037] = 32'h8be854dc;
    ram_cell[   35038] = 32'hdc4b4148;
    ram_cell[   35039] = 32'h005a0e8a;
    ram_cell[   35040] = 32'h9d44e41f;
    ram_cell[   35041] = 32'h58833a4c;
    ram_cell[   35042] = 32'hf145fc0d;
    ram_cell[   35043] = 32'h516567c0;
    ram_cell[   35044] = 32'h49235a67;
    ram_cell[   35045] = 32'h2e1cefd9;
    ram_cell[   35046] = 32'hb0cd04ea;
    ram_cell[   35047] = 32'hce18ee85;
    ram_cell[   35048] = 32'hc650e0dd;
    ram_cell[   35049] = 32'h022a3ba5;
    ram_cell[   35050] = 32'h2bb2e6d1;
    ram_cell[   35051] = 32'h35a10222;
    ram_cell[   35052] = 32'h4b01ae84;
    ram_cell[   35053] = 32'h8be256cc;
    ram_cell[   35054] = 32'h3d86f337;
    ram_cell[   35055] = 32'h70447b76;
    ram_cell[   35056] = 32'h55e0cba1;
    ram_cell[   35057] = 32'h35a9000c;
    ram_cell[   35058] = 32'hed4ff0b3;
    ram_cell[   35059] = 32'h1a0ef279;
    ram_cell[   35060] = 32'h2b79d4c4;
    ram_cell[   35061] = 32'h72d47f03;
    ram_cell[   35062] = 32'he93b421c;
    ram_cell[   35063] = 32'h1cbeaed9;
    ram_cell[   35064] = 32'h43c181de;
    ram_cell[   35065] = 32'hc3162f5d;
    ram_cell[   35066] = 32'hafd69e30;
    ram_cell[   35067] = 32'h90717184;
    ram_cell[   35068] = 32'hc6e49b91;
    ram_cell[   35069] = 32'h3813a5db;
    ram_cell[   35070] = 32'h0fee6b48;
    ram_cell[   35071] = 32'h4c9d021d;
    ram_cell[   35072] = 32'h15bc262d;
    ram_cell[   35073] = 32'h291e2c12;
    ram_cell[   35074] = 32'h53afe5b0;
    ram_cell[   35075] = 32'ha5aac07b;
    ram_cell[   35076] = 32'h1f831a15;
    ram_cell[   35077] = 32'he6cc3069;
    ram_cell[   35078] = 32'h224d2472;
    ram_cell[   35079] = 32'h74774b1b;
    ram_cell[   35080] = 32'hd5e3e797;
    ram_cell[   35081] = 32'h07ed99a3;
    ram_cell[   35082] = 32'hdf1b2fce;
    ram_cell[   35083] = 32'ha5d56213;
    ram_cell[   35084] = 32'hc2dde083;
    ram_cell[   35085] = 32'hab638e4a;
    ram_cell[   35086] = 32'h0bb1da0c;
    ram_cell[   35087] = 32'h25ca4e16;
    ram_cell[   35088] = 32'h7b14ce0f;
    ram_cell[   35089] = 32'h8a7579ac;
    ram_cell[   35090] = 32'h6783b504;
    ram_cell[   35091] = 32'h5960a0be;
    ram_cell[   35092] = 32'h0ea64e66;
    ram_cell[   35093] = 32'h6971749b;
    ram_cell[   35094] = 32'h5f0bc8ce;
    ram_cell[   35095] = 32'h312b0cc0;
    ram_cell[   35096] = 32'hdc164495;
    ram_cell[   35097] = 32'h5cc35034;
    ram_cell[   35098] = 32'ha594e185;
    ram_cell[   35099] = 32'h465e76e5;
    ram_cell[   35100] = 32'h2bd8a3e0;
    ram_cell[   35101] = 32'h5dbf60f2;
    ram_cell[   35102] = 32'h64515c34;
    ram_cell[   35103] = 32'hd9f5c918;
    ram_cell[   35104] = 32'h2f72f2a1;
    ram_cell[   35105] = 32'h57f33f76;
    ram_cell[   35106] = 32'hfa881cb2;
    ram_cell[   35107] = 32'h559fbeee;
    ram_cell[   35108] = 32'h35829915;
    ram_cell[   35109] = 32'h4e2c4c91;
    ram_cell[   35110] = 32'h02c80002;
    ram_cell[   35111] = 32'h9766da9d;
    ram_cell[   35112] = 32'hd573eae7;
    ram_cell[   35113] = 32'h33687f83;
    ram_cell[   35114] = 32'h275b38c2;
    ram_cell[   35115] = 32'hf7f2dd27;
    ram_cell[   35116] = 32'hd10d50ac;
    ram_cell[   35117] = 32'hd3d98245;
    ram_cell[   35118] = 32'hce21248d;
    ram_cell[   35119] = 32'haae1cc0f;
    ram_cell[   35120] = 32'hb404290c;
    ram_cell[   35121] = 32'hd6b2e716;
    ram_cell[   35122] = 32'hd24c69ce;
    ram_cell[   35123] = 32'h60c66f60;
    ram_cell[   35124] = 32'h28948b1d;
    ram_cell[   35125] = 32'hf79504db;
    ram_cell[   35126] = 32'h3cc24069;
    ram_cell[   35127] = 32'hf83f030a;
    ram_cell[   35128] = 32'h754d64cb;
    ram_cell[   35129] = 32'h30f5960a;
    ram_cell[   35130] = 32'hc4902ca9;
    ram_cell[   35131] = 32'h2f3aeaf1;
    ram_cell[   35132] = 32'h38732cc4;
    ram_cell[   35133] = 32'h725266bc;
    ram_cell[   35134] = 32'hbad273fd;
    ram_cell[   35135] = 32'h27a13d78;
    ram_cell[   35136] = 32'h48558669;
    ram_cell[   35137] = 32'ha93d5eb2;
    ram_cell[   35138] = 32'h46023c3b;
    ram_cell[   35139] = 32'h0898197a;
    ram_cell[   35140] = 32'h8d208525;
    ram_cell[   35141] = 32'h0f294490;
    ram_cell[   35142] = 32'h6fa00827;
    ram_cell[   35143] = 32'h53875eae;
    ram_cell[   35144] = 32'hd09e5a4a;
    ram_cell[   35145] = 32'h56191f8a;
    ram_cell[   35146] = 32'h2e9ba88e;
    ram_cell[   35147] = 32'h3aa47272;
    ram_cell[   35148] = 32'h11508d02;
    ram_cell[   35149] = 32'h7dc406dc;
    ram_cell[   35150] = 32'h72c62529;
    ram_cell[   35151] = 32'h25d8812d;
    ram_cell[   35152] = 32'h5e5b7463;
    ram_cell[   35153] = 32'h42110372;
    ram_cell[   35154] = 32'h4dd5b4cd;
    ram_cell[   35155] = 32'hf151523f;
    ram_cell[   35156] = 32'h37686a80;
    ram_cell[   35157] = 32'hde4602ac;
    ram_cell[   35158] = 32'h2da55eef;
    ram_cell[   35159] = 32'h4e057783;
    ram_cell[   35160] = 32'hc8cf0532;
    ram_cell[   35161] = 32'had14be76;
    ram_cell[   35162] = 32'h0054b6a6;
    ram_cell[   35163] = 32'h89bcc6cc;
    ram_cell[   35164] = 32'hb246b8de;
    ram_cell[   35165] = 32'hddc80954;
    ram_cell[   35166] = 32'hc1a30081;
    ram_cell[   35167] = 32'h0b2635cb;
    ram_cell[   35168] = 32'hb5deb4b6;
    ram_cell[   35169] = 32'h441d95c1;
    ram_cell[   35170] = 32'h61789347;
    ram_cell[   35171] = 32'h12f09b32;
    ram_cell[   35172] = 32'h04a6aa5d;
    ram_cell[   35173] = 32'h81564aef;
    ram_cell[   35174] = 32'hc64eded7;
    ram_cell[   35175] = 32'h50840f5a;
    ram_cell[   35176] = 32'he1cab531;
    ram_cell[   35177] = 32'hc18c7679;
    ram_cell[   35178] = 32'h018330ed;
    ram_cell[   35179] = 32'ha1df5fd6;
    ram_cell[   35180] = 32'h7660b3aa;
    ram_cell[   35181] = 32'h90f87ab0;
    ram_cell[   35182] = 32'hbbffdcac;
    ram_cell[   35183] = 32'h80b868b6;
    ram_cell[   35184] = 32'h1de387ab;
    ram_cell[   35185] = 32'h0647d087;
    ram_cell[   35186] = 32'h8cba6bd6;
    ram_cell[   35187] = 32'h74dd7582;
    ram_cell[   35188] = 32'hdbbd4c48;
    ram_cell[   35189] = 32'h64a820f7;
    ram_cell[   35190] = 32'hf3b41097;
    ram_cell[   35191] = 32'he9bb3b9b;
    ram_cell[   35192] = 32'h34b7586a;
    ram_cell[   35193] = 32'hda67cef1;
    ram_cell[   35194] = 32'he363e403;
    ram_cell[   35195] = 32'h242022f2;
    ram_cell[   35196] = 32'hc8fd342f;
    ram_cell[   35197] = 32'h1b5c9f11;
    ram_cell[   35198] = 32'h8628279e;
    ram_cell[   35199] = 32'h0dea8a87;
    ram_cell[   35200] = 32'h36d0f735;
    ram_cell[   35201] = 32'h4749b96d;
    ram_cell[   35202] = 32'hf49d9abd;
    ram_cell[   35203] = 32'h5d1bb595;
    ram_cell[   35204] = 32'h9451b99c;
    ram_cell[   35205] = 32'hc1bf2c6a;
    ram_cell[   35206] = 32'h08e27671;
    ram_cell[   35207] = 32'h4a551deb;
    ram_cell[   35208] = 32'h9d2e3448;
    ram_cell[   35209] = 32'ha1072b9d;
    ram_cell[   35210] = 32'h029f3b26;
    ram_cell[   35211] = 32'h52902da5;
    ram_cell[   35212] = 32'he022e58f;
    ram_cell[   35213] = 32'h67dc0768;
    ram_cell[   35214] = 32'hbd19e64e;
    ram_cell[   35215] = 32'h2ee261ca;
    ram_cell[   35216] = 32'hfc2fd0fb;
    ram_cell[   35217] = 32'ha8397fc1;
    ram_cell[   35218] = 32'h5a30f936;
    ram_cell[   35219] = 32'h41d62e92;
    ram_cell[   35220] = 32'h045f9772;
    ram_cell[   35221] = 32'h66a4b9ac;
    ram_cell[   35222] = 32'hf9116ff6;
    ram_cell[   35223] = 32'h33017008;
    ram_cell[   35224] = 32'h38de1f1a;
    ram_cell[   35225] = 32'h3cfa30e7;
    ram_cell[   35226] = 32'h290467f3;
    ram_cell[   35227] = 32'hf5ad6598;
    ram_cell[   35228] = 32'h1e6da350;
    ram_cell[   35229] = 32'hb77023f1;
    ram_cell[   35230] = 32'hd27c38ec;
    ram_cell[   35231] = 32'hd8bb37cd;
    ram_cell[   35232] = 32'he2b17276;
    ram_cell[   35233] = 32'hf9d53b03;
    ram_cell[   35234] = 32'h30f001c4;
    ram_cell[   35235] = 32'h12e92675;
    ram_cell[   35236] = 32'ha118be95;
    ram_cell[   35237] = 32'hb7eca55d;
    ram_cell[   35238] = 32'h22cb63ec;
    ram_cell[   35239] = 32'h3ec1241a;
    ram_cell[   35240] = 32'hfc1ccf2c;
    ram_cell[   35241] = 32'h73b0bf9f;
    ram_cell[   35242] = 32'h436fc077;
    ram_cell[   35243] = 32'h4b699ae4;
    ram_cell[   35244] = 32'h8fd85db0;
    ram_cell[   35245] = 32'h41b3c750;
    ram_cell[   35246] = 32'h04b3dd4c;
    ram_cell[   35247] = 32'hf124184c;
    ram_cell[   35248] = 32'h3f7bc703;
    ram_cell[   35249] = 32'hafa42060;
    ram_cell[   35250] = 32'h26eec12b;
    ram_cell[   35251] = 32'h209a0365;
    ram_cell[   35252] = 32'h874e5471;
    ram_cell[   35253] = 32'habd931ea;
    ram_cell[   35254] = 32'h68254110;
    ram_cell[   35255] = 32'h140b1263;
    ram_cell[   35256] = 32'h5cb805b6;
    ram_cell[   35257] = 32'h5ec30c68;
    ram_cell[   35258] = 32'hcd28975d;
    ram_cell[   35259] = 32'h87697b5d;
    ram_cell[   35260] = 32'h28bd8c4a;
    ram_cell[   35261] = 32'h6dff9a99;
    ram_cell[   35262] = 32'h63194ea0;
    ram_cell[   35263] = 32'hac536f03;
    ram_cell[   35264] = 32'h12a61185;
    ram_cell[   35265] = 32'h8902772c;
    ram_cell[   35266] = 32'h19aecc8e;
    ram_cell[   35267] = 32'h99954d59;
    ram_cell[   35268] = 32'hb73bd7f4;
    ram_cell[   35269] = 32'h8a9cc290;
    ram_cell[   35270] = 32'hc883f8ff;
    ram_cell[   35271] = 32'h54aa6f30;
    ram_cell[   35272] = 32'h71f41c14;
    ram_cell[   35273] = 32'h1cfdb86f;
    ram_cell[   35274] = 32'he3eb09ae;
    ram_cell[   35275] = 32'hb3d128eb;
    ram_cell[   35276] = 32'hd8f1a135;
    ram_cell[   35277] = 32'h62d9d94c;
    ram_cell[   35278] = 32'h5b7da4fa;
    ram_cell[   35279] = 32'hd32c6657;
    ram_cell[   35280] = 32'he2513843;
    ram_cell[   35281] = 32'h9f13c46d;
    ram_cell[   35282] = 32'hce8adbb7;
    ram_cell[   35283] = 32'h1ddbffe6;
    ram_cell[   35284] = 32'h137106ec;
    ram_cell[   35285] = 32'hd6c537cf;
    ram_cell[   35286] = 32'h68be2b58;
    ram_cell[   35287] = 32'h6cafd919;
    ram_cell[   35288] = 32'h01c881d1;
    ram_cell[   35289] = 32'hc0733fbf;
    ram_cell[   35290] = 32'hf836f669;
    ram_cell[   35291] = 32'h1fc37e62;
    ram_cell[   35292] = 32'h19d5a551;
    ram_cell[   35293] = 32'hb5eff935;
    ram_cell[   35294] = 32'he07e6eff;
    ram_cell[   35295] = 32'h8cb5384a;
    ram_cell[   35296] = 32'h1c500b18;
    ram_cell[   35297] = 32'h52901c13;
    ram_cell[   35298] = 32'hc6efb111;
    ram_cell[   35299] = 32'h82218c04;
    ram_cell[   35300] = 32'ha3066c4f;
    ram_cell[   35301] = 32'h723b4e5c;
    ram_cell[   35302] = 32'h75e467ba;
    ram_cell[   35303] = 32'h829bfa69;
    ram_cell[   35304] = 32'hcb4d0866;
    ram_cell[   35305] = 32'h31979cd5;
    ram_cell[   35306] = 32'h39e61ab3;
    ram_cell[   35307] = 32'hd18a64bf;
    ram_cell[   35308] = 32'h5e0b1f83;
    ram_cell[   35309] = 32'hc01a63d2;
    ram_cell[   35310] = 32'h9ed23304;
    ram_cell[   35311] = 32'hccf3d002;
    ram_cell[   35312] = 32'h7fc7ed76;
    ram_cell[   35313] = 32'h48115dab;
    ram_cell[   35314] = 32'h6c780b7a;
    ram_cell[   35315] = 32'h4f5bef42;
    ram_cell[   35316] = 32'h48969983;
    ram_cell[   35317] = 32'h5101b062;
    ram_cell[   35318] = 32'hd5fcad37;
    ram_cell[   35319] = 32'he96cd06f;
    ram_cell[   35320] = 32'hd356166f;
    ram_cell[   35321] = 32'hb01b47e1;
    ram_cell[   35322] = 32'h0b5ae5cc;
    ram_cell[   35323] = 32'h06b0edb6;
    ram_cell[   35324] = 32'h66975db8;
    ram_cell[   35325] = 32'hf1f327b9;
    ram_cell[   35326] = 32'h30f4188c;
    ram_cell[   35327] = 32'hc161df58;
    ram_cell[   35328] = 32'hdddbb9c3;
    ram_cell[   35329] = 32'h35efde13;
    ram_cell[   35330] = 32'h9a7d7da7;
    ram_cell[   35331] = 32'h048355d5;
    ram_cell[   35332] = 32'h27aaed4e;
    ram_cell[   35333] = 32'hdd5972bd;
    ram_cell[   35334] = 32'h1f96130f;
    ram_cell[   35335] = 32'h99a95746;
    ram_cell[   35336] = 32'h0ee58c32;
    ram_cell[   35337] = 32'h3b4bfc70;
    ram_cell[   35338] = 32'h2e960bb9;
    ram_cell[   35339] = 32'h421b7950;
    ram_cell[   35340] = 32'h46e7a5b1;
    ram_cell[   35341] = 32'hd17c0a3a;
    ram_cell[   35342] = 32'h8cba5b00;
    ram_cell[   35343] = 32'hf6f7092d;
    ram_cell[   35344] = 32'h905e38dc;
    ram_cell[   35345] = 32'h5ec7869e;
    ram_cell[   35346] = 32'hb8f2a012;
    ram_cell[   35347] = 32'hfcf35c12;
    ram_cell[   35348] = 32'h8b3bd51e;
    ram_cell[   35349] = 32'hd203a46b;
    ram_cell[   35350] = 32'h8a6dbc9c;
    ram_cell[   35351] = 32'h098668a9;
    ram_cell[   35352] = 32'h48c64df7;
    ram_cell[   35353] = 32'h2d4a5da2;
    ram_cell[   35354] = 32'he47ff20a;
    ram_cell[   35355] = 32'h0750cda7;
    ram_cell[   35356] = 32'hedb79b5b;
    ram_cell[   35357] = 32'h6d2148c9;
    ram_cell[   35358] = 32'hacc0372d;
    ram_cell[   35359] = 32'h8641198b;
    ram_cell[   35360] = 32'h6072ce79;
    ram_cell[   35361] = 32'h108bcac8;
    ram_cell[   35362] = 32'hd763d7b1;
    ram_cell[   35363] = 32'hb6c80d00;
    ram_cell[   35364] = 32'hd64ba17e;
    ram_cell[   35365] = 32'h87cb8de9;
    ram_cell[   35366] = 32'h7fecfdc0;
    ram_cell[   35367] = 32'h3a20863f;
    ram_cell[   35368] = 32'h2977b651;
    ram_cell[   35369] = 32'h32c5e42e;
    ram_cell[   35370] = 32'h6ae6238a;
    ram_cell[   35371] = 32'h8ae962a1;
    ram_cell[   35372] = 32'h7ca50148;
    ram_cell[   35373] = 32'h34cb44c7;
    ram_cell[   35374] = 32'h835dcf98;
    ram_cell[   35375] = 32'h213b3831;
    ram_cell[   35376] = 32'h66766a55;
    ram_cell[   35377] = 32'h398d7f06;
    ram_cell[   35378] = 32'hfe86ddad;
    ram_cell[   35379] = 32'hef8412bb;
    ram_cell[   35380] = 32'h00a97a2e;
    ram_cell[   35381] = 32'h0f5bd06d;
    ram_cell[   35382] = 32'hcc0d11fd;
    ram_cell[   35383] = 32'h8b8d03ae;
    ram_cell[   35384] = 32'h2c7a421c;
    ram_cell[   35385] = 32'h9034f913;
    ram_cell[   35386] = 32'h4cfb2f7e;
    ram_cell[   35387] = 32'hd5c581f7;
    ram_cell[   35388] = 32'hdb7a1f55;
    ram_cell[   35389] = 32'h559a609b;
    ram_cell[   35390] = 32'hf59ef15b;
    ram_cell[   35391] = 32'h5da03008;
    ram_cell[   35392] = 32'h8d2251dc;
    ram_cell[   35393] = 32'h83d14089;
    ram_cell[   35394] = 32'h64d7d5d9;
    ram_cell[   35395] = 32'h858f386c;
    ram_cell[   35396] = 32'hfc45d0a5;
    ram_cell[   35397] = 32'h6fc31d9f;
    ram_cell[   35398] = 32'hd7ec0b22;
    ram_cell[   35399] = 32'h68185a40;
    ram_cell[   35400] = 32'h96a61348;
    ram_cell[   35401] = 32'hc39991f7;
    ram_cell[   35402] = 32'h9d5aefac;
    ram_cell[   35403] = 32'h281ca26a;
    ram_cell[   35404] = 32'h43099dcb;
    ram_cell[   35405] = 32'h4b0bfab8;
    ram_cell[   35406] = 32'h32180b24;
    ram_cell[   35407] = 32'h7dab3c63;
    ram_cell[   35408] = 32'hc60e7707;
    ram_cell[   35409] = 32'h85f75099;
    ram_cell[   35410] = 32'h508eb3ae;
    ram_cell[   35411] = 32'h3e90b64e;
    ram_cell[   35412] = 32'hf6b6b254;
    ram_cell[   35413] = 32'he0cb6169;
    ram_cell[   35414] = 32'h876c6bbb;
    ram_cell[   35415] = 32'h6ead61d1;
    ram_cell[   35416] = 32'h6a2e16f7;
    ram_cell[   35417] = 32'hcc3a9f7f;
    ram_cell[   35418] = 32'h890bf314;
    ram_cell[   35419] = 32'hb2735dd0;
    ram_cell[   35420] = 32'he4198603;
    ram_cell[   35421] = 32'h96467959;
    ram_cell[   35422] = 32'hb4b77461;
    ram_cell[   35423] = 32'ha6fe3aaa;
    ram_cell[   35424] = 32'h9ef18085;
    ram_cell[   35425] = 32'h1071d7eb;
    ram_cell[   35426] = 32'hab8d97be;
    ram_cell[   35427] = 32'hc80153f4;
    ram_cell[   35428] = 32'h3e2bd3d3;
    ram_cell[   35429] = 32'h2f4ea5c2;
    ram_cell[   35430] = 32'he068165c;
    ram_cell[   35431] = 32'h37e2a4a4;
    ram_cell[   35432] = 32'hf335ebac;
    ram_cell[   35433] = 32'h80dbab63;
    ram_cell[   35434] = 32'h28dc183f;
    ram_cell[   35435] = 32'h2dd056b8;
    ram_cell[   35436] = 32'h682337ed;
    ram_cell[   35437] = 32'hf6cb6d60;
    ram_cell[   35438] = 32'h534e47de;
    ram_cell[   35439] = 32'hf1b9c855;
    ram_cell[   35440] = 32'h90c81216;
    ram_cell[   35441] = 32'hc9b3aba1;
    ram_cell[   35442] = 32'h1aedcce9;
    ram_cell[   35443] = 32'he7ed5757;
    ram_cell[   35444] = 32'h42b08052;
    ram_cell[   35445] = 32'h68e70799;
    ram_cell[   35446] = 32'hf142a928;
    ram_cell[   35447] = 32'h8c1c76d8;
    ram_cell[   35448] = 32'h0fe9a410;
    ram_cell[   35449] = 32'h964d5e56;
    ram_cell[   35450] = 32'hdca054f0;
    ram_cell[   35451] = 32'hbad80bfb;
    ram_cell[   35452] = 32'h85b89696;
    ram_cell[   35453] = 32'h2688569f;
    ram_cell[   35454] = 32'h6d85da37;
    ram_cell[   35455] = 32'h308ed3f3;
    ram_cell[   35456] = 32'h08befb61;
    ram_cell[   35457] = 32'h86820be7;
    ram_cell[   35458] = 32'hb7624593;
    ram_cell[   35459] = 32'h63ea7c95;
    ram_cell[   35460] = 32'hfdf2ceed;
    ram_cell[   35461] = 32'h387a4882;
    ram_cell[   35462] = 32'h4c38f544;
    ram_cell[   35463] = 32'hf05c4809;
    ram_cell[   35464] = 32'h8cb9ee8b;
    ram_cell[   35465] = 32'h027b10b6;
    ram_cell[   35466] = 32'h6a610d23;
    ram_cell[   35467] = 32'h101182fe;
    ram_cell[   35468] = 32'h95d65a5e;
    ram_cell[   35469] = 32'hf57cf21f;
    ram_cell[   35470] = 32'h96c1a107;
    ram_cell[   35471] = 32'hfbf3c116;
    ram_cell[   35472] = 32'h0226f7c6;
    ram_cell[   35473] = 32'h8adcdef9;
    ram_cell[   35474] = 32'h22e2545b;
    ram_cell[   35475] = 32'h740eaa48;
    ram_cell[   35476] = 32'h23bf9a0d;
    ram_cell[   35477] = 32'hcef5c880;
    ram_cell[   35478] = 32'hb25e26b1;
    ram_cell[   35479] = 32'h387b2983;
    ram_cell[   35480] = 32'h752e3086;
    ram_cell[   35481] = 32'hbeb73737;
    ram_cell[   35482] = 32'h98e914ea;
    ram_cell[   35483] = 32'haf85213a;
    ram_cell[   35484] = 32'h29b4ff56;
    ram_cell[   35485] = 32'h88cf2114;
    ram_cell[   35486] = 32'ha8e7c72f;
    ram_cell[   35487] = 32'h8c41938c;
    ram_cell[   35488] = 32'h731f0118;
    ram_cell[   35489] = 32'h86ebbf21;
    ram_cell[   35490] = 32'hc062d1c2;
    ram_cell[   35491] = 32'h406eba5c;
    ram_cell[   35492] = 32'h3ecad8ea;
    ram_cell[   35493] = 32'h32b9c30e;
    ram_cell[   35494] = 32'h98d36d4c;
    ram_cell[   35495] = 32'h30a370a3;
    ram_cell[   35496] = 32'h69397aeb;
    ram_cell[   35497] = 32'h0dc2da26;
    ram_cell[   35498] = 32'ha9f6bd7d;
    ram_cell[   35499] = 32'h79cc871d;
    ram_cell[   35500] = 32'hcba32708;
    ram_cell[   35501] = 32'h29333a9e;
    ram_cell[   35502] = 32'h7e01f279;
    ram_cell[   35503] = 32'hb30dd929;
    ram_cell[   35504] = 32'h1c2e844d;
    ram_cell[   35505] = 32'h258e49ea;
    ram_cell[   35506] = 32'h10f3d264;
    ram_cell[   35507] = 32'h57ee8451;
    ram_cell[   35508] = 32'h07391244;
    ram_cell[   35509] = 32'hb2477e38;
    ram_cell[   35510] = 32'h7577a861;
    ram_cell[   35511] = 32'h140f720b;
    ram_cell[   35512] = 32'ha430e58c;
    ram_cell[   35513] = 32'h8b1390d6;
    ram_cell[   35514] = 32'h2fc5557b;
    ram_cell[   35515] = 32'h5d86a668;
    ram_cell[   35516] = 32'h65514b4e;
    ram_cell[   35517] = 32'h25dd7b1d;
    ram_cell[   35518] = 32'hab6a3d95;
    ram_cell[   35519] = 32'h27ae0f91;
    ram_cell[   35520] = 32'h977e90a0;
    ram_cell[   35521] = 32'hdc2dbc96;
    ram_cell[   35522] = 32'h6734ca58;
    ram_cell[   35523] = 32'h7077e274;
    ram_cell[   35524] = 32'ha89321c8;
    ram_cell[   35525] = 32'h0693e7df;
    ram_cell[   35526] = 32'h9340de57;
    ram_cell[   35527] = 32'haa274b08;
    ram_cell[   35528] = 32'h765bc37d;
    ram_cell[   35529] = 32'h6e8e8cd6;
    ram_cell[   35530] = 32'h6bdeb054;
    ram_cell[   35531] = 32'h3d1e6ab8;
    ram_cell[   35532] = 32'h742da448;
    ram_cell[   35533] = 32'haf998bac;
    ram_cell[   35534] = 32'h1eb0dd47;
    ram_cell[   35535] = 32'h2251f01b;
    ram_cell[   35536] = 32'h94051ef8;
    ram_cell[   35537] = 32'hfca26069;
    ram_cell[   35538] = 32'hc8f3bf01;
    ram_cell[   35539] = 32'hf60c0860;
    ram_cell[   35540] = 32'hc196d79a;
    ram_cell[   35541] = 32'hb43718be;
    ram_cell[   35542] = 32'h5bc4c66a;
    ram_cell[   35543] = 32'hef24396d;
    ram_cell[   35544] = 32'he438db70;
    ram_cell[   35545] = 32'h77bd6d4a;
    ram_cell[   35546] = 32'hf65e2f4a;
    ram_cell[   35547] = 32'h9c9b162e;
    ram_cell[   35548] = 32'h222be4c6;
    ram_cell[   35549] = 32'h1354c671;
    ram_cell[   35550] = 32'h2d1a37dd;
    ram_cell[   35551] = 32'h3862f397;
    ram_cell[   35552] = 32'h25499fa6;
    ram_cell[   35553] = 32'hffbe0b1c;
    ram_cell[   35554] = 32'hb4a80a17;
    ram_cell[   35555] = 32'h096beb23;
    ram_cell[   35556] = 32'had5e0764;
    ram_cell[   35557] = 32'h450a4280;
    ram_cell[   35558] = 32'hadafa1d9;
    ram_cell[   35559] = 32'h8f82f07c;
    ram_cell[   35560] = 32'he7a233ae;
    ram_cell[   35561] = 32'h12312d18;
    ram_cell[   35562] = 32'h777fef98;
    ram_cell[   35563] = 32'h315d77f5;
    ram_cell[   35564] = 32'h3eaced01;
    ram_cell[   35565] = 32'h753d0b16;
    ram_cell[   35566] = 32'h3e8971e7;
    ram_cell[   35567] = 32'hd9d26aa8;
    ram_cell[   35568] = 32'h4976abe4;
    ram_cell[   35569] = 32'h9709bd6c;
    ram_cell[   35570] = 32'hcf8a54ed;
    ram_cell[   35571] = 32'hfb31fd78;
    ram_cell[   35572] = 32'h8661aabe;
    ram_cell[   35573] = 32'hc6ef6de6;
    ram_cell[   35574] = 32'h3a4e5082;
    ram_cell[   35575] = 32'h5b83b5ef;
    ram_cell[   35576] = 32'hfe8c5a6c;
    ram_cell[   35577] = 32'h3b6c8fbb;
    ram_cell[   35578] = 32'haa8eae70;
    ram_cell[   35579] = 32'hb3191f56;
    ram_cell[   35580] = 32'h03374b32;
    ram_cell[   35581] = 32'hcdf08435;
    ram_cell[   35582] = 32'ha34d8d91;
    ram_cell[   35583] = 32'h68e5326f;
    ram_cell[   35584] = 32'h65f54229;
    ram_cell[   35585] = 32'h4fa307fc;
    ram_cell[   35586] = 32'hcd6ce499;
    ram_cell[   35587] = 32'hf52a4886;
    ram_cell[   35588] = 32'h64de8a54;
    ram_cell[   35589] = 32'hdb4487bf;
    ram_cell[   35590] = 32'h9ad35b02;
    ram_cell[   35591] = 32'h86e4c002;
    ram_cell[   35592] = 32'h9ecfc234;
    ram_cell[   35593] = 32'hbd8bf6cd;
    ram_cell[   35594] = 32'h5e201faf;
    ram_cell[   35595] = 32'h576925cc;
    ram_cell[   35596] = 32'h9706fad0;
    ram_cell[   35597] = 32'hb3b6f4da;
    ram_cell[   35598] = 32'h26810d0f;
    ram_cell[   35599] = 32'h979474b0;
    ram_cell[   35600] = 32'hff7ed148;
    ram_cell[   35601] = 32'h08f094a7;
    ram_cell[   35602] = 32'h87489845;
    ram_cell[   35603] = 32'h476872b0;
    ram_cell[   35604] = 32'h38366615;
    ram_cell[   35605] = 32'hecfaf43b;
    ram_cell[   35606] = 32'hff3be517;
    ram_cell[   35607] = 32'h3fad3c06;
    ram_cell[   35608] = 32'h9d52017b;
    ram_cell[   35609] = 32'h9ed1f6a6;
    ram_cell[   35610] = 32'hc566146b;
    ram_cell[   35611] = 32'h567d578f;
    ram_cell[   35612] = 32'h065c945f;
    ram_cell[   35613] = 32'h41661b00;
    ram_cell[   35614] = 32'h0846b0f3;
    ram_cell[   35615] = 32'he80847e5;
    ram_cell[   35616] = 32'h583f11d8;
    ram_cell[   35617] = 32'he2a1464e;
    ram_cell[   35618] = 32'h520e6783;
    ram_cell[   35619] = 32'h14bdc0c9;
    ram_cell[   35620] = 32'h015a76a1;
    ram_cell[   35621] = 32'h204b32db;
    ram_cell[   35622] = 32'hb0810c4a;
    ram_cell[   35623] = 32'he9042c3c;
    ram_cell[   35624] = 32'hd151f185;
    ram_cell[   35625] = 32'hef4af0b1;
    ram_cell[   35626] = 32'h04a78de4;
    ram_cell[   35627] = 32'h4f44403b;
    ram_cell[   35628] = 32'h2d8f6e1a;
    ram_cell[   35629] = 32'h34d9f6ad;
    ram_cell[   35630] = 32'h091479b5;
    ram_cell[   35631] = 32'h53f3111c;
    ram_cell[   35632] = 32'hde0dbac5;
    ram_cell[   35633] = 32'h71812d79;
    ram_cell[   35634] = 32'hd275160e;
    ram_cell[   35635] = 32'h8b817dcf;
    ram_cell[   35636] = 32'h5d11cfd2;
    ram_cell[   35637] = 32'h0540425a;
    ram_cell[   35638] = 32'hc0615603;
    ram_cell[   35639] = 32'h743539f5;
    ram_cell[   35640] = 32'ha9bba282;
    ram_cell[   35641] = 32'ha53ee2ef;
    ram_cell[   35642] = 32'he2dd5a19;
    ram_cell[   35643] = 32'ha6fda69b;
    ram_cell[   35644] = 32'h36ae2ace;
    ram_cell[   35645] = 32'h718bb94e;
    ram_cell[   35646] = 32'hd3125d83;
    ram_cell[   35647] = 32'h07e7e62e;
    ram_cell[   35648] = 32'ha606f3ba;
    ram_cell[   35649] = 32'hf90c0557;
    ram_cell[   35650] = 32'h6f6d19df;
    ram_cell[   35651] = 32'h31584150;
    ram_cell[   35652] = 32'hd1bfe464;
    ram_cell[   35653] = 32'h2b2321f6;
    ram_cell[   35654] = 32'hc33fa81b;
    ram_cell[   35655] = 32'h4441d49b;
    ram_cell[   35656] = 32'hd7500781;
    ram_cell[   35657] = 32'hddc93ab4;
    ram_cell[   35658] = 32'h53f3df57;
    ram_cell[   35659] = 32'hac591432;
    ram_cell[   35660] = 32'hb3b1d7f6;
    ram_cell[   35661] = 32'h00c296b8;
    ram_cell[   35662] = 32'h1f42f355;
    ram_cell[   35663] = 32'he1281569;
    ram_cell[   35664] = 32'hf0a8c48d;
    ram_cell[   35665] = 32'hbf002de8;
    ram_cell[   35666] = 32'h8bb420df;
    ram_cell[   35667] = 32'hd8eee141;
    ram_cell[   35668] = 32'ha6783a06;
    ram_cell[   35669] = 32'h199303a1;
    ram_cell[   35670] = 32'he4bbfceb;
    ram_cell[   35671] = 32'hb310c28a;
    ram_cell[   35672] = 32'h0b6e9579;
    ram_cell[   35673] = 32'h2753039b;
    ram_cell[   35674] = 32'h82ac129e;
    ram_cell[   35675] = 32'h21b6acf6;
    ram_cell[   35676] = 32'hcfcced7d;
    ram_cell[   35677] = 32'hd0d5eeff;
    ram_cell[   35678] = 32'h6c376895;
    ram_cell[   35679] = 32'h923234f3;
    ram_cell[   35680] = 32'ha28d7c3e;
    ram_cell[   35681] = 32'hefba0f46;
    ram_cell[   35682] = 32'h5a56f239;
    ram_cell[   35683] = 32'h63e25c09;
    ram_cell[   35684] = 32'h3485f29e;
    ram_cell[   35685] = 32'ha4cdbe02;
    ram_cell[   35686] = 32'h6ff32993;
    ram_cell[   35687] = 32'hd210dc7f;
    ram_cell[   35688] = 32'hb040bf3b;
    ram_cell[   35689] = 32'h864f6a5e;
    ram_cell[   35690] = 32'hff251307;
    ram_cell[   35691] = 32'hb976f0f7;
    ram_cell[   35692] = 32'ha69fe5ff;
    ram_cell[   35693] = 32'hc11348ba;
    ram_cell[   35694] = 32'h9a0befa3;
    ram_cell[   35695] = 32'hf42769c8;
    ram_cell[   35696] = 32'hc92048c8;
    ram_cell[   35697] = 32'h82f43d29;
    ram_cell[   35698] = 32'h55660c28;
    ram_cell[   35699] = 32'h96ebbc3b;
    ram_cell[   35700] = 32'h39cf1ed3;
    ram_cell[   35701] = 32'hf82c26eb;
    ram_cell[   35702] = 32'h8c5ac234;
    ram_cell[   35703] = 32'h08f8d9ed;
    ram_cell[   35704] = 32'h617c99cf;
    ram_cell[   35705] = 32'hef7753bb;
    ram_cell[   35706] = 32'h6ce3fe56;
    ram_cell[   35707] = 32'he35ee0a6;
    ram_cell[   35708] = 32'h1b257496;
    ram_cell[   35709] = 32'h7eb4236e;
    ram_cell[   35710] = 32'h95ac0946;
    ram_cell[   35711] = 32'he84e8d7e;
    ram_cell[   35712] = 32'h64e065d0;
    ram_cell[   35713] = 32'hfb8086a1;
    ram_cell[   35714] = 32'h606cace6;
    ram_cell[   35715] = 32'h9cc7949d;
    ram_cell[   35716] = 32'h76756e34;
    ram_cell[   35717] = 32'hf02caa73;
    ram_cell[   35718] = 32'h214fb364;
    ram_cell[   35719] = 32'hbbf48876;
    ram_cell[   35720] = 32'h552e097c;
    ram_cell[   35721] = 32'h95c11cd1;
    ram_cell[   35722] = 32'h7342f9cf;
    ram_cell[   35723] = 32'h75badd3b;
    ram_cell[   35724] = 32'hb6e84c78;
    ram_cell[   35725] = 32'h37a064e9;
    ram_cell[   35726] = 32'h9d7b7945;
    ram_cell[   35727] = 32'heebea205;
    ram_cell[   35728] = 32'h65c9336a;
    ram_cell[   35729] = 32'h800b47ef;
    ram_cell[   35730] = 32'hbab117a4;
    ram_cell[   35731] = 32'h6821b787;
    ram_cell[   35732] = 32'h250c1989;
    ram_cell[   35733] = 32'h7abc4d15;
    ram_cell[   35734] = 32'h285ad394;
    ram_cell[   35735] = 32'h621d6ec6;
    ram_cell[   35736] = 32'he21e450a;
    ram_cell[   35737] = 32'hffbeab66;
    ram_cell[   35738] = 32'h7028d300;
    ram_cell[   35739] = 32'h576090fc;
    ram_cell[   35740] = 32'hf8b8f82e;
    ram_cell[   35741] = 32'h8d5ee4e4;
    ram_cell[   35742] = 32'h84016454;
    ram_cell[   35743] = 32'hdbc0d333;
    ram_cell[   35744] = 32'h3ab014db;
    ram_cell[   35745] = 32'hcf5cd11b;
    ram_cell[   35746] = 32'h5a8fc292;
    ram_cell[   35747] = 32'h41dd25e6;
    ram_cell[   35748] = 32'hf9a8bdc1;
    ram_cell[   35749] = 32'h88120da8;
    ram_cell[   35750] = 32'h7e41c2b6;
    ram_cell[   35751] = 32'h25b7172f;
    ram_cell[   35752] = 32'hb3d56cb4;
    ram_cell[   35753] = 32'h7f75c9fd;
    ram_cell[   35754] = 32'h1d04ac23;
    ram_cell[   35755] = 32'h38aa6abd;
    ram_cell[   35756] = 32'hdf25749e;
    ram_cell[   35757] = 32'h70bedf2c;
    ram_cell[   35758] = 32'hfc6fd22e;
    ram_cell[   35759] = 32'he9ddaa14;
    ram_cell[   35760] = 32'h4fd1a144;
    ram_cell[   35761] = 32'h97ff72c3;
    ram_cell[   35762] = 32'h57fbb354;
    ram_cell[   35763] = 32'h12e8e053;
    ram_cell[   35764] = 32'h1c18a9da;
    ram_cell[   35765] = 32'h50d9b7bc;
    ram_cell[   35766] = 32'ha96128dc;
    ram_cell[   35767] = 32'h9e2e732b;
    ram_cell[   35768] = 32'hb29a32d4;
    ram_cell[   35769] = 32'h88436ba9;
    ram_cell[   35770] = 32'he829b0f3;
    ram_cell[   35771] = 32'hc2bbccb3;
    ram_cell[   35772] = 32'h12562eba;
    ram_cell[   35773] = 32'h4741b2db;
    ram_cell[   35774] = 32'hd8813af2;
    ram_cell[   35775] = 32'h5958b296;
    ram_cell[   35776] = 32'h49091f99;
    ram_cell[   35777] = 32'hb6617f02;
    ram_cell[   35778] = 32'h7c03ba85;
    ram_cell[   35779] = 32'hbabdd14b;
    ram_cell[   35780] = 32'hc202377b;
    ram_cell[   35781] = 32'h897f41c6;
    ram_cell[   35782] = 32'h24026f9b;
    ram_cell[   35783] = 32'h2a0e5640;
    ram_cell[   35784] = 32'hec4009fc;
    ram_cell[   35785] = 32'hf88dc212;
    ram_cell[   35786] = 32'h3381ed40;
    ram_cell[   35787] = 32'h51f9e7d4;
    ram_cell[   35788] = 32'hfa0795e7;
    ram_cell[   35789] = 32'h496d2a9d;
    ram_cell[   35790] = 32'h5f5b8081;
    ram_cell[   35791] = 32'hf54a2ba2;
    ram_cell[   35792] = 32'he4213211;
    ram_cell[   35793] = 32'hdc6ceea9;
    ram_cell[   35794] = 32'h4f09642d;
    ram_cell[   35795] = 32'h74ed99f3;
    ram_cell[   35796] = 32'h5cf9b54b;
    ram_cell[   35797] = 32'h382007a1;
    ram_cell[   35798] = 32'h9040c842;
    ram_cell[   35799] = 32'hc37c3022;
    ram_cell[   35800] = 32'hdfb51a9f;
    ram_cell[   35801] = 32'h5f856bdb;
    ram_cell[   35802] = 32'h0f9f73de;
    ram_cell[   35803] = 32'h483e58e7;
    ram_cell[   35804] = 32'hd4e9f8a6;
    ram_cell[   35805] = 32'h1be72aa4;
    ram_cell[   35806] = 32'h60d952c2;
    ram_cell[   35807] = 32'h7f063e65;
    ram_cell[   35808] = 32'hdb4bf11f;
    ram_cell[   35809] = 32'h46545e38;
    ram_cell[   35810] = 32'hba03b97b;
    ram_cell[   35811] = 32'h2dbb9351;
    ram_cell[   35812] = 32'h58df4cf2;
    ram_cell[   35813] = 32'h52a2b4e5;
    ram_cell[   35814] = 32'hea633aa8;
    ram_cell[   35815] = 32'hbd8a2e11;
    ram_cell[   35816] = 32'hdd07c7dc;
    ram_cell[   35817] = 32'h155e0ded;
    ram_cell[   35818] = 32'hbc7fb041;
    ram_cell[   35819] = 32'he1e530f9;
    ram_cell[   35820] = 32'ha795419e;
    ram_cell[   35821] = 32'he10d40c8;
    ram_cell[   35822] = 32'hdde76234;
    ram_cell[   35823] = 32'ha2254365;
    ram_cell[   35824] = 32'hc756810c;
    ram_cell[   35825] = 32'h64d5532e;
    ram_cell[   35826] = 32'h84ed2ac2;
    ram_cell[   35827] = 32'h41cd131d;
    ram_cell[   35828] = 32'hd25a6ca2;
    ram_cell[   35829] = 32'h4da68f8e;
    ram_cell[   35830] = 32'h93a04d26;
    ram_cell[   35831] = 32'h21451657;
    ram_cell[   35832] = 32'h968cdde7;
    ram_cell[   35833] = 32'hb9fb3743;
    ram_cell[   35834] = 32'h82fdbbdb;
    ram_cell[   35835] = 32'hb4072712;
    ram_cell[   35836] = 32'h2495445b;
    ram_cell[   35837] = 32'hd7ad8125;
    ram_cell[   35838] = 32'h1fb07ef7;
    ram_cell[   35839] = 32'h872ec8d3;
    ram_cell[   35840] = 32'h0b7636ca;
    ram_cell[   35841] = 32'h50b4a568;
    ram_cell[   35842] = 32'haf5b0798;
    ram_cell[   35843] = 32'hf10eaec5;
    ram_cell[   35844] = 32'hbc7b4daf;
    ram_cell[   35845] = 32'hfc8f8873;
    ram_cell[   35846] = 32'hf29285b5;
    ram_cell[   35847] = 32'h0f011ec5;
    ram_cell[   35848] = 32'h7c1ce9dd;
    ram_cell[   35849] = 32'h55f909cd;
    ram_cell[   35850] = 32'h5828cc0f;
    ram_cell[   35851] = 32'hb4970947;
    ram_cell[   35852] = 32'hd4b8d56a;
    ram_cell[   35853] = 32'heb3e53dc;
    ram_cell[   35854] = 32'h818e39e8;
    ram_cell[   35855] = 32'hd92ac098;
    ram_cell[   35856] = 32'h06fd58f7;
    ram_cell[   35857] = 32'hc25c4c7a;
    ram_cell[   35858] = 32'hd91f1c05;
    ram_cell[   35859] = 32'h0895573a;
    ram_cell[   35860] = 32'h59fcd5e7;
    ram_cell[   35861] = 32'hc0224f9d;
    ram_cell[   35862] = 32'he630f832;
    ram_cell[   35863] = 32'h2d9ba919;
    ram_cell[   35864] = 32'h665d26ad;
    ram_cell[   35865] = 32'h49e7a5b3;
    ram_cell[   35866] = 32'ha648924d;
    ram_cell[   35867] = 32'hb75aa6ae;
    ram_cell[   35868] = 32'h18c92a30;
    ram_cell[   35869] = 32'h2bd3bc98;
    ram_cell[   35870] = 32'he67dc91c;
    ram_cell[   35871] = 32'h830b4aa4;
    ram_cell[   35872] = 32'ha6e23a50;
    ram_cell[   35873] = 32'hf962b715;
    ram_cell[   35874] = 32'h78ada1ca;
    ram_cell[   35875] = 32'he3f5cb1a;
    ram_cell[   35876] = 32'hf8d2cbc1;
    ram_cell[   35877] = 32'h7aa0543c;
    ram_cell[   35878] = 32'h4bbf11c7;
    ram_cell[   35879] = 32'hf13145e1;
    ram_cell[   35880] = 32'hed0d5bfb;
    ram_cell[   35881] = 32'h7ffbedf7;
    ram_cell[   35882] = 32'h155df809;
    ram_cell[   35883] = 32'h1b0e3680;
    ram_cell[   35884] = 32'h1ad3777c;
    ram_cell[   35885] = 32'h51db9c43;
    ram_cell[   35886] = 32'h98e85a02;
    ram_cell[   35887] = 32'h2f03fb87;
    ram_cell[   35888] = 32'hb7fa2b4b;
    ram_cell[   35889] = 32'hf889d2f3;
    ram_cell[   35890] = 32'he8a91788;
    ram_cell[   35891] = 32'h08e16aa4;
    ram_cell[   35892] = 32'h124dbb47;
    ram_cell[   35893] = 32'h0a0276a1;
    ram_cell[   35894] = 32'h13ec6078;
    ram_cell[   35895] = 32'h351a1d42;
    ram_cell[   35896] = 32'h8656b395;
    ram_cell[   35897] = 32'h01e87b44;
    ram_cell[   35898] = 32'hf4f08e62;
    ram_cell[   35899] = 32'h25085108;
    ram_cell[   35900] = 32'hc8f4f897;
    ram_cell[   35901] = 32'hb0cd8fbb;
    ram_cell[   35902] = 32'h0433019c;
    ram_cell[   35903] = 32'h6614364a;
    ram_cell[   35904] = 32'h5906f17b;
    ram_cell[   35905] = 32'h52c8624d;
    ram_cell[   35906] = 32'hd9a5a380;
    ram_cell[   35907] = 32'h47f2519c;
    ram_cell[   35908] = 32'hfaba209b;
    ram_cell[   35909] = 32'h333ff53b;
    ram_cell[   35910] = 32'h791dac11;
    ram_cell[   35911] = 32'h8b13ee8d;
    ram_cell[   35912] = 32'ha0d879e0;
    ram_cell[   35913] = 32'h99b4e089;
    ram_cell[   35914] = 32'h9f38dd20;
    ram_cell[   35915] = 32'hacc4a5b5;
    ram_cell[   35916] = 32'h96dfc258;
    ram_cell[   35917] = 32'h6650d7c6;
    ram_cell[   35918] = 32'h59836f50;
    ram_cell[   35919] = 32'h6c9acb96;
    ram_cell[   35920] = 32'h4baaaeb7;
    ram_cell[   35921] = 32'h1dde056c;
    ram_cell[   35922] = 32'h54844e14;
    ram_cell[   35923] = 32'h463384cc;
    ram_cell[   35924] = 32'hc866c49e;
    ram_cell[   35925] = 32'h3baf67b9;
    ram_cell[   35926] = 32'h72c623b9;
    ram_cell[   35927] = 32'he318daa0;
    ram_cell[   35928] = 32'h5fc5f45e;
    ram_cell[   35929] = 32'h8fecb71e;
    ram_cell[   35930] = 32'h5393337b;
    ram_cell[   35931] = 32'he8d68914;
    ram_cell[   35932] = 32'hac2c78a6;
    ram_cell[   35933] = 32'hb0b2b99b;
    ram_cell[   35934] = 32'h14b6348a;
    ram_cell[   35935] = 32'hd4f235aa;
    ram_cell[   35936] = 32'h7847f08c;
    ram_cell[   35937] = 32'h2f0a606d;
    ram_cell[   35938] = 32'hf09d1d9c;
    ram_cell[   35939] = 32'h230ed927;
    ram_cell[   35940] = 32'h9820122b;
    ram_cell[   35941] = 32'h51b89deb;
    ram_cell[   35942] = 32'h1d427950;
    ram_cell[   35943] = 32'hbdc7b9eb;
    ram_cell[   35944] = 32'h98f4b2e5;
    ram_cell[   35945] = 32'h404172a5;
    ram_cell[   35946] = 32'h9ebcea87;
    ram_cell[   35947] = 32'hba9feef8;
    ram_cell[   35948] = 32'h7f9a4adb;
    ram_cell[   35949] = 32'hff734b77;
    ram_cell[   35950] = 32'h38f1e07e;
    ram_cell[   35951] = 32'h0b3c27a3;
    ram_cell[   35952] = 32'h80b3dec2;
    ram_cell[   35953] = 32'h81dd05b2;
    ram_cell[   35954] = 32'hbee05b1f;
    ram_cell[   35955] = 32'hbdf5c3fa;
    ram_cell[   35956] = 32'h9447ea2a;
    ram_cell[   35957] = 32'h6ebc7448;
    ram_cell[   35958] = 32'h3e3b4ffd;
    ram_cell[   35959] = 32'h27ef1116;
    ram_cell[   35960] = 32'h64b27ddd;
    ram_cell[   35961] = 32'h4c1bc918;
    ram_cell[   35962] = 32'hbd9a8ff1;
    ram_cell[   35963] = 32'hdddf9835;
    ram_cell[   35964] = 32'h2e00851c;
    ram_cell[   35965] = 32'hbbf7f226;
    ram_cell[   35966] = 32'hf8666f1e;
    ram_cell[   35967] = 32'h444dc961;
    ram_cell[   35968] = 32'h447bfa02;
    ram_cell[   35969] = 32'h0839736e;
    ram_cell[   35970] = 32'h37002e62;
    ram_cell[   35971] = 32'hc99c7611;
    ram_cell[   35972] = 32'h7a0b93d0;
    ram_cell[   35973] = 32'h1b2b7d0b;
    ram_cell[   35974] = 32'hcd89e732;
    ram_cell[   35975] = 32'hd1e30060;
    ram_cell[   35976] = 32'h79c96090;
    ram_cell[   35977] = 32'hf55790ff;
    ram_cell[   35978] = 32'hcc805a2c;
    ram_cell[   35979] = 32'h758110ea;
    ram_cell[   35980] = 32'h43f7a8f7;
    ram_cell[   35981] = 32'h749e7397;
    ram_cell[   35982] = 32'h9146b966;
    ram_cell[   35983] = 32'h96a30d43;
    ram_cell[   35984] = 32'h12c6130d;
    ram_cell[   35985] = 32'h11e68ef0;
    ram_cell[   35986] = 32'hd57c1c76;
    ram_cell[   35987] = 32'hda62ba0f;
    ram_cell[   35988] = 32'h090bab41;
    ram_cell[   35989] = 32'hca2c1824;
    ram_cell[   35990] = 32'hd5d48354;
    ram_cell[   35991] = 32'hbeed38e0;
    ram_cell[   35992] = 32'h8e8e4f88;
    ram_cell[   35993] = 32'ha63168a3;
    ram_cell[   35994] = 32'he065e329;
    ram_cell[   35995] = 32'h855081eb;
    ram_cell[   35996] = 32'h19a0aaf1;
    ram_cell[   35997] = 32'h23b8fc5f;
    ram_cell[   35998] = 32'hc522a73c;
    ram_cell[   35999] = 32'h533143e2;
    ram_cell[   36000] = 32'h25a08403;
    ram_cell[   36001] = 32'hb428a363;
    ram_cell[   36002] = 32'hc4eb77a4;
    ram_cell[   36003] = 32'h2cac8875;
    ram_cell[   36004] = 32'hd43cb669;
    ram_cell[   36005] = 32'hbf83cc83;
    ram_cell[   36006] = 32'hbef7152d;
    ram_cell[   36007] = 32'hf0cf6c3f;
    ram_cell[   36008] = 32'h14f5d94a;
    ram_cell[   36009] = 32'h120db304;
    ram_cell[   36010] = 32'hd5b814a4;
    ram_cell[   36011] = 32'h36fccb4d;
    ram_cell[   36012] = 32'h107c8f1f;
    ram_cell[   36013] = 32'h6ea8e411;
    ram_cell[   36014] = 32'hfbd62dec;
    ram_cell[   36015] = 32'h8d937ffa;
    ram_cell[   36016] = 32'h329c90bc;
    ram_cell[   36017] = 32'haffe7bf8;
    ram_cell[   36018] = 32'h8c465ae6;
    ram_cell[   36019] = 32'hc046bf50;
    ram_cell[   36020] = 32'h15d7e6d9;
    ram_cell[   36021] = 32'hff42e27f;
    ram_cell[   36022] = 32'hb1f9f756;
    ram_cell[   36023] = 32'hf9e24b3c;
    ram_cell[   36024] = 32'hc04d21d0;
    ram_cell[   36025] = 32'h178e90aa;
    ram_cell[   36026] = 32'h3da2e737;
    ram_cell[   36027] = 32'h2b7bc84e;
    ram_cell[   36028] = 32'h8c4fb0ae;
    ram_cell[   36029] = 32'h46695771;
    ram_cell[   36030] = 32'hf2c1e962;
    ram_cell[   36031] = 32'h8fe7bd10;
    ram_cell[   36032] = 32'h5e6a3c4e;
    ram_cell[   36033] = 32'h87eabb1e;
    ram_cell[   36034] = 32'hd855d7fd;
    ram_cell[   36035] = 32'hb745f9c4;
    ram_cell[   36036] = 32'he0af08ab;
    ram_cell[   36037] = 32'h0b7596d8;
    ram_cell[   36038] = 32'hb320be7d;
    ram_cell[   36039] = 32'h19eb7876;
    ram_cell[   36040] = 32'ha84e6183;
    ram_cell[   36041] = 32'hbe9db4bf;
    ram_cell[   36042] = 32'h13c08322;
    ram_cell[   36043] = 32'h416b0556;
    ram_cell[   36044] = 32'h4bf095a1;
    ram_cell[   36045] = 32'had400781;
    ram_cell[   36046] = 32'h9f1b7d77;
    ram_cell[   36047] = 32'h720a8058;
    ram_cell[   36048] = 32'hd9869b79;
    ram_cell[   36049] = 32'h7aad77ab;
    ram_cell[   36050] = 32'h74c5bfc7;
    ram_cell[   36051] = 32'h175154be;
    ram_cell[   36052] = 32'h54995a3b;
    ram_cell[   36053] = 32'he5d0547f;
    ram_cell[   36054] = 32'hdfc28acd;
    ram_cell[   36055] = 32'he9a798f7;
    ram_cell[   36056] = 32'h9a6ac796;
    ram_cell[   36057] = 32'h52b81f51;
    ram_cell[   36058] = 32'hbb804f7a;
    ram_cell[   36059] = 32'hd2ddada2;
    ram_cell[   36060] = 32'hfabbc2f6;
    ram_cell[   36061] = 32'h771cc813;
    ram_cell[   36062] = 32'hd75947f9;
    ram_cell[   36063] = 32'hfe4e048f;
    ram_cell[   36064] = 32'hf5b35d7e;
    ram_cell[   36065] = 32'h131199d4;
    ram_cell[   36066] = 32'hcc1869a4;
    ram_cell[   36067] = 32'h0849293b;
    ram_cell[   36068] = 32'hff6dfcc4;
    ram_cell[   36069] = 32'h5efba03b;
    ram_cell[   36070] = 32'h9b60ad9e;
    ram_cell[   36071] = 32'h37e454ac;
    ram_cell[   36072] = 32'h64450f2b;
    ram_cell[   36073] = 32'h2e318161;
    ram_cell[   36074] = 32'hde54faca;
    ram_cell[   36075] = 32'h28efef00;
    ram_cell[   36076] = 32'ha5c2ae62;
    ram_cell[   36077] = 32'h0a93627c;
    ram_cell[   36078] = 32'hf805f5dd;
    ram_cell[   36079] = 32'h4113fd6c;
    ram_cell[   36080] = 32'h9503fc5e;
    ram_cell[   36081] = 32'hd8f459bf;
    ram_cell[   36082] = 32'hab8c8da0;
    ram_cell[   36083] = 32'h9b0dff7c;
    ram_cell[   36084] = 32'hcb0fdf32;
    ram_cell[   36085] = 32'h9ebdbfd5;
    ram_cell[   36086] = 32'h6e36b78c;
    ram_cell[   36087] = 32'h6a5e6f17;
    ram_cell[   36088] = 32'h9530c4dd;
    ram_cell[   36089] = 32'h236c2ce3;
    ram_cell[   36090] = 32'h6dfef176;
    ram_cell[   36091] = 32'h5f7fdc6f;
    ram_cell[   36092] = 32'h5c02319b;
    ram_cell[   36093] = 32'h090521f8;
    ram_cell[   36094] = 32'h72c84c6e;
    ram_cell[   36095] = 32'ha4feb512;
    ram_cell[   36096] = 32'h38a009c9;
    ram_cell[   36097] = 32'h43f09817;
    ram_cell[   36098] = 32'hb00fa528;
    ram_cell[   36099] = 32'hb9250baf;
    ram_cell[   36100] = 32'ha4400d3a;
    ram_cell[   36101] = 32'h6acc7738;
    ram_cell[   36102] = 32'h384d8545;
    ram_cell[   36103] = 32'h91707138;
    ram_cell[   36104] = 32'h5da18207;
    ram_cell[   36105] = 32'h0dec8ae0;
    ram_cell[   36106] = 32'h3a9f0e64;
    ram_cell[   36107] = 32'h902b82a4;
    ram_cell[   36108] = 32'hbe325ce0;
    ram_cell[   36109] = 32'h54a22f45;
    ram_cell[   36110] = 32'h2f3807b3;
    ram_cell[   36111] = 32'h562945f0;
    ram_cell[   36112] = 32'h7a50b014;
    ram_cell[   36113] = 32'hf6e461ed;
    ram_cell[   36114] = 32'hac78bcaf;
    ram_cell[   36115] = 32'h7e548a66;
    ram_cell[   36116] = 32'he7e0035c;
    ram_cell[   36117] = 32'hfc2eeaef;
    ram_cell[   36118] = 32'h7da1f385;
    ram_cell[   36119] = 32'ha657ef1c;
    ram_cell[   36120] = 32'hc110f431;
    ram_cell[   36121] = 32'h270f4d00;
    ram_cell[   36122] = 32'h1088eff9;
    ram_cell[   36123] = 32'h1a6d9232;
    ram_cell[   36124] = 32'hda4e3bbb;
    ram_cell[   36125] = 32'h59f746cf;
    ram_cell[   36126] = 32'h21bef19d;
    ram_cell[   36127] = 32'h1e75f384;
    ram_cell[   36128] = 32'hdeab279e;
    ram_cell[   36129] = 32'h44910d9b;
    ram_cell[   36130] = 32'he055cbb2;
    ram_cell[   36131] = 32'ha587cb16;
    ram_cell[   36132] = 32'hd50e0a67;
    ram_cell[   36133] = 32'h992ffc87;
    ram_cell[   36134] = 32'h97e6fc01;
    ram_cell[   36135] = 32'he47e0cb0;
    ram_cell[   36136] = 32'ha5a62c51;
    ram_cell[   36137] = 32'ha62c3e42;
    ram_cell[   36138] = 32'hc94b1e82;
    ram_cell[   36139] = 32'he376332b;
    ram_cell[   36140] = 32'hac252479;
    ram_cell[   36141] = 32'h882c87af;
    ram_cell[   36142] = 32'hc79346df;
    ram_cell[   36143] = 32'h0b88425d;
    ram_cell[   36144] = 32'h7ff7a87e;
    ram_cell[   36145] = 32'hb983b645;
    ram_cell[   36146] = 32'hf67fbaad;
    ram_cell[   36147] = 32'hd948914f;
    ram_cell[   36148] = 32'h9661df54;
    ram_cell[   36149] = 32'h9571b5cd;
    ram_cell[   36150] = 32'hd7945c85;
    ram_cell[   36151] = 32'hef396086;
    ram_cell[   36152] = 32'hc9ac994e;
    ram_cell[   36153] = 32'h03dab8bf;
    ram_cell[   36154] = 32'h734e7e9a;
    ram_cell[   36155] = 32'ha55c58b3;
    ram_cell[   36156] = 32'h98b3b465;
    ram_cell[   36157] = 32'h1f473e0d;
    ram_cell[   36158] = 32'h0bc5b1f4;
    ram_cell[   36159] = 32'h978a8619;
    ram_cell[   36160] = 32'h7d40f7fa;
    ram_cell[   36161] = 32'h46a914ba;
    ram_cell[   36162] = 32'h23aa71b2;
    ram_cell[   36163] = 32'ha4894666;
    ram_cell[   36164] = 32'h2e3c2339;
    ram_cell[   36165] = 32'h122cfc17;
    ram_cell[   36166] = 32'h91776e54;
    ram_cell[   36167] = 32'hbeecab82;
    ram_cell[   36168] = 32'hf716c4a1;
    ram_cell[   36169] = 32'hf99299dc;
    ram_cell[   36170] = 32'h65fa529a;
    ram_cell[   36171] = 32'ha6d10647;
    ram_cell[   36172] = 32'hc03bd7bf;
    ram_cell[   36173] = 32'h9e6885c6;
    ram_cell[   36174] = 32'h4b94fb2f;
    ram_cell[   36175] = 32'h4ad5155f;
    ram_cell[   36176] = 32'he66583cd;
    ram_cell[   36177] = 32'hf7adfaa0;
    ram_cell[   36178] = 32'hfc6743b3;
    ram_cell[   36179] = 32'h3e2ef72d;
    ram_cell[   36180] = 32'h711b847a;
    ram_cell[   36181] = 32'hc4741d32;
    ram_cell[   36182] = 32'h5fbbdb93;
    ram_cell[   36183] = 32'he2864330;
    ram_cell[   36184] = 32'h3975fe9a;
    ram_cell[   36185] = 32'h0b0565b9;
    ram_cell[   36186] = 32'h9f84fbdd;
    ram_cell[   36187] = 32'h50bbb172;
    ram_cell[   36188] = 32'hb1facbef;
    ram_cell[   36189] = 32'hfeb12d5f;
    ram_cell[   36190] = 32'hce90b401;
    ram_cell[   36191] = 32'h0b62e85f;
    ram_cell[   36192] = 32'h06c81108;
    ram_cell[   36193] = 32'h45bcc86b;
    ram_cell[   36194] = 32'h2f01ad8e;
    ram_cell[   36195] = 32'h6dc70d89;
    ram_cell[   36196] = 32'head4f49c;
    ram_cell[   36197] = 32'h8207fde2;
    ram_cell[   36198] = 32'h3a205e33;
    ram_cell[   36199] = 32'hdbe89e11;
    ram_cell[   36200] = 32'h0ea12eb5;
    ram_cell[   36201] = 32'h8db6938d;
    ram_cell[   36202] = 32'h8f68b3fd;
    ram_cell[   36203] = 32'h836b6a2a;
    ram_cell[   36204] = 32'h669dade3;
    ram_cell[   36205] = 32'h57b9b08c;
    ram_cell[   36206] = 32'hdd0e0cea;
    ram_cell[   36207] = 32'hc25ee441;
    ram_cell[   36208] = 32'h2e38beac;
    ram_cell[   36209] = 32'he1c3b69c;
    ram_cell[   36210] = 32'h4c97cd75;
    ram_cell[   36211] = 32'h1b933b9d;
    ram_cell[   36212] = 32'h11f2c70c;
    ram_cell[   36213] = 32'h7d02c48e;
    ram_cell[   36214] = 32'h3ca531f8;
    ram_cell[   36215] = 32'h575c5166;
    ram_cell[   36216] = 32'h334355ac;
    ram_cell[   36217] = 32'ha41579a7;
    ram_cell[   36218] = 32'h7646bd37;
    ram_cell[   36219] = 32'h599eceaa;
    ram_cell[   36220] = 32'h9b7e7dce;
    ram_cell[   36221] = 32'h1055d6f4;
    ram_cell[   36222] = 32'h9e5bc59e;
    ram_cell[   36223] = 32'hee91e9d1;
    ram_cell[   36224] = 32'h3789041c;
    ram_cell[   36225] = 32'h07ad3972;
    ram_cell[   36226] = 32'h58da3384;
    ram_cell[   36227] = 32'h69241922;
    ram_cell[   36228] = 32'h576a036b;
    ram_cell[   36229] = 32'h9bfd3aa2;
    ram_cell[   36230] = 32'ha3ae4989;
    ram_cell[   36231] = 32'hc320ea55;
    ram_cell[   36232] = 32'h27ae2179;
    ram_cell[   36233] = 32'hbd726450;
    ram_cell[   36234] = 32'h346124fc;
    ram_cell[   36235] = 32'h6f600669;
    ram_cell[   36236] = 32'h7e1c84f2;
    ram_cell[   36237] = 32'hb132befe;
    ram_cell[   36238] = 32'h5f58c8ed;
    ram_cell[   36239] = 32'hdeb1075a;
    ram_cell[   36240] = 32'h4e463cb1;
    ram_cell[   36241] = 32'hf866e148;
    ram_cell[   36242] = 32'hb1934f3d;
    ram_cell[   36243] = 32'h2f1576de;
    ram_cell[   36244] = 32'h17ce1dbd;
    ram_cell[   36245] = 32'hdab69874;
    ram_cell[   36246] = 32'hc3571d46;
    ram_cell[   36247] = 32'h65349c28;
    ram_cell[   36248] = 32'hf14d79a6;
    ram_cell[   36249] = 32'hee1961fe;
    ram_cell[   36250] = 32'hbdef78da;
    ram_cell[   36251] = 32'hfbfea532;
    ram_cell[   36252] = 32'h61852e89;
    ram_cell[   36253] = 32'hf4d355ce;
    ram_cell[   36254] = 32'h30203c18;
    ram_cell[   36255] = 32'ha4b82e9d;
    ram_cell[   36256] = 32'h80338a29;
    ram_cell[   36257] = 32'h6a6dad0e;
    ram_cell[   36258] = 32'h36f6dcac;
    ram_cell[   36259] = 32'hefac3799;
    ram_cell[   36260] = 32'h3a2e7a37;
    ram_cell[   36261] = 32'h5d5006ca;
    ram_cell[   36262] = 32'h4fb8fdeb;
    ram_cell[   36263] = 32'ha42fa1ef;
    ram_cell[   36264] = 32'h3f231f91;
    ram_cell[   36265] = 32'h37cfe7d5;
    ram_cell[   36266] = 32'h2ffd56e0;
    ram_cell[   36267] = 32'h036783a2;
    ram_cell[   36268] = 32'hd89a6b59;
    ram_cell[   36269] = 32'h8f34db15;
    ram_cell[   36270] = 32'h674845a6;
    ram_cell[   36271] = 32'h9cb8acff;
    ram_cell[   36272] = 32'hd0321c60;
    ram_cell[   36273] = 32'h3ce97e19;
    ram_cell[   36274] = 32'haef73883;
    ram_cell[   36275] = 32'hd3c4629d;
    ram_cell[   36276] = 32'ha37f323d;
    ram_cell[   36277] = 32'h48993e4d;
    ram_cell[   36278] = 32'h313085f6;
    ram_cell[   36279] = 32'hbcf8140e;
    ram_cell[   36280] = 32'hc414f358;
    ram_cell[   36281] = 32'h5fe52bb6;
    ram_cell[   36282] = 32'h4f95c1ab;
    ram_cell[   36283] = 32'h12577b5a;
    ram_cell[   36284] = 32'h7fc00e2d;
    ram_cell[   36285] = 32'h2f8bbd56;
    ram_cell[   36286] = 32'h639cd2a7;
    ram_cell[   36287] = 32'h5a4d7ef2;
    ram_cell[   36288] = 32'h194770b3;
    ram_cell[   36289] = 32'hccb0deaf;
    ram_cell[   36290] = 32'h9e9e884a;
    ram_cell[   36291] = 32'h61bd9784;
    ram_cell[   36292] = 32'h2f50ae5f;
    ram_cell[   36293] = 32'ha34cd351;
    ram_cell[   36294] = 32'hab03f0b8;
    ram_cell[   36295] = 32'hf6ba6b91;
    ram_cell[   36296] = 32'h7e981a4e;
    ram_cell[   36297] = 32'h1c4b098a;
    ram_cell[   36298] = 32'h0a9d98a3;
    ram_cell[   36299] = 32'hfe481985;
    ram_cell[   36300] = 32'hffe5326f;
    ram_cell[   36301] = 32'hfd5a2307;
    ram_cell[   36302] = 32'ha1fd3ecd;
    ram_cell[   36303] = 32'he55adb78;
    ram_cell[   36304] = 32'h08689d5b;
    ram_cell[   36305] = 32'h47e45f5e;
    ram_cell[   36306] = 32'h0177981e;
    ram_cell[   36307] = 32'h9381bc05;
    ram_cell[   36308] = 32'h791e570f;
    ram_cell[   36309] = 32'h882b8f67;
    ram_cell[   36310] = 32'h784842c4;
    ram_cell[   36311] = 32'h8c66599e;
    ram_cell[   36312] = 32'hc76c94e0;
    ram_cell[   36313] = 32'h5ed759b0;
    ram_cell[   36314] = 32'haeb9ce6a;
    ram_cell[   36315] = 32'h0ae78fc6;
    ram_cell[   36316] = 32'h86145f39;
    ram_cell[   36317] = 32'hec0d69a1;
    ram_cell[   36318] = 32'h51d9df44;
    ram_cell[   36319] = 32'h4c8de89e;
    ram_cell[   36320] = 32'hc3069704;
    ram_cell[   36321] = 32'h3cc591ac;
    ram_cell[   36322] = 32'hc44845bd;
    ram_cell[   36323] = 32'hf3b5a6c1;
    ram_cell[   36324] = 32'hc7135e62;
    ram_cell[   36325] = 32'hce8b6f0e;
    ram_cell[   36326] = 32'h1e80d9d2;
    ram_cell[   36327] = 32'hcfdf8646;
    ram_cell[   36328] = 32'h0378ff61;
    ram_cell[   36329] = 32'h4b0b69e8;
    ram_cell[   36330] = 32'h143733a6;
    ram_cell[   36331] = 32'h623acc01;
    ram_cell[   36332] = 32'h643158f8;
    ram_cell[   36333] = 32'h734588cd;
    ram_cell[   36334] = 32'had5c6ea6;
    ram_cell[   36335] = 32'h97717a05;
    ram_cell[   36336] = 32'h14489c0e;
    ram_cell[   36337] = 32'h58f9f873;
    ram_cell[   36338] = 32'h12c954fa;
    ram_cell[   36339] = 32'h55c3bacb;
    ram_cell[   36340] = 32'h9cf520e3;
    ram_cell[   36341] = 32'h945ac0f0;
    ram_cell[   36342] = 32'h25485ae6;
    ram_cell[   36343] = 32'h3ffdde9c;
    ram_cell[   36344] = 32'h1b617cbb;
    ram_cell[   36345] = 32'hf5343d36;
    ram_cell[   36346] = 32'h2db0e588;
    ram_cell[   36347] = 32'h6aa7dec1;
    ram_cell[   36348] = 32'hd10c7ced;
    ram_cell[   36349] = 32'h223f1c8c;
    ram_cell[   36350] = 32'h1d975840;
    ram_cell[   36351] = 32'hdcb896f3;
    ram_cell[   36352] = 32'ha6b27c2a;
    ram_cell[   36353] = 32'h18750d8a;
    ram_cell[   36354] = 32'hdb91026c;
    ram_cell[   36355] = 32'h5d7e9c09;
    ram_cell[   36356] = 32'h89b4ce31;
    ram_cell[   36357] = 32'hb695840c;
    ram_cell[   36358] = 32'h7b9fb89d;
    ram_cell[   36359] = 32'ha450e58c;
    ram_cell[   36360] = 32'he9fb423f;
    ram_cell[   36361] = 32'h04f97540;
    ram_cell[   36362] = 32'h68e4d466;
    ram_cell[   36363] = 32'h5264239d;
    ram_cell[   36364] = 32'he33abc56;
    ram_cell[   36365] = 32'hee7be308;
    ram_cell[   36366] = 32'h2ae7c7ab;
    ram_cell[   36367] = 32'hdfb03198;
    ram_cell[   36368] = 32'h351da2d3;
    ram_cell[   36369] = 32'he8fd8fef;
    ram_cell[   36370] = 32'hcb8041ed;
    ram_cell[   36371] = 32'h35c1ca4d;
    ram_cell[   36372] = 32'h7a2ac569;
    ram_cell[   36373] = 32'h0d9e47b9;
    ram_cell[   36374] = 32'ha7300f76;
    ram_cell[   36375] = 32'hdfe21431;
    ram_cell[   36376] = 32'h6c256891;
    ram_cell[   36377] = 32'h975c818b;
    ram_cell[   36378] = 32'he9b977ee;
    ram_cell[   36379] = 32'ha75f3d41;
    ram_cell[   36380] = 32'h93241fc1;
    ram_cell[   36381] = 32'h8fc0d497;
    ram_cell[   36382] = 32'h6178b7a1;
    ram_cell[   36383] = 32'h5cfe54ff;
    ram_cell[   36384] = 32'h6e6efb6a;
    ram_cell[   36385] = 32'hb67f9081;
    ram_cell[   36386] = 32'h21e190d7;
    ram_cell[   36387] = 32'h0789ec4b;
    ram_cell[   36388] = 32'h28c99c69;
    ram_cell[   36389] = 32'h6547233a;
    ram_cell[   36390] = 32'hb29c7871;
    ram_cell[   36391] = 32'hdd3cceaa;
    ram_cell[   36392] = 32'h4d70a47d;
    ram_cell[   36393] = 32'h4197b1c2;
    ram_cell[   36394] = 32'ha4ef7cb7;
    ram_cell[   36395] = 32'hfe642d69;
    ram_cell[   36396] = 32'hc6dab12c;
    ram_cell[   36397] = 32'h851ca1d9;
    ram_cell[   36398] = 32'h02233043;
    ram_cell[   36399] = 32'h2cab12eb;
    ram_cell[   36400] = 32'h12bfa32e;
    ram_cell[   36401] = 32'h0bcfbe9d;
    ram_cell[   36402] = 32'hb337a389;
    ram_cell[   36403] = 32'hf3273403;
    ram_cell[   36404] = 32'hb96ad0ef;
    ram_cell[   36405] = 32'h72154f81;
    ram_cell[   36406] = 32'h7af3506e;
    ram_cell[   36407] = 32'h5f1c26fe;
    ram_cell[   36408] = 32'hd4f19031;
    ram_cell[   36409] = 32'h875fcb92;
    ram_cell[   36410] = 32'h36474338;
    ram_cell[   36411] = 32'h14a94310;
    ram_cell[   36412] = 32'h72cd610f;
    ram_cell[   36413] = 32'h544ec809;
    ram_cell[   36414] = 32'h21a4ffa0;
    ram_cell[   36415] = 32'h9dc513aa;
    ram_cell[   36416] = 32'h474f381c;
    ram_cell[   36417] = 32'h019a22a5;
    ram_cell[   36418] = 32'h20c5af62;
    ram_cell[   36419] = 32'hc770a155;
    ram_cell[   36420] = 32'h93a1e886;
    ram_cell[   36421] = 32'hfb55c825;
    ram_cell[   36422] = 32'h7b70ca24;
    ram_cell[   36423] = 32'haeaa61d7;
    ram_cell[   36424] = 32'h7b5679ef;
    ram_cell[   36425] = 32'h6156ac00;
    ram_cell[   36426] = 32'h50915f38;
    ram_cell[   36427] = 32'hca449d6e;
    ram_cell[   36428] = 32'h196c656b;
    ram_cell[   36429] = 32'hd3c8a6c7;
    ram_cell[   36430] = 32'he2bc4c11;
    ram_cell[   36431] = 32'h4ee1bd8f;
    ram_cell[   36432] = 32'h717e28d9;
    ram_cell[   36433] = 32'hf32cd2c5;
    ram_cell[   36434] = 32'hd6109715;
    ram_cell[   36435] = 32'hd4c283f6;
    ram_cell[   36436] = 32'he46aefcb;
    ram_cell[   36437] = 32'h1e4b365d;
    ram_cell[   36438] = 32'hf999f1bf;
    ram_cell[   36439] = 32'h80f654ec;
    ram_cell[   36440] = 32'h73685ad2;
    ram_cell[   36441] = 32'h13f9e832;
    ram_cell[   36442] = 32'h508b754c;
    ram_cell[   36443] = 32'h9950a7b9;
    ram_cell[   36444] = 32'h7b673465;
    ram_cell[   36445] = 32'h54e5f132;
    ram_cell[   36446] = 32'h562ca97d;
    ram_cell[   36447] = 32'h7401d356;
    ram_cell[   36448] = 32'hbfd9ec84;
    ram_cell[   36449] = 32'hae635b30;
    ram_cell[   36450] = 32'h4a1b921f;
    ram_cell[   36451] = 32'h66c2b209;
    ram_cell[   36452] = 32'h477888c3;
    ram_cell[   36453] = 32'h85f39254;
    ram_cell[   36454] = 32'h4fcbb8fa;
    ram_cell[   36455] = 32'hb5c6a933;
    ram_cell[   36456] = 32'h13860d46;
    ram_cell[   36457] = 32'h47334320;
    ram_cell[   36458] = 32'heaeadfb6;
    ram_cell[   36459] = 32'hfc917125;
    ram_cell[   36460] = 32'h765d82e5;
    ram_cell[   36461] = 32'hddc4a91d;
    ram_cell[   36462] = 32'h07c3e717;
    ram_cell[   36463] = 32'h3fa93b84;
    ram_cell[   36464] = 32'hd145c373;
    ram_cell[   36465] = 32'hf48ef693;
    ram_cell[   36466] = 32'h04abf87d;
    ram_cell[   36467] = 32'h0fe94573;
    ram_cell[   36468] = 32'h912cd82e;
    ram_cell[   36469] = 32'h01d7c04b;
    ram_cell[   36470] = 32'h0818277d;
    ram_cell[   36471] = 32'h01f0a053;
    ram_cell[   36472] = 32'hded0b5ba;
    ram_cell[   36473] = 32'h1ffb56af;
    ram_cell[   36474] = 32'h0b5e2409;
    ram_cell[   36475] = 32'ha2726cb2;
    ram_cell[   36476] = 32'hec9ccb39;
    ram_cell[   36477] = 32'h6268b4c1;
    ram_cell[   36478] = 32'hd1982611;
    ram_cell[   36479] = 32'h820c5f44;
    ram_cell[   36480] = 32'he4115228;
    ram_cell[   36481] = 32'h8d19d1c4;
    ram_cell[   36482] = 32'hb0397e6c;
    ram_cell[   36483] = 32'h731f7db7;
    ram_cell[   36484] = 32'hc02d199a;
    ram_cell[   36485] = 32'h9ab7782f;
    ram_cell[   36486] = 32'h6dc50989;
    ram_cell[   36487] = 32'h97915001;
    ram_cell[   36488] = 32'hee244f3a;
    ram_cell[   36489] = 32'h7aa2e940;
    ram_cell[   36490] = 32'hb273f45e;
    ram_cell[   36491] = 32'h3673870b;
    ram_cell[   36492] = 32'hf8cfda51;
    ram_cell[   36493] = 32'h5e8fa913;
    ram_cell[   36494] = 32'h4d834c84;
    ram_cell[   36495] = 32'h962c21f3;
    ram_cell[   36496] = 32'hdab054ae;
    ram_cell[   36497] = 32'hb3c532b1;
    ram_cell[   36498] = 32'hf8ca309a;
    ram_cell[   36499] = 32'h2d81df6d;
    ram_cell[   36500] = 32'h6ae17c01;
    ram_cell[   36501] = 32'h06c4015e;
    ram_cell[   36502] = 32'he4609afb;
    ram_cell[   36503] = 32'h02432234;
    ram_cell[   36504] = 32'h9ee73e1e;
    ram_cell[   36505] = 32'h7d291a42;
    ram_cell[   36506] = 32'h7aa2309e;
    ram_cell[   36507] = 32'hc12943eb;
    ram_cell[   36508] = 32'h806bca46;
    ram_cell[   36509] = 32'h562c9881;
    ram_cell[   36510] = 32'hf31739b7;
    ram_cell[   36511] = 32'hf7b5892a;
    ram_cell[   36512] = 32'hbd1e7e4e;
    ram_cell[   36513] = 32'hc72f0ef3;
    ram_cell[   36514] = 32'h4edb6482;
    ram_cell[   36515] = 32'h0f18fc71;
    ram_cell[   36516] = 32'h383a1aac;
    ram_cell[   36517] = 32'he422a6a1;
    ram_cell[   36518] = 32'h78b35cbc;
    ram_cell[   36519] = 32'ha2621fcd;
    ram_cell[   36520] = 32'h488e8141;
    ram_cell[   36521] = 32'h026ad001;
    ram_cell[   36522] = 32'h634af0e5;
    ram_cell[   36523] = 32'h8adacf56;
    ram_cell[   36524] = 32'h2df6635a;
    ram_cell[   36525] = 32'h91011550;
    ram_cell[   36526] = 32'h38d42de7;
    ram_cell[   36527] = 32'h97b583ee;
    ram_cell[   36528] = 32'h77697a42;
    ram_cell[   36529] = 32'h3913481b;
    ram_cell[   36530] = 32'h4c47f87d;
    ram_cell[   36531] = 32'hbcbe0ef6;
    ram_cell[   36532] = 32'hef1309aa;
    ram_cell[   36533] = 32'h9aaa78d4;
    ram_cell[   36534] = 32'h0892ca9b;
    ram_cell[   36535] = 32'h7d3a1262;
    ram_cell[   36536] = 32'h4b199687;
    ram_cell[   36537] = 32'hca1a0a07;
    ram_cell[   36538] = 32'h8275e7af;
    ram_cell[   36539] = 32'h9e0d4397;
    ram_cell[   36540] = 32'h8bdd7896;
    ram_cell[   36541] = 32'hd122b6b6;
    ram_cell[   36542] = 32'h49ec6b05;
    ram_cell[   36543] = 32'hf80fe4c9;
    ram_cell[   36544] = 32'hdb29d25d;
    ram_cell[   36545] = 32'h5c39b42e;
    ram_cell[   36546] = 32'hc5890956;
    ram_cell[   36547] = 32'h01299f96;
    ram_cell[   36548] = 32'h0f7ca3f4;
    ram_cell[   36549] = 32'h1e71a71a;
    ram_cell[   36550] = 32'hc225b4e2;
    ram_cell[   36551] = 32'hdce6e857;
    ram_cell[   36552] = 32'hddba60c0;
    ram_cell[   36553] = 32'h778a429b;
    ram_cell[   36554] = 32'h3976d12c;
    ram_cell[   36555] = 32'ha2358fe5;
    ram_cell[   36556] = 32'haa5565fe;
    ram_cell[   36557] = 32'h254ffd69;
    ram_cell[   36558] = 32'hf7ee0349;
    ram_cell[   36559] = 32'h83b86c51;
    ram_cell[   36560] = 32'h2fc90a2a;
    ram_cell[   36561] = 32'h4c0bd012;
    ram_cell[   36562] = 32'h9f40d53f;
    ram_cell[   36563] = 32'hbee7ac57;
    ram_cell[   36564] = 32'hc56fcbc6;
    ram_cell[   36565] = 32'hf9c46182;
    ram_cell[   36566] = 32'h5793b87b;
    ram_cell[   36567] = 32'hb37e2ec5;
    ram_cell[   36568] = 32'h286201eb;
    ram_cell[   36569] = 32'hdb5afd91;
    ram_cell[   36570] = 32'h3c08d88c;
    ram_cell[   36571] = 32'h2faa8877;
    ram_cell[   36572] = 32'h9b56f0e3;
    ram_cell[   36573] = 32'h2d42d056;
    ram_cell[   36574] = 32'h48d1b457;
    ram_cell[   36575] = 32'heae77247;
    ram_cell[   36576] = 32'h68c19f06;
    ram_cell[   36577] = 32'h26f58977;
    ram_cell[   36578] = 32'h20a5799d;
    ram_cell[   36579] = 32'hd2fed687;
    ram_cell[   36580] = 32'h7993b11e;
    ram_cell[   36581] = 32'hf8d30887;
    ram_cell[   36582] = 32'h2f2e8c0b;
    ram_cell[   36583] = 32'h3401c68f;
    ram_cell[   36584] = 32'haa9b1441;
    ram_cell[   36585] = 32'h9b37f754;
    ram_cell[   36586] = 32'h303838f4;
    ram_cell[   36587] = 32'hbb253c18;
    ram_cell[   36588] = 32'h81d9145e;
    ram_cell[   36589] = 32'hc3bf0828;
    ram_cell[   36590] = 32'hf2bb97b7;
    ram_cell[   36591] = 32'hb34ca15e;
    ram_cell[   36592] = 32'h1afeda51;
    ram_cell[   36593] = 32'hacf245c9;
    ram_cell[   36594] = 32'hf7041f27;
    ram_cell[   36595] = 32'h1736aa0a;
    ram_cell[   36596] = 32'h58513f92;
    ram_cell[   36597] = 32'h657a5ee9;
    ram_cell[   36598] = 32'he462f8c9;
    ram_cell[   36599] = 32'h86dfa8df;
    ram_cell[   36600] = 32'hfe6ec992;
    ram_cell[   36601] = 32'h2be02dcb;
    ram_cell[   36602] = 32'h90cac685;
    ram_cell[   36603] = 32'h80ce40d4;
    ram_cell[   36604] = 32'h16946797;
    ram_cell[   36605] = 32'h7dd3dd08;
    ram_cell[   36606] = 32'hb99e4cbe;
    ram_cell[   36607] = 32'h7a897a60;
    ram_cell[   36608] = 32'he1dba132;
    ram_cell[   36609] = 32'h0a43ceb1;
    ram_cell[   36610] = 32'h27245e66;
    ram_cell[   36611] = 32'he167ecb4;
    ram_cell[   36612] = 32'h5e453796;
    ram_cell[   36613] = 32'h7887561d;
    ram_cell[   36614] = 32'h82e77f38;
    ram_cell[   36615] = 32'h49db3e39;
    ram_cell[   36616] = 32'h03523eac;
    ram_cell[   36617] = 32'h33fe52c0;
    ram_cell[   36618] = 32'hba48832e;
    ram_cell[   36619] = 32'h536e2a2d;
    ram_cell[   36620] = 32'hfd091ce8;
    ram_cell[   36621] = 32'h3758886b;
    ram_cell[   36622] = 32'he69a554d;
    ram_cell[   36623] = 32'h4b3be386;
    ram_cell[   36624] = 32'h7047895f;
    ram_cell[   36625] = 32'h6cecd05a;
    ram_cell[   36626] = 32'h3485e696;
    ram_cell[   36627] = 32'h5e6a0af4;
    ram_cell[   36628] = 32'ha7d3b0f7;
    ram_cell[   36629] = 32'h91f6390e;
    ram_cell[   36630] = 32'h97f25401;
    ram_cell[   36631] = 32'he11ae762;
    ram_cell[   36632] = 32'h10dd9bf1;
    ram_cell[   36633] = 32'h419d55c4;
    ram_cell[   36634] = 32'h58f9a5e9;
    ram_cell[   36635] = 32'hfb1d99da;
    ram_cell[   36636] = 32'hf2652210;
    ram_cell[   36637] = 32'h38fce42a;
    ram_cell[   36638] = 32'h9154b7dd;
    ram_cell[   36639] = 32'hdec119e7;
    ram_cell[   36640] = 32'hd38ac1b5;
    ram_cell[   36641] = 32'hcd5ee89b;
    ram_cell[   36642] = 32'h9cb6ae8d;
    ram_cell[   36643] = 32'hf25eea1d;
    ram_cell[   36644] = 32'h78c4c5f1;
    ram_cell[   36645] = 32'h947ae60e;
    ram_cell[   36646] = 32'h880e3514;
    ram_cell[   36647] = 32'hb6addcb4;
    ram_cell[   36648] = 32'hf9774a7c;
    ram_cell[   36649] = 32'h56f4c086;
    ram_cell[   36650] = 32'h7ad8e10a;
    ram_cell[   36651] = 32'hbed29a04;
    ram_cell[   36652] = 32'hba320130;
    ram_cell[   36653] = 32'h845f4afe;
    ram_cell[   36654] = 32'hd2e8752a;
    ram_cell[   36655] = 32'hffa699ed;
    ram_cell[   36656] = 32'h7b84a444;
    ram_cell[   36657] = 32'h1cd9d7b9;
    ram_cell[   36658] = 32'h2bbc5425;
    ram_cell[   36659] = 32'h25d994ab;
    ram_cell[   36660] = 32'h587c62ec;
    ram_cell[   36661] = 32'hba00c00f;
    ram_cell[   36662] = 32'ha10a90ba;
    ram_cell[   36663] = 32'hfbdd366e;
    ram_cell[   36664] = 32'hc4ab81af;
    ram_cell[   36665] = 32'h84f75b8d;
    ram_cell[   36666] = 32'hea255cb7;
    ram_cell[   36667] = 32'h178da5d4;
    ram_cell[   36668] = 32'h0e22f524;
    ram_cell[   36669] = 32'h13c86b41;
    ram_cell[   36670] = 32'h794af2d0;
    ram_cell[   36671] = 32'h570ab536;
    ram_cell[   36672] = 32'h4cb71431;
    ram_cell[   36673] = 32'h32d28f64;
    ram_cell[   36674] = 32'heb23bf8e;
    ram_cell[   36675] = 32'h9755d1a9;
    ram_cell[   36676] = 32'h8646c62c;
    ram_cell[   36677] = 32'h0653cd50;
    ram_cell[   36678] = 32'h7bc8ebc5;
    ram_cell[   36679] = 32'ha7ab3ce8;
    ram_cell[   36680] = 32'hbc313379;
    ram_cell[   36681] = 32'hae38b0b7;
    ram_cell[   36682] = 32'hef88d111;
    ram_cell[   36683] = 32'h0c74f85f;
    ram_cell[   36684] = 32'hcebf39c1;
    ram_cell[   36685] = 32'h1f3fa5d0;
    ram_cell[   36686] = 32'hecc7abd4;
    ram_cell[   36687] = 32'hf1900e30;
    ram_cell[   36688] = 32'hea990d88;
    ram_cell[   36689] = 32'h56f60c6e;
    ram_cell[   36690] = 32'h8244ce9f;
    ram_cell[   36691] = 32'h8c2f679d;
    ram_cell[   36692] = 32'h737bb649;
    ram_cell[   36693] = 32'h8c8b1d4f;
    ram_cell[   36694] = 32'hc9781e72;
    ram_cell[   36695] = 32'he3aefd69;
    ram_cell[   36696] = 32'h58d20764;
    ram_cell[   36697] = 32'h81a4dac9;
    ram_cell[   36698] = 32'hf95b319c;
    ram_cell[   36699] = 32'hb80f39d6;
    ram_cell[   36700] = 32'h29380769;
    ram_cell[   36701] = 32'h725f1eda;
    ram_cell[   36702] = 32'h0a973ded;
    ram_cell[   36703] = 32'h04d91829;
    ram_cell[   36704] = 32'h0bc753af;
    ram_cell[   36705] = 32'hdcbb7eda;
    ram_cell[   36706] = 32'hdcdb2318;
    ram_cell[   36707] = 32'h861d1f21;
    ram_cell[   36708] = 32'hf36f0f0e;
    ram_cell[   36709] = 32'h603f0daa;
    ram_cell[   36710] = 32'h37d5f571;
    ram_cell[   36711] = 32'h260ba11d;
    ram_cell[   36712] = 32'h1eaa18fb;
    ram_cell[   36713] = 32'ha4b5802b;
    ram_cell[   36714] = 32'he7932810;
    ram_cell[   36715] = 32'h93bb1005;
    ram_cell[   36716] = 32'hd9a89f27;
    ram_cell[   36717] = 32'hd3ebe84c;
    ram_cell[   36718] = 32'h4c0297e3;
    ram_cell[   36719] = 32'hf2300346;
    ram_cell[   36720] = 32'h27145fd8;
    ram_cell[   36721] = 32'h5297b046;
    ram_cell[   36722] = 32'h65ddf18a;
    ram_cell[   36723] = 32'hf09111cc;
    ram_cell[   36724] = 32'he94e9b39;
    ram_cell[   36725] = 32'h5b62e4bd;
    ram_cell[   36726] = 32'hc5145ca5;
    ram_cell[   36727] = 32'hec692b83;
    ram_cell[   36728] = 32'h1ac70e6b;
    ram_cell[   36729] = 32'h9a510238;
    ram_cell[   36730] = 32'hba80fc2e;
    ram_cell[   36731] = 32'haa4e6363;
    ram_cell[   36732] = 32'h97d24804;
    ram_cell[   36733] = 32'hf0890c0b;
    ram_cell[   36734] = 32'h1d0910a0;
    ram_cell[   36735] = 32'hbb354e1f;
    ram_cell[   36736] = 32'h52065df7;
    ram_cell[   36737] = 32'h0f5ed9c8;
    ram_cell[   36738] = 32'h5c17f575;
    ram_cell[   36739] = 32'h6c5e3f40;
    ram_cell[   36740] = 32'h4e0e9e7a;
    ram_cell[   36741] = 32'ha4491c35;
    ram_cell[   36742] = 32'h3d02de7e;
    ram_cell[   36743] = 32'hfd8b492a;
    ram_cell[   36744] = 32'h80b35e2a;
    ram_cell[   36745] = 32'h95904fa4;
    ram_cell[   36746] = 32'hb4150157;
    ram_cell[   36747] = 32'hfac00ec9;
    ram_cell[   36748] = 32'hddcf45b2;
    ram_cell[   36749] = 32'h356db952;
    ram_cell[   36750] = 32'h0b664771;
    ram_cell[   36751] = 32'h303b0a21;
    ram_cell[   36752] = 32'h66fdeb70;
    ram_cell[   36753] = 32'hcfc25103;
    ram_cell[   36754] = 32'h873335e6;
    ram_cell[   36755] = 32'h68dbed2a;
    ram_cell[   36756] = 32'he9d95143;
    ram_cell[   36757] = 32'ha5fc0431;
    ram_cell[   36758] = 32'ha6ce21f0;
    ram_cell[   36759] = 32'hf89f5097;
    ram_cell[   36760] = 32'h7597fa37;
    ram_cell[   36761] = 32'hc3555601;
    ram_cell[   36762] = 32'hbd964575;
    ram_cell[   36763] = 32'h2de78b9c;
    ram_cell[   36764] = 32'he36f48da;
    ram_cell[   36765] = 32'he4cf4e1f;
    ram_cell[   36766] = 32'h6784a9c2;
    ram_cell[   36767] = 32'hb155bc6d;
    ram_cell[   36768] = 32'h5c2b79a3;
    ram_cell[   36769] = 32'heb42a738;
    ram_cell[   36770] = 32'hc47b2920;
    ram_cell[   36771] = 32'h8caee874;
    ram_cell[   36772] = 32'hbd51f1c6;
    ram_cell[   36773] = 32'h9ffae39f;
    ram_cell[   36774] = 32'h78343579;
    ram_cell[   36775] = 32'h602049cf;
    ram_cell[   36776] = 32'hfb52341e;
    ram_cell[   36777] = 32'h60b4ea46;
    ram_cell[   36778] = 32'h1d0c6d92;
    ram_cell[   36779] = 32'h544a2241;
    ram_cell[   36780] = 32'h7fe50a48;
    ram_cell[   36781] = 32'h69c10afb;
    ram_cell[   36782] = 32'h0ece3e24;
    ram_cell[   36783] = 32'hdfa5fcc3;
    ram_cell[   36784] = 32'h5837c4ad;
    ram_cell[   36785] = 32'hd6bc8905;
    ram_cell[   36786] = 32'hffdfccea;
    ram_cell[   36787] = 32'h4eff99c6;
    ram_cell[   36788] = 32'h21b72afd;
    ram_cell[   36789] = 32'h9acbd354;
    ram_cell[   36790] = 32'h2171e933;
    ram_cell[   36791] = 32'hf3970938;
    ram_cell[   36792] = 32'h0cb25d1e;
    ram_cell[   36793] = 32'h04d61653;
    ram_cell[   36794] = 32'h02ba8762;
    ram_cell[   36795] = 32'h6a705d61;
    ram_cell[   36796] = 32'h9127945b;
    ram_cell[   36797] = 32'hf2552174;
    ram_cell[   36798] = 32'h89b5c005;
    ram_cell[   36799] = 32'h15981c2f;
    ram_cell[   36800] = 32'h5063c019;
    ram_cell[   36801] = 32'hcdc6e2ab;
    ram_cell[   36802] = 32'hb88e950c;
    ram_cell[   36803] = 32'h75ea3474;
    ram_cell[   36804] = 32'he22ba287;
    ram_cell[   36805] = 32'h63495195;
    ram_cell[   36806] = 32'hd3841911;
    ram_cell[   36807] = 32'hb99471e4;
    ram_cell[   36808] = 32'h7fa6601f;
    ram_cell[   36809] = 32'he8614d67;
    ram_cell[   36810] = 32'h92f98ed5;
    ram_cell[   36811] = 32'h3740aa7a;
    ram_cell[   36812] = 32'h3538bf98;
    ram_cell[   36813] = 32'h4cc93a28;
    ram_cell[   36814] = 32'hfb65d72f;
    ram_cell[   36815] = 32'h2c2c80b3;
    ram_cell[   36816] = 32'hcbc6556c;
    ram_cell[   36817] = 32'ha138a36e;
    ram_cell[   36818] = 32'hbdc841e9;
    ram_cell[   36819] = 32'h9c24bbf8;
    ram_cell[   36820] = 32'h075814bd;
    ram_cell[   36821] = 32'h62b11423;
    ram_cell[   36822] = 32'head4c908;
    ram_cell[   36823] = 32'hab6dad4a;
    ram_cell[   36824] = 32'h49f930fc;
    ram_cell[   36825] = 32'h9fef81de;
    ram_cell[   36826] = 32'h51973735;
    ram_cell[   36827] = 32'h5c49f47c;
    ram_cell[   36828] = 32'ha21394f1;
    ram_cell[   36829] = 32'h742b7311;
    ram_cell[   36830] = 32'h580c9f9b;
    ram_cell[   36831] = 32'hd9bfb496;
    ram_cell[   36832] = 32'hed615290;
    ram_cell[   36833] = 32'hb6094d90;
    ram_cell[   36834] = 32'h8d19cd47;
    ram_cell[   36835] = 32'h63f5a07b;
    ram_cell[   36836] = 32'ha9180501;
    ram_cell[   36837] = 32'heaf4490a;
    ram_cell[   36838] = 32'h0a8db073;
    ram_cell[   36839] = 32'h53fbbafa;
    ram_cell[   36840] = 32'h90109fd7;
    ram_cell[   36841] = 32'hfa5f1d46;
    ram_cell[   36842] = 32'h2843b23a;
    ram_cell[   36843] = 32'h34860eef;
    ram_cell[   36844] = 32'hab36a150;
    ram_cell[   36845] = 32'hda6e3c2c;
    ram_cell[   36846] = 32'hb58a1489;
    ram_cell[   36847] = 32'hf8b06f67;
    ram_cell[   36848] = 32'h5c018d2c;
    ram_cell[   36849] = 32'ha89d31f9;
    ram_cell[   36850] = 32'h1f7849fa;
    ram_cell[   36851] = 32'h2ffc5914;
    ram_cell[   36852] = 32'h84c69866;
    ram_cell[   36853] = 32'h3cd81add;
    ram_cell[   36854] = 32'he296fa19;
    ram_cell[   36855] = 32'h7510cb55;
    ram_cell[   36856] = 32'h85aa1d88;
    ram_cell[   36857] = 32'h09c501f0;
    ram_cell[   36858] = 32'hb63e6dcc;
    ram_cell[   36859] = 32'h5ad8119a;
    ram_cell[   36860] = 32'h34f60c7c;
    ram_cell[   36861] = 32'h620ba7b1;
    ram_cell[   36862] = 32'h635c821e;
    ram_cell[   36863] = 32'h2bb961b0;
    ram_cell[   36864] = 32'h662e5d01;
    ram_cell[   36865] = 32'h240c9f4f;
    ram_cell[   36866] = 32'h6b909408;
    ram_cell[   36867] = 32'hf773689f;
    ram_cell[   36868] = 32'h31f426b7;
    ram_cell[   36869] = 32'h00b41d90;
    ram_cell[   36870] = 32'h659a8ab1;
    ram_cell[   36871] = 32'h1c2e39f7;
    ram_cell[   36872] = 32'hd7d18ae0;
    ram_cell[   36873] = 32'ha36f71c2;
    ram_cell[   36874] = 32'h5dd2ae97;
    ram_cell[   36875] = 32'hbe8c9f24;
    ram_cell[   36876] = 32'h5cfafceb;
    ram_cell[   36877] = 32'hff3a8cdf;
    ram_cell[   36878] = 32'hdb888f60;
    ram_cell[   36879] = 32'h4700d380;
    ram_cell[   36880] = 32'h7210f32a;
    ram_cell[   36881] = 32'hdbca36d8;
    ram_cell[   36882] = 32'h4a26eb8e;
    ram_cell[   36883] = 32'hfcebd640;
    ram_cell[   36884] = 32'hb4ddb9fc;
    ram_cell[   36885] = 32'h1660164c;
    ram_cell[   36886] = 32'h8289ab16;
    ram_cell[   36887] = 32'h8b776d6e;
    ram_cell[   36888] = 32'he309064e;
    ram_cell[   36889] = 32'h6c4310b8;
    ram_cell[   36890] = 32'h65b8ab13;
    ram_cell[   36891] = 32'hb6bcd287;
    ram_cell[   36892] = 32'h66098fcc;
    ram_cell[   36893] = 32'h90785e99;
    ram_cell[   36894] = 32'hbeef4a6c;
    ram_cell[   36895] = 32'h480f8e0b;
    ram_cell[   36896] = 32'hd7ca0ed5;
    ram_cell[   36897] = 32'hfa21f20c;
    ram_cell[   36898] = 32'hb5987dec;
    ram_cell[   36899] = 32'h420e81e6;
    ram_cell[   36900] = 32'h0ff39fb8;
    ram_cell[   36901] = 32'h5c5905b0;
    ram_cell[   36902] = 32'h546718c2;
    ram_cell[   36903] = 32'h3c743dbb;
    ram_cell[   36904] = 32'h24176264;
    ram_cell[   36905] = 32'hf8e736a6;
    ram_cell[   36906] = 32'h77235d76;
    ram_cell[   36907] = 32'h94304c50;
    ram_cell[   36908] = 32'hca556ebc;
    ram_cell[   36909] = 32'h2bdba2ef;
    ram_cell[   36910] = 32'hd3e7b6ed;
    ram_cell[   36911] = 32'h67eda3d7;
    ram_cell[   36912] = 32'h89fcabbf;
    ram_cell[   36913] = 32'hfad727f3;
    ram_cell[   36914] = 32'hf3578404;
    ram_cell[   36915] = 32'h2a522cc3;
    ram_cell[   36916] = 32'ha5a0bf56;
    ram_cell[   36917] = 32'h04c9858d;
    ram_cell[   36918] = 32'hfdc568fb;
    ram_cell[   36919] = 32'h26642179;
    ram_cell[   36920] = 32'h1346cab6;
    ram_cell[   36921] = 32'h7664485c;
    ram_cell[   36922] = 32'h01821a5d;
    ram_cell[   36923] = 32'h90a4e3ed;
    ram_cell[   36924] = 32'h7b6061be;
    ram_cell[   36925] = 32'h9bd042ed;
    ram_cell[   36926] = 32'h345a58aa;
    ram_cell[   36927] = 32'hdfba419e;
    ram_cell[   36928] = 32'h720fadd9;
    ram_cell[   36929] = 32'h1fa71414;
    ram_cell[   36930] = 32'h59f3a6e9;
    ram_cell[   36931] = 32'h6b84992c;
    ram_cell[   36932] = 32'h6f589b67;
    ram_cell[   36933] = 32'h499bae31;
    ram_cell[   36934] = 32'h68f14693;
    ram_cell[   36935] = 32'ha86d0720;
    ram_cell[   36936] = 32'hc7aa846a;
    ram_cell[   36937] = 32'hc922c095;
    ram_cell[   36938] = 32'h4ae1869f;
    ram_cell[   36939] = 32'h1d8d0458;
    ram_cell[   36940] = 32'hcc9f9ac3;
    ram_cell[   36941] = 32'h460c6bb5;
    ram_cell[   36942] = 32'hd6a3d35e;
    ram_cell[   36943] = 32'hd168d485;
    ram_cell[   36944] = 32'h003fd1a8;
    ram_cell[   36945] = 32'h637c6dba;
    ram_cell[   36946] = 32'h4b9a250f;
    ram_cell[   36947] = 32'h0dd50fee;
    ram_cell[   36948] = 32'hf7d6bece;
    ram_cell[   36949] = 32'h904efb8d;
    ram_cell[   36950] = 32'hdb0d7730;
    ram_cell[   36951] = 32'h091c5ae6;
    ram_cell[   36952] = 32'h7624298a;
    ram_cell[   36953] = 32'h8f8e1dc8;
    ram_cell[   36954] = 32'h1904e46e;
    ram_cell[   36955] = 32'h174ae63e;
    ram_cell[   36956] = 32'h4b969aa9;
    ram_cell[   36957] = 32'haab4c879;
    ram_cell[   36958] = 32'haf1c63c7;
    ram_cell[   36959] = 32'h68ce62a4;
    ram_cell[   36960] = 32'h68a67a51;
    ram_cell[   36961] = 32'h43b6edf7;
    ram_cell[   36962] = 32'h5998f0a8;
    ram_cell[   36963] = 32'h49f7b204;
    ram_cell[   36964] = 32'hb59aaa2a;
    ram_cell[   36965] = 32'h37880326;
    ram_cell[   36966] = 32'h903abd53;
    ram_cell[   36967] = 32'h8063b53f;
    ram_cell[   36968] = 32'h8eca400b;
    ram_cell[   36969] = 32'heb45adf6;
    ram_cell[   36970] = 32'hef15b939;
    ram_cell[   36971] = 32'he6bc346f;
    ram_cell[   36972] = 32'h9e8c8ec0;
    ram_cell[   36973] = 32'h4fe5945b;
    ram_cell[   36974] = 32'h5ce90b53;
    ram_cell[   36975] = 32'hc92a78f9;
    ram_cell[   36976] = 32'h01f93988;
    ram_cell[   36977] = 32'ha16f0f04;
    ram_cell[   36978] = 32'hb6cd929e;
    ram_cell[   36979] = 32'h99b59e58;
    ram_cell[   36980] = 32'ha6a71b7d;
    ram_cell[   36981] = 32'h8cf9ad45;
    ram_cell[   36982] = 32'hdc6b3254;
    ram_cell[   36983] = 32'h7b42fca4;
    ram_cell[   36984] = 32'hf39709a4;
    ram_cell[   36985] = 32'h77566c47;
    ram_cell[   36986] = 32'h4d01175b;
    ram_cell[   36987] = 32'h3e857cad;
    ram_cell[   36988] = 32'h13b0a4fa;
    ram_cell[   36989] = 32'hb8d0a798;
    ram_cell[   36990] = 32'h12c5af75;
    ram_cell[   36991] = 32'h6c77c9b4;
    ram_cell[   36992] = 32'had4f13b9;
    ram_cell[   36993] = 32'h320136cb;
    ram_cell[   36994] = 32'h466f4b63;
    ram_cell[   36995] = 32'ha8b44b3e;
    ram_cell[   36996] = 32'hdcbefe0c;
    ram_cell[   36997] = 32'h8d87a273;
    ram_cell[   36998] = 32'h7d1eb8fa;
    ram_cell[   36999] = 32'hcb51b72d;
    ram_cell[   37000] = 32'h12500935;
    ram_cell[   37001] = 32'h8dfc696a;
    ram_cell[   37002] = 32'h9ae75edf;
    ram_cell[   37003] = 32'hb09f81c5;
    ram_cell[   37004] = 32'hb3b1a9ad;
    ram_cell[   37005] = 32'hc74c3385;
    ram_cell[   37006] = 32'h342644bd;
    ram_cell[   37007] = 32'hbf24a398;
    ram_cell[   37008] = 32'hcb903047;
    ram_cell[   37009] = 32'h4b97980c;
    ram_cell[   37010] = 32'hd0da9957;
    ram_cell[   37011] = 32'h9152f149;
    ram_cell[   37012] = 32'h8b55d7c1;
    ram_cell[   37013] = 32'h484addd1;
    ram_cell[   37014] = 32'h98a2a82b;
    ram_cell[   37015] = 32'he64a3e29;
    ram_cell[   37016] = 32'h36bda4b7;
    ram_cell[   37017] = 32'had1ef5be;
    ram_cell[   37018] = 32'he14706fe;
    ram_cell[   37019] = 32'h23fd5af1;
    ram_cell[   37020] = 32'hf1e44622;
    ram_cell[   37021] = 32'hf8556b58;
    ram_cell[   37022] = 32'h21f3e7ae;
    ram_cell[   37023] = 32'hf41d9890;
    ram_cell[   37024] = 32'h5932c6f7;
    ram_cell[   37025] = 32'h6d4614d7;
    ram_cell[   37026] = 32'h5ee04c8d;
    ram_cell[   37027] = 32'h0bbf675c;
    ram_cell[   37028] = 32'h2240ad17;
    ram_cell[   37029] = 32'h2574834d;
    ram_cell[   37030] = 32'hc1ac8707;
    ram_cell[   37031] = 32'h82dca21c;
    ram_cell[   37032] = 32'h76d998bf;
    ram_cell[   37033] = 32'h46e4043d;
    ram_cell[   37034] = 32'hb1f0b356;
    ram_cell[   37035] = 32'h0312fc01;
    ram_cell[   37036] = 32'h92b82c46;
    ram_cell[   37037] = 32'h3252f679;
    ram_cell[   37038] = 32'hcaccc1d7;
    ram_cell[   37039] = 32'hfc03aba2;
    ram_cell[   37040] = 32'hc61be73a;
    ram_cell[   37041] = 32'hb51ca2b1;
    ram_cell[   37042] = 32'h0b331e78;
    ram_cell[   37043] = 32'h9c3cebd8;
    ram_cell[   37044] = 32'hff86ebb0;
    ram_cell[   37045] = 32'h3afe868d;
    ram_cell[   37046] = 32'h4a43338e;
    ram_cell[   37047] = 32'h0a9fa089;
    ram_cell[   37048] = 32'hebf70efc;
    ram_cell[   37049] = 32'h55a3afed;
    ram_cell[   37050] = 32'h38ae6f11;
    ram_cell[   37051] = 32'hd397a908;
    ram_cell[   37052] = 32'h852aa222;
    ram_cell[   37053] = 32'hdb0ea1b7;
    ram_cell[   37054] = 32'h60718cb9;
    ram_cell[   37055] = 32'hd055bf8f;
    ram_cell[   37056] = 32'h1d960063;
    ram_cell[   37057] = 32'hf9c51829;
    ram_cell[   37058] = 32'h2d428b56;
    ram_cell[   37059] = 32'h44951dd4;
    ram_cell[   37060] = 32'h0fc37a2f;
    ram_cell[   37061] = 32'hf6ff6f88;
    ram_cell[   37062] = 32'h988f7f96;
    ram_cell[   37063] = 32'h52ea4fc9;
    ram_cell[   37064] = 32'hcd358559;
    ram_cell[   37065] = 32'hc874a3c5;
    ram_cell[   37066] = 32'h4d8ebd4b;
    ram_cell[   37067] = 32'h90cf99ee;
    ram_cell[   37068] = 32'hf3fe38f8;
    ram_cell[   37069] = 32'h6772006b;
    ram_cell[   37070] = 32'heaa1cc07;
    ram_cell[   37071] = 32'h437d392d;
    ram_cell[   37072] = 32'haaf62305;
    ram_cell[   37073] = 32'h6a87e09b;
    ram_cell[   37074] = 32'h70736ed5;
    ram_cell[   37075] = 32'heabcfb50;
    ram_cell[   37076] = 32'hb5f7ec0c;
    ram_cell[   37077] = 32'h6c6f6c79;
    ram_cell[   37078] = 32'h45b745eb;
    ram_cell[   37079] = 32'hac1f6b34;
    ram_cell[   37080] = 32'h7567fedd;
    ram_cell[   37081] = 32'h77d3544f;
    ram_cell[   37082] = 32'h00b8131a;
    ram_cell[   37083] = 32'h33d4abdb;
    ram_cell[   37084] = 32'hb8544c35;
    ram_cell[   37085] = 32'h63060a42;
    ram_cell[   37086] = 32'h0f25f2d1;
    ram_cell[   37087] = 32'h04778b59;
    ram_cell[   37088] = 32'hf13c9f06;
    ram_cell[   37089] = 32'h2bdbc74d;
    ram_cell[   37090] = 32'h53d87110;
    ram_cell[   37091] = 32'h38863e86;
    ram_cell[   37092] = 32'h0ce09418;
    ram_cell[   37093] = 32'h430d10b5;
    ram_cell[   37094] = 32'h8c1a7a43;
    ram_cell[   37095] = 32'h411fe79f;
    ram_cell[   37096] = 32'h6379e45a;
    ram_cell[   37097] = 32'h09eed8fa;
    ram_cell[   37098] = 32'hc132d3cc;
    ram_cell[   37099] = 32'h1c14a8ee;
    ram_cell[   37100] = 32'hda59180b;
    ram_cell[   37101] = 32'hb0dc9017;
    ram_cell[   37102] = 32'h810a9f8a;
    ram_cell[   37103] = 32'h3021e888;
    ram_cell[   37104] = 32'hc4f91ae0;
    ram_cell[   37105] = 32'h4e73cb51;
    ram_cell[   37106] = 32'hca19f74b;
    ram_cell[   37107] = 32'h9ef51ee1;
    ram_cell[   37108] = 32'h930acb2b;
    ram_cell[   37109] = 32'h842e151b;
    ram_cell[   37110] = 32'h4427e136;
    ram_cell[   37111] = 32'hff873ad0;
    ram_cell[   37112] = 32'h90d66111;
    ram_cell[   37113] = 32'hac20e535;
    ram_cell[   37114] = 32'hb909355d;
    ram_cell[   37115] = 32'hd5c53ab8;
    ram_cell[   37116] = 32'haf5b1a28;
    ram_cell[   37117] = 32'h0a922bb1;
    ram_cell[   37118] = 32'h74ab0ad4;
    ram_cell[   37119] = 32'h6e9f93cf;
    ram_cell[   37120] = 32'h49fdd1fd;
    ram_cell[   37121] = 32'h0827c4e4;
    ram_cell[   37122] = 32'h54057732;
    ram_cell[   37123] = 32'h32dc5692;
    ram_cell[   37124] = 32'hd50fba87;
    ram_cell[   37125] = 32'h20be3fa6;
    ram_cell[   37126] = 32'h69a838a8;
    ram_cell[   37127] = 32'h0128a5aa;
    ram_cell[   37128] = 32'h9485e7a9;
    ram_cell[   37129] = 32'h2cdcf541;
    ram_cell[   37130] = 32'h4d189393;
    ram_cell[   37131] = 32'h2e029d26;
    ram_cell[   37132] = 32'h51a062e6;
    ram_cell[   37133] = 32'h59ff1e33;
    ram_cell[   37134] = 32'hcb2a5059;
    ram_cell[   37135] = 32'ha4859b4b;
    ram_cell[   37136] = 32'h746c42d0;
    ram_cell[   37137] = 32'hdd87fb91;
    ram_cell[   37138] = 32'h53eb2bb2;
    ram_cell[   37139] = 32'h93aea9bc;
    ram_cell[   37140] = 32'h109ce06f;
    ram_cell[   37141] = 32'h2ee419ee;
    ram_cell[   37142] = 32'h6f16d6a4;
    ram_cell[   37143] = 32'haf5e8edb;
    ram_cell[   37144] = 32'h9b7e4330;
    ram_cell[   37145] = 32'h1f375829;
    ram_cell[   37146] = 32'h4c8599cc;
    ram_cell[   37147] = 32'h487536d6;
    ram_cell[   37148] = 32'h777afd4c;
    ram_cell[   37149] = 32'hc68a9d0c;
    ram_cell[   37150] = 32'h3fd84037;
    ram_cell[   37151] = 32'he8ffb0c4;
    ram_cell[   37152] = 32'he9d16e54;
    ram_cell[   37153] = 32'hf57ef097;
    ram_cell[   37154] = 32'h1b25d7b2;
    ram_cell[   37155] = 32'h126f0a18;
    ram_cell[   37156] = 32'haf090536;
    ram_cell[   37157] = 32'h190847ae;
    ram_cell[   37158] = 32'he6ddd45f;
    ram_cell[   37159] = 32'h94a0031f;
    ram_cell[   37160] = 32'h09e7d2e1;
    ram_cell[   37161] = 32'hb6c28277;
    ram_cell[   37162] = 32'h8c16e9b0;
    ram_cell[   37163] = 32'h0c25c491;
    ram_cell[   37164] = 32'h9989a963;
    ram_cell[   37165] = 32'he27ccfe2;
    ram_cell[   37166] = 32'h5d671b25;
    ram_cell[   37167] = 32'he6a49fc0;
    ram_cell[   37168] = 32'h60c55681;
    ram_cell[   37169] = 32'h485d3882;
    ram_cell[   37170] = 32'h1541f1f3;
    ram_cell[   37171] = 32'hec6bf945;
    ram_cell[   37172] = 32'h751263ac;
    ram_cell[   37173] = 32'h43bba6a3;
    ram_cell[   37174] = 32'h565acb64;
    ram_cell[   37175] = 32'h08a046cb;
    ram_cell[   37176] = 32'h08ffd66e;
    ram_cell[   37177] = 32'h73a91c7f;
    ram_cell[   37178] = 32'h833cb823;
    ram_cell[   37179] = 32'h2b167dda;
    ram_cell[   37180] = 32'h98ea4537;
    ram_cell[   37181] = 32'h897c06de;
    ram_cell[   37182] = 32'he35903f3;
    ram_cell[   37183] = 32'hdb0ebdc9;
    ram_cell[   37184] = 32'h5909a684;
    ram_cell[   37185] = 32'ha5f416f4;
    ram_cell[   37186] = 32'h2301c33b;
    ram_cell[   37187] = 32'he8bb61bb;
    ram_cell[   37188] = 32'h0d10600c;
    ram_cell[   37189] = 32'ha2c4ed38;
    ram_cell[   37190] = 32'h17b56cbd;
    ram_cell[   37191] = 32'hfc1f15e4;
    ram_cell[   37192] = 32'hf9d3ff21;
    ram_cell[   37193] = 32'h673010c8;
    ram_cell[   37194] = 32'h6f27e3df;
    ram_cell[   37195] = 32'hfbb56972;
    ram_cell[   37196] = 32'h6b52da30;
    ram_cell[   37197] = 32'h9f4208b0;
    ram_cell[   37198] = 32'h843c4c08;
    ram_cell[   37199] = 32'h012044b8;
    ram_cell[   37200] = 32'h2fa60d13;
    ram_cell[   37201] = 32'he4cf5767;
    ram_cell[   37202] = 32'he2ad988a;
    ram_cell[   37203] = 32'hc2cd3ead;
    ram_cell[   37204] = 32'hbaee89c6;
    ram_cell[   37205] = 32'h92e6bcb0;
    ram_cell[   37206] = 32'h2203cecd;
    ram_cell[   37207] = 32'h3149edf1;
    ram_cell[   37208] = 32'h390ff5cd;
    ram_cell[   37209] = 32'h804949f9;
    ram_cell[   37210] = 32'h543b9d12;
    ram_cell[   37211] = 32'haf15292f;
    ram_cell[   37212] = 32'hc8d12fae;
    ram_cell[   37213] = 32'h9c215491;
    ram_cell[   37214] = 32'hda99de1c;
    ram_cell[   37215] = 32'he0f73dce;
    ram_cell[   37216] = 32'ha81878ec;
    ram_cell[   37217] = 32'h62fa58c5;
    ram_cell[   37218] = 32'h23a996ce;
    ram_cell[   37219] = 32'h6d723742;
    ram_cell[   37220] = 32'h5b14689f;
    ram_cell[   37221] = 32'hf9a7d3fd;
    ram_cell[   37222] = 32'hf879d927;
    ram_cell[   37223] = 32'h4675871d;
    ram_cell[   37224] = 32'h8d6fa89e;
    ram_cell[   37225] = 32'h2ee43b87;
    ram_cell[   37226] = 32'haefa2548;
    ram_cell[   37227] = 32'h590c6e25;
    ram_cell[   37228] = 32'hc0b7c68e;
    ram_cell[   37229] = 32'h5a9c9215;
    ram_cell[   37230] = 32'h0513eec8;
    ram_cell[   37231] = 32'h75e4d858;
    ram_cell[   37232] = 32'ha9b9d265;
    ram_cell[   37233] = 32'h0cc6e988;
    ram_cell[   37234] = 32'h416520ae;
    ram_cell[   37235] = 32'h2fc8f3e4;
    ram_cell[   37236] = 32'h7d433c66;
    ram_cell[   37237] = 32'h680882e8;
    ram_cell[   37238] = 32'h9b9442dd;
    ram_cell[   37239] = 32'h3313212a;
    ram_cell[   37240] = 32'hdaf2853c;
    ram_cell[   37241] = 32'hacffd5fe;
    ram_cell[   37242] = 32'h607b707d;
    ram_cell[   37243] = 32'hb18a37d8;
    ram_cell[   37244] = 32'h20aac4c7;
    ram_cell[   37245] = 32'h83634e4f;
    ram_cell[   37246] = 32'h1be4039e;
    ram_cell[   37247] = 32'ha66f4f4a;
    ram_cell[   37248] = 32'hbc7ae68b;
    ram_cell[   37249] = 32'hb695076c;
    ram_cell[   37250] = 32'hb69d7bbe;
    ram_cell[   37251] = 32'he47f4dde;
    ram_cell[   37252] = 32'hbc42c476;
    ram_cell[   37253] = 32'h5fe9d63d;
    ram_cell[   37254] = 32'h1920f96a;
    ram_cell[   37255] = 32'h658a5f02;
    ram_cell[   37256] = 32'h1660f9e4;
    ram_cell[   37257] = 32'hc93c5b12;
    ram_cell[   37258] = 32'he937adc0;
    ram_cell[   37259] = 32'hc0640aa5;
    ram_cell[   37260] = 32'hab86c60f;
    ram_cell[   37261] = 32'hd96d31c5;
    ram_cell[   37262] = 32'h57cf3d7f;
    ram_cell[   37263] = 32'hc5c298de;
    ram_cell[   37264] = 32'h88d6db9c;
    ram_cell[   37265] = 32'h10f6042b;
    ram_cell[   37266] = 32'hab4a19d3;
    ram_cell[   37267] = 32'h1e01d0ae;
    ram_cell[   37268] = 32'h4f7be529;
    ram_cell[   37269] = 32'h0bed3055;
    ram_cell[   37270] = 32'h6c3826f9;
    ram_cell[   37271] = 32'h37dd68dd;
    ram_cell[   37272] = 32'hba83d668;
    ram_cell[   37273] = 32'hfba5fe94;
    ram_cell[   37274] = 32'hb6a8b68c;
    ram_cell[   37275] = 32'hd91ee84e;
    ram_cell[   37276] = 32'hd6d62fa2;
    ram_cell[   37277] = 32'hbbf72f50;
    ram_cell[   37278] = 32'h6d121b93;
    ram_cell[   37279] = 32'ha81bf767;
    ram_cell[   37280] = 32'hc1a9354d;
    ram_cell[   37281] = 32'h13644517;
    ram_cell[   37282] = 32'hd929e4a7;
    ram_cell[   37283] = 32'h242ac07f;
    ram_cell[   37284] = 32'h950a1741;
    ram_cell[   37285] = 32'h8a1556ae;
    ram_cell[   37286] = 32'h2a95f0bb;
    ram_cell[   37287] = 32'hc4592f25;
    ram_cell[   37288] = 32'hd2db589a;
    ram_cell[   37289] = 32'hed135741;
    ram_cell[   37290] = 32'h99336e52;
    ram_cell[   37291] = 32'hadd0aa83;
    ram_cell[   37292] = 32'h706d1b51;
    ram_cell[   37293] = 32'h4203cffd;
    ram_cell[   37294] = 32'h5ed1f457;
    ram_cell[   37295] = 32'h76d1846d;
    ram_cell[   37296] = 32'h1f946980;
    ram_cell[   37297] = 32'h40eecaa6;
    ram_cell[   37298] = 32'h13bc4f53;
    ram_cell[   37299] = 32'hdeb86070;
    ram_cell[   37300] = 32'h6bb15d61;
    ram_cell[   37301] = 32'hfe5f2a3c;
    ram_cell[   37302] = 32'h7e009861;
    ram_cell[   37303] = 32'h115b9ea1;
    ram_cell[   37304] = 32'hd57b7d97;
    ram_cell[   37305] = 32'h3134aa7a;
    ram_cell[   37306] = 32'h9f08421d;
    ram_cell[   37307] = 32'hd96f469e;
    ram_cell[   37308] = 32'h0b9024f8;
    ram_cell[   37309] = 32'h47bea526;
    ram_cell[   37310] = 32'h0e7fe5fe;
    ram_cell[   37311] = 32'h7dcedc2d;
    ram_cell[   37312] = 32'h2fa2d371;
    ram_cell[   37313] = 32'hbbfb4973;
    ram_cell[   37314] = 32'h7030f5e2;
    ram_cell[   37315] = 32'h3d3af6d3;
    ram_cell[   37316] = 32'h0664779b;
    ram_cell[   37317] = 32'h0f1950f2;
    ram_cell[   37318] = 32'h7af2d265;
    ram_cell[   37319] = 32'h0c07df1b;
    ram_cell[   37320] = 32'ha96daae3;
    ram_cell[   37321] = 32'hbdbed698;
    ram_cell[   37322] = 32'hff753670;
    ram_cell[   37323] = 32'h00887c64;
    ram_cell[   37324] = 32'h5131bc38;
    ram_cell[   37325] = 32'hd1d0d65d;
    ram_cell[   37326] = 32'h7fd71dfb;
    ram_cell[   37327] = 32'h4a5b6558;
    ram_cell[   37328] = 32'hb1dc6daa;
    ram_cell[   37329] = 32'hf93d65f6;
    ram_cell[   37330] = 32'h13077f08;
    ram_cell[   37331] = 32'hd2bab67a;
    ram_cell[   37332] = 32'h6248a1a6;
    ram_cell[   37333] = 32'h4c2ebe29;
    ram_cell[   37334] = 32'h9788daeb;
    ram_cell[   37335] = 32'hb6f54a52;
    ram_cell[   37336] = 32'hd1ee9475;
    ram_cell[   37337] = 32'h1937f174;
    ram_cell[   37338] = 32'h25eb8e4c;
    ram_cell[   37339] = 32'h1772177e;
    ram_cell[   37340] = 32'h936eaf69;
    ram_cell[   37341] = 32'hb2bd9df4;
    ram_cell[   37342] = 32'h2ca854eb;
    ram_cell[   37343] = 32'he21f2dfc;
    ram_cell[   37344] = 32'h76ddc3f3;
    ram_cell[   37345] = 32'h92b0aab6;
    ram_cell[   37346] = 32'h2af7b75b;
    ram_cell[   37347] = 32'ha23f2910;
    ram_cell[   37348] = 32'h4ef01efc;
    ram_cell[   37349] = 32'hc8279fac;
    ram_cell[   37350] = 32'h3c1d8bdb;
    ram_cell[   37351] = 32'h4e52db71;
    ram_cell[   37352] = 32'hf1de302d;
    ram_cell[   37353] = 32'hf83891cc;
    ram_cell[   37354] = 32'hb4a48396;
    ram_cell[   37355] = 32'he75f4180;
    ram_cell[   37356] = 32'h99edf1d7;
    ram_cell[   37357] = 32'he45679d3;
    ram_cell[   37358] = 32'h2b3cf85e;
    ram_cell[   37359] = 32'hf9e3e7d9;
    ram_cell[   37360] = 32'h6bc1d948;
    ram_cell[   37361] = 32'h88f3eeeb;
    ram_cell[   37362] = 32'hb499e1a8;
    ram_cell[   37363] = 32'hf3565af1;
    ram_cell[   37364] = 32'h7f1608ec;
    ram_cell[   37365] = 32'h9c2b4a4a;
    ram_cell[   37366] = 32'h3696963c;
    ram_cell[   37367] = 32'h1146ff12;
    ram_cell[   37368] = 32'hb45ce465;
    ram_cell[   37369] = 32'hc5004bad;
    ram_cell[   37370] = 32'hcf87176c;
    ram_cell[   37371] = 32'h8acb4411;
    ram_cell[   37372] = 32'h3d56bb9e;
    ram_cell[   37373] = 32'h13a96ca2;
    ram_cell[   37374] = 32'h7bde5dd6;
    ram_cell[   37375] = 32'h9939b250;
    ram_cell[   37376] = 32'h1b1bc70e;
    ram_cell[   37377] = 32'ha249d1d6;
    ram_cell[   37378] = 32'h40b6e3e0;
    ram_cell[   37379] = 32'h0edc7895;
    ram_cell[   37380] = 32'haaf9dc19;
    ram_cell[   37381] = 32'h20e21656;
    ram_cell[   37382] = 32'h107b081e;
    ram_cell[   37383] = 32'hd2446984;
    ram_cell[   37384] = 32'h347492fe;
    ram_cell[   37385] = 32'h5b8cf257;
    ram_cell[   37386] = 32'h2a4f05a7;
    ram_cell[   37387] = 32'h3fec9531;
    ram_cell[   37388] = 32'ha684acad;
    ram_cell[   37389] = 32'h6ca732ba;
    ram_cell[   37390] = 32'hbbdd38f2;
    ram_cell[   37391] = 32'hcb17ade2;
    ram_cell[   37392] = 32'hfdbb6a64;
    ram_cell[   37393] = 32'h377418c9;
    ram_cell[   37394] = 32'hf9c78bb3;
    ram_cell[   37395] = 32'h6c61800d;
    ram_cell[   37396] = 32'hdb96848f;
    ram_cell[   37397] = 32'hd91b8b0f;
    ram_cell[   37398] = 32'h069aa548;
    ram_cell[   37399] = 32'h3a56fa55;
    ram_cell[   37400] = 32'he3f0299b;
    ram_cell[   37401] = 32'hc93dd513;
    ram_cell[   37402] = 32'h1a5746cd;
    ram_cell[   37403] = 32'hb0600a70;
    ram_cell[   37404] = 32'h49426929;
    ram_cell[   37405] = 32'hf155818d;
    ram_cell[   37406] = 32'h429bf922;
    ram_cell[   37407] = 32'hf53ea08f;
    ram_cell[   37408] = 32'h4ddef9d3;
    ram_cell[   37409] = 32'hc181555c;
    ram_cell[   37410] = 32'h962e7a7f;
    ram_cell[   37411] = 32'hf50af3a9;
    ram_cell[   37412] = 32'h50bc24ae;
    ram_cell[   37413] = 32'h2a0d2ddf;
    ram_cell[   37414] = 32'h1afc6d80;
    ram_cell[   37415] = 32'h70b4bf39;
    ram_cell[   37416] = 32'h99fe352f;
    ram_cell[   37417] = 32'h8b0a3a16;
    ram_cell[   37418] = 32'h007308e3;
    ram_cell[   37419] = 32'h11f6d576;
    ram_cell[   37420] = 32'hb6238065;
    ram_cell[   37421] = 32'h4c234e4e;
    ram_cell[   37422] = 32'h66d2043e;
    ram_cell[   37423] = 32'h1e1b9974;
    ram_cell[   37424] = 32'h060eb9f8;
    ram_cell[   37425] = 32'h734fb01b;
    ram_cell[   37426] = 32'h1fd81ceb;
    ram_cell[   37427] = 32'h61810c7c;
    ram_cell[   37428] = 32'h8700a33c;
    ram_cell[   37429] = 32'hd44c56a6;
    ram_cell[   37430] = 32'h9bf9d73f;
    ram_cell[   37431] = 32'hc286a614;
    ram_cell[   37432] = 32'h59acf255;
    ram_cell[   37433] = 32'hd4bd76d4;
    ram_cell[   37434] = 32'h0ffb2299;
    ram_cell[   37435] = 32'h16402aa0;
    ram_cell[   37436] = 32'he9860b32;
    ram_cell[   37437] = 32'haa448405;
    ram_cell[   37438] = 32'h3313dad0;
    ram_cell[   37439] = 32'h97e72810;
    ram_cell[   37440] = 32'hc1a9ebe5;
    ram_cell[   37441] = 32'h16105186;
    ram_cell[   37442] = 32'h52b77af7;
    ram_cell[   37443] = 32'he6e13e18;
    ram_cell[   37444] = 32'h4d557b9f;
    ram_cell[   37445] = 32'h9cbd8b2a;
    ram_cell[   37446] = 32'h6100a84d;
    ram_cell[   37447] = 32'hbb8d06fc;
    ram_cell[   37448] = 32'h324fed7d;
    ram_cell[   37449] = 32'h1ad7b221;
    ram_cell[   37450] = 32'h88b0dce3;
    ram_cell[   37451] = 32'h8d5904c8;
    ram_cell[   37452] = 32'h61a58ac6;
    ram_cell[   37453] = 32'h2ae1b214;
    ram_cell[   37454] = 32'hf47e8f8a;
    ram_cell[   37455] = 32'ha2b88d1d;
    ram_cell[   37456] = 32'hf6fe561a;
    ram_cell[   37457] = 32'hb093246a;
    ram_cell[   37458] = 32'h8b7d6a35;
    ram_cell[   37459] = 32'h2d3f9436;
    ram_cell[   37460] = 32'hafa581dc;
    ram_cell[   37461] = 32'h33dcd6c2;
    ram_cell[   37462] = 32'h5e5941da;
    ram_cell[   37463] = 32'h5af97696;
    ram_cell[   37464] = 32'ha733a2bf;
    ram_cell[   37465] = 32'h2c9f9843;
    ram_cell[   37466] = 32'hf8266058;
    ram_cell[   37467] = 32'ha8a4ea62;
    ram_cell[   37468] = 32'hb48b71be;
    ram_cell[   37469] = 32'hc674f28a;
    ram_cell[   37470] = 32'h21fbbdaf;
    ram_cell[   37471] = 32'h55d46075;
    ram_cell[   37472] = 32'hc5155288;
    ram_cell[   37473] = 32'h6c1851f7;
    ram_cell[   37474] = 32'hfe5a60ba;
    ram_cell[   37475] = 32'h99452cd9;
    ram_cell[   37476] = 32'h2f7aa699;
    ram_cell[   37477] = 32'h6ac66b2f;
    ram_cell[   37478] = 32'h86fce883;
    ram_cell[   37479] = 32'h7bb48800;
    ram_cell[   37480] = 32'he00dc711;
    ram_cell[   37481] = 32'hb4f1a464;
    ram_cell[   37482] = 32'h6770ae75;
    ram_cell[   37483] = 32'h37a68d2c;
    ram_cell[   37484] = 32'ha9a8a886;
    ram_cell[   37485] = 32'h890c7497;
    ram_cell[   37486] = 32'hb4ea4095;
    ram_cell[   37487] = 32'hc5342c15;
    ram_cell[   37488] = 32'hb038b65e;
    ram_cell[   37489] = 32'h60e718a5;
    ram_cell[   37490] = 32'ha0284500;
    ram_cell[   37491] = 32'h36c07d60;
    ram_cell[   37492] = 32'hdd463401;
    ram_cell[   37493] = 32'haf4f0b6a;
    ram_cell[   37494] = 32'h4520cd7a;
    ram_cell[   37495] = 32'ha9e0a405;
    ram_cell[   37496] = 32'h2b771b24;
    ram_cell[   37497] = 32'h35a3fc26;
    ram_cell[   37498] = 32'hbac272cf;
    ram_cell[   37499] = 32'h0a830f07;
    ram_cell[   37500] = 32'hbf4a015a;
    ram_cell[   37501] = 32'hbe21a6a5;
    ram_cell[   37502] = 32'h1c5a590a;
    ram_cell[   37503] = 32'h07dde8a0;
    ram_cell[   37504] = 32'h92b5cc04;
    ram_cell[   37505] = 32'h82af15e2;
    ram_cell[   37506] = 32'hef512267;
    ram_cell[   37507] = 32'h716de9ef;
    ram_cell[   37508] = 32'h2e0038bb;
    ram_cell[   37509] = 32'h4c3c0855;
    ram_cell[   37510] = 32'h6ed829ff;
    ram_cell[   37511] = 32'h66151dca;
    ram_cell[   37512] = 32'hd54d5e77;
    ram_cell[   37513] = 32'h282356ab;
    ram_cell[   37514] = 32'h16a3b9cd;
    ram_cell[   37515] = 32'h90d4fdc7;
    ram_cell[   37516] = 32'h9f3c72af;
    ram_cell[   37517] = 32'h8d982913;
    ram_cell[   37518] = 32'h2e0c7659;
    ram_cell[   37519] = 32'heb8535cf;
    ram_cell[   37520] = 32'h5a48bd4d;
    ram_cell[   37521] = 32'h560da4fc;
    ram_cell[   37522] = 32'h0f827c5d;
    ram_cell[   37523] = 32'hfe2fdaec;
    ram_cell[   37524] = 32'hd57232b6;
    ram_cell[   37525] = 32'hdaaea8e2;
    ram_cell[   37526] = 32'h86419400;
    ram_cell[   37527] = 32'h81ef4227;
    ram_cell[   37528] = 32'hf460ce42;
    ram_cell[   37529] = 32'h0dd8e2a0;
    ram_cell[   37530] = 32'h45ea1443;
    ram_cell[   37531] = 32'h2215695e;
    ram_cell[   37532] = 32'h1ab3b522;
    ram_cell[   37533] = 32'hf9d326fa;
    ram_cell[   37534] = 32'h77bf88c2;
    ram_cell[   37535] = 32'hfb3226b6;
    ram_cell[   37536] = 32'h209211ee;
    ram_cell[   37537] = 32'h37264ec9;
    ram_cell[   37538] = 32'h6d9220c5;
    ram_cell[   37539] = 32'h7308fce2;
    ram_cell[   37540] = 32'h923f05f3;
    ram_cell[   37541] = 32'h719e9b11;
    ram_cell[   37542] = 32'h280d71c1;
    ram_cell[   37543] = 32'h8d94d850;
    ram_cell[   37544] = 32'h4b221823;
    ram_cell[   37545] = 32'hb2e43e55;
    ram_cell[   37546] = 32'hc4b59255;
    ram_cell[   37547] = 32'h002d2c3b;
    ram_cell[   37548] = 32'h41be7969;
    ram_cell[   37549] = 32'h15b8233d;
    ram_cell[   37550] = 32'ha50af3cf;
    ram_cell[   37551] = 32'h61d29828;
    ram_cell[   37552] = 32'h753fcab6;
    ram_cell[   37553] = 32'h85be86c5;
    ram_cell[   37554] = 32'hca593fef;
    ram_cell[   37555] = 32'hd316cd5f;
    ram_cell[   37556] = 32'hd1b35f6b;
    ram_cell[   37557] = 32'h83585776;
    ram_cell[   37558] = 32'h5bd0286a;
    ram_cell[   37559] = 32'hc82c801e;
    ram_cell[   37560] = 32'h8517b871;
    ram_cell[   37561] = 32'h543ce09e;
    ram_cell[   37562] = 32'h017435e8;
    ram_cell[   37563] = 32'h7c83e2a7;
    ram_cell[   37564] = 32'h03b7bbc0;
    ram_cell[   37565] = 32'hd588f7b7;
    ram_cell[   37566] = 32'h3d89aa4f;
    ram_cell[   37567] = 32'h6aca36b6;
    ram_cell[   37568] = 32'hcb2e63e4;
    ram_cell[   37569] = 32'hf6f276b7;
    ram_cell[   37570] = 32'h91305b58;
    ram_cell[   37571] = 32'h4ee9c0b2;
    ram_cell[   37572] = 32'h84d5cfbe;
    ram_cell[   37573] = 32'hf43cc539;
    ram_cell[   37574] = 32'hd4e7d033;
    ram_cell[   37575] = 32'h23b28d37;
    ram_cell[   37576] = 32'h83ba6e40;
    ram_cell[   37577] = 32'h3bc5b4f3;
    ram_cell[   37578] = 32'hebfe5242;
    ram_cell[   37579] = 32'h154927e2;
    ram_cell[   37580] = 32'hda405e6c;
    ram_cell[   37581] = 32'ha34c6fe4;
    ram_cell[   37582] = 32'hf740a306;
    ram_cell[   37583] = 32'hf2e411ba;
    ram_cell[   37584] = 32'h99e7c516;
    ram_cell[   37585] = 32'h6bc1db40;
    ram_cell[   37586] = 32'hfb1bae48;
    ram_cell[   37587] = 32'h2f6205b8;
    ram_cell[   37588] = 32'h2c7bcdd2;
    ram_cell[   37589] = 32'h98bcc2eb;
    ram_cell[   37590] = 32'hc5b2574d;
    ram_cell[   37591] = 32'h16b320be;
    ram_cell[   37592] = 32'h8fd6cb2f;
    ram_cell[   37593] = 32'hd54e8bbc;
    ram_cell[   37594] = 32'hc562acd3;
    ram_cell[   37595] = 32'h22de4b6d;
    ram_cell[   37596] = 32'h0c41ce0a;
    ram_cell[   37597] = 32'h6112235d;
    ram_cell[   37598] = 32'h7a661895;
    ram_cell[   37599] = 32'h269573c9;
    ram_cell[   37600] = 32'hac27a5ac;
    ram_cell[   37601] = 32'he7778a7f;
    ram_cell[   37602] = 32'h27c62372;
    ram_cell[   37603] = 32'h9437f0fb;
    ram_cell[   37604] = 32'haf974cd7;
    ram_cell[   37605] = 32'h4255f225;
    ram_cell[   37606] = 32'h91628c47;
    ram_cell[   37607] = 32'hbbba8a95;
    ram_cell[   37608] = 32'h36df3c7c;
    ram_cell[   37609] = 32'h204945e8;
    ram_cell[   37610] = 32'hfd655af6;
    ram_cell[   37611] = 32'h73c750dc;
    ram_cell[   37612] = 32'h78313e1d;
    ram_cell[   37613] = 32'h8b8a2fcf;
    ram_cell[   37614] = 32'hc9177f67;
    ram_cell[   37615] = 32'he67e9868;
    ram_cell[   37616] = 32'ha58078c6;
    ram_cell[   37617] = 32'h081c764e;
    ram_cell[   37618] = 32'h6276cceb;
    ram_cell[   37619] = 32'hcc1663a6;
    ram_cell[   37620] = 32'hff87d3a0;
    ram_cell[   37621] = 32'he6c16025;
    ram_cell[   37622] = 32'ha6538438;
    ram_cell[   37623] = 32'h6ecf6a34;
    ram_cell[   37624] = 32'h893771cd;
    ram_cell[   37625] = 32'heee7bfdd;
    ram_cell[   37626] = 32'he4d2cdd3;
    ram_cell[   37627] = 32'h0c30f068;
    ram_cell[   37628] = 32'h90c7efa0;
    ram_cell[   37629] = 32'h1f966a18;
    ram_cell[   37630] = 32'h3bbfc5f3;
    ram_cell[   37631] = 32'h37b1a83a;
    ram_cell[   37632] = 32'h216950ba;
    ram_cell[   37633] = 32'h1cd18f56;
    ram_cell[   37634] = 32'h160e4f85;
    ram_cell[   37635] = 32'h4fcdb37f;
    ram_cell[   37636] = 32'hf1ae9aa7;
    ram_cell[   37637] = 32'h1f82ebec;
    ram_cell[   37638] = 32'h0064c462;
    ram_cell[   37639] = 32'h8feec71a;
    ram_cell[   37640] = 32'hfbe5aecc;
    ram_cell[   37641] = 32'h58fb9c0d;
    ram_cell[   37642] = 32'h3343b24f;
    ram_cell[   37643] = 32'hff09bfc6;
    ram_cell[   37644] = 32'hadfaa5dc;
    ram_cell[   37645] = 32'h9e003a2e;
    ram_cell[   37646] = 32'h2e8c825b;
    ram_cell[   37647] = 32'h6d928065;
    ram_cell[   37648] = 32'h4f3fc88a;
    ram_cell[   37649] = 32'ha44de7dd;
    ram_cell[   37650] = 32'h8f76e8d9;
    ram_cell[   37651] = 32'h50e73ba3;
    ram_cell[   37652] = 32'h6ef6abfd;
    ram_cell[   37653] = 32'h21d740f6;
    ram_cell[   37654] = 32'h79f7a9aa;
    ram_cell[   37655] = 32'hcce02bd7;
    ram_cell[   37656] = 32'hb96561b6;
    ram_cell[   37657] = 32'h66448750;
    ram_cell[   37658] = 32'h667df2ed;
    ram_cell[   37659] = 32'h5d431c68;
    ram_cell[   37660] = 32'hdd4c2234;
    ram_cell[   37661] = 32'h9993e900;
    ram_cell[   37662] = 32'hddb2a8cc;
    ram_cell[   37663] = 32'h5d0ef888;
    ram_cell[   37664] = 32'hc408133e;
    ram_cell[   37665] = 32'h8242ece3;
    ram_cell[   37666] = 32'h2486fe83;
    ram_cell[   37667] = 32'haed96e02;
    ram_cell[   37668] = 32'ha2d69e1e;
    ram_cell[   37669] = 32'hf8218495;
    ram_cell[   37670] = 32'hd1f926cb;
    ram_cell[   37671] = 32'h5b959540;
    ram_cell[   37672] = 32'he088b7a0;
    ram_cell[   37673] = 32'h3a83ad36;
    ram_cell[   37674] = 32'heffc8d19;
    ram_cell[   37675] = 32'ha11ceea8;
    ram_cell[   37676] = 32'hc60025b5;
    ram_cell[   37677] = 32'hf493324b;
    ram_cell[   37678] = 32'h2ad163ea;
    ram_cell[   37679] = 32'ha92cb2d2;
    ram_cell[   37680] = 32'h873af76e;
    ram_cell[   37681] = 32'h0f7e15ee;
    ram_cell[   37682] = 32'h872578d9;
    ram_cell[   37683] = 32'hf8a9fbc6;
    ram_cell[   37684] = 32'hd8caea5c;
    ram_cell[   37685] = 32'h9449a390;
    ram_cell[   37686] = 32'h1c9afb5b;
    ram_cell[   37687] = 32'h10ac7f49;
    ram_cell[   37688] = 32'h188c473c;
    ram_cell[   37689] = 32'ha1213c8f;
    ram_cell[   37690] = 32'ha53476fc;
    ram_cell[   37691] = 32'ha031d2b7;
    ram_cell[   37692] = 32'h93b6e259;
    ram_cell[   37693] = 32'hf0e8d429;
    ram_cell[   37694] = 32'h883516d3;
    ram_cell[   37695] = 32'h61bac4cf;
    ram_cell[   37696] = 32'h4ea77967;
    ram_cell[   37697] = 32'h7f95e63c;
    ram_cell[   37698] = 32'h6bbff779;
    ram_cell[   37699] = 32'hfd24c3b6;
    ram_cell[   37700] = 32'h90a00499;
    ram_cell[   37701] = 32'ha2cd3a98;
    ram_cell[   37702] = 32'h822905a4;
    ram_cell[   37703] = 32'h2b46377f;
    ram_cell[   37704] = 32'hbad85b42;
    ram_cell[   37705] = 32'h94f90698;
    ram_cell[   37706] = 32'h454ad7ec;
    ram_cell[   37707] = 32'h32d8739d;
    ram_cell[   37708] = 32'he113cdd6;
    ram_cell[   37709] = 32'hfd71ae71;
    ram_cell[   37710] = 32'h9bf123f7;
    ram_cell[   37711] = 32'h618206e7;
    ram_cell[   37712] = 32'h41f3ecdd;
    ram_cell[   37713] = 32'h17edb23a;
    ram_cell[   37714] = 32'h16ca00a3;
    ram_cell[   37715] = 32'h4fc0d589;
    ram_cell[   37716] = 32'h35a4d534;
    ram_cell[   37717] = 32'h3e0bec01;
    ram_cell[   37718] = 32'hfa430aeb;
    ram_cell[   37719] = 32'h5b23a12d;
    ram_cell[   37720] = 32'h00b9cdb9;
    ram_cell[   37721] = 32'hf02d1829;
    ram_cell[   37722] = 32'h0457ae76;
    ram_cell[   37723] = 32'hddea3b6f;
    ram_cell[   37724] = 32'h1437454d;
    ram_cell[   37725] = 32'hd937124c;
    ram_cell[   37726] = 32'h6f25927d;
    ram_cell[   37727] = 32'hedeccfa5;
    ram_cell[   37728] = 32'ha948f3f7;
    ram_cell[   37729] = 32'h820e8ad4;
    ram_cell[   37730] = 32'h00805da9;
    ram_cell[   37731] = 32'h537d9a9b;
    ram_cell[   37732] = 32'h3529e51e;
    ram_cell[   37733] = 32'ha6a5c62f;
    ram_cell[   37734] = 32'h134f2a4b;
    ram_cell[   37735] = 32'hd78e95c7;
    ram_cell[   37736] = 32'hc4c9a02b;
    ram_cell[   37737] = 32'h5ada8384;
    ram_cell[   37738] = 32'hbe01c7ea;
    ram_cell[   37739] = 32'h5151d937;
    ram_cell[   37740] = 32'h61104b11;
    ram_cell[   37741] = 32'h66e1cf17;
    ram_cell[   37742] = 32'h0c318368;
    ram_cell[   37743] = 32'h80a92b72;
    ram_cell[   37744] = 32'hbe56a8ce;
    ram_cell[   37745] = 32'hdd248cd0;
    ram_cell[   37746] = 32'hbb6e539f;
    ram_cell[   37747] = 32'h36eacb5c;
    ram_cell[   37748] = 32'h426f3303;
    ram_cell[   37749] = 32'hce6d19a4;
    ram_cell[   37750] = 32'h0f6d645f;
    ram_cell[   37751] = 32'h9af7aed6;
    ram_cell[   37752] = 32'h67d97645;
    ram_cell[   37753] = 32'h52d61f1e;
    ram_cell[   37754] = 32'h9236a7dd;
    ram_cell[   37755] = 32'h9fd5f627;
    ram_cell[   37756] = 32'hf74b9086;
    ram_cell[   37757] = 32'hd37e01f7;
    ram_cell[   37758] = 32'h0fb28531;
    ram_cell[   37759] = 32'hdee12729;
    ram_cell[   37760] = 32'h0c3b6f3a;
    ram_cell[   37761] = 32'hf7d7e637;
    ram_cell[   37762] = 32'he4701903;
    ram_cell[   37763] = 32'h9fea9d8e;
    ram_cell[   37764] = 32'h7ca8c414;
    ram_cell[   37765] = 32'h85bfb696;
    ram_cell[   37766] = 32'hb54f39f1;
    ram_cell[   37767] = 32'hbceb4bba;
    ram_cell[   37768] = 32'h788bbd4b;
    ram_cell[   37769] = 32'h539f2b34;
    ram_cell[   37770] = 32'h3b16f754;
    ram_cell[   37771] = 32'ha21a5f75;
    ram_cell[   37772] = 32'h335c9210;
    ram_cell[   37773] = 32'he38a39e7;
    ram_cell[   37774] = 32'h784ecfab;
    ram_cell[   37775] = 32'h1e02324b;
    ram_cell[   37776] = 32'hc47c3957;
    ram_cell[   37777] = 32'ha87a17bd;
    ram_cell[   37778] = 32'ha9b82d02;
    ram_cell[   37779] = 32'h57fa72d5;
    ram_cell[   37780] = 32'hec0e3130;
    ram_cell[   37781] = 32'h4bab69aa;
    ram_cell[   37782] = 32'h46aeed07;
    ram_cell[   37783] = 32'ha60a17f8;
    ram_cell[   37784] = 32'ha064c201;
    ram_cell[   37785] = 32'h360a3e56;
    ram_cell[   37786] = 32'h7a38b424;
    ram_cell[   37787] = 32'h2d399e11;
    ram_cell[   37788] = 32'h9f5e74aa;
    ram_cell[   37789] = 32'h9c46505f;
    ram_cell[   37790] = 32'h89232c73;
    ram_cell[   37791] = 32'h6ff2a1eb;
    ram_cell[   37792] = 32'h1f1f195e;
    ram_cell[   37793] = 32'hf09205a7;
    ram_cell[   37794] = 32'h84d6e7c5;
    ram_cell[   37795] = 32'h33d0962a;
    ram_cell[   37796] = 32'h397d8b31;
    ram_cell[   37797] = 32'h97a37ba2;
    ram_cell[   37798] = 32'h7694eb52;
    ram_cell[   37799] = 32'hd16d55a5;
    ram_cell[   37800] = 32'h69b97eff;
    ram_cell[   37801] = 32'he5a23e48;
    ram_cell[   37802] = 32'h5a560a44;
    ram_cell[   37803] = 32'h3ed83e6b;
    ram_cell[   37804] = 32'hec6059dd;
    ram_cell[   37805] = 32'h5df69844;
    ram_cell[   37806] = 32'he27ae952;
    ram_cell[   37807] = 32'h4026c1fb;
    ram_cell[   37808] = 32'h10a0a9c0;
    ram_cell[   37809] = 32'h00eaa104;
    ram_cell[   37810] = 32'hb4fbdd6a;
    ram_cell[   37811] = 32'hb5d8b2a6;
    ram_cell[   37812] = 32'h52836f93;
    ram_cell[   37813] = 32'hf1a0f6c4;
    ram_cell[   37814] = 32'h22b8e157;
    ram_cell[   37815] = 32'h244448b3;
    ram_cell[   37816] = 32'h7039afeb;
    ram_cell[   37817] = 32'h424c0ef4;
    ram_cell[   37818] = 32'h95b5f1ed;
    ram_cell[   37819] = 32'hf3fe9880;
    ram_cell[   37820] = 32'h9ba1ef8d;
    ram_cell[   37821] = 32'hd80cb7e9;
    ram_cell[   37822] = 32'ha2738603;
    ram_cell[   37823] = 32'h350d6299;
    ram_cell[   37824] = 32'ha4e7b8c9;
    ram_cell[   37825] = 32'hd7a9d5b3;
    ram_cell[   37826] = 32'haaff62fb;
    ram_cell[   37827] = 32'hf71e943b;
    ram_cell[   37828] = 32'h9164fb2a;
    ram_cell[   37829] = 32'h4af406fa;
    ram_cell[   37830] = 32'h9d4c47ec;
    ram_cell[   37831] = 32'hf7090f74;
    ram_cell[   37832] = 32'hb3349d08;
    ram_cell[   37833] = 32'h07ddec2a;
    ram_cell[   37834] = 32'hf999f8c6;
    ram_cell[   37835] = 32'h6a9d655d;
    ram_cell[   37836] = 32'h01badeb7;
    ram_cell[   37837] = 32'h4008b320;
    ram_cell[   37838] = 32'h0941c302;
    ram_cell[   37839] = 32'h0a810833;
    ram_cell[   37840] = 32'h5680c670;
    ram_cell[   37841] = 32'h2c7445a3;
    ram_cell[   37842] = 32'h27bf293b;
    ram_cell[   37843] = 32'hb80a8482;
    ram_cell[   37844] = 32'h7886819a;
    ram_cell[   37845] = 32'hdc11c13f;
    ram_cell[   37846] = 32'he64b3593;
    ram_cell[   37847] = 32'h023de077;
    ram_cell[   37848] = 32'hb5bf537b;
    ram_cell[   37849] = 32'h98b2bc80;
    ram_cell[   37850] = 32'hde6b67a1;
    ram_cell[   37851] = 32'h86df740f;
    ram_cell[   37852] = 32'h7f7a48f7;
    ram_cell[   37853] = 32'h01cd43d7;
    ram_cell[   37854] = 32'h2d2862bc;
    ram_cell[   37855] = 32'h0afbde27;
    ram_cell[   37856] = 32'h78eee63c;
    ram_cell[   37857] = 32'hb6536489;
    ram_cell[   37858] = 32'h25e0c571;
    ram_cell[   37859] = 32'h55b7fa92;
    ram_cell[   37860] = 32'h82b6a6bc;
    ram_cell[   37861] = 32'hb7c448f0;
    ram_cell[   37862] = 32'h6d0ada83;
    ram_cell[   37863] = 32'h92eca30e;
    ram_cell[   37864] = 32'h5bf5681b;
    ram_cell[   37865] = 32'h7a5fc2f7;
    ram_cell[   37866] = 32'h2db43896;
    ram_cell[   37867] = 32'h727dbd55;
    ram_cell[   37868] = 32'h7ea549d5;
    ram_cell[   37869] = 32'ha87ccef0;
    ram_cell[   37870] = 32'hb9d7f93b;
    ram_cell[   37871] = 32'h4652fb1c;
    ram_cell[   37872] = 32'hc48a8d68;
    ram_cell[   37873] = 32'hf66351d8;
    ram_cell[   37874] = 32'hfe1ced24;
    ram_cell[   37875] = 32'h48247824;
    ram_cell[   37876] = 32'h7793f706;
    ram_cell[   37877] = 32'h93a2bad3;
    ram_cell[   37878] = 32'hd3412a77;
    ram_cell[   37879] = 32'h8d781f16;
    ram_cell[   37880] = 32'hce907d82;
    ram_cell[   37881] = 32'h6e9cd235;
    ram_cell[   37882] = 32'hb4149a9d;
    ram_cell[   37883] = 32'h0085742c;
    ram_cell[   37884] = 32'h89070422;
    ram_cell[   37885] = 32'h54af2e80;
    ram_cell[   37886] = 32'h488b6993;
    ram_cell[   37887] = 32'h823b7a09;
    ram_cell[   37888] = 32'ha262ce57;
    ram_cell[   37889] = 32'hac680a56;
    ram_cell[   37890] = 32'h378328e5;
    ram_cell[   37891] = 32'h9e7a2847;
    ram_cell[   37892] = 32'h14510996;
    ram_cell[   37893] = 32'h0b4d69f5;
    ram_cell[   37894] = 32'hcb4c1d2c;
    ram_cell[   37895] = 32'h29402f47;
    ram_cell[   37896] = 32'h2828636b;
    ram_cell[   37897] = 32'h94bb3c4c;
    ram_cell[   37898] = 32'h66e3bc4f;
    ram_cell[   37899] = 32'h07f2cfb2;
    ram_cell[   37900] = 32'hbc356910;
    ram_cell[   37901] = 32'h6df177a9;
    ram_cell[   37902] = 32'h2bda36c5;
    ram_cell[   37903] = 32'h3a9f8f03;
    ram_cell[   37904] = 32'hc6326754;
    ram_cell[   37905] = 32'ha9cf88dd;
    ram_cell[   37906] = 32'h47260c2a;
    ram_cell[   37907] = 32'hd3513859;
    ram_cell[   37908] = 32'hf017eda8;
    ram_cell[   37909] = 32'h74a35caf;
    ram_cell[   37910] = 32'h0768a9ef;
    ram_cell[   37911] = 32'h4f1d8ced;
    ram_cell[   37912] = 32'he70ee6c3;
    ram_cell[   37913] = 32'h0291d6f7;
    ram_cell[   37914] = 32'h3f79515d;
    ram_cell[   37915] = 32'h0884134e;
    ram_cell[   37916] = 32'hb35840ac;
    ram_cell[   37917] = 32'h1d3533d3;
    ram_cell[   37918] = 32'hf50aab32;
    ram_cell[   37919] = 32'h1ec56dc3;
    ram_cell[   37920] = 32'habe29f62;
    ram_cell[   37921] = 32'h19108c86;
    ram_cell[   37922] = 32'h5a0bfa95;
    ram_cell[   37923] = 32'hfebea50e;
    ram_cell[   37924] = 32'h542787cc;
    ram_cell[   37925] = 32'hd5cb95bd;
    ram_cell[   37926] = 32'hedd20db0;
    ram_cell[   37927] = 32'h5434b914;
    ram_cell[   37928] = 32'h477d715c;
    ram_cell[   37929] = 32'h9bc3ef93;
    ram_cell[   37930] = 32'h85326f0a;
    ram_cell[   37931] = 32'he17a816d;
    ram_cell[   37932] = 32'hfe133bd6;
    ram_cell[   37933] = 32'h1dde270a;
    ram_cell[   37934] = 32'h0ab92e36;
    ram_cell[   37935] = 32'ha672d145;
    ram_cell[   37936] = 32'hc3166b7b;
    ram_cell[   37937] = 32'h124d8e12;
    ram_cell[   37938] = 32'hcbc2f289;
    ram_cell[   37939] = 32'h5e092c7c;
    ram_cell[   37940] = 32'hf16eb611;
    ram_cell[   37941] = 32'h8bd10242;
    ram_cell[   37942] = 32'hbf9c06b7;
    ram_cell[   37943] = 32'he60b8d45;
    ram_cell[   37944] = 32'hf8cbd1a8;
    ram_cell[   37945] = 32'hea53bd3e;
    ram_cell[   37946] = 32'hcb252bac;
    ram_cell[   37947] = 32'h050f55e6;
    ram_cell[   37948] = 32'h8540335c;
    ram_cell[   37949] = 32'hff12f8d7;
    ram_cell[   37950] = 32'hbbad0d62;
    ram_cell[   37951] = 32'hd03a4cf2;
    ram_cell[   37952] = 32'hb013e685;
    ram_cell[   37953] = 32'h9830e1b4;
    ram_cell[   37954] = 32'hc17e8129;
    ram_cell[   37955] = 32'h24eaf3ea;
    ram_cell[   37956] = 32'h069a9195;
    ram_cell[   37957] = 32'hcd17aa1d;
    ram_cell[   37958] = 32'h331915d2;
    ram_cell[   37959] = 32'hb5f2d01a;
    ram_cell[   37960] = 32'hb88c6d55;
    ram_cell[   37961] = 32'h2571bc64;
    ram_cell[   37962] = 32'h7117a88c;
    ram_cell[   37963] = 32'he7cdb283;
    ram_cell[   37964] = 32'hb79c670b;
    ram_cell[   37965] = 32'hf61002a4;
    ram_cell[   37966] = 32'h6ebf38c7;
    ram_cell[   37967] = 32'hb09ef42f;
    ram_cell[   37968] = 32'h753707c5;
    ram_cell[   37969] = 32'he50cb39a;
    ram_cell[   37970] = 32'h295c3777;
    ram_cell[   37971] = 32'hcb99f58c;
    ram_cell[   37972] = 32'h86ce8356;
    ram_cell[   37973] = 32'h8bf07753;
    ram_cell[   37974] = 32'h45e32bca;
    ram_cell[   37975] = 32'h84cd19d2;
    ram_cell[   37976] = 32'h747237bf;
    ram_cell[   37977] = 32'h281ae74e;
    ram_cell[   37978] = 32'h880f22c5;
    ram_cell[   37979] = 32'h10e7a5e2;
    ram_cell[   37980] = 32'h71845171;
    ram_cell[   37981] = 32'h6253965f;
    ram_cell[   37982] = 32'he50e330f;
    ram_cell[   37983] = 32'h306f4826;
    ram_cell[   37984] = 32'he8255c00;
    ram_cell[   37985] = 32'h8eef8aef;
    ram_cell[   37986] = 32'h6ed97ae4;
    ram_cell[   37987] = 32'hce6ac351;
    ram_cell[   37988] = 32'hfca1bbbf;
    ram_cell[   37989] = 32'h780c0143;
    ram_cell[   37990] = 32'h225ba87f;
    ram_cell[   37991] = 32'hcf8f907e;
    ram_cell[   37992] = 32'h6134926d;
    ram_cell[   37993] = 32'hebe3022a;
    ram_cell[   37994] = 32'hb1f474b1;
    ram_cell[   37995] = 32'hb8e79e5e;
    ram_cell[   37996] = 32'hd0af29f5;
    ram_cell[   37997] = 32'hb4d84b89;
    ram_cell[   37998] = 32'h6a63b059;
    ram_cell[   37999] = 32'h1390bb1e;
    ram_cell[   38000] = 32'h9dac0235;
    ram_cell[   38001] = 32'h6ec0648a;
    ram_cell[   38002] = 32'ha70ee9dc;
    ram_cell[   38003] = 32'hb8325874;
    ram_cell[   38004] = 32'hdbad322b;
    ram_cell[   38005] = 32'h8bea0000;
    ram_cell[   38006] = 32'h1cf4aaa5;
    ram_cell[   38007] = 32'haa29309e;
    ram_cell[   38008] = 32'hf1a1b12d;
    ram_cell[   38009] = 32'h46595d2f;
    ram_cell[   38010] = 32'h313e5bec;
    ram_cell[   38011] = 32'hca2e2032;
    ram_cell[   38012] = 32'h11e76d05;
    ram_cell[   38013] = 32'h6d649b87;
    ram_cell[   38014] = 32'h686c4603;
    ram_cell[   38015] = 32'h34a80381;
    ram_cell[   38016] = 32'he0d7fb49;
    ram_cell[   38017] = 32'hdb5e762a;
    ram_cell[   38018] = 32'h295fc490;
    ram_cell[   38019] = 32'h80bb28e8;
    ram_cell[   38020] = 32'heaeb1087;
    ram_cell[   38021] = 32'h18f703d6;
    ram_cell[   38022] = 32'h9bb86118;
    ram_cell[   38023] = 32'h08c2fb54;
    ram_cell[   38024] = 32'h2fd9fef4;
    ram_cell[   38025] = 32'hc82e9817;
    ram_cell[   38026] = 32'h176e6f27;
    ram_cell[   38027] = 32'hf1cb118c;
    ram_cell[   38028] = 32'h691fc4a0;
    ram_cell[   38029] = 32'h75fe562d;
    ram_cell[   38030] = 32'hf4761ed3;
    ram_cell[   38031] = 32'h1d9ccefd;
    ram_cell[   38032] = 32'h19576bca;
    ram_cell[   38033] = 32'hdaec81b7;
    ram_cell[   38034] = 32'ha7322433;
    ram_cell[   38035] = 32'habc9c252;
    ram_cell[   38036] = 32'h49230c3e;
    ram_cell[   38037] = 32'hb928fe88;
    ram_cell[   38038] = 32'h442265c5;
    ram_cell[   38039] = 32'hba4f90ed;
    ram_cell[   38040] = 32'h482a4a4e;
    ram_cell[   38041] = 32'h3e76d3ec;
    ram_cell[   38042] = 32'h29d2fe09;
    ram_cell[   38043] = 32'hc271995c;
    ram_cell[   38044] = 32'h8728f0a6;
    ram_cell[   38045] = 32'h5abd958b;
    ram_cell[   38046] = 32'h6d442aea;
    ram_cell[   38047] = 32'ha794a1da;
    ram_cell[   38048] = 32'hfc837e4e;
    ram_cell[   38049] = 32'h1ac98255;
    ram_cell[   38050] = 32'h37b0f9c7;
    ram_cell[   38051] = 32'h4639160c;
    ram_cell[   38052] = 32'h308fbbe6;
    ram_cell[   38053] = 32'h6b46d787;
    ram_cell[   38054] = 32'h4beec2b5;
    ram_cell[   38055] = 32'h1f1f71f3;
    ram_cell[   38056] = 32'h178d2596;
    ram_cell[   38057] = 32'h18be9650;
    ram_cell[   38058] = 32'haadabb1d;
    ram_cell[   38059] = 32'h94cf16ee;
    ram_cell[   38060] = 32'h030ea7a2;
    ram_cell[   38061] = 32'h7ba4ca5f;
    ram_cell[   38062] = 32'h90755404;
    ram_cell[   38063] = 32'hcd44e343;
    ram_cell[   38064] = 32'h7be7b0fa;
    ram_cell[   38065] = 32'h7d35bc2b;
    ram_cell[   38066] = 32'he741b64c;
    ram_cell[   38067] = 32'h77edab63;
    ram_cell[   38068] = 32'hecb6a11a;
    ram_cell[   38069] = 32'hb0663153;
    ram_cell[   38070] = 32'hf66a84c8;
    ram_cell[   38071] = 32'hef18b5c4;
    ram_cell[   38072] = 32'h96d58814;
    ram_cell[   38073] = 32'h282442a5;
    ram_cell[   38074] = 32'he4241dec;
    ram_cell[   38075] = 32'ha59c539f;
    ram_cell[   38076] = 32'hbe3aa14b;
    ram_cell[   38077] = 32'hcbf2636e;
    ram_cell[   38078] = 32'heed41c17;
    ram_cell[   38079] = 32'haa8009c9;
    ram_cell[   38080] = 32'ha1909f9d;
    ram_cell[   38081] = 32'h36636a8e;
    ram_cell[   38082] = 32'h6a62be72;
    ram_cell[   38083] = 32'hed1a671b;
    ram_cell[   38084] = 32'hec52ef20;
    ram_cell[   38085] = 32'h858758b3;
    ram_cell[   38086] = 32'h05be6539;
    ram_cell[   38087] = 32'h94b1ec85;
    ram_cell[   38088] = 32'hd90f6815;
    ram_cell[   38089] = 32'he40137cf;
    ram_cell[   38090] = 32'h492201a8;
    ram_cell[   38091] = 32'h4d0516a3;
    ram_cell[   38092] = 32'hade13ea8;
    ram_cell[   38093] = 32'h78010310;
    ram_cell[   38094] = 32'h6e613c55;
    ram_cell[   38095] = 32'hdaedd884;
    ram_cell[   38096] = 32'he7de33af;
    ram_cell[   38097] = 32'h355f80b1;
    ram_cell[   38098] = 32'h562c0282;
    ram_cell[   38099] = 32'hd804e3b2;
    ram_cell[   38100] = 32'h5b1b1433;
    ram_cell[   38101] = 32'hf1c5cd90;
    ram_cell[   38102] = 32'hac9836e5;
    ram_cell[   38103] = 32'h9d3c3bfd;
    ram_cell[   38104] = 32'hbf1d570e;
    ram_cell[   38105] = 32'hf60c05e8;
    ram_cell[   38106] = 32'hda04573f;
    ram_cell[   38107] = 32'h28481aeb;
    ram_cell[   38108] = 32'h7907d276;
    ram_cell[   38109] = 32'h9be8f015;
    ram_cell[   38110] = 32'h7c04a8be;
    ram_cell[   38111] = 32'ha768d3ea;
    ram_cell[   38112] = 32'h6abaefbe;
    ram_cell[   38113] = 32'h5a8b37be;
    ram_cell[   38114] = 32'hcf3cb9f7;
    ram_cell[   38115] = 32'h7d1b0fe9;
    ram_cell[   38116] = 32'h64688a1e;
    ram_cell[   38117] = 32'hbb7d1f0e;
    ram_cell[   38118] = 32'hc86e7927;
    ram_cell[   38119] = 32'he613f008;
    ram_cell[   38120] = 32'h2e2b87f3;
    ram_cell[   38121] = 32'hd5c19dc1;
    ram_cell[   38122] = 32'ha50a88e3;
    ram_cell[   38123] = 32'h588998cf;
    ram_cell[   38124] = 32'hce22e8f1;
    ram_cell[   38125] = 32'h80057852;
    ram_cell[   38126] = 32'h06a3880b;
    ram_cell[   38127] = 32'hc0d603cf;
    ram_cell[   38128] = 32'h5caeb5b5;
    ram_cell[   38129] = 32'hbcb9ef76;
    ram_cell[   38130] = 32'h046242d7;
    ram_cell[   38131] = 32'h7a01303c;
    ram_cell[   38132] = 32'hc12d5851;
    ram_cell[   38133] = 32'hfb163468;
    ram_cell[   38134] = 32'hb3f53ac1;
    ram_cell[   38135] = 32'h517ce1cc;
    ram_cell[   38136] = 32'h18f56b88;
    ram_cell[   38137] = 32'h2194e6e2;
    ram_cell[   38138] = 32'hcb3d01ad;
    ram_cell[   38139] = 32'h975a5e05;
    ram_cell[   38140] = 32'h42eea67f;
    ram_cell[   38141] = 32'h90ae13a1;
    ram_cell[   38142] = 32'h563e43a9;
    ram_cell[   38143] = 32'h2d3df696;
    ram_cell[   38144] = 32'hc51cbc0f;
    ram_cell[   38145] = 32'h445bf8a0;
    ram_cell[   38146] = 32'hf9fa0ad6;
    ram_cell[   38147] = 32'h5c1c188b;
    ram_cell[   38148] = 32'h60586997;
    ram_cell[   38149] = 32'h2679c6ff;
    ram_cell[   38150] = 32'h3ab09c5e;
    ram_cell[   38151] = 32'hacdde2ea;
    ram_cell[   38152] = 32'h5dff77b7;
    ram_cell[   38153] = 32'h1863c162;
    ram_cell[   38154] = 32'hf9be03a4;
    ram_cell[   38155] = 32'h4fac8d91;
    ram_cell[   38156] = 32'h771b956d;
    ram_cell[   38157] = 32'h28eb6d63;
    ram_cell[   38158] = 32'hea9162ac;
    ram_cell[   38159] = 32'h60b5b045;
    ram_cell[   38160] = 32'ha54a5381;
    ram_cell[   38161] = 32'h8a575b21;
    ram_cell[   38162] = 32'h0d0404d5;
    ram_cell[   38163] = 32'h61f4ae9a;
    ram_cell[   38164] = 32'h17637e47;
    ram_cell[   38165] = 32'hf82ea2c0;
    ram_cell[   38166] = 32'h3024c535;
    ram_cell[   38167] = 32'h5f826b69;
    ram_cell[   38168] = 32'h2011b562;
    ram_cell[   38169] = 32'h76f060af;
    ram_cell[   38170] = 32'hd5a32279;
    ram_cell[   38171] = 32'h06cb748e;
    ram_cell[   38172] = 32'h1fe64336;
    ram_cell[   38173] = 32'hd0e8cd90;
    ram_cell[   38174] = 32'hf5eb88ff;
    ram_cell[   38175] = 32'hab03fecd;
    ram_cell[   38176] = 32'h8bba2116;
    ram_cell[   38177] = 32'hba57b4b3;
    ram_cell[   38178] = 32'hd47ca5e0;
    ram_cell[   38179] = 32'h998b553c;
    ram_cell[   38180] = 32'h9932acce;
    ram_cell[   38181] = 32'hacc29dda;
    ram_cell[   38182] = 32'h93f6f52f;
    ram_cell[   38183] = 32'h1dbbd362;
    ram_cell[   38184] = 32'hc7d3ea9f;
    ram_cell[   38185] = 32'h5d1cf59e;
    ram_cell[   38186] = 32'h6a475d13;
    ram_cell[   38187] = 32'hcbda9c05;
    ram_cell[   38188] = 32'he77a9b44;
    ram_cell[   38189] = 32'h902c1f3c;
    ram_cell[   38190] = 32'h79c64a3f;
    ram_cell[   38191] = 32'h9b2baf0b;
    ram_cell[   38192] = 32'h3f7b783a;
    ram_cell[   38193] = 32'h1e651472;
    ram_cell[   38194] = 32'hd58572e6;
    ram_cell[   38195] = 32'h32443424;
    ram_cell[   38196] = 32'hdaa1f4dc;
    ram_cell[   38197] = 32'h86f1b242;
    ram_cell[   38198] = 32'h243631ac;
    ram_cell[   38199] = 32'h095d9356;
    ram_cell[   38200] = 32'hdd81b7d7;
    ram_cell[   38201] = 32'h3ecb8911;
    ram_cell[   38202] = 32'hba226453;
    ram_cell[   38203] = 32'h6dcf7a4e;
    ram_cell[   38204] = 32'h86e564d3;
    ram_cell[   38205] = 32'h7568605e;
    ram_cell[   38206] = 32'hc72238ec;
    ram_cell[   38207] = 32'h2e4ec95a;
    ram_cell[   38208] = 32'h84bafc6d;
    ram_cell[   38209] = 32'h34b9e234;
    ram_cell[   38210] = 32'h48859b16;
    ram_cell[   38211] = 32'h42ec28c5;
    ram_cell[   38212] = 32'h3b079f79;
    ram_cell[   38213] = 32'ha28503f4;
    ram_cell[   38214] = 32'ha86369c7;
    ram_cell[   38215] = 32'hda6db661;
    ram_cell[   38216] = 32'h33e5d1ed;
    ram_cell[   38217] = 32'h71fa5fdf;
    ram_cell[   38218] = 32'h47ea7060;
    ram_cell[   38219] = 32'h084a0664;
    ram_cell[   38220] = 32'he9803f25;
    ram_cell[   38221] = 32'h7697beab;
    ram_cell[   38222] = 32'h4437f627;
    ram_cell[   38223] = 32'ha2721b59;
    ram_cell[   38224] = 32'h404ae8c1;
    ram_cell[   38225] = 32'h4b5bca59;
    ram_cell[   38226] = 32'h1095092d;
    ram_cell[   38227] = 32'h4be44f94;
    ram_cell[   38228] = 32'h8c1deb06;
    ram_cell[   38229] = 32'hadc8542e;
    ram_cell[   38230] = 32'h766c5bec;
    ram_cell[   38231] = 32'h1f38bc23;
    ram_cell[   38232] = 32'h5f27365a;
    ram_cell[   38233] = 32'hce7e6afe;
    ram_cell[   38234] = 32'h840b708e;
    ram_cell[   38235] = 32'hb27006af;
    ram_cell[   38236] = 32'hb4562e91;
    ram_cell[   38237] = 32'ha6bf4302;
    ram_cell[   38238] = 32'h4a945ee9;
    ram_cell[   38239] = 32'h5f9cb67e;
    ram_cell[   38240] = 32'hfcb51eba;
    ram_cell[   38241] = 32'h1042e7fc;
    ram_cell[   38242] = 32'h49d76cf7;
    ram_cell[   38243] = 32'he4e4e877;
    ram_cell[   38244] = 32'h93f7ace7;
    ram_cell[   38245] = 32'hc3e96884;
    ram_cell[   38246] = 32'h87bf8c3a;
    ram_cell[   38247] = 32'h466285e5;
    ram_cell[   38248] = 32'hfa0e90de;
    ram_cell[   38249] = 32'h90419aea;
    ram_cell[   38250] = 32'h5d947ef4;
    ram_cell[   38251] = 32'h1ee81aed;
    ram_cell[   38252] = 32'hd94e7b5e;
    ram_cell[   38253] = 32'h8acf14ac;
    ram_cell[   38254] = 32'he24d5638;
    ram_cell[   38255] = 32'he3f2bb2f;
    ram_cell[   38256] = 32'h56d245c7;
    ram_cell[   38257] = 32'hb661be32;
    ram_cell[   38258] = 32'h943ddb2c;
    ram_cell[   38259] = 32'h5983b1ec;
    ram_cell[   38260] = 32'h2524fdda;
    ram_cell[   38261] = 32'h7ac2cc72;
    ram_cell[   38262] = 32'h25b4f436;
    ram_cell[   38263] = 32'hd3aa1d2a;
    ram_cell[   38264] = 32'hf42aa805;
    ram_cell[   38265] = 32'h2060214a;
    ram_cell[   38266] = 32'h8c14bd4a;
    ram_cell[   38267] = 32'h24d98a74;
    ram_cell[   38268] = 32'hf34c6710;
    ram_cell[   38269] = 32'he6122062;
    ram_cell[   38270] = 32'hdf4f61d3;
    ram_cell[   38271] = 32'h17d95cc1;
    ram_cell[   38272] = 32'ha66ad7f3;
    ram_cell[   38273] = 32'ha305b5f5;
    ram_cell[   38274] = 32'h2e96088a;
    ram_cell[   38275] = 32'h5e75614e;
    ram_cell[   38276] = 32'h0c1d4315;
    ram_cell[   38277] = 32'h27944cb8;
    ram_cell[   38278] = 32'h32ae72c4;
    ram_cell[   38279] = 32'h5342c66b;
    ram_cell[   38280] = 32'hc0ad8d63;
    ram_cell[   38281] = 32'he95d9c2c;
    ram_cell[   38282] = 32'h23b3662f;
    ram_cell[   38283] = 32'h9511a007;
    ram_cell[   38284] = 32'h6858f6c9;
    ram_cell[   38285] = 32'hb3e0c1f0;
    ram_cell[   38286] = 32'h86ddb90c;
    ram_cell[   38287] = 32'hf2695935;
    ram_cell[   38288] = 32'h9bef08ed;
    ram_cell[   38289] = 32'hf6dcc746;
    ram_cell[   38290] = 32'h4edf298c;
    ram_cell[   38291] = 32'hb652505d;
    ram_cell[   38292] = 32'hfefeb3d9;
    ram_cell[   38293] = 32'heb0c4015;
    ram_cell[   38294] = 32'h5cce2d4d;
    ram_cell[   38295] = 32'hab9db028;
    ram_cell[   38296] = 32'hcf176223;
    ram_cell[   38297] = 32'h8e8df202;
    ram_cell[   38298] = 32'h0f0521ea;
    ram_cell[   38299] = 32'h6324b2ac;
    ram_cell[   38300] = 32'hc59800bd;
    ram_cell[   38301] = 32'h850cd22a;
    ram_cell[   38302] = 32'hf588b146;
    ram_cell[   38303] = 32'h23e2685b;
    ram_cell[   38304] = 32'h49555f51;
    ram_cell[   38305] = 32'h9e5dc06b;
    ram_cell[   38306] = 32'hefb45916;
    ram_cell[   38307] = 32'hd44ffd71;
    ram_cell[   38308] = 32'h27c9149a;
    ram_cell[   38309] = 32'hccb1b53a;
    ram_cell[   38310] = 32'h6eb1bb37;
    ram_cell[   38311] = 32'h5dc772ed;
    ram_cell[   38312] = 32'h30a3d99a;
    ram_cell[   38313] = 32'h37350f16;
    ram_cell[   38314] = 32'h5d7a660c;
    ram_cell[   38315] = 32'h7d245ffb;
    ram_cell[   38316] = 32'hfc9e4fb9;
    ram_cell[   38317] = 32'hbcb3959e;
    ram_cell[   38318] = 32'h031b8925;
    ram_cell[   38319] = 32'h21e0e443;
    ram_cell[   38320] = 32'hff4379ae;
    ram_cell[   38321] = 32'h1a2277dd;
    ram_cell[   38322] = 32'h9862a6f3;
    ram_cell[   38323] = 32'ha8eb72e6;
    ram_cell[   38324] = 32'h954b1620;
    ram_cell[   38325] = 32'hbd93fc29;
    ram_cell[   38326] = 32'hba69c13a;
    ram_cell[   38327] = 32'hedbb91de;
    ram_cell[   38328] = 32'hdec71aca;
    ram_cell[   38329] = 32'h7ccba26f;
    ram_cell[   38330] = 32'hd82924cd;
    ram_cell[   38331] = 32'hc4021987;
    ram_cell[   38332] = 32'hde5a2b68;
    ram_cell[   38333] = 32'h54a9d692;
    ram_cell[   38334] = 32'he1d12fd9;
    ram_cell[   38335] = 32'h13f30ecf;
    ram_cell[   38336] = 32'h66d8ba26;
    ram_cell[   38337] = 32'hb2aa18cb;
    ram_cell[   38338] = 32'h17b6fbec;
    ram_cell[   38339] = 32'h224b3c24;
    ram_cell[   38340] = 32'h34ecd0ae;
    ram_cell[   38341] = 32'h80541101;
    ram_cell[   38342] = 32'ha03b377c;
    ram_cell[   38343] = 32'hed2fc8b0;
    ram_cell[   38344] = 32'hd07b71b2;
    ram_cell[   38345] = 32'h08345551;
    ram_cell[   38346] = 32'h11380746;
    ram_cell[   38347] = 32'hc4a13072;
    ram_cell[   38348] = 32'h23cadb8e;
    ram_cell[   38349] = 32'h189bea0f;
    ram_cell[   38350] = 32'h993a849a;
    ram_cell[   38351] = 32'h70bf7b6b;
    ram_cell[   38352] = 32'hbf458304;
    ram_cell[   38353] = 32'hcf939acf;
    ram_cell[   38354] = 32'h80275691;
    ram_cell[   38355] = 32'ha3df62af;
    ram_cell[   38356] = 32'h0e53eae8;
    ram_cell[   38357] = 32'hb9857111;
    ram_cell[   38358] = 32'hd7b9f8d5;
    ram_cell[   38359] = 32'h9b84db43;
    ram_cell[   38360] = 32'h3dc1eb1f;
    ram_cell[   38361] = 32'hf98ea32f;
    ram_cell[   38362] = 32'h5a79fa7b;
    ram_cell[   38363] = 32'hbb8555d3;
    ram_cell[   38364] = 32'h7cd87929;
    ram_cell[   38365] = 32'h78339631;
    ram_cell[   38366] = 32'h1f19f9e1;
    ram_cell[   38367] = 32'hadaa6c76;
    ram_cell[   38368] = 32'hf6a0886c;
    ram_cell[   38369] = 32'h544066c8;
    ram_cell[   38370] = 32'hcc98e111;
    ram_cell[   38371] = 32'h00cf84ba;
    ram_cell[   38372] = 32'he1905fba;
    ram_cell[   38373] = 32'h2bcc6503;
    ram_cell[   38374] = 32'h8593b2f9;
    ram_cell[   38375] = 32'h67fbbdf8;
    ram_cell[   38376] = 32'h8c0609af;
    ram_cell[   38377] = 32'h00b9a6d7;
    ram_cell[   38378] = 32'h9df44908;
    ram_cell[   38379] = 32'h5483d950;
    ram_cell[   38380] = 32'h7411a3e7;
    ram_cell[   38381] = 32'h9270baf1;
    ram_cell[   38382] = 32'h588352dc;
    ram_cell[   38383] = 32'h7b32e152;
    ram_cell[   38384] = 32'h1f9e8d34;
    ram_cell[   38385] = 32'hbd51b451;
    ram_cell[   38386] = 32'hb551eb01;
    ram_cell[   38387] = 32'h333a616e;
    ram_cell[   38388] = 32'h40b5c782;
    ram_cell[   38389] = 32'h24fbc657;
    ram_cell[   38390] = 32'h830eeb47;
    ram_cell[   38391] = 32'h60a8a78d;
    ram_cell[   38392] = 32'hd1df8658;
    ram_cell[   38393] = 32'h82f2aa99;
    ram_cell[   38394] = 32'he53d82ff;
    ram_cell[   38395] = 32'h6ee98f94;
    ram_cell[   38396] = 32'h8939f6a0;
    ram_cell[   38397] = 32'hbef410f8;
    ram_cell[   38398] = 32'h4e83e061;
    ram_cell[   38399] = 32'he5194f1a;
    ram_cell[   38400] = 32'hbbe54771;
    ram_cell[   38401] = 32'h91f57231;
    ram_cell[   38402] = 32'hdad8ebe7;
    ram_cell[   38403] = 32'he44d881c;
    ram_cell[   38404] = 32'h790942de;
    ram_cell[   38405] = 32'h6773ce97;
    ram_cell[   38406] = 32'hdff21ea0;
    ram_cell[   38407] = 32'h762a9a5c;
    ram_cell[   38408] = 32'hf7465af0;
    ram_cell[   38409] = 32'h7bf95a3f;
    ram_cell[   38410] = 32'h84fabba4;
    ram_cell[   38411] = 32'hdec38f57;
    ram_cell[   38412] = 32'ha32bf2cb;
    ram_cell[   38413] = 32'hc1fbb858;
    ram_cell[   38414] = 32'hef267a63;
    ram_cell[   38415] = 32'he23f2aed;
    ram_cell[   38416] = 32'he4df7973;
    ram_cell[   38417] = 32'hdf57b895;
    ram_cell[   38418] = 32'he4c0f248;
    ram_cell[   38419] = 32'h0e203daa;
    ram_cell[   38420] = 32'h8afc528a;
    ram_cell[   38421] = 32'h11c1936f;
    ram_cell[   38422] = 32'hc9954227;
    ram_cell[   38423] = 32'h5ebb85da;
    ram_cell[   38424] = 32'h193dd8e1;
    ram_cell[   38425] = 32'h83a33463;
    ram_cell[   38426] = 32'hb7e6103a;
    ram_cell[   38427] = 32'hbad7ad73;
    ram_cell[   38428] = 32'h723299af;
    ram_cell[   38429] = 32'h606cb2ee;
    ram_cell[   38430] = 32'h51821980;
    ram_cell[   38431] = 32'h6e8fb85f;
    ram_cell[   38432] = 32'h8c4b937e;
    ram_cell[   38433] = 32'h30947222;
    ram_cell[   38434] = 32'h01026006;
    ram_cell[   38435] = 32'h6e48ab22;
    ram_cell[   38436] = 32'hdfccdfbe;
    ram_cell[   38437] = 32'hb51b6406;
    ram_cell[   38438] = 32'h9b730302;
    ram_cell[   38439] = 32'h5a610c1f;
    ram_cell[   38440] = 32'hee0394a0;
    ram_cell[   38441] = 32'h12d92ad7;
    ram_cell[   38442] = 32'hf7948bab;
    ram_cell[   38443] = 32'hb230f77c;
    ram_cell[   38444] = 32'h338c82b6;
    ram_cell[   38445] = 32'h610ff339;
    ram_cell[   38446] = 32'h9d3bebf2;
    ram_cell[   38447] = 32'h2d07bcb4;
    ram_cell[   38448] = 32'h58baef8e;
    ram_cell[   38449] = 32'h97da1608;
    ram_cell[   38450] = 32'h8652aa6d;
    ram_cell[   38451] = 32'hcdead085;
    ram_cell[   38452] = 32'h1dbacae6;
    ram_cell[   38453] = 32'hcf9ca1e3;
    ram_cell[   38454] = 32'h9f7dbc6f;
    ram_cell[   38455] = 32'ha34c7016;
    ram_cell[   38456] = 32'h4da05dc7;
    ram_cell[   38457] = 32'h04fac65e;
    ram_cell[   38458] = 32'h0274f93c;
    ram_cell[   38459] = 32'he62f7d66;
    ram_cell[   38460] = 32'h17becaaa;
    ram_cell[   38461] = 32'h5cf4da6e;
    ram_cell[   38462] = 32'h4edf1577;
    ram_cell[   38463] = 32'h803e6b29;
    ram_cell[   38464] = 32'h9c60da63;
    ram_cell[   38465] = 32'hc1493c1f;
    ram_cell[   38466] = 32'ha069eac7;
    ram_cell[   38467] = 32'h93de39cc;
    ram_cell[   38468] = 32'hefbbb73a;
    ram_cell[   38469] = 32'h97d84758;
    ram_cell[   38470] = 32'hcd357f5f;
    ram_cell[   38471] = 32'h29117c4b;
    ram_cell[   38472] = 32'hd0f39435;
    ram_cell[   38473] = 32'heb026a0b;
    ram_cell[   38474] = 32'h3d91a340;
    ram_cell[   38475] = 32'h74b94b35;
    ram_cell[   38476] = 32'h0b2f6e26;
    ram_cell[   38477] = 32'h8e72036e;
    ram_cell[   38478] = 32'hed7eaf6d;
    ram_cell[   38479] = 32'hc1297452;
    ram_cell[   38480] = 32'h9957e1b0;
    ram_cell[   38481] = 32'h920c640b;
    ram_cell[   38482] = 32'h9251f9f7;
    ram_cell[   38483] = 32'hb8392b9e;
    ram_cell[   38484] = 32'hde04f35b;
    ram_cell[   38485] = 32'ha8630eb9;
    ram_cell[   38486] = 32'h0d997ee7;
    ram_cell[   38487] = 32'h0be94d36;
    ram_cell[   38488] = 32'h657fdc5b;
    ram_cell[   38489] = 32'h959b69de;
    ram_cell[   38490] = 32'hc391fb53;
    ram_cell[   38491] = 32'he4265b2a;
    ram_cell[   38492] = 32'hfceeee21;
    ram_cell[   38493] = 32'h1263aa33;
    ram_cell[   38494] = 32'h2b73a77b;
    ram_cell[   38495] = 32'h0c45c978;
    ram_cell[   38496] = 32'ha89a1e93;
    ram_cell[   38497] = 32'h992fb7ef;
    ram_cell[   38498] = 32'h80068520;
    ram_cell[   38499] = 32'hdaf128ca;
    ram_cell[   38500] = 32'h2b26e03b;
    ram_cell[   38501] = 32'hecc93aab;
    ram_cell[   38502] = 32'h7784b774;
    ram_cell[   38503] = 32'ha2009a87;
    ram_cell[   38504] = 32'hbed155e0;
    ram_cell[   38505] = 32'ha4aeb337;
    ram_cell[   38506] = 32'hb9750ecc;
    ram_cell[   38507] = 32'hdfe35679;
    ram_cell[   38508] = 32'hc5f085c8;
    ram_cell[   38509] = 32'h1b4120a3;
    ram_cell[   38510] = 32'hfee953eb;
    ram_cell[   38511] = 32'h23109537;
    ram_cell[   38512] = 32'hd8ebb5ca;
    ram_cell[   38513] = 32'h94acd8fc;
    ram_cell[   38514] = 32'h9f127a52;
    ram_cell[   38515] = 32'hda42e52f;
    ram_cell[   38516] = 32'hec46f4a8;
    ram_cell[   38517] = 32'hdc98674b;
    ram_cell[   38518] = 32'h2f0d2414;
    ram_cell[   38519] = 32'hedbc65c2;
    ram_cell[   38520] = 32'h74487ee0;
    ram_cell[   38521] = 32'h3567baec;
    ram_cell[   38522] = 32'hd802edb0;
    ram_cell[   38523] = 32'h022b9194;
    ram_cell[   38524] = 32'h90bd7729;
    ram_cell[   38525] = 32'hde37ab97;
    ram_cell[   38526] = 32'h3d44c329;
    ram_cell[   38527] = 32'h951dc3ff;
    ram_cell[   38528] = 32'h110f639e;
    ram_cell[   38529] = 32'hf182e9e0;
    ram_cell[   38530] = 32'h4c589deb;
    ram_cell[   38531] = 32'h936a6aa7;
    ram_cell[   38532] = 32'h6385ccaf;
    ram_cell[   38533] = 32'h7129696a;
    ram_cell[   38534] = 32'hafa0ad13;
    ram_cell[   38535] = 32'h6446c75b;
    ram_cell[   38536] = 32'hf7e6f923;
    ram_cell[   38537] = 32'hf4e76348;
    ram_cell[   38538] = 32'h4e0a9c5d;
    ram_cell[   38539] = 32'h73a888a2;
    ram_cell[   38540] = 32'ha12096fd;
    ram_cell[   38541] = 32'h8195bc5b;
    ram_cell[   38542] = 32'h81b71026;
    ram_cell[   38543] = 32'h724be47f;
    ram_cell[   38544] = 32'hd0674db7;
    ram_cell[   38545] = 32'h9dd390dd;
    ram_cell[   38546] = 32'h61333798;
    ram_cell[   38547] = 32'hf7e280f3;
    ram_cell[   38548] = 32'h89df7191;
    ram_cell[   38549] = 32'h2f5ce393;
    ram_cell[   38550] = 32'hb00704e9;
    ram_cell[   38551] = 32'h97ee04ce;
    ram_cell[   38552] = 32'h75068607;
    ram_cell[   38553] = 32'h637671a8;
    ram_cell[   38554] = 32'hc7120378;
    ram_cell[   38555] = 32'h83c68779;
    ram_cell[   38556] = 32'hc3ea11da;
    ram_cell[   38557] = 32'h411b44c1;
    ram_cell[   38558] = 32'h9705abff;
    ram_cell[   38559] = 32'hd0c9a577;
    ram_cell[   38560] = 32'h44fddb02;
    ram_cell[   38561] = 32'h60342d2a;
    ram_cell[   38562] = 32'h9d824afd;
    ram_cell[   38563] = 32'hf2da77c9;
    ram_cell[   38564] = 32'hdb9b8e5b;
    ram_cell[   38565] = 32'h15bd19fc;
    ram_cell[   38566] = 32'h404f8538;
    ram_cell[   38567] = 32'ha43823a2;
    ram_cell[   38568] = 32'h1691a43a;
    ram_cell[   38569] = 32'hb2a0c8f9;
    ram_cell[   38570] = 32'h9b6890c3;
    ram_cell[   38571] = 32'h7b1ce2a5;
    ram_cell[   38572] = 32'h54d3afd6;
    ram_cell[   38573] = 32'hd19e0839;
    ram_cell[   38574] = 32'he8345e53;
    ram_cell[   38575] = 32'h6e604362;
    ram_cell[   38576] = 32'h2e000ab5;
    ram_cell[   38577] = 32'h1a63f661;
    ram_cell[   38578] = 32'h0146374e;
    ram_cell[   38579] = 32'h5826d93d;
    ram_cell[   38580] = 32'h5bfb7a6d;
    ram_cell[   38581] = 32'he16a2ec8;
    ram_cell[   38582] = 32'h7571a558;
    ram_cell[   38583] = 32'h9cfc9579;
    ram_cell[   38584] = 32'h338f3d0f;
    ram_cell[   38585] = 32'h916656cd;
    ram_cell[   38586] = 32'h0bcba8d5;
    ram_cell[   38587] = 32'h4fbab61b;
    ram_cell[   38588] = 32'h16d4b6cf;
    ram_cell[   38589] = 32'hbaca7b21;
    ram_cell[   38590] = 32'hb96db2a1;
    ram_cell[   38591] = 32'hababee18;
    ram_cell[   38592] = 32'h2c25b09e;
    ram_cell[   38593] = 32'hcb036d2a;
    ram_cell[   38594] = 32'ha5d4ccc0;
    ram_cell[   38595] = 32'hdb5a71c8;
    ram_cell[   38596] = 32'hb18aaeae;
    ram_cell[   38597] = 32'h04861494;
    ram_cell[   38598] = 32'hb1ac40a0;
    ram_cell[   38599] = 32'h21b16010;
    ram_cell[   38600] = 32'hbbe821b8;
    ram_cell[   38601] = 32'hd4f62c64;
    ram_cell[   38602] = 32'h6b69e328;
    ram_cell[   38603] = 32'h4902f669;
    ram_cell[   38604] = 32'h8657a6f0;
    ram_cell[   38605] = 32'hc584722b;
    ram_cell[   38606] = 32'h051605a4;
    ram_cell[   38607] = 32'h50ff188b;
    ram_cell[   38608] = 32'hccd0f783;
    ram_cell[   38609] = 32'h07aa4d96;
    ram_cell[   38610] = 32'h5042827c;
    ram_cell[   38611] = 32'h8b349e9e;
    ram_cell[   38612] = 32'h3f6607f2;
    ram_cell[   38613] = 32'h6f6b62f4;
    ram_cell[   38614] = 32'hf05f6052;
    ram_cell[   38615] = 32'h3d303599;
    ram_cell[   38616] = 32'h64b19f1e;
    ram_cell[   38617] = 32'hcce79a54;
    ram_cell[   38618] = 32'h31730c65;
    ram_cell[   38619] = 32'hcc442d5f;
    ram_cell[   38620] = 32'h0af7c264;
    ram_cell[   38621] = 32'hd90e32c4;
    ram_cell[   38622] = 32'hfd89fd80;
    ram_cell[   38623] = 32'hec416b14;
    ram_cell[   38624] = 32'hc1cc1089;
    ram_cell[   38625] = 32'h8c1f79a1;
    ram_cell[   38626] = 32'h0f3e7a84;
    ram_cell[   38627] = 32'hd32e78a9;
    ram_cell[   38628] = 32'h60ae514e;
    ram_cell[   38629] = 32'h36c55a7a;
    ram_cell[   38630] = 32'h4ae94efa;
    ram_cell[   38631] = 32'hfbb14a08;
    ram_cell[   38632] = 32'h896ac170;
    ram_cell[   38633] = 32'h69369480;
    ram_cell[   38634] = 32'h841c0bf4;
    ram_cell[   38635] = 32'h5a3787e6;
    ram_cell[   38636] = 32'h5a731d84;
    ram_cell[   38637] = 32'h68c02f7d;
    ram_cell[   38638] = 32'hfbef210d;
    ram_cell[   38639] = 32'h88588730;
    ram_cell[   38640] = 32'h103f401d;
    ram_cell[   38641] = 32'h20659e89;
    ram_cell[   38642] = 32'h14999db6;
    ram_cell[   38643] = 32'hfb1a81ac;
    ram_cell[   38644] = 32'heba5b7e5;
    ram_cell[   38645] = 32'h7c24c1e3;
    ram_cell[   38646] = 32'h0491c524;
    ram_cell[   38647] = 32'hbbbe6745;
    ram_cell[   38648] = 32'h11f338a7;
    ram_cell[   38649] = 32'hec64b5fd;
    ram_cell[   38650] = 32'h392036dc;
    ram_cell[   38651] = 32'hd5d318a4;
    ram_cell[   38652] = 32'h95eefb8a;
    ram_cell[   38653] = 32'h27d56540;
    ram_cell[   38654] = 32'hf4424bf9;
    ram_cell[   38655] = 32'hcadf3472;
    ram_cell[   38656] = 32'h80cedf30;
    ram_cell[   38657] = 32'h878da20c;
    ram_cell[   38658] = 32'h9ce85219;
    ram_cell[   38659] = 32'h55bd6dca;
    ram_cell[   38660] = 32'hbdbc2ce5;
    ram_cell[   38661] = 32'h4bb2412e;
    ram_cell[   38662] = 32'h97916df1;
    ram_cell[   38663] = 32'hdeec941e;
    ram_cell[   38664] = 32'h998f4518;
    ram_cell[   38665] = 32'heec7521f;
    ram_cell[   38666] = 32'h2c587795;
    ram_cell[   38667] = 32'h8c64c78b;
    ram_cell[   38668] = 32'h1af6c94c;
    ram_cell[   38669] = 32'h6fdb05fc;
    ram_cell[   38670] = 32'h3d4e8292;
    ram_cell[   38671] = 32'hc03310e0;
    ram_cell[   38672] = 32'h1fad4aa7;
    ram_cell[   38673] = 32'h0f65dad4;
    ram_cell[   38674] = 32'hec06e169;
    ram_cell[   38675] = 32'hd367de3b;
    ram_cell[   38676] = 32'h8752e8e3;
    ram_cell[   38677] = 32'hae0e26e4;
    ram_cell[   38678] = 32'h9faf105a;
    ram_cell[   38679] = 32'hb8a1baf0;
    ram_cell[   38680] = 32'hca98de9a;
    ram_cell[   38681] = 32'hd7c13944;
    ram_cell[   38682] = 32'h6f859037;
    ram_cell[   38683] = 32'h82410b08;
    ram_cell[   38684] = 32'he283cc3c;
    ram_cell[   38685] = 32'hf0173c2c;
    ram_cell[   38686] = 32'h890ca40c;
    ram_cell[   38687] = 32'h9bbf4dc4;
    ram_cell[   38688] = 32'h178c00d0;
    ram_cell[   38689] = 32'hb0316e3f;
    ram_cell[   38690] = 32'hf0564c03;
    ram_cell[   38691] = 32'hdab14f86;
    ram_cell[   38692] = 32'he88c81fb;
    ram_cell[   38693] = 32'hcc036baa;
    ram_cell[   38694] = 32'h45e7ee3d;
    ram_cell[   38695] = 32'hc94b6c3d;
    ram_cell[   38696] = 32'h099ab51e;
    ram_cell[   38697] = 32'h6e2a1c84;
    ram_cell[   38698] = 32'hf3901237;
    ram_cell[   38699] = 32'h9f55772c;
    ram_cell[   38700] = 32'h168db85f;
    ram_cell[   38701] = 32'hcf20dcf8;
    ram_cell[   38702] = 32'h80306ad5;
    ram_cell[   38703] = 32'h0b27aea9;
    ram_cell[   38704] = 32'h68def7d6;
    ram_cell[   38705] = 32'h3ed73d75;
    ram_cell[   38706] = 32'h12df8bc7;
    ram_cell[   38707] = 32'hce7292fb;
    ram_cell[   38708] = 32'h0e3d7cd8;
    ram_cell[   38709] = 32'he0ed6666;
    ram_cell[   38710] = 32'h60e22eb3;
    ram_cell[   38711] = 32'hc2945087;
    ram_cell[   38712] = 32'h8624d220;
    ram_cell[   38713] = 32'h5d39f06b;
    ram_cell[   38714] = 32'h74889965;
    ram_cell[   38715] = 32'h334fd0a1;
    ram_cell[   38716] = 32'h433e0d62;
    ram_cell[   38717] = 32'h68589f9c;
    ram_cell[   38718] = 32'h6931625d;
    ram_cell[   38719] = 32'h72740236;
    ram_cell[   38720] = 32'h1c52cba6;
    ram_cell[   38721] = 32'h8583591d;
    ram_cell[   38722] = 32'hcb16823f;
    ram_cell[   38723] = 32'h00d11968;
    ram_cell[   38724] = 32'hedb023f3;
    ram_cell[   38725] = 32'h71c67cd8;
    ram_cell[   38726] = 32'hd88decef;
    ram_cell[   38727] = 32'hcdcb033c;
    ram_cell[   38728] = 32'h682e6b22;
    ram_cell[   38729] = 32'h9df33c67;
    ram_cell[   38730] = 32'hc2f6eca2;
    ram_cell[   38731] = 32'h404b4863;
    ram_cell[   38732] = 32'h70b73f1d;
    ram_cell[   38733] = 32'h85b51714;
    ram_cell[   38734] = 32'hcee2c8e9;
    ram_cell[   38735] = 32'h4fa931ee;
    ram_cell[   38736] = 32'had4210f4;
    ram_cell[   38737] = 32'hd6269f7a;
    ram_cell[   38738] = 32'ha60b825b;
    ram_cell[   38739] = 32'hc9cb5b85;
    ram_cell[   38740] = 32'h67d3c598;
    ram_cell[   38741] = 32'h41bf4028;
    ram_cell[   38742] = 32'hf1f95095;
    ram_cell[   38743] = 32'hca0d877a;
    ram_cell[   38744] = 32'h24d23921;
    ram_cell[   38745] = 32'hb1d269be;
    ram_cell[   38746] = 32'h698f52bf;
    ram_cell[   38747] = 32'h21d0b668;
    ram_cell[   38748] = 32'h6c18edbf;
    ram_cell[   38749] = 32'h902edafb;
    ram_cell[   38750] = 32'hf6dfb9b2;
    ram_cell[   38751] = 32'h772d8e36;
    ram_cell[   38752] = 32'h7f2b8c22;
    ram_cell[   38753] = 32'hb2d0a4ce;
    ram_cell[   38754] = 32'h2abfea1e;
    ram_cell[   38755] = 32'h62946905;
    ram_cell[   38756] = 32'hc47f0673;
    ram_cell[   38757] = 32'h64c6131a;
    ram_cell[   38758] = 32'ha89e1f56;
    ram_cell[   38759] = 32'h1be3f28e;
    ram_cell[   38760] = 32'ha69e3ce3;
    ram_cell[   38761] = 32'hd6d5d7e6;
    ram_cell[   38762] = 32'h45fe09d4;
    ram_cell[   38763] = 32'h90037ad5;
    ram_cell[   38764] = 32'h58b8e88c;
    ram_cell[   38765] = 32'h75905f7f;
    ram_cell[   38766] = 32'h98cfd767;
    ram_cell[   38767] = 32'h72c406ed;
    ram_cell[   38768] = 32'h0a800c34;
    ram_cell[   38769] = 32'h54649504;
    ram_cell[   38770] = 32'ha79b5db9;
    ram_cell[   38771] = 32'h2a2951b2;
    ram_cell[   38772] = 32'hdaf2fff9;
    ram_cell[   38773] = 32'h4003f91a;
    ram_cell[   38774] = 32'h919494bf;
    ram_cell[   38775] = 32'h1afaa0b4;
    ram_cell[   38776] = 32'h02f1c6c8;
    ram_cell[   38777] = 32'h269f5a20;
    ram_cell[   38778] = 32'h638a95a1;
    ram_cell[   38779] = 32'h262116b2;
    ram_cell[   38780] = 32'h486a3222;
    ram_cell[   38781] = 32'h91185380;
    ram_cell[   38782] = 32'h1c2aef37;
    ram_cell[   38783] = 32'h81c8c8f1;
    ram_cell[   38784] = 32'h1aa50e49;
    ram_cell[   38785] = 32'h34bc9ad1;
    ram_cell[   38786] = 32'h55c249d1;
    ram_cell[   38787] = 32'h558869f8;
    ram_cell[   38788] = 32'he177146b;
    ram_cell[   38789] = 32'hd7f79fa5;
    ram_cell[   38790] = 32'h09fb0d7c;
    ram_cell[   38791] = 32'h1a35f016;
    ram_cell[   38792] = 32'h1c2c2264;
    ram_cell[   38793] = 32'h6fcc7d12;
    ram_cell[   38794] = 32'h423327d2;
    ram_cell[   38795] = 32'h991e422f;
    ram_cell[   38796] = 32'hc8a0152b;
    ram_cell[   38797] = 32'h3fcd01bc;
    ram_cell[   38798] = 32'h388dcd30;
    ram_cell[   38799] = 32'h96dc9a39;
    ram_cell[   38800] = 32'he7ed36dd;
    ram_cell[   38801] = 32'hdf5410c4;
    ram_cell[   38802] = 32'h701f222a;
    ram_cell[   38803] = 32'h4c2c5508;
    ram_cell[   38804] = 32'h74baa5b8;
    ram_cell[   38805] = 32'haca462cb;
    ram_cell[   38806] = 32'h2af51c4d;
    ram_cell[   38807] = 32'h5ae5cb91;
    ram_cell[   38808] = 32'h3c4bf4b3;
    ram_cell[   38809] = 32'h5c1cc97f;
    ram_cell[   38810] = 32'he51f5ada;
    ram_cell[   38811] = 32'h375f7720;
    ram_cell[   38812] = 32'h20242269;
    ram_cell[   38813] = 32'h88343dd9;
    ram_cell[   38814] = 32'h8dfe91f1;
    ram_cell[   38815] = 32'h7a95cbe5;
    ram_cell[   38816] = 32'hac50a83f;
    ram_cell[   38817] = 32'hda0bd81d;
    ram_cell[   38818] = 32'h1f981508;
    ram_cell[   38819] = 32'hbf60f0f0;
    ram_cell[   38820] = 32'had6b373b;
    ram_cell[   38821] = 32'h6807fe43;
    ram_cell[   38822] = 32'h6ff89d11;
    ram_cell[   38823] = 32'h944d7b77;
    ram_cell[   38824] = 32'hfb7f0bde;
    ram_cell[   38825] = 32'hc27f305c;
    ram_cell[   38826] = 32'h81ccfb70;
    ram_cell[   38827] = 32'hdedba746;
    ram_cell[   38828] = 32'h4bb25549;
    ram_cell[   38829] = 32'h4105e332;
    ram_cell[   38830] = 32'heb119df5;
    ram_cell[   38831] = 32'h555d35a8;
    ram_cell[   38832] = 32'hce8f8fc4;
    ram_cell[   38833] = 32'h8cf73c1b;
    ram_cell[   38834] = 32'heced772e;
    ram_cell[   38835] = 32'h7816f2fd;
    ram_cell[   38836] = 32'h783d1d06;
    ram_cell[   38837] = 32'hb7eb2ef3;
    ram_cell[   38838] = 32'h0ce6653e;
    ram_cell[   38839] = 32'h26f0f615;
    ram_cell[   38840] = 32'h6a577010;
    ram_cell[   38841] = 32'h7dbb6f8f;
    ram_cell[   38842] = 32'h63db6508;
    ram_cell[   38843] = 32'hb707086d;
    ram_cell[   38844] = 32'h6d5c94a2;
    ram_cell[   38845] = 32'he0053532;
    ram_cell[   38846] = 32'h30f43aa3;
    ram_cell[   38847] = 32'h518415dc;
    ram_cell[   38848] = 32'h071d1766;
    ram_cell[   38849] = 32'h26a2c91c;
    ram_cell[   38850] = 32'h08633379;
    ram_cell[   38851] = 32'hafc4991e;
    ram_cell[   38852] = 32'h4eaad0e0;
    ram_cell[   38853] = 32'h85bef2aa;
    ram_cell[   38854] = 32'h5d77cdc5;
    ram_cell[   38855] = 32'h1f4a725b;
    ram_cell[   38856] = 32'h9cadc504;
    ram_cell[   38857] = 32'hd82e4db9;
    ram_cell[   38858] = 32'h0c688256;
    ram_cell[   38859] = 32'h38186c70;
    ram_cell[   38860] = 32'h49360671;
    ram_cell[   38861] = 32'hcec5d758;
    ram_cell[   38862] = 32'ha57de6cd;
    ram_cell[   38863] = 32'h3aaa7801;
    ram_cell[   38864] = 32'hf2c933af;
    ram_cell[   38865] = 32'h1f3c146f;
    ram_cell[   38866] = 32'hc716e83c;
    ram_cell[   38867] = 32'h27e9dacb;
    ram_cell[   38868] = 32'h54a5e6b3;
    ram_cell[   38869] = 32'hbf43215e;
    ram_cell[   38870] = 32'h388d25d0;
    ram_cell[   38871] = 32'hc72750ae;
    ram_cell[   38872] = 32'h066f7a31;
    ram_cell[   38873] = 32'h40cd3a3d;
    ram_cell[   38874] = 32'h3fc28553;
    ram_cell[   38875] = 32'h27926f5e;
    ram_cell[   38876] = 32'h829ce256;
    ram_cell[   38877] = 32'h3e2b6bb1;
    ram_cell[   38878] = 32'he9337d64;
    ram_cell[   38879] = 32'hf7c92b26;
    ram_cell[   38880] = 32'ha05276e9;
    ram_cell[   38881] = 32'hfcef43f1;
    ram_cell[   38882] = 32'h4f4833d6;
    ram_cell[   38883] = 32'heb0f9208;
    ram_cell[   38884] = 32'hf09c26fa;
    ram_cell[   38885] = 32'hd8480a57;
    ram_cell[   38886] = 32'h781434cd;
    ram_cell[   38887] = 32'he0bb5b12;
    ram_cell[   38888] = 32'h1f84c289;
    ram_cell[   38889] = 32'h81627f99;
    ram_cell[   38890] = 32'h6f97b25e;
    ram_cell[   38891] = 32'h075404b6;
    ram_cell[   38892] = 32'h6f69d9d9;
    ram_cell[   38893] = 32'h71737a2b;
    ram_cell[   38894] = 32'h8e99dd80;
    ram_cell[   38895] = 32'h16054a61;
    ram_cell[   38896] = 32'h5cdc3286;
    ram_cell[   38897] = 32'hd94423c4;
    ram_cell[   38898] = 32'h450abeee;
    ram_cell[   38899] = 32'h1f19867d;
    ram_cell[   38900] = 32'hd580eecb;
    ram_cell[   38901] = 32'h921145d3;
    ram_cell[   38902] = 32'h01797829;
    ram_cell[   38903] = 32'h9f5607db;
    ram_cell[   38904] = 32'he6fc5e6f;
    ram_cell[   38905] = 32'h1ee630a9;
    ram_cell[   38906] = 32'h92abf8f9;
    ram_cell[   38907] = 32'hb074226b;
    ram_cell[   38908] = 32'h22db3d2b;
    ram_cell[   38909] = 32'hd58e05e2;
    ram_cell[   38910] = 32'he9334886;
    ram_cell[   38911] = 32'hf52ff1d9;
    ram_cell[   38912] = 32'h4d575e79;
    ram_cell[   38913] = 32'hce030454;
    ram_cell[   38914] = 32'h8be0f8e6;
    ram_cell[   38915] = 32'h25254165;
    ram_cell[   38916] = 32'h39c38213;
    ram_cell[   38917] = 32'he601b811;
    ram_cell[   38918] = 32'h47be8984;
    ram_cell[   38919] = 32'hf709949a;
    ram_cell[   38920] = 32'he08c2212;
    ram_cell[   38921] = 32'h424c9409;
    ram_cell[   38922] = 32'h48566d60;
    ram_cell[   38923] = 32'h76b336b8;
    ram_cell[   38924] = 32'h95c66caf;
    ram_cell[   38925] = 32'hcf2579d2;
    ram_cell[   38926] = 32'h3eeb1d84;
    ram_cell[   38927] = 32'hc3c5bd07;
    ram_cell[   38928] = 32'hdd43db7d;
    ram_cell[   38929] = 32'h763cbfef;
    ram_cell[   38930] = 32'hfd30748c;
    ram_cell[   38931] = 32'he8a6097b;
    ram_cell[   38932] = 32'h6b7a24ec;
    ram_cell[   38933] = 32'hcdcd8dc6;
    ram_cell[   38934] = 32'h30f726d2;
    ram_cell[   38935] = 32'h6b9d55cc;
    ram_cell[   38936] = 32'hf5a792c0;
    ram_cell[   38937] = 32'h2d14d852;
    ram_cell[   38938] = 32'h8a7b0b8a;
    ram_cell[   38939] = 32'h40fef521;
    ram_cell[   38940] = 32'h0fd10cbb;
    ram_cell[   38941] = 32'h6353e1ba;
    ram_cell[   38942] = 32'hc0835205;
    ram_cell[   38943] = 32'h36ebe340;
    ram_cell[   38944] = 32'h465c895b;
    ram_cell[   38945] = 32'hc366a3ce;
    ram_cell[   38946] = 32'h03a10e5c;
    ram_cell[   38947] = 32'hd9f2e20b;
    ram_cell[   38948] = 32'h7e7b81cd;
    ram_cell[   38949] = 32'h6d5b95ef;
    ram_cell[   38950] = 32'h941f28f4;
    ram_cell[   38951] = 32'h26ffcc17;
    ram_cell[   38952] = 32'hab4a2d64;
    ram_cell[   38953] = 32'hbc96839c;
    ram_cell[   38954] = 32'hba4cc9e0;
    ram_cell[   38955] = 32'hda32362d;
    ram_cell[   38956] = 32'hc15f1e5c;
    ram_cell[   38957] = 32'ha9542f4a;
    ram_cell[   38958] = 32'hd1f52638;
    ram_cell[   38959] = 32'h3dac2065;
    ram_cell[   38960] = 32'hd5ca3779;
    ram_cell[   38961] = 32'hdfc6ff3c;
    ram_cell[   38962] = 32'h82923f66;
    ram_cell[   38963] = 32'h01f3ed32;
    ram_cell[   38964] = 32'h04061fdf;
    ram_cell[   38965] = 32'hd0394b74;
    ram_cell[   38966] = 32'hc435cce6;
    ram_cell[   38967] = 32'hcf35f376;
    ram_cell[   38968] = 32'h0a5acb39;
    ram_cell[   38969] = 32'hdff48143;
    ram_cell[   38970] = 32'h3ed8ba38;
    ram_cell[   38971] = 32'h13948a82;
    ram_cell[   38972] = 32'h37823a58;
    ram_cell[   38973] = 32'h5ad865a9;
    ram_cell[   38974] = 32'h94b7b5fb;
    ram_cell[   38975] = 32'hf67e35da;
    ram_cell[   38976] = 32'h74828688;
    ram_cell[   38977] = 32'h096233d2;
    ram_cell[   38978] = 32'h86f97e3c;
    ram_cell[   38979] = 32'h486702fa;
    ram_cell[   38980] = 32'h0e1bede6;
    ram_cell[   38981] = 32'h69e73c1f;
    ram_cell[   38982] = 32'h985fce00;
    ram_cell[   38983] = 32'h80fcfca4;
    ram_cell[   38984] = 32'h6d55fbaa;
    ram_cell[   38985] = 32'h9badc362;
    ram_cell[   38986] = 32'h4022278a;
    ram_cell[   38987] = 32'h7067ac40;
    ram_cell[   38988] = 32'h30a922c5;
    ram_cell[   38989] = 32'haaeae58a;
    ram_cell[   38990] = 32'h5b3a7f7f;
    ram_cell[   38991] = 32'h202c126a;
    ram_cell[   38992] = 32'he864425b;
    ram_cell[   38993] = 32'h8cdb5a55;
    ram_cell[   38994] = 32'had6ca364;
    ram_cell[   38995] = 32'h2b890161;
    ram_cell[   38996] = 32'hb4a2f6f5;
    ram_cell[   38997] = 32'h1f124adc;
    ram_cell[   38998] = 32'h0d6a2e11;
    ram_cell[   38999] = 32'hfbe9a223;
    ram_cell[   39000] = 32'he9480631;
    ram_cell[   39001] = 32'h1bd03d06;
    ram_cell[   39002] = 32'hfa2537c3;
    ram_cell[   39003] = 32'hbb443160;
    ram_cell[   39004] = 32'he9951e40;
    ram_cell[   39005] = 32'h4c0312d9;
    ram_cell[   39006] = 32'hb6a8fa74;
    ram_cell[   39007] = 32'hbb9e4580;
    ram_cell[   39008] = 32'h3dbee3fa;
    ram_cell[   39009] = 32'h8a0d7f43;
    ram_cell[   39010] = 32'hd6bcded0;
    ram_cell[   39011] = 32'hb9193e20;
    ram_cell[   39012] = 32'h593608d8;
    ram_cell[   39013] = 32'h4aa83929;
    ram_cell[   39014] = 32'hf178bbf3;
    ram_cell[   39015] = 32'h42bd46b2;
    ram_cell[   39016] = 32'ha616c5d3;
    ram_cell[   39017] = 32'hd389b4a1;
    ram_cell[   39018] = 32'h8a3ea6c4;
    ram_cell[   39019] = 32'h0b76c0ef;
    ram_cell[   39020] = 32'h5a3756b9;
    ram_cell[   39021] = 32'h3332227e;
    ram_cell[   39022] = 32'h1a312006;
    ram_cell[   39023] = 32'h58e06686;
    ram_cell[   39024] = 32'hdbd3e193;
    ram_cell[   39025] = 32'h48e2a293;
    ram_cell[   39026] = 32'h98e5dc93;
    ram_cell[   39027] = 32'h59901749;
    ram_cell[   39028] = 32'h73169500;
    ram_cell[   39029] = 32'h3d96013f;
    ram_cell[   39030] = 32'h7b36196a;
    ram_cell[   39031] = 32'h1c69d116;
    ram_cell[   39032] = 32'h0c1bdd1a;
    ram_cell[   39033] = 32'h899c2aa2;
    ram_cell[   39034] = 32'h1fb0025e;
    ram_cell[   39035] = 32'hbdcdf343;
    ram_cell[   39036] = 32'h819e93bb;
    ram_cell[   39037] = 32'hed4446c5;
    ram_cell[   39038] = 32'h9a79a9d3;
    ram_cell[   39039] = 32'ha9c76d90;
    ram_cell[   39040] = 32'h86ddc042;
    ram_cell[   39041] = 32'h069e8e5a;
    ram_cell[   39042] = 32'h000b6c67;
    ram_cell[   39043] = 32'h4a2b3275;
    ram_cell[   39044] = 32'hf5e2181a;
    ram_cell[   39045] = 32'h26a56edc;
    ram_cell[   39046] = 32'h734bd9c6;
    ram_cell[   39047] = 32'hb375e4cb;
    ram_cell[   39048] = 32'hce753b96;
    ram_cell[   39049] = 32'he5cb1305;
    ram_cell[   39050] = 32'h96563df9;
    ram_cell[   39051] = 32'h97d92ae4;
    ram_cell[   39052] = 32'h1acaa899;
    ram_cell[   39053] = 32'h62962b0a;
    ram_cell[   39054] = 32'hc3bfd932;
    ram_cell[   39055] = 32'hec0b4c2d;
    ram_cell[   39056] = 32'h2fcf5190;
    ram_cell[   39057] = 32'ha8fb790b;
    ram_cell[   39058] = 32'h35d593cf;
    ram_cell[   39059] = 32'h94deb4cf;
    ram_cell[   39060] = 32'hbe59b0a9;
    ram_cell[   39061] = 32'hb7ef26b8;
    ram_cell[   39062] = 32'h5315154d;
    ram_cell[   39063] = 32'hca107517;
    ram_cell[   39064] = 32'hb87dcb76;
    ram_cell[   39065] = 32'h0df4f4de;
    ram_cell[   39066] = 32'hd926f12a;
    ram_cell[   39067] = 32'heec4bb89;
    ram_cell[   39068] = 32'h84d60186;
    ram_cell[   39069] = 32'hb3bce76e;
    ram_cell[   39070] = 32'hbd914164;
    ram_cell[   39071] = 32'h14ed09e5;
    ram_cell[   39072] = 32'h2ff20dee;
    ram_cell[   39073] = 32'h142d0350;
    ram_cell[   39074] = 32'hadcf55c2;
    ram_cell[   39075] = 32'hd42069c1;
    ram_cell[   39076] = 32'h60cf8427;
    ram_cell[   39077] = 32'hc8f9f504;
    ram_cell[   39078] = 32'hf9202433;
    ram_cell[   39079] = 32'h7de4d188;
    ram_cell[   39080] = 32'h1fe584ea;
    ram_cell[   39081] = 32'hefb050b9;
    ram_cell[   39082] = 32'hc9ff686d;
    ram_cell[   39083] = 32'h8ddc6702;
    ram_cell[   39084] = 32'hf4fb8ca2;
    ram_cell[   39085] = 32'ha7940958;
    ram_cell[   39086] = 32'hd7505461;
    ram_cell[   39087] = 32'h1d0b8759;
    ram_cell[   39088] = 32'h7d0b3648;
    ram_cell[   39089] = 32'h685193cb;
    ram_cell[   39090] = 32'hc496a2ad;
    ram_cell[   39091] = 32'h7ff6d1b7;
    ram_cell[   39092] = 32'h556df71b;
    ram_cell[   39093] = 32'hbebfba49;
    ram_cell[   39094] = 32'h250e1145;
    ram_cell[   39095] = 32'h9a6bc748;
    ram_cell[   39096] = 32'h79aaa84d;
    ram_cell[   39097] = 32'h34c6ed4c;
    ram_cell[   39098] = 32'h45180eb0;
    ram_cell[   39099] = 32'h354db98b;
    ram_cell[   39100] = 32'hba6f4da8;
    ram_cell[   39101] = 32'h3ea2f97e;
    ram_cell[   39102] = 32'hcc53b85b;
    ram_cell[   39103] = 32'h1bdf16bf;
    ram_cell[   39104] = 32'h24ae9d12;
    ram_cell[   39105] = 32'hcff4db0a;
    ram_cell[   39106] = 32'hae7cdc6a;
    ram_cell[   39107] = 32'h6430a402;
    ram_cell[   39108] = 32'h6d951db2;
    ram_cell[   39109] = 32'h47d2c80f;
    ram_cell[   39110] = 32'h60968240;
    ram_cell[   39111] = 32'hdbca2035;
    ram_cell[   39112] = 32'hf8363073;
    ram_cell[   39113] = 32'h6f3cf295;
    ram_cell[   39114] = 32'hcec222da;
    ram_cell[   39115] = 32'h147a8fac;
    ram_cell[   39116] = 32'h0ab12e81;
    ram_cell[   39117] = 32'ha3715e54;
    ram_cell[   39118] = 32'h578f289f;
    ram_cell[   39119] = 32'h39e8bbc9;
    ram_cell[   39120] = 32'h24cd50ea;
    ram_cell[   39121] = 32'hcdf84be6;
    ram_cell[   39122] = 32'h6b7e949f;
    ram_cell[   39123] = 32'hf8163476;
    ram_cell[   39124] = 32'hff3a18e7;
    ram_cell[   39125] = 32'hbc4650e9;
    ram_cell[   39126] = 32'h85ce3833;
    ram_cell[   39127] = 32'h997b3c19;
    ram_cell[   39128] = 32'h1953102d;
    ram_cell[   39129] = 32'hfb5defd4;
    ram_cell[   39130] = 32'hf697dc6f;
    ram_cell[   39131] = 32'h53317293;
    ram_cell[   39132] = 32'h69b3e8a8;
    ram_cell[   39133] = 32'h440c6da4;
    ram_cell[   39134] = 32'h348490a5;
    ram_cell[   39135] = 32'hdbb67cc4;
    ram_cell[   39136] = 32'hb8942f1a;
    ram_cell[   39137] = 32'h0656bc7f;
    ram_cell[   39138] = 32'h1505bc72;
    ram_cell[   39139] = 32'h87c0f482;
    ram_cell[   39140] = 32'h07238347;
    ram_cell[   39141] = 32'h6e4a8926;
    ram_cell[   39142] = 32'h3d5383f5;
    ram_cell[   39143] = 32'h7a1ff9e1;
    ram_cell[   39144] = 32'hd65eff69;
    ram_cell[   39145] = 32'h1336b76d;
    ram_cell[   39146] = 32'h22315072;
    ram_cell[   39147] = 32'h43d55429;
    ram_cell[   39148] = 32'h027b286f;
    ram_cell[   39149] = 32'hf41712b4;
    ram_cell[   39150] = 32'hb0a7caf8;
    ram_cell[   39151] = 32'h02d8fedb;
    ram_cell[   39152] = 32'h056dfdc0;
    ram_cell[   39153] = 32'h64b8ff03;
    ram_cell[   39154] = 32'h9489e837;
    ram_cell[   39155] = 32'h00e25375;
    ram_cell[   39156] = 32'h4c6f968f;
    ram_cell[   39157] = 32'hb53728aa;
    ram_cell[   39158] = 32'h26970d58;
    ram_cell[   39159] = 32'hdf27dfed;
    ram_cell[   39160] = 32'h007f904c;
    ram_cell[   39161] = 32'h2d7669d0;
    ram_cell[   39162] = 32'hbb07c79f;
    ram_cell[   39163] = 32'h477d4351;
    ram_cell[   39164] = 32'h4d3bd627;
    ram_cell[   39165] = 32'h992d0930;
    ram_cell[   39166] = 32'h23260b40;
    ram_cell[   39167] = 32'hae144b2b;
    ram_cell[   39168] = 32'h940c35c0;
    ram_cell[   39169] = 32'h4a57fccb;
    ram_cell[   39170] = 32'h9ed49bb5;
    ram_cell[   39171] = 32'h86d69eac;
    ram_cell[   39172] = 32'hd19e9c0e;
    ram_cell[   39173] = 32'hfd4e07a0;
    ram_cell[   39174] = 32'he57c4cfb;
    ram_cell[   39175] = 32'h3718557a;
    ram_cell[   39176] = 32'hd3b81e3c;
    ram_cell[   39177] = 32'hf49a2712;
    ram_cell[   39178] = 32'hffff781c;
    ram_cell[   39179] = 32'h6a77cd17;
    ram_cell[   39180] = 32'h0ff867e3;
    ram_cell[   39181] = 32'h18f7221c;
    ram_cell[   39182] = 32'h1a3207e6;
    ram_cell[   39183] = 32'hdeb66c88;
    ram_cell[   39184] = 32'h0c548118;
    ram_cell[   39185] = 32'h272c5da4;
    ram_cell[   39186] = 32'h98b9e22f;
    ram_cell[   39187] = 32'h4db5285d;
    ram_cell[   39188] = 32'h7c37930b;
    ram_cell[   39189] = 32'h9db2f637;
    ram_cell[   39190] = 32'hbb5686bd;
    ram_cell[   39191] = 32'h037b3e3c;
    ram_cell[   39192] = 32'h80780038;
    ram_cell[   39193] = 32'ha3081007;
    ram_cell[   39194] = 32'h58e0bddd;
    ram_cell[   39195] = 32'h5cd9be98;
    ram_cell[   39196] = 32'h5470048b;
    ram_cell[   39197] = 32'h37d91b03;
    ram_cell[   39198] = 32'h6f37693a;
    ram_cell[   39199] = 32'hef828126;
    ram_cell[   39200] = 32'h558eacd9;
    ram_cell[   39201] = 32'h445eb27f;
    ram_cell[   39202] = 32'hf81adb66;
    ram_cell[   39203] = 32'hfb17fc6b;
    ram_cell[   39204] = 32'hc594a91b;
    ram_cell[   39205] = 32'h922ed758;
    ram_cell[   39206] = 32'hbc5b74d6;
    ram_cell[   39207] = 32'h9ff21c0b;
    ram_cell[   39208] = 32'hb20efdd2;
    ram_cell[   39209] = 32'h9b49af71;
    ram_cell[   39210] = 32'h3d8b3701;
    ram_cell[   39211] = 32'h69ef40bf;
    ram_cell[   39212] = 32'hf83b67d7;
    ram_cell[   39213] = 32'h287fe16f;
    ram_cell[   39214] = 32'hfeb58f4a;
    ram_cell[   39215] = 32'hf89f868c;
    ram_cell[   39216] = 32'h7673ad19;
    ram_cell[   39217] = 32'hcadec70c;
    ram_cell[   39218] = 32'h8ac44b42;
    ram_cell[   39219] = 32'hbd53307c;
    ram_cell[   39220] = 32'h27c629f9;
    ram_cell[   39221] = 32'hb3fd0b2f;
    ram_cell[   39222] = 32'h1a852f2f;
    ram_cell[   39223] = 32'h8e2e2f83;
    ram_cell[   39224] = 32'he18b967d;
    ram_cell[   39225] = 32'h9a847978;
    ram_cell[   39226] = 32'h7602cb72;
    ram_cell[   39227] = 32'h0f53fb28;
    ram_cell[   39228] = 32'h9e72f29e;
    ram_cell[   39229] = 32'hb10ebc4e;
    ram_cell[   39230] = 32'h8bfb9b81;
    ram_cell[   39231] = 32'hf81b9602;
    ram_cell[   39232] = 32'h61189a4f;
    ram_cell[   39233] = 32'hdba8114c;
    ram_cell[   39234] = 32'h7b833ae7;
    ram_cell[   39235] = 32'hc9fad50e;
    ram_cell[   39236] = 32'hcd950528;
    ram_cell[   39237] = 32'h8479683d;
    ram_cell[   39238] = 32'h07eb59dd;
    ram_cell[   39239] = 32'h1d1f035e;
    ram_cell[   39240] = 32'hddf41968;
    ram_cell[   39241] = 32'hdf346133;
    ram_cell[   39242] = 32'hbb60f094;
    ram_cell[   39243] = 32'hdc80fe82;
    ram_cell[   39244] = 32'h234fa26d;
    ram_cell[   39245] = 32'h70bc1e37;
    ram_cell[   39246] = 32'hfe623b2c;
    ram_cell[   39247] = 32'h46ddd65e;
    ram_cell[   39248] = 32'haae88ec8;
    ram_cell[   39249] = 32'h3d04b697;
    ram_cell[   39250] = 32'h7b9fe342;
    ram_cell[   39251] = 32'h023d5b3c;
    ram_cell[   39252] = 32'hd69467b6;
    ram_cell[   39253] = 32'ha99b40eb;
    ram_cell[   39254] = 32'h60858103;
    ram_cell[   39255] = 32'hc7e55ff6;
    ram_cell[   39256] = 32'h0e27fc9c;
    ram_cell[   39257] = 32'h1b65a320;
    ram_cell[   39258] = 32'h0ce27f07;
    ram_cell[   39259] = 32'hb4c0c8aa;
    ram_cell[   39260] = 32'h2947cb40;
    ram_cell[   39261] = 32'h848cd230;
    ram_cell[   39262] = 32'h015e3bc6;
    ram_cell[   39263] = 32'h62b7f276;
    ram_cell[   39264] = 32'h247f0d00;
    ram_cell[   39265] = 32'h51c2e97b;
    ram_cell[   39266] = 32'h46d15a53;
    ram_cell[   39267] = 32'h5cf6dc0c;
    ram_cell[   39268] = 32'hd42221b2;
    ram_cell[   39269] = 32'h8eab1b1e;
    ram_cell[   39270] = 32'h819c71c2;
    ram_cell[   39271] = 32'h0b220dc1;
    ram_cell[   39272] = 32'h129dc113;
    ram_cell[   39273] = 32'he2bd2612;
    ram_cell[   39274] = 32'hecf55af7;
    ram_cell[   39275] = 32'h4dc65aff;
    ram_cell[   39276] = 32'h2f857069;
    ram_cell[   39277] = 32'h2aea41c9;
    ram_cell[   39278] = 32'hd118268c;
    ram_cell[   39279] = 32'hcb6dda2c;
    ram_cell[   39280] = 32'h05d21613;
    ram_cell[   39281] = 32'h6c9edeb2;
    ram_cell[   39282] = 32'h29c7138c;
    ram_cell[   39283] = 32'h6f44a7be;
    ram_cell[   39284] = 32'h95cc09cd;
    ram_cell[   39285] = 32'haf76edfa;
    ram_cell[   39286] = 32'h15fc5723;
    ram_cell[   39287] = 32'h86ff5b29;
    ram_cell[   39288] = 32'h48ade4c1;
    ram_cell[   39289] = 32'h205b40e8;
    ram_cell[   39290] = 32'h89efd63c;
    ram_cell[   39291] = 32'hffeabd7f;
    ram_cell[   39292] = 32'h6643317c;
    ram_cell[   39293] = 32'he9155aa4;
    ram_cell[   39294] = 32'h3dc22be9;
    ram_cell[   39295] = 32'h8bdd5a16;
    ram_cell[   39296] = 32'hce324232;
    ram_cell[   39297] = 32'h93824cb1;
    ram_cell[   39298] = 32'h04e3c5af;
    ram_cell[   39299] = 32'hf1cf666e;
    ram_cell[   39300] = 32'h71cf1170;
    ram_cell[   39301] = 32'hda316112;
    ram_cell[   39302] = 32'h7cabe28a;
    ram_cell[   39303] = 32'h2e06648c;
    ram_cell[   39304] = 32'h7bf9d48e;
    ram_cell[   39305] = 32'hc6214200;
    ram_cell[   39306] = 32'h31dfc0b1;
    ram_cell[   39307] = 32'h7f40a321;
    ram_cell[   39308] = 32'h7c9a6a0a;
    ram_cell[   39309] = 32'hddefb903;
    ram_cell[   39310] = 32'h3bf93912;
    ram_cell[   39311] = 32'ha8672511;
    ram_cell[   39312] = 32'h3e4130ad;
    ram_cell[   39313] = 32'h4b5d44b1;
    ram_cell[   39314] = 32'h167af2d2;
    ram_cell[   39315] = 32'hdb4645d1;
    ram_cell[   39316] = 32'h47eb0192;
    ram_cell[   39317] = 32'hcf1c82fb;
    ram_cell[   39318] = 32'h05265eb3;
    ram_cell[   39319] = 32'h724e5a60;
    ram_cell[   39320] = 32'h022406b0;
    ram_cell[   39321] = 32'h483189a3;
    ram_cell[   39322] = 32'h7cf71455;
    ram_cell[   39323] = 32'h213ec8d1;
    ram_cell[   39324] = 32'h41ea90ec;
    ram_cell[   39325] = 32'h16cbd26d;
    ram_cell[   39326] = 32'h344a7d1d;
    ram_cell[   39327] = 32'h672dd45f;
    ram_cell[   39328] = 32'heaf23ce7;
    ram_cell[   39329] = 32'h13439ed2;
    ram_cell[   39330] = 32'h7143397c;
    ram_cell[   39331] = 32'h78f27204;
    ram_cell[   39332] = 32'h8056eedc;
    ram_cell[   39333] = 32'hc55a089c;
    ram_cell[   39334] = 32'h2aaa9dbc;
    ram_cell[   39335] = 32'h0d6581df;
    ram_cell[   39336] = 32'hc7debaab;
    ram_cell[   39337] = 32'h0e3f39ce;
    ram_cell[   39338] = 32'hca02c820;
    ram_cell[   39339] = 32'hca693681;
    ram_cell[   39340] = 32'h8f028a94;
    ram_cell[   39341] = 32'hd814024f;
    ram_cell[   39342] = 32'h5aa8ac77;
    ram_cell[   39343] = 32'h35faa159;
    ram_cell[   39344] = 32'h98284af9;
    ram_cell[   39345] = 32'hf5a36ae3;
    ram_cell[   39346] = 32'h5ee14528;
    ram_cell[   39347] = 32'heb6bbac4;
    ram_cell[   39348] = 32'h30eb7904;
    ram_cell[   39349] = 32'h9ae76b24;
    ram_cell[   39350] = 32'hca41bafa;
    ram_cell[   39351] = 32'h7c75f90b;
    ram_cell[   39352] = 32'h21ed78e9;
    ram_cell[   39353] = 32'h298e42a4;
    ram_cell[   39354] = 32'h117d5b23;
    ram_cell[   39355] = 32'h42f6d1a0;
    ram_cell[   39356] = 32'h3aafcd8b;
    ram_cell[   39357] = 32'hf78a62b1;
    ram_cell[   39358] = 32'h1cf21025;
    ram_cell[   39359] = 32'h64496d9b;
    ram_cell[   39360] = 32'h5f423e4e;
    ram_cell[   39361] = 32'hc387feb2;
    ram_cell[   39362] = 32'h54821413;
    ram_cell[   39363] = 32'h9ba81896;
    ram_cell[   39364] = 32'h717b6f26;
    ram_cell[   39365] = 32'h5490f282;
    ram_cell[   39366] = 32'h015c0f40;
    ram_cell[   39367] = 32'hfbbdce64;
    ram_cell[   39368] = 32'h787adc8f;
    ram_cell[   39369] = 32'h786eaaac;
    ram_cell[   39370] = 32'hd5fa06ce;
    ram_cell[   39371] = 32'ha6ffd7cd;
    ram_cell[   39372] = 32'h8c1df07d;
    ram_cell[   39373] = 32'h09a0fa8b;
    ram_cell[   39374] = 32'h4ac5931c;
    ram_cell[   39375] = 32'h6323f1f5;
    ram_cell[   39376] = 32'heee06d3a;
    ram_cell[   39377] = 32'haf7fb0d2;
    ram_cell[   39378] = 32'he414e989;
    ram_cell[   39379] = 32'h21881c5b;
    ram_cell[   39380] = 32'h29dd3ce3;
    ram_cell[   39381] = 32'hf500d471;
    ram_cell[   39382] = 32'h1692e63f;
    ram_cell[   39383] = 32'hc4857338;
    ram_cell[   39384] = 32'h269cfe6c;
    ram_cell[   39385] = 32'hbea8627d;
    ram_cell[   39386] = 32'hfe9bb73f;
    ram_cell[   39387] = 32'hd2a9cf4b;
    ram_cell[   39388] = 32'hd23d058a;
    ram_cell[   39389] = 32'h8191287f;
    ram_cell[   39390] = 32'h447f8cb5;
    ram_cell[   39391] = 32'h8961071a;
    ram_cell[   39392] = 32'hca2950d1;
    ram_cell[   39393] = 32'hadbf9312;
    ram_cell[   39394] = 32'h65bfd68d;
    ram_cell[   39395] = 32'ha4b836e3;
    ram_cell[   39396] = 32'h1c1637ae;
    ram_cell[   39397] = 32'h093d1ea9;
    ram_cell[   39398] = 32'he3e01cb9;
    ram_cell[   39399] = 32'hdb53d4ad;
    ram_cell[   39400] = 32'h4a871117;
    ram_cell[   39401] = 32'h29bc6878;
    ram_cell[   39402] = 32'h0c43fc3b;
    ram_cell[   39403] = 32'h24f9e588;
    ram_cell[   39404] = 32'h25daae6d;
    ram_cell[   39405] = 32'h8a3f9708;
    ram_cell[   39406] = 32'h51f1fcc7;
    ram_cell[   39407] = 32'h6075572c;
    ram_cell[   39408] = 32'h0a9c47e4;
    ram_cell[   39409] = 32'hdce77191;
    ram_cell[   39410] = 32'h4f30636b;
    ram_cell[   39411] = 32'h5f427950;
    ram_cell[   39412] = 32'he4492818;
    ram_cell[   39413] = 32'hdb089866;
    ram_cell[   39414] = 32'h8da9cbe4;
    ram_cell[   39415] = 32'hbf12adcd;
    ram_cell[   39416] = 32'h53276c03;
    ram_cell[   39417] = 32'h0b63fa83;
    ram_cell[   39418] = 32'h350bb381;
    ram_cell[   39419] = 32'h7d569538;
    ram_cell[   39420] = 32'h7044d927;
    ram_cell[   39421] = 32'he6e38461;
    ram_cell[   39422] = 32'h4e0f8ae7;
    ram_cell[   39423] = 32'h154b6266;
    ram_cell[   39424] = 32'h7846856f;
    ram_cell[   39425] = 32'he41b2df4;
    ram_cell[   39426] = 32'h42779fb4;
    ram_cell[   39427] = 32'h22c89801;
    ram_cell[   39428] = 32'hdc3f8567;
    ram_cell[   39429] = 32'h3e471900;
    ram_cell[   39430] = 32'h3aaf6608;
    ram_cell[   39431] = 32'h576992a5;
    ram_cell[   39432] = 32'h24c2cb17;
    ram_cell[   39433] = 32'hd7f47e0b;
    ram_cell[   39434] = 32'hf7953804;
    ram_cell[   39435] = 32'h0ba5c980;
    ram_cell[   39436] = 32'hbf4e4f03;
    ram_cell[   39437] = 32'h0a0be65a;
    ram_cell[   39438] = 32'ha3b63c5f;
    ram_cell[   39439] = 32'hb7450e68;
    ram_cell[   39440] = 32'h806dfc97;
    ram_cell[   39441] = 32'h1e3dcd8a;
    ram_cell[   39442] = 32'h41478a72;
    ram_cell[   39443] = 32'ha8700093;
    ram_cell[   39444] = 32'h6ad989c3;
    ram_cell[   39445] = 32'h8657b4e4;
    ram_cell[   39446] = 32'he7d4b73a;
    ram_cell[   39447] = 32'h2f62a32e;
    ram_cell[   39448] = 32'h24c45823;
    ram_cell[   39449] = 32'h396ad3c1;
    ram_cell[   39450] = 32'hd17e1dfd;
    ram_cell[   39451] = 32'h8c005b91;
    ram_cell[   39452] = 32'h0e445f63;
    ram_cell[   39453] = 32'h1a03c915;
    ram_cell[   39454] = 32'hc23304e6;
    ram_cell[   39455] = 32'h2dda3867;
    ram_cell[   39456] = 32'he171d0cd;
    ram_cell[   39457] = 32'h16f32507;
    ram_cell[   39458] = 32'he4ead2e1;
    ram_cell[   39459] = 32'h6e7ac3f7;
    ram_cell[   39460] = 32'hc4257f09;
    ram_cell[   39461] = 32'hcd228ae1;
    ram_cell[   39462] = 32'h6dfda165;
    ram_cell[   39463] = 32'hd8d523bd;
    ram_cell[   39464] = 32'h91b9dd8f;
    ram_cell[   39465] = 32'h466b7c11;
    ram_cell[   39466] = 32'h930ac06f;
    ram_cell[   39467] = 32'h79385b5e;
    ram_cell[   39468] = 32'hd1801f42;
    ram_cell[   39469] = 32'hbafed901;
    ram_cell[   39470] = 32'h9ce8387b;
    ram_cell[   39471] = 32'h762521a1;
    ram_cell[   39472] = 32'h789586b9;
    ram_cell[   39473] = 32'h61c36316;
    ram_cell[   39474] = 32'h28d054bb;
    ram_cell[   39475] = 32'he6b68b98;
    ram_cell[   39476] = 32'h3f5b3d5a;
    ram_cell[   39477] = 32'h0e002b57;
    ram_cell[   39478] = 32'h8ae9b1b0;
    ram_cell[   39479] = 32'hd8bde041;
    ram_cell[   39480] = 32'hc1d98ef8;
    ram_cell[   39481] = 32'hb50db59e;
    ram_cell[   39482] = 32'h5af71ca2;
    ram_cell[   39483] = 32'hd593c767;
    ram_cell[   39484] = 32'hc97e1f63;
    ram_cell[   39485] = 32'h08a8b878;
    ram_cell[   39486] = 32'h8afd9f8d;
    ram_cell[   39487] = 32'hc1a64aea;
    ram_cell[   39488] = 32'hf14c4f37;
    ram_cell[   39489] = 32'h4b0bf290;
    ram_cell[   39490] = 32'hc97d920b;
    ram_cell[   39491] = 32'h75a1ce62;
    ram_cell[   39492] = 32'hd1c8f6c8;
    ram_cell[   39493] = 32'he6bf652f;
    ram_cell[   39494] = 32'he4044c3c;
    ram_cell[   39495] = 32'h50cde6e7;
    ram_cell[   39496] = 32'h4e841d48;
    ram_cell[   39497] = 32'h8c4531c8;
    ram_cell[   39498] = 32'hdf4cbd04;
    ram_cell[   39499] = 32'heb22de4a;
    ram_cell[   39500] = 32'h821724c5;
    ram_cell[   39501] = 32'hcefe7919;
    ram_cell[   39502] = 32'h89924a6d;
    ram_cell[   39503] = 32'h58c61e7c;
    ram_cell[   39504] = 32'h586c2035;
    ram_cell[   39505] = 32'h0f77180e;
    ram_cell[   39506] = 32'h4c168962;
    ram_cell[   39507] = 32'he45bd032;
    ram_cell[   39508] = 32'hb4750ad8;
    ram_cell[   39509] = 32'h85a9983e;
    ram_cell[   39510] = 32'h32906c99;
    ram_cell[   39511] = 32'h51a2e03c;
    ram_cell[   39512] = 32'h21875bcd;
    ram_cell[   39513] = 32'hf0168962;
    ram_cell[   39514] = 32'haa418cb7;
    ram_cell[   39515] = 32'h0f6152a5;
    ram_cell[   39516] = 32'h3d5bdc1a;
    ram_cell[   39517] = 32'h81355e13;
    ram_cell[   39518] = 32'h4c7b68bf;
    ram_cell[   39519] = 32'h33a4244c;
    ram_cell[   39520] = 32'h15d27736;
    ram_cell[   39521] = 32'h1dec163f;
    ram_cell[   39522] = 32'h0fbc0ded;
    ram_cell[   39523] = 32'h955ffd47;
    ram_cell[   39524] = 32'h3a662422;
    ram_cell[   39525] = 32'hcbb9c2ec;
    ram_cell[   39526] = 32'h7683952b;
    ram_cell[   39527] = 32'hb12c4563;
    ram_cell[   39528] = 32'he98ea612;
    ram_cell[   39529] = 32'h870535fd;
    ram_cell[   39530] = 32'h5419a2c7;
    ram_cell[   39531] = 32'h90c613d4;
    ram_cell[   39532] = 32'h39df2c33;
    ram_cell[   39533] = 32'h07c837a0;
    ram_cell[   39534] = 32'h3ea3ea53;
    ram_cell[   39535] = 32'hd942e3dd;
    ram_cell[   39536] = 32'h67f034d4;
    ram_cell[   39537] = 32'h2510f5ea;
    ram_cell[   39538] = 32'h7961812a;
    ram_cell[   39539] = 32'hbd784b38;
    ram_cell[   39540] = 32'he0d59136;
    ram_cell[   39541] = 32'hac847dbc;
    ram_cell[   39542] = 32'hdb7292ee;
    ram_cell[   39543] = 32'h514db577;
    ram_cell[   39544] = 32'hf55f589d;
    ram_cell[   39545] = 32'hcefe89e8;
    ram_cell[   39546] = 32'h6252019f;
    ram_cell[   39547] = 32'h1f0d6ee3;
    ram_cell[   39548] = 32'h96066e28;
    ram_cell[   39549] = 32'hd9265657;
    ram_cell[   39550] = 32'he0d48fb8;
    ram_cell[   39551] = 32'hd392998c;
    ram_cell[   39552] = 32'h9473578e;
    ram_cell[   39553] = 32'hed2f0abb;
    ram_cell[   39554] = 32'h6daada84;
    ram_cell[   39555] = 32'h4f9984fd;
    ram_cell[   39556] = 32'h86a908e8;
    ram_cell[   39557] = 32'h492102e0;
    ram_cell[   39558] = 32'hafc73476;
    ram_cell[   39559] = 32'h77a9f079;
    ram_cell[   39560] = 32'h9fdb35e2;
    ram_cell[   39561] = 32'h414f9fa9;
    ram_cell[   39562] = 32'h838ba39f;
    ram_cell[   39563] = 32'h75feccba;
    ram_cell[   39564] = 32'hb5da5072;
    ram_cell[   39565] = 32'h45807193;
    ram_cell[   39566] = 32'hdd783d14;
    ram_cell[   39567] = 32'h75a2429a;
    ram_cell[   39568] = 32'h00396e83;
    ram_cell[   39569] = 32'hc1e7666f;
    ram_cell[   39570] = 32'h1147b089;
    ram_cell[   39571] = 32'hfbcac937;
    ram_cell[   39572] = 32'hf96ee945;
    ram_cell[   39573] = 32'h72dbdd10;
    ram_cell[   39574] = 32'hcd4c4e42;
    ram_cell[   39575] = 32'h84e7db06;
    ram_cell[   39576] = 32'ha298cc81;
    ram_cell[   39577] = 32'hd06c7c85;
    ram_cell[   39578] = 32'h4e91ea95;
    ram_cell[   39579] = 32'h944ecadc;
    ram_cell[   39580] = 32'hcafed161;
    ram_cell[   39581] = 32'h687379c0;
    ram_cell[   39582] = 32'hb03e647a;
    ram_cell[   39583] = 32'h81ce9b98;
    ram_cell[   39584] = 32'h127da55f;
    ram_cell[   39585] = 32'h74a3d85e;
    ram_cell[   39586] = 32'h29680402;
    ram_cell[   39587] = 32'h5ed75e6c;
    ram_cell[   39588] = 32'h380ee534;
    ram_cell[   39589] = 32'hd43ecc5b;
    ram_cell[   39590] = 32'h06f63899;
    ram_cell[   39591] = 32'ha31eacd6;
    ram_cell[   39592] = 32'h297319cb;
    ram_cell[   39593] = 32'h637d24db;
    ram_cell[   39594] = 32'hbdf444b1;
    ram_cell[   39595] = 32'h6942baba;
    ram_cell[   39596] = 32'h551c2a7f;
    ram_cell[   39597] = 32'h09dc2b19;
    ram_cell[   39598] = 32'h55bcfcbc;
    ram_cell[   39599] = 32'h250cfa1c;
    ram_cell[   39600] = 32'h23250ab9;
    ram_cell[   39601] = 32'hdd8385d6;
    ram_cell[   39602] = 32'hce368c13;
    ram_cell[   39603] = 32'hd7b1ff68;
    ram_cell[   39604] = 32'h2cf4efee;
    ram_cell[   39605] = 32'h920409c3;
    ram_cell[   39606] = 32'h7a0cc1e6;
    ram_cell[   39607] = 32'he1e48b4b;
    ram_cell[   39608] = 32'h62a2eb87;
    ram_cell[   39609] = 32'he7ee5e80;
    ram_cell[   39610] = 32'h01d418b9;
    ram_cell[   39611] = 32'h66ec10f5;
    ram_cell[   39612] = 32'h9e55e8ff;
    ram_cell[   39613] = 32'hafaf1862;
    ram_cell[   39614] = 32'hf8b3c730;
    ram_cell[   39615] = 32'h268d9afd;
    ram_cell[   39616] = 32'h2fb3a922;
    ram_cell[   39617] = 32'hb2e31b69;
    ram_cell[   39618] = 32'h6ba2547e;
    ram_cell[   39619] = 32'hd91d8911;
    ram_cell[   39620] = 32'he4bd2c88;
    ram_cell[   39621] = 32'h2b733743;
    ram_cell[   39622] = 32'hd60032e7;
    ram_cell[   39623] = 32'he38a1e66;
    ram_cell[   39624] = 32'h94428705;
    ram_cell[   39625] = 32'hf15b1ed6;
    ram_cell[   39626] = 32'he24015d7;
    ram_cell[   39627] = 32'h8b6b4f1d;
    ram_cell[   39628] = 32'hffbb6e2e;
    ram_cell[   39629] = 32'hb5b1072b;
    ram_cell[   39630] = 32'had5a1d48;
    ram_cell[   39631] = 32'h5d8a9ee8;
    ram_cell[   39632] = 32'h9cb06600;
    ram_cell[   39633] = 32'h85138ce9;
    ram_cell[   39634] = 32'he87a8452;
    ram_cell[   39635] = 32'hac3bfa38;
    ram_cell[   39636] = 32'ha58b76ee;
    ram_cell[   39637] = 32'hb9f6d1cd;
    ram_cell[   39638] = 32'hf475b78e;
    ram_cell[   39639] = 32'h426c48d4;
    ram_cell[   39640] = 32'h3abf2c11;
    ram_cell[   39641] = 32'h6c5b3f64;
    ram_cell[   39642] = 32'hd7f3dfb9;
    ram_cell[   39643] = 32'h9418ba6c;
    ram_cell[   39644] = 32'hab9f4404;
    ram_cell[   39645] = 32'h8172ec7f;
    ram_cell[   39646] = 32'h18d8cc16;
    ram_cell[   39647] = 32'h6ab1b938;
    ram_cell[   39648] = 32'hef40c3b6;
    ram_cell[   39649] = 32'h98e3c157;
    ram_cell[   39650] = 32'h57ed75d4;
    ram_cell[   39651] = 32'h2194c5dd;
    ram_cell[   39652] = 32'hfaad5a74;
    ram_cell[   39653] = 32'h75bac251;
    ram_cell[   39654] = 32'hd1b04f86;
    ram_cell[   39655] = 32'h841a9ea6;
    ram_cell[   39656] = 32'h54f98efd;
    ram_cell[   39657] = 32'h3c3920ae;
    ram_cell[   39658] = 32'hd3864d18;
    ram_cell[   39659] = 32'hca5e181f;
    ram_cell[   39660] = 32'h7c140b1a;
    ram_cell[   39661] = 32'h6fcd0051;
    ram_cell[   39662] = 32'hc3565bab;
    ram_cell[   39663] = 32'h19d8107c;
    ram_cell[   39664] = 32'h0310cf16;
    ram_cell[   39665] = 32'h99ad671d;
    ram_cell[   39666] = 32'h938b203e;
    ram_cell[   39667] = 32'h9c665a24;
    ram_cell[   39668] = 32'h681fb650;
    ram_cell[   39669] = 32'h17cc0d39;
    ram_cell[   39670] = 32'h3b3ad78a;
    ram_cell[   39671] = 32'h97e59496;
    ram_cell[   39672] = 32'hbb378296;
    ram_cell[   39673] = 32'h32212c47;
    ram_cell[   39674] = 32'h16b7fac2;
    ram_cell[   39675] = 32'h30c7a4e3;
    ram_cell[   39676] = 32'h89d44760;
    ram_cell[   39677] = 32'h8c0e2b17;
    ram_cell[   39678] = 32'hc08017e1;
    ram_cell[   39679] = 32'h849da2cd;
    ram_cell[   39680] = 32'h75a7ba21;
    ram_cell[   39681] = 32'hb9fba018;
    ram_cell[   39682] = 32'h4f836fb4;
    ram_cell[   39683] = 32'he4870d2f;
    ram_cell[   39684] = 32'ha88db356;
    ram_cell[   39685] = 32'h6aa91d3d;
    ram_cell[   39686] = 32'hf482a1b5;
    ram_cell[   39687] = 32'h005443e2;
    ram_cell[   39688] = 32'hc269a0d2;
    ram_cell[   39689] = 32'h1bb26a3a;
    ram_cell[   39690] = 32'hbfe18549;
    ram_cell[   39691] = 32'h42ce987e;
    ram_cell[   39692] = 32'h44af941c;
    ram_cell[   39693] = 32'h447ee8d7;
    ram_cell[   39694] = 32'h25e409df;
    ram_cell[   39695] = 32'h93439167;
    ram_cell[   39696] = 32'hb254c79e;
    ram_cell[   39697] = 32'hfe26225a;
    ram_cell[   39698] = 32'h67ee7b27;
    ram_cell[   39699] = 32'h7317ab81;
    ram_cell[   39700] = 32'hc6ec3856;
    ram_cell[   39701] = 32'hfe87e2fd;
    ram_cell[   39702] = 32'h573625a1;
    ram_cell[   39703] = 32'hd663422f;
    ram_cell[   39704] = 32'hd101d8f2;
    ram_cell[   39705] = 32'h4437151d;
    ram_cell[   39706] = 32'h76f81290;
    ram_cell[   39707] = 32'h4529fa3b;
    ram_cell[   39708] = 32'h3b2dc98a;
    ram_cell[   39709] = 32'h5ea335b6;
    ram_cell[   39710] = 32'he77a0106;
    ram_cell[   39711] = 32'h84c38a45;
    ram_cell[   39712] = 32'h66ab573f;
    ram_cell[   39713] = 32'h68e500e1;
    ram_cell[   39714] = 32'hedea50d6;
    ram_cell[   39715] = 32'hc079c0e6;
    ram_cell[   39716] = 32'h4305b79b;
    ram_cell[   39717] = 32'h3f1cd719;
    ram_cell[   39718] = 32'h49750b36;
    ram_cell[   39719] = 32'h34d98557;
    ram_cell[   39720] = 32'he9bb9ba4;
    ram_cell[   39721] = 32'h3c832a1f;
    ram_cell[   39722] = 32'h0b6bb405;
    ram_cell[   39723] = 32'he1274ccf;
    ram_cell[   39724] = 32'hae09112f;
    ram_cell[   39725] = 32'h2e91b20a;
    ram_cell[   39726] = 32'hc17028db;
    ram_cell[   39727] = 32'he860cdd2;
    ram_cell[   39728] = 32'h3bc10ea9;
    ram_cell[   39729] = 32'h6ec3b1f5;
    ram_cell[   39730] = 32'h3d9d17e8;
    ram_cell[   39731] = 32'ha8d110e0;
    ram_cell[   39732] = 32'hd8e0b416;
    ram_cell[   39733] = 32'h412e9f70;
    ram_cell[   39734] = 32'hd3b74e41;
    ram_cell[   39735] = 32'hf9f610ab;
    ram_cell[   39736] = 32'h6ab664a2;
    ram_cell[   39737] = 32'ha84a30c9;
    ram_cell[   39738] = 32'hb5fcdbaa;
    ram_cell[   39739] = 32'h13901362;
    ram_cell[   39740] = 32'ha9f02a6b;
    ram_cell[   39741] = 32'h33e61c00;
    ram_cell[   39742] = 32'h12b5fa02;
    ram_cell[   39743] = 32'h96e4b2ba;
    ram_cell[   39744] = 32'h613141ee;
    ram_cell[   39745] = 32'h4daf6a29;
    ram_cell[   39746] = 32'h2122083f;
    ram_cell[   39747] = 32'h0d459baa;
    ram_cell[   39748] = 32'h68e63c96;
    ram_cell[   39749] = 32'h77fc2846;
    ram_cell[   39750] = 32'h95dbdfd4;
    ram_cell[   39751] = 32'h7325af0b;
    ram_cell[   39752] = 32'h4db36118;
    ram_cell[   39753] = 32'hc461d899;
    ram_cell[   39754] = 32'hb22c1ef2;
    ram_cell[   39755] = 32'he2278815;
    ram_cell[   39756] = 32'h156e2f1b;
    ram_cell[   39757] = 32'h9bc069e8;
    ram_cell[   39758] = 32'hc58ddb17;
    ram_cell[   39759] = 32'haf3ba495;
    ram_cell[   39760] = 32'h3751f18d;
    ram_cell[   39761] = 32'h55a1ee5d;
    ram_cell[   39762] = 32'h67120042;
    ram_cell[   39763] = 32'h1ee32f17;
    ram_cell[   39764] = 32'h60f08b03;
    ram_cell[   39765] = 32'h4a9f4571;
    ram_cell[   39766] = 32'hc09fc38e;
    ram_cell[   39767] = 32'hb56e01b7;
    ram_cell[   39768] = 32'hf77c975f;
    ram_cell[   39769] = 32'h129f421e;
    ram_cell[   39770] = 32'h79b169ed;
    ram_cell[   39771] = 32'h66d6a170;
    ram_cell[   39772] = 32'h0c17f8a9;
    ram_cell[   39773] = 32'hdd58ff55;
    ram_cell[   39774] = 32'h8ee7a658;
    ram_cell[   39775] = 32'h142e5e5d;
    ram_cell[   39776] = 32'h70085c9b;
    ram_cell[   39777] = 32'hcc74248c;
    ram_cell[   39778] = 32'h1750a28f;
    ram_cell[   39779] = 32'h0b8de1c9;
    ram_cell[   39780] = 32'hf335d20f;
    ram_cell[   39781] = 32'h1e7feb99;
    ram_cell[   39782] = 32'hbad9fb5d;
    ram_cell[   39783] = 32'hb056642f;
    ram_cell[   39784] = 32'h70c79e62;
    ram_cell[   39785] = 32'h45cd531d;
    ram_cell[   39786] = 32'ha442f154;
    ram_cell[   39787] = 32'hb3480af6;
    ram_cell[   39788] = 32'h1168ef35;
    ram_cell[   39789] = 32'h539e53bd;
    ram_cell[   39790] = 32'h50bf4edc;
    ram_cell[   39791] = 32'h822edf92;
    ram_cell[   39792] = 32'h83f160cb;
    ram_cell[   39793] = 32'ha5bce44c;
    ram_cell[   39794] = 32'hab6174fa;
    ram_cell[   39795] = 32'he7e79df5;
    ram_cell[   39796] = 32'h81d326ed;
    ram_cell[   39797] = 32'h733f09ff;
    ram_cell[   39798] = 32'h1fff42ae;
    ram_cell[   39799] = 32'h7d4fd5a8;
    ram_cell[   39800] = 32'h4e9cf9bf;
    ram_cell[   39801] = 32'h5a441666;
    ram_cell[   39802] = 32'h45f07f8e;
    ram_cell[   39803] = 32'h2d7df5ad;
    ram_cell[   39804] = 32'h373ff1fa;
    ram_cell[   39805] = 32'h7f34cf69;
    ram_cell[   39806] = 32'h082ea793;
    ram_cell[   39807] = 32'h6badefab;
    ram_cell[   39808] = 32'hc1561aba;
    ram_cell[   39809] = 32'h6baa728e;
    ram_cell[   39810] = 32'h09c3899b;
    ram_cell[   39811] = 32'h2766498b;
    ram_cell[   39812] = 32'haefeced9;
    ram_cell[   39813] = 32'h73c396cd;
    ram_cell[   39814] = 32'h97bbd5f1;
    ram_cell[   39815] = 32'had43c8a3;
    ram_cell[   39816] = 32'h8949ed16;
    ram_cell[   39817] = 32'h633755a6;
    ram_cell[   39818] = 32'ha9547127;
    ram_cell[   39819] = 32'h6916649f;
    ram_cell[   39820] = 32'h87ea14ea;
    ram_cell[   39821] = 32'h3bf5604d;
    ram_cell[   39822] = 32'h64c8c7d9;
    ram_cell[   39823] = 32'hd8fc8750;
    ram_cell[   39824] = 32'h62dd8181;
    ram_cell[   39825] = 32'hea4b99b7;
    ram_cell[   39826] = 32'h30363ff8;
    ram_cell[   39827] = 32'hb085c48a;
    ram_cell[   39828] = 32'h0f6ecf21;
    ram_cell[   39829] = 32'h84ab2f77;
    ram_cell[   39830] = 32'hb3c6e8d2;
    ram_cell[   39831] = 32'hd095c3d5;
    ram_cell[   39832] = 32'h20922c6d;
    ram_cell[   39833] = 32'h6671c947;
    ram_cell[   39834] = 32'h719e2525;
    ram_cell[   39835] = 32'hbae011b9;
    ram_cell[   39836] = 32'h1a46b699;
    ram_cell[   39837] = 32'ha29210eb;
    ram_cell[   39838] = 32'hb4faa803;
    ram_cell[   39839] = 32'h03299046;
    ram_cell[   39840] = 32'h5902a0e3;
    ram_cell[   39841] = 32'hde0c9a39;
    ram_cell[   39842] = 32'h50cf2fd2;
    ram_cell[   39843] = 32'h57b37313;
    ram_cell[   39844] = 32'h575314da;
    ram_cell[   39845] = 32'h589917b7;
    ram_cell[   39846] = 32'h3300cebf;
    ram_cell[   39847] = 32'hf724dffc;
    ram_cell[   39848] = 32'h87042843;
    ram_cell[   39849] = 32'h50285671;
    ram_cell[   39850] = 32'h6fad25c5;
    ram_cell[   39851] = 32'h223e9273;
    ram_cell[   39852] = 32'h0c29182c;
    ram_cell[   39853] = 32'h3a9a1fef;
    ram_cell[   39854] = 32'h53eb6e5d;
    ram_cell[   39855] = 32'h0a28598f;
    ram_cell[   39856] = 32'ha04541fd;
    ram_cell[   39857] = 32'hcbbc36ea;
    ram_cell[   39858] = 32'h09bb5dd8;
    ram_cell[   39859] = 32'he95dcc1b;
    ram_cell[   39860] = 32'hd79dc45d;
    ram_cell[   39861] = 32'hfb2d3edb;
    ram_cell[   39862] = 32'hc7d7e482;
    ram_cell[   39863] = 32'hca4a4ba0;
    ram_cell[   39864] = 32'h025c67de;
    ram_cell[   39865] = 32'h814ef04d;
    ram_cell[   39866] = 32'hc26260ef;
    ram_cell[   39867] = 32'he08efb53;
    ram_cell[   39868] = 32'hd4a893b4;
    ram_cell[   39869] = 32'he8d54fb8;
    ram_cell[   39870] = 32'h61577493;
    ram_cell[   39871] = 32'h9bc31eaf;
    ram_cell[   39872] = 32'h80938d15;
    ram_cell[   39873] = 32'h6a6d189d;
    ram_cell[   39874] = 32'hb8ebfae1;
    ram_cell[   39875] = 32'h6776cdc6;
    ram_cell[   39876] = 32'hc904b462;
    ram_cell[   39877] = 32'h728a31e6;
    ram_cell[   39878] = 32'hb1d0e816;
    ram_cell[   39879] = 32'hcbf1e031;
    ram_cell[   39880] = 32'h2c4fda5e;
    ram_cell[   39881] = 32'he6c1414b;
    ram_cell[   39882] = 32'hd54989e6;
    ram_cell[   39883] = 32'h0fb562f0;
    ram_cell[   39884] = 32'hec9504bb;
    ram_cell[   39885] = 32'ha44070e9;
    ram_cell[   39886] = 32'h176e9eae;
    ram_cell[   39887] = 32'h0c8f6bae;
    ram_cell[   39888] = 32'h100499ee;
    ram_cell[   39889] = 32'h3f920760;
    ram_cell[   39890] = 32'h85fd14c1;
    ram_cell[   39891] = 32'h84a6acdb;
    ram_cell[   39892] = 32'h1007248f;
    ram_cell[   39893] = 32'h0687cfd4;
    ram_cell[   39894] = 32'he39c02be;
    ram_cell[   39895] = 32'h56659181;
    ram_cell[   39896] = 32'h3c0f9ec2;
    ram_cell[   39897] = 32'hf9b67bce;
    ram_cell[   39898] = 32'h6c925bc7;
    ram_cell[   39899] = 32'h4da2d0e4;
    ram_cell[   39900] = 32'h5eccef01;
    ram_cell[   39901] = 32'hd5dd0cfa;
    ram_cell[   39902] = 32'hf90295f7;
    ram_cell[   39903] = 32'h9af714be;
    ram_cell[   39904] = 32'h329d5d65;
    ram_cell[   39905] = 32'hcb7e49da;
    ram_cell[   39906] = 32'h2db0bbdb;
    ram_cell[   39907] = 32'h2b678be4;
    ram_cell[   39908] = 32'h34ce5eed;
    ram_cell[   39909] = 32'h29142011;
    ram_cell[   39910] = 32'hec2ec65a;
    ram_cell[   39911] = 32'h48cefa66;
    ram_cell[   39912] = 32'hb783bcd9;
    ram_cell[   39913] = 32'h966cb193;
    ram_cell[   39914] = 32'h793188a7;
    ram_cell[   39915] = 32'h29f9e313;
    ram_cell[   39916] = 32'ha23bd9b4;
    ram_cell[   39917] = 32'h456ebfca;
    ram_cell[   39918] = 32'h51fdbe9d;
    ram_cell[   39919] = 32'h23f1e1f4;
    ram_cell[   39920] = 32'h591dc888;
    ram_cell[   39921] = 32'he23a3c7c;
    ram_cell[   39922] = 32'h2fa55fed;
    ram_cell[   39923] = 32'h3994c9a8;
    ram_cell[   39924] = 32'h18016f87;
    ram_cell[   39925] = 32'hb0bc7a38;
    ram_cell[   39926] = 32'h7448ff16;
    ram_cell[   39927] = 32'hb3565e82;
    ram_cell[   39928] = 32'h4556be8f;
    ram_cell[   39929] = 32'h07b9c363;
    ram_cell[   39930] = 32'h8b3b7c8d;
    ram_cell[   39931] = 32'h2436066d;
    ram_cell[   39932] = 32'h262909f8;
    ram_cell[   39933] = 32'h7ace57f5;
    ram_cell[   39934] = 32'hf6b16c0e;
    ram_cell[   39935] = 32'h89f621d9;
    ram_cell[   39936] = 32'h1eca5d19;
    ram_cell[   39937] = 32'hb12d6abb;
    ram_cell[   39938] = 32'hb0eff0ad;
    ram_cell[   39939] = 32'hd117f113;
    ram_cell[   39940] = 32'haf83adcc;
    ram_cell[   39941] = 32'h53de9b13;
    ram_cell[   39942] = 32'h396fc57d;
    ram_cell[   39943] = 32'h17889446;
    ram_cell[   39944] = 32'h62b788cd;
    ram_cell[   39945] = 32'hbc6fca88;
    ram_cell[   39946] = 32'h68ab41aa;
    ram_cell[   39947] = 32'hd7a528b0;
    ram_cell[   39948] = 32'h1ae25b7a;
    ram_cell[   39949] = 32'h61222235;
    ram_cell[   39950] = 32'h59e83b87;
    ram_cell[   39951] = 32'h9d60dd7f;
    ram_cell[   39952] = 32'h22aeccbe;
    ram_cell[   39953] = 32'h84c64178;
    ram_cell[   39954] = 32'h7aa01d0d;
    ram_cell[   39955] = 32'h143d1dae;
    ram_cell[   39956] = 32'h1ee10383;
    ram_cell[   39957] = 32'h9f24cfa2;
    ram_cell[   39958] = 32'hb7b5ee4a;
    ram_cell[   39959] = 32'h1199abb0;
    ram_cell[   39960] = 32'he8b97bdf;
    ram_cell[   39961] = 32'h27d34403;
    ram_cell[   39962] = 32'h57763728;
    ram_cell[   39963] = 32'h27621950;
    ram_cell[   39964] = 32'h2563f28b;
    ram_cell[   39965] = 32'h7888f94b;
    ram_cell[   39966] = 32'hbbc0cdc0;
    ram_cell[   39967] = 32'h5eaf47eb;
    ram_cell[   39968] = 32'h41a055ac;
    ram_cell[   39969] = 32'h39aa6e87;
    ram_cell[   39970] = 32'ha8bbb20c;
    ram_cell[   39971] = 32'h898dce15;
    ram_cell[   39972] = 32'hc088819e;
    ram_cell[   39973] = 32'h24cd2706;
    ram_cell[   39974] = 32'h0918ddba;
    ram_cell[   39975] = 32'h6da09807;
    ram_cell[   39976] = 32'h616e99c2;
    ram_cell[   39977] = 32'hab303163;
    ram_cell[   39978] = 32'h11c2f026;
    ram_cell[   39979] = 32'ha0ade4f0;
    ram_cell[   39980] = 32'hf5129b53;
    ram_cell[   39981] = 32'h0e7c55ad;
    ram_cell[   39982] = 32'hbdc56cc6;
    ram_cell[   39983] = 32'h581f6b0a;
    ram_cell[   39984] = 32'h0af40670;
    ram_cell[   39985] = 32'h988ac830;
    ram_cell[   39986] = 32'h7e279b6a;
    ram_cell[   39987] = 32'h18043822;
    ram_cell[   39988] = 32'h8a63f08e;
    ram_cell[   39989] = 32'h8c483441;
    ram_cell[   39990] = 32'h09ea5738;
    ram_cell[   39991] = 32'hc9df9e2e;
    ram_cell[   39992] = 32'haa736f37;
    ram_cell[   39993] = 32'he20b1a73;
    ram_cell[   39994] = 32'h0db414e8;
    ram_cell[   39995] = 32'h6bd982d9;
    ram_cell[   39996] = 32'h5648ad4b;
    ram_cell[   39997] = 32'h38d13e85;
    ram_cell[   39998] = 32'hba79b6a8;
    ram_cell[   39999] = 32'h652f8059;
    ram_cell[   40000] = 32'hc14f16c8;
    ram_cell[   40001] = 32'h4b788206;
    ram_cell[   40002] = 32'h015ee4e7;
    ram_cell[   40003] = 32'h1dc28406;
    ram_cell[   40004] = 32'h5a47867f;
    ram_cell[   40005] = 32'h786dca4d;
    ram_cell[   40006] = 32'heeeee4fe;
    ram_cell[   40007] = 32'hf36807f5;
    ram_cell[   40008] = 32'hc0470966;
    ram_cell[   40009] = 32'h007db370;
    ram_cell[   40010] = 32'h796e7f08;
    ram_cell[   40011] = 32'hd7ef7100;
    ram_cell[   40012] = 32'h24667c76;
    ram_cell[   40013] = 32'h6a7d5560;
    ram_cell[   40014] = 32'ha3fba25b;
    ram_cell[   40015] = 32'h9a87e0c0;
    ram_cell[   40016] = 32'h5a9ae56e;
    ram_cell[   40017] = 32'hd37a4dab;
    ram_cell[   40018] = 32'h34bb00be;
    ram_cell[   40019] = 32'h7449fcd7;
    ram_cell[   40020] = 32'h78c8fd95;
    ram_cell[   40021] = 32'hbfcfcca3;
    ram_cell[   40022] = 32'hc2cc924d;
    ram_cell[   40023] = 32'hb921f28a;
    ram_cell[   40024] = 32'h893fe4c8;
    ram_cell[   40025] = 32'h842d803f;
    ram_cell[   40026] = 32'hc9f3d7ad;
    ram_cell[   40027] = 32'h7958a744;
    ram_cell[   40028] = 32'h590ffb15;
    ram_cell[   40029] = 32'h7b99737b;
    ram_cell[   40030] = 32'hcc690e1d;
    ram_cell[   40031] = 32'h1ff40b3a;
    ram_cell[   40032] = 32'hfe8a1087;
    ram_cell[   40033] = 32'h277b02b8;
    ram_cell[   40034] = 32'h05a39f1d;
    ram_cell[   40035] = 32'hdf093136;
    ram_cell[   40036] = 32'he9b2f5de;
    ram_cell[   40037] = 32'h103feaf4;
    ram_cell[   40038] = 32'hbb4592f6;
    ram_cell[   40039] = 32'h00d74a4b;
    ram_cell[   40040] = 32'he9ae1188;
    ram_cell[   40041] = 32'haaf3ef78;
    ram_cell[   40042] = 32'he77855d1;
    ram_cell[   40043] = 32'h1648654c;
    ram_cell[   40044] = 32'h9abbf8bc;
    ram_cell[   40045] = 32'h5fa90415;
    ram_cell[   40046] = 32'h65aeb6c7;
    ram_cell[   40047] = 32'h1615ce9e;
    ram_cell[   40048] = 32'hde791acc;
    ram_cell[   40049] = 32'h52d0997a;
    ram_cell[   40050] = 32'hc2daea12;
    ram_cell[   40051] = 32'h63cdde37;
    ram_cell[   40052] = 32'h6dde0d57;
    ram_cell[   40053] = 32'he9002d39;
    ram_cell[   40054] = 32'h16ebeb6e;
    ram_cell[   40055] = 32'hd30960d0;
    ram_cell[   40056] = 32'h946de19f;
    ram_cell[   40057] = 32'h161afcf2;
    ram_cell[   40058] = 32'hfdfe89ac;
    ram_cell[   40059] = 32'ha8737c50;
    ram_cell[   40060] = 32'h18105f37;
    ram_cell[   40061] = 32'hafe9aee0;
    ram_cell[   40062] = 32'h7435b588;
    ram_cell[   40063] = 32'h1178350d;
    ram_cell[   40064] = 32'hcb71ef32;
    ram_cell[   40065] = 32'h9b089ee6;
    ram_cell[   40066] = 32'hcb42d2dc;
    ram_cell[   40067] = 32'h31f47740;
    ram_cell[   40068] = 32'h1c2f8239;
    ram_cell[   40069] = 32'h89bfe35f;
    ram_cell[   40070] = 32'h9b8f27dd;
    ram_cell[   40071] = 32'hf50f6f0d;
    ram_cell[   40072] = 32'h72ceb831;
    ram_cell[   40073] = 32'h40d332a7;
    ram_cell[   40074] = 32'h7fb49121;
    ram_cell[   40075] = 32'h71c96b57;
    ram_cell[   40076] = 32'ha6e0f041;
    ram_cell[   40077] = 32'h00ce7e46;
    ram_cell[   40078] = 32'h1a33f5cd;
    ram_cell[   40079] = 32'h8e1c3f6a;
    ram_cell[   40080] = 32'h73ee3bb6;
    ram_cell[   40081] = 32'hac10a895;
    ram_cell[   40082] = 32'hc386491c;
    ram_cell[   40083] = 32'h0a1299e5;
    ram_cell[   40084] = 32'h7a39c993;
    ram_cell[   40085] = 32'hdd42cd05;
    ram_cell[   40086] = 32'h6ce55350;
    ram_cell[   40087] = 32'he34ac26f;
    ram_cell[   40088] = 32'hd9ae5a6c;
    ram_cell[   40089] = 32'hf512d75d;
    ram_cell[   40090] = 32'h73653995;
    ram_cell[   40091] = 32'h23453ba8;
    ram_cell[   40092] = 32'he736f1db;
    ram_cell[   40093] = 32'ha8d97bc4;
    ram_cell[   40094] = 32'h096b0c13;
    ram_cell[   40095] = 32'h044a2ee0;
    ram_cell[   40096] = 32'hceec51ec;
    ram_cell[   40097] = 32'h11dea368;
    ram_cell[   40098] = 32'hc869560a;
    ram_cell[   40099] = 32'h064118fd;
    ram_cell[   40100] = 32'h107d6547;
    ram_cell[   40101] = 32'h10bbb9c0;
    ram_cell[   40102] = 32'h86c2ea23;
    ram_cell[   40103] = 32'h800aa629;
    ram_cell[   40104] = 32'h6c27adf9;
    ram_cell[   40105] = 32'h34a3bf66;
    ram_cell[   40106] = 32'hc91f1b45;
    ram_cell[   40107] = 32'he55658a6;
    ram_cell[   40108] = 32'he4faeb23;
    ram_cell[   40109] = 32'hb194acb2;
    ram_cell[   40110] = 32'hd0b80324;
    ram_cell[   40111] = 32'he14d7aaa;
    ram_cell[   40112] = 32'h52b65a81;
    ram_cell[   40113] = 32'h975274f8;
    ram_cell[   40114] = 32'h483b1c0a;
    ram_cell[   40115] = 32'h824a84ee;
    ram_cell[   40116] = 32'hfcc72a52;
    ram_cell[   40117] = 32'h7311692d;
    ram_cell[   40118] = 32'h79570204;
    ram_cell[   40119] = 32'h22f56536;
    ram_cell[   40120] = 32'h98cd4a07;
    ram_cell[   40121] = 32'h44944653;
    ram_cell[   40122] = 32'h51be0940;
    ram_cell[   40123] = 32'h3db7b67a;
    ram_cell[   40124] = 32'hbb990de5;
    ram_cell[   40125] = 32'habc0666e;
    ram_cell[   40126] = 32'h9f36264b;
    ram_cell[   40127] = 32'ha343d367;
    ram_cell[   40128] = 32'h44671559;
    ram_cell[   40129] = 32'hbdd47f77;
    ram_cell[   40130] = 32'hb716de1b;
    ram_cell[   40131] = 32'hff2f0f6a;
    ram_cell[   40132] = 32'h5cfbecca;
    ram_cell[   40133] = 32'hcf29ca22;
    ram_cell[   40134] = 32'h324bd05b;
    ram_cell[   40135] = 32'h8f6e4dfa;
    ram_cell[   40136] = 32'hdaefaa76;
    ram_cell[   40137] = 32'h17c773a5;
    ram_cell[   40138] = 32'h09ff2ca3;
    ram_cell[   40139] = 32'h8105b941;
    ram_cell[   40140] = 32'h2fc0d057;
    ram_cell[   40141] = 32'h17495819;
    ram_cell[   40142] = 32'hcc2213a0;
    ram_cell[   40143] = 32'h65a0a8f4;
    ram_cell[   40144] = 32'h7ef193ae;
    ram_cell[   40145] = 32'h498aa89f;
    ram_cell[   40146] = 32'h2cb684bf;
    ram_cell[   40147] = 32'h660b80a2;
    ram_cell[   40148] = 32'hcde0e866;
    ram_cell[   40149] = 32'h0eabfa70;
    ram_cell[   40150] = 32'h265bb685;
    ram_cell[   40151] = 32'h61cfff9e;
    ram_cell[   40152] = 32'h3fc210e2;
    ram_cell[   40153] = 32'hbfe0cadc;
    ram_cell[   40154] = 32'hf8f2974d;
    ram_cell[   40155] = 32'h24f7242d;
    ram_cell[   40156] = 32'h02fd92f8;
    ram_cell[   40157] = 32'hb0a67e05;
    ram_cell[   40158] = 32'h0c7b7f14;
    ram_cell[   40159] = 32'h58b96077;
    ram_cell[   40160] = 32'ha3347e91;
    ram_cell[   40161] = 32'h13d581e7;
    ram_cell[   40162] = 32'h520b5ee6;
    ram_cell[   40163] = 32'h7d617e71;
    ram_cell[   40164] = 32'hf55542a5;
    ram_cell[   40165] = 32'h9d8fa5d3;
    ram_cell[   40166] = 32'h84b6f8f3;
    ram_cell[   40167] = 32'hc6aa9e4f;
    ram_cell[   40168] = 32'h8b03aacd;
    ram_cell[   40169] = 32'h84d8f1eb;
    ram_cell[   40170] = 32'h5933933e;
    ram_cell[   40171] = 32'h7d27b180;
    ram_cell[   40172] = 32'h3a05ebb2;
    ram_cell[   40173] = 32'hf6249079;
    ram_cell[   40174] = 32'hbd295775;
    ram_cell[   40175] = 32'he5a1171a;
    ram_cell[   40176] = 32'h83b4b8a0;
    ram_cell[   40177] = 32'h1ecae43d;
    ram_cell[   40178] = 32'h9fb13280;
    ram_cell[   40179] = 32'h240b710f;
    ram_cell[   40180] = 32'ha45c040e;
    ram_cell[   40181] = 32'h15049cfe;
    ram_cell[   40182] = 32'h85ac993b;
    ram_cell[   40183] = 32'h76e40cce;
    ram_cell[   40184] = 32'h75cb74c2;
    ram_cell[   40185] = 32'h1577aa32;
    ram_cell[   40186] = 32'h2d092506;
    ram_cell[   40187] = 32'h0c21f401;
    ram_cell[   40188] = 32'h737c21d5;
    ram_cell[   40189] = 32'hce98ffbf;
    ram_cell[   40190] = 32'h643194b7;
    ram_cell[   40191] = 32'hba1e73f2;
    ram_cell[   40192] = 32'h1e00b618;
    ram_cell[   40193] = 32'h3ef67235;
    ram_cell[   40194] = 32'h2f858b2b;
    ram_cell[   40195] = 32'ha700362d;
    ram_cell[   40196] = 32'h1768ef0c;
    ram_cell[   40197] = 32'h13b55516;
    ram_cell[   40198] = 32'h810166cb;
    ram_cell[   40199] = 32'hbb3e836f;
    ram_cell[   40200] = 32'h3a539010;
    ram_cell[   40201] = 32'h87de5494;
    ram_cell[   40202] = 32'h4666173b;
    ram_cell[   40203] = 32'ha8085ae2;
    ram_cell[   40204] = 32'h9ab4e52a;
    ram_cell[   40205] = 32'hd307f882;
    ram_cell[   40206] = 32'h75ebd207;
    ram_cell[   40207] = 32'h3d183e65;
    ram_cell[   40208] = 32'h30ba2440;
    ram_cell[   40209] = 32'hd19ca856;
    ram_cell[   40210] = 32'h74700544;
    ram_cell[   40211] = 32'h1aa1a264;
    ram_cell[   40212] = 32'h65fb95c4;
    ram_cell[   40213] = 32'h61086809;
    ram_cell[   40214] = 32'hfd35b9de;
    ram_cell[   40215] = 32'h51254a61;
    ram_cell[   40216] = 32'hdd07f4ab;
    ram_cell[   40217] = 32'h7b812b29;
    ram_cell[   40218] = 32'hfbf4d53d;
    ram_cell[   40219] = 32'h7faf682d;
    ram_cell[   40220] = 32'h6c12d7c4;
    ram_cell[   40221] = 32'he482b783;
    ram_cell[   40222] = 32'hb8f2b71d;
    ram_cell[   40223] = 32'h4bc56bad;
    ram_cell[   40224] = 32'h501f919a;
    ram_cell[   40225] = 32'ha881d29d;
    ram_cell[   40226] = 32'h55a387a1;
    ram_cell[   40227] = 32'he0082fe5;
    ram_cell[   40228] = 32'h1117e811;
    ram_cell[   40229] = 32'h77d6cac5;
    ram_cell[   40230] = 32'h2f5f7bfd;
    ram_cell[   40231] = 32'h3fa7efb8;
    ram_cell[   40232] = 32'h03ea1296;
    ram_cell[   40233] = 32'h07708c84;
    ram_cell[   40234] = 32'h36e5ddbb;
    ram_cell[   40235] = 32'h352a4bbe;
    ram_cell[   40236] = 32'h288f0b9f;
    ram_cell[   40237] = 32'hc3132db4;
    ram_cell[   40238] = 32'ha7c3ba29;
    ram_cell[   40239] = 32'h47c7b48f;
    ram_cell[   40240] = 32'h8fcf3940;
    ram_cell[   40241] = 32'hc49386fb;
    ram_cell[   40242] = 32'hed22040c;
    ram_cell[   40243] = 32'h13774b3d;
    ram_cell[   40244] = 32'h856cb94d;
    ram_cell[   40245] = 32'hf6a979b3;
    ram_cell[   40246] = 32'h08569bb9;
    ram_cell[   40247] = 32'ha5d47d72;
    ram_cell[   40248] = 32'h95c45cae;
    ram_cell[   40249] = 32'hef0e77a7;
    ram_cell[   40250] = 32'he01b4df4;
    ram_cell[   40251] = 32'hddaf85a6;
    ram_cell[   40252] = 32'hd81eaf70;
    ram_cell[   40253] = 32'h2f54f25b;
    ram_cell[   40254] = 32'h1fcb22b2;
    ram_cell[   40255] = 32'he62c35ca;
    ram_cell[   40256] = 32'he6cc7c8b;
    ram_cell[   40257] = 32'hecef9dd6;
    ram_cell[   40258] = 32'h413f98bb;
    ram_cell[   40259] = 32'h418a90e3;
    ram_cell[   40260] = 32'h9043cd45;
    ram_cell[   40261] = 32'haf6fe53e;
    ram_cell[   40262] = 32'hd4e91c66;
    ram_cell[   40263] = 32'ha3636674;
    ram_cell[   40264] = 32'hceeae44d;
    ram_cell[   40265] = 32'h223a3c60;
    ram_cell[   40266] = 32'hef69898a;
    ram_cell[   40267] = 32'h8a9d9d51;
    ram_cell[   40268] = 32'h01bad160;
    ram_cell[   40269] = 32'h47bebab2;
    ram_cell[   40270] = 32'h620a8a7f;
    ram_cell[   40271] = 32'h99d191b7;
    ram_cell[   40272] = 32'hec9160ee;
    ram_cell[   40273] = 32'heb219399;
    ram_cell[   40274] = 32'he76bbf46;
    ram_cell[   40275] = 32'hb8144b3e;
    ram_cell[   40276] = 32'h48334fa1;
    ram_cell[   40277] = 32'h43f12a1c;
    ram_cell[   40278] = 32'he6eadd56;
    ram_cell[   40279] = 32'hc4d29e1a;
    ram_cell[   40280] = 32'h7409cef8;
    ram_cell[   40281] = 32'h90fc0d7d;
    ram_cell[   40282] = 32'hdb65e31a;
    ram_cell[   40283] = 32'h4e645af2;
    ram_cell[   40284] = 32'h0704708a;
    ram_cell[   40285] = 32'h90bc0a3c;
    ram_cell[   40286] = 32'he05312d5;
    ram_cell[   40287] = 32'h94a59244;
    ram_cell[   40288] = 32'hb98dae50;
    ram_cell[   40289] = 32'h00fd5eb1;
    ram_cell[   40290] = 32'hdaad1ddf;
    ram_cell[   40291] = 32'h885de959;
    ram_cell[   40292] = 32'hda4c7b7c;
    ram_cell[   40293] = 32'h719c123b;
    ram_cell[   40294] = 32'h608047c9;
    ram_cell[   40295] = 32'hb89fa0c8;
    ram_cell[   40296] = 32'ha070bf1a;
    ram_cell[   40297] = 32'h6e24d085;
    ram_cell[   40298] = 32'h2a4354ac;
    ram_cell[   40299] = 32'hf3e4f86e;
    ram_cell[   40300] = 32'hcce40221;
    ram_cell[   40301] = 32'h3f9ab3b4;
    ram_cell[   40302] = 32'h198c6138;
    ram_cell[   40303] = 32'h7900afab;
    ram_cell[   40304] = 32'hfbce3f40;
    ram_cell[   40305] = 32'h20bddaa4;
    ram_cell[   40306] = 32'hcce7c3c1;
    ram_cell[   40307] = 32'h3f28cf02;
    ram_cell[   40308] = 32'h3d7cef77;
    ram_cell[   40309] = 32'h265550bb;
    ram_cell[   40310] = 32'hf861d071;
    ram_cell[   40311] = 32'h4ce66749;
    ram_cell[   40312] = 32'h055f4995;
    ram_cell[   40313] = 32'h80869503;
    ram_cell[   40314] = 32'hf128ba4d;
    ram_cell[   40315] = 32'he056016f;
    ram_cell[   40316] = 32'he31cb83a;
    ram_cell[   40317] = 32'h6413ea34;
    ram_cell[   40318] = 32'h3eb23554;
    ram_cell[   40319] = 32'hf46da264;
    ram_cell[   40320] = 32'h4faa6d11;
    ram_cell[   40321] = 32'h81630e18;
    ram_cell[   40322] = 32'hf5fe102e;
    ram_cell[   40323] = 32'h08bf1af4;
    ram_cell[   40324] = 32'h51d3eedc;
    ram_cell[   40325] = 32'hb89ea615;
    ram_cell[   40326] = 32'hf58d0538;
    ram_cell[   40327] = 32'h7f9b47ab;
    ram_cell[   40328] = 32'hdf9bcf8a;
    ram_cell[   40329] = 32'h90c2d4ba;
    ram_cell[   40330] = 32'hd57c7bd9;
    ram_cell[   40331] = 32'h9c8b1fbf;
    ram_cell[   40332] = 32'h70fd582a;
    ram_cell[   40333] = 32'hecb0c04e;
    ram_cell[   40334] = 32'h1090c0d1;
    ram_cell[   40335] = 32'h35cdd948;
    ram_cell[   40336] = 32'hb4defe12;
    ram_cell[   40337] = 32'h9f131d05;
    ram_cell[   40338] = 32'h38e18803;
    ram_cell[   40339] = 32'hf89d70aa;
    ram_cell[   40340] = 32'hbb55708f;
    ram_cell[   40341] = 32'h7dcc7642;
    ram_cell[   40342] = 32'h6280a761;
    ram_cell[   40343] = 32'hfacf6dbb;
    ram_cell[   40344] = 32'hdbb8c7b3;
    ram_cell[   40345] = 32'h8ab53336;
    ram_cell[   40346] = 32'h152e457d;
    ram_cell[   40347] = 32'h2ec1abc5;
    ram_cell[   40348] = 32'hf2d333fe;
    ram_cell[   40349] = 32'heace7331;
    ram_cell[   40350] = 32'h79bb83ec;
    ram_cell[   40351] = 32'hfef0f502;
    ram_cell[   40352] = 32'h2eeabbae;
    ram_cell[   40353] = 32'h9015dc3f;
    ram_cell[   40354] = 32'h81b0e480;
    ram_cell[   40355] = 32'h8fd27de2;
    ram_cell[   40356] = 32'hdcc4d509;
    ram_cell[   40357] = 32'he06594e4;
    ram_cell[   40358] = 32'h596d3a03;
    ram_cell[   40359] = 32'ha6154b1b;
    ram_cell[   40360] = 32'h8a5e1128;
    ram_cell[   40361] = 32'hcabae096;
    ram_cell[   40362] = 32'hadfd2064;
    ram_cell[   40363] = 32'hffd672dc;
    ram_cell[   40364] = 32'hb3ea2370;
    ram_cell[   40365] = 32'h1f696d0a;
    ram_cell[   40366] = 32'h34e0aed6;
    ram_cell[   40367] = 32'h1b546ea6;
    ram_cell[   40368] = 32'hf71b7e82;
    ram_cell[   40369] = 32'h27a4e92f;
    ram_cell[   40370] = 32'hecd006d6;
    ram_cell[   40371] = 32'hc39e1549;
    ram_cell[   40372] = 32'he4985a9b;
    ram_cell[   40373] = 32'hdda178c7;
    ram_cell[   40374] = 32'h5c9c66da;
    ram_cell[   40375] = 32'heb664f20;
    ram_cell[   40376] = 32'h4d40fe6a;
    ram_cell[   40377] = 32'hef564331;
    ram_cell[   40378] = 32'hf444e88c;
    ram_cell[   40379] = 32'h82041ba4;
    ram_cell[   40380] = 32'h1d294717;
    ram_cell[   40381] = 32'hdae4e61d;
    ram_cell[   40382] = 32'h355072e1;
    ram_cell[   40383] = 32'haf977eba;
    ram_cell[   40384] = 32'hfc8693df;
    ram_cell[   40385] = 32'h52bfa3f3;
    ram_cell[   40386] = 32'h94234ff9;
    ram_cell[   40387] = 32'h76812405;
    ram_cell[   40388] = 32'hd0ceebbf;
    ram_cell[   40389] = 32'h7e27f2d7;
    ram_cell[   40390] = 32'hd9667d53;
    ram_cell[   40391] = 32'h6f2cbf58;
    ram_cell[   40392] = 32'h4c93fcaa;
    ram_cell[   40393] = 32'h143ebe8c;
    ram_cell[   40394] = 32'hee62a6f2;
    ram_cell[   40395] = 32'h8de7b6c5;
    ram_cell[   40396] = 32'hedbec567;
    ram_cell[   40397] = 32'h24479209;
    ram_cell[   40398] = 32'h67501817;
    ram_cell[   40399] = 32'h87439b8f;
    ram_cell[   40400] = 32'h9b7e5f1b;
    ram_cell[   40401] = 32'h1eb3c4dc;
    ram_cell[   40402] = 32'h46db7f9b;
    ram_cell[   40403] = 32'ha76f2845;
    ram_cell[   40404] = 32'h10b04696;
    ram_cell[   40405] = 32'h218d1db5;
    ram_cell[   40406] = 32'h29d527c4;
    ram_cell[   40407] = 32'he8402dbe;
    ram_cell[   40408] = 32'h7fe9dbf2;
    ram_cell[   40409] = 32'ha9d9e53e;
    ram_cell[   40410] = 32'h6bba9b7a;
    ram_cell[   40411] = 32'hfedac020;
    ram_cell[   40412] = 32'h5865bff4;
    ram_cell[   40413] = 32'he9d3897e;
    ram_cell[   40414] = 32'h10e735b9;
    ram_cell[   40415] = 32'h8b192b10;
    ram_cell[   40416] = 32'hfbbccb2f;
    ram_cell[   40417] = 32'h60307363;
    ram_cell[   40418] = 32'hfe3195a9;
    ram_cell[   40419] = 32'h354d2581;
    ram_cell[   40420] = 32'ha53d56d1;
    ram_cell[   40421] = 32'hf198c067;
    ram_cell[   40422] = 32'h93632c0f;
    ram_cell[   40423] = 32'h885be22b;
    ram_cell[   40424] = 32'hd7354f13;
    ram_cell[   40425] = 32'h1f897e2c;
    ram_cell[   40426] = 32'he0531427;
    ram_cell[   40427] = 32'h5a9759b6;
    ram_cell[   40428] = 32'h48700910;
    ram_cell[   40429] = 32'h3d5e66a3;
    ram_cell[   40430] = 32'hcfa9d1a7;
    ram_cell[   40431] = 32'hb8967861;
    ram_cell[   40432] = 32'h1035d315;
    ram_cell[   40433] = 32'h434735f4;
    ram_cell[   40434] = 32'h9548ed96;
    ram_cell[   40435] = 32'hee70989e;
    ram_cell[   40436] = 32'he8f6bba4;
    ram_cell[   40437] = 32'h67bb5306;
    ram_cell[   40438] = 32'h218e8a77;
    ram_cell[   40439] = 32'h400b86a0;
    ram_cell[   40440] = 32'h0f1903d5;
    ram_cell[   40441] = 32'h9a216184;
    ram_cell[   40442] = 32'he1d92184;
    ram_cell[   40443] = 32'h2e0b1d12;
    ram_cell[   40444] = 32'h53694697;
    ram_cell[   40445] = 32'ha5bdfd4f;
    ram_cell[   40446] = 32'hd55d0172;
    ram_cell[   40447] = 32'h53fc9ffc;
    ram_cell[   40448] = 32'h9a6a70a6;
    ram_cell[   40449] = 32'h214181a0;
    ram_cell[   40450] = 32'h1c708e68;
    ram_cell[   40451] = 32'h4a2ea159;
    ram_cell[   40452] = 32'h345f081d;
    ram_cell[   40453] = 32'h92d7592d;
    ram_cell[   40454] = 32'h463fc787;
    ram_cell[   40455] = 32'h1e17dd91;
    ram_cell[   40456] = 32'h133f52ff;
    ram_cell[   40457] = 32'hc8752dea;
    ram_cell[   40458] = 32'hed14e21c;
    ram_cell[   40459] = 32'h56b04853;
    ram_cell[   40460] = 32'h936ae64b;
    ram_cell[   40461] = 32'hb0dc98d7;
    ram_cell[   40462] = 32'h73df8a35;
    ram_cell[   40463] = 32'h72debad6;
    ram_cell[   40464] = 32'h59a5d13a;
    ram_cell[   40465] = 32'hdfccec27;
    ram_cell[   40466] = 32'hba861c80;
    ram_cell[   40467] = 32'h87e1e4e4;
    ram_cell[   40468] = 32'h17a72721;
    ram_cell[   40469] = 32'h5f410133;
    ram_cell[   40470] = 32'hd979a09d;
    ram_cell[   40471] = 32'h0fb35359;
    ram_cell[   40472] = 32'h5db84db8;
    ram_cell[   40473] = 32'hf6561b8e;
    ram_cell[   40474] = 32'hf2465ab8;
    ram_cell[   40475] = 32'h8ce92bfb;
    ram_cell[   40476] = 32'h0d629347;
    ram_cell[   40477] = 32'h19e91916;
    ram_cell[   40478] = 32'h5870a3b3;
    ram_cell[   40479] = 32'h156208b4;
    ram_cell[   40480] = 32'hf7663e95;
    ram_cell[   40481] = 32'hb4370879;
    ram_cell[   40482] = 32'h99108710;
    ram_cell[   40483] = 32'h76c58a89;
    ram_cell[   40484] = 32'h064d77f9;
    ram_cell[   40485] = 32'h35d8223e;
    ram_cell[   40486] = 32'hfccb681b;
    ram_cell[   40487] = 32'hf1da7d01;
    ram_cell[   40488] = 32'h46825083;
    ram_cell[   40489] = 32'hea4d85e0;
    ram_cell[   40490] = 32'h58411677;
    ram_cell[   40491] = 32'hc7c23a9b;
    ram_cell[   40492] = 32'h40e3f76e;
    ram_cell[   40493] = 32'h9d14a643;
    ram_cell[   40494] = 32'h8d0e9622;
    ram_cell[   40495] = 32'hc2f0f017;
    ram_cell[   40496] = 32'h84fe5f66;
    ram_cell[   40497] = 32'h71a22862;
    ram_cell[   40498] = 32'h8d3b2825;
    ram_cell[   40499] = 32'h47e802a8;
    ram_cell[   40500] = 32'hb360e294;
    ram_cell[   40501] = 32'h6f1c63bc;
    ram_cell[   40502] = 32'hb6fc8424;
    ram_cell[   40503] = 32'h00295af8;
    ram_cell[   40504] = 32'h50dc291e;
    ram_cell[   40505] = 32'h5ee49b59;
    ram_cell[   40506] = 32'hc425227f;
    ram_cell[   40507] = 32'h5bcc66f7;
    ram_cell[   40508] = 32'h054bc464;
    ram_cell[   40509] = 32'h989a8e36;
    ram_cell[   40510] = 32'h788908b3;
    ram_cell[   40511] = 32'hd36f615b;
    ram_cell[   40512] = 32'he838dea9;
    ram_cell[   40513] = 32'h33f06562;
    ram_cell[   40514] = 32'hc354a5c0;
    ram_cell[   40515] = 32'h6447daf7;
    ram_cell[   40516] = 32'h2515b197;
    ram_cell[   40517] = 32'h622a9807;
    ram_cell[   40518] = 32'h37670204;
    ram_cell[   40519] = 32'h6bd3177f;
    ram_cell[   40520] = 32'hbf5cd47c;
    ram_cell[   40521] = 32'h6d2ddd58;
    ram_cell[   40522] = 32'h4a7e2830;
    ram_cell[   40523] = 32'ha37c7844;
    ram_cell[   40524] = 32'h704c2261;
    ram_cell[   40525] = 32'h5510ddc0;
    ram_cell[   40526] = 32'hb887ed07;
    ram_cell[   40527] = 32'h00b23f14;
    ram_cell[   40528] = 32'hc6055492;
    ram_cell[   40529] = 32'h8f5c70cb;
    ram_cell[   40530] = 32'hdfb151cf;
    ram_cell[   40531] = 32'hbcfa51d3;
    ram_cell[   40532] = 32'h718419e2;
    ram_cell[   40533] = 32'h32d47106;
    ram_cell[   40534] = 32'h7f1e160d;
    ram_cell[   40535] = 32'h328afc7d;
    ram_cell[   40536] = 32'hb321cbb6;
    ram_cell[   40537] = 32'h1479eede;
    ram_cell[   40538] = 32'h6c17dcd0;
    ram_cell[   40539] = 32'hd15f5114;
    ram_cell[   40540] = 32'h33702dbe;
    ram_cell[   40541] = 32'hb5d0e993;
    ram_cell[   40542] = 32'h583b8364;
    ram_cell[   40543] = 32'h73f81813;
    ram_cell[   40544] = 32'h21e50c01;
    ram_cell[   40545] = 32'hd92b9a2a;
    ram_cell[   40546] = 32'h3d509c20;
    ram_cell[   40547] = 32'ha5f87fc9;
    ram_cell[   40548] = 32'h3f32ba8e;
    ram_cell[   40549] = 32'h86abeada;
    ram_cell[   40550] = 32'hb1e20f77;
    ram_cell[   40551] = 32'hb203603c;
    ram_cell[   40552] = 32'hcdcefe92;
    ram_cell[   40553] = 32'hf713a97a;
    ram_cell[   40554] = 32'h0b1b846c;
    ram_cell[   40555] = 32'h8c5ff025;
    ram_cell[   40556] = 32'hee16cb5d;
    ram_cell[   40557] = 32'h33ed0657;
    ram_cell[   40558] = 32'h81531e70;
    ram_cell[   40559] = 32'h3eddb164;
    ram_cell[   40560] = 32'hb5fc6f8d;
    ram_cell[   40561] = 32'h921e617a;
    ram_cell[   40562] = 32'h3cffcb07;
    ram_cell[   40563] = 32'h0da11394;
    ram_cell[   40564] = 32'h523fc214;
    ram_cell[   40565] = 32'h5ac59d96;
    ram_cell[   40566] = 32'h7be8b73f;
    ram_cell[   40567] = 32'h7ce2c867;
    ram_cell[   40568] = 32'he0de0406;
    ram_cell[   40569] = 32'h56c4e83f;
    ram_cell[   40570] = 32'h32edd1a4;
    ram_cell[   40571] = 32'hc81899d3;
    ram_cell[   40572] = 32'ha279274a;
    ram_cell[   40573] = 32'h48fed640;
    ram_cell[   40574] = 32'hf665baab;
    ram_cell[   40575] = 32'h3691fc62;
    ram_cell[   40576] = 32'he21dbe13;
    ram_cell[   40577] = 32'h0f26bd06;
    ram_cell[   40578] = 32'h10224381;
    ram_cell[   40579] = 32'h47549ac4;
    ram_cell[   40580] = 32'h13d08f4e;
    ram_cell[   40581] = 32'h2d780485;
    ram_cell[   40582] = 32'ha688e0a8;
    ram_cell[   40583] = 32'h56f94a21;
    ram_cell[   40584] = 32'hfae68c89;
    ram_cell[   40585] = 32'hfea0ede9;
    ram_cell[   40586] = 32'h0be7d8d9;
    ram_cell[   40587] = 32'h77ae3bdc;
    ram_cell[   40588] = 32'h79dea692;
    ram_cell[   40589] = 32'h854cceb9;
    ram_cell[   40590] = 32'ha2dcbfa5;
    ram_cell[   40591] = 32'hce969281;
    ram_cell[   40592] = 32'h9bed7d59;
    ram_cell[   40593] = 32'h8f52f60e;
    ram_cell[   40594] = 32'hb61598dc;
    ram_cell[   40595] = 32'h7c886fa9;
    ram_cell[   40596] = 32'hecc6f56c;
    ram_cell[   40597] = 32'h60cb72ab;
    ram_cell[   40598] = 32'h3c8e4a36;
    ram_cell[   40599] = 32'h842bb7a9;
    ram_cell[   40600] = 32'h0102633d;
    ram_cell[   40601] = 32'he80abe80;
    ram_cell[   40602] = 32'h9a781fa3;
    ram_cell[   40603] = 32'h00ec74fd;
    ram_cell[   40604] = 32'h1fa8a04d;
    ram_cell[   40605] = 32'h8ad82ee8;
    ram_cell[   40606] = 32'hfad2b7e5;
    ram_cell[   40607] = 32'h361659e1;
    ram_cell[   40608] = 32'h2990ae46;
    ram_cell[   40609] = 32'h38e2184f;
    ram_cell[   40610] = 32'h74e5068a;
    ram_cell[   40611] = 32'h9c228da1;
    ram_cell[   40612] = 32'h63029291;
    ram_cell[   40613] = 32'hef0edd79;
    ram_cell[   40614] = 32'h8c0f8bba;
    ram_cell[   40615] = 32'h6cafe3b3;
    ram_cell[   40616] = 32'h7c08dc88;
    ram_cell[   40617] = 32'h758fae4d;
    ram_cell[   40618] = 32'h406dc797;
    ram_cell[   40619] = 32'h63d19134;
    ram_cell[   40620] = 32'h49fc4a3f;
    ram_cell[   40621] = 32'he37a9740;
    ram_cell[   40622] = 32'h2a039e71;
    ram_cell[   40623] = 32'h17497e8f;
    ram_cell[   40624] = 32'h83774fdc;
    ram_cell[   40625] = 32'hb34fb6c3;
    ram_cell[   40626] = 32'h688d3b8c;
    ram_cell[   40627] = 32'h8390b1c7;
    ram_cell[   40628] = 32'h0030c3b9;
    ram_cell[   40629] = 32'h9c2cf65c;
    ram_cell[   40630] = 32'ha18bc570;
    ram_cell[   40631] = 32'h615253be;
    ram_cell[   40632] = 32'h27b3ee18;
    ram_cell[   40633] = 32'h44498df1;
    ram_cell[   40634] = 32'h592b9e80;
    ram_cell[   40635] = 32'hf062492a;
    ram_cell[   40636] = 32'h0166de67;
    ram_cell[   40637] = 32'h06a3f955;
    ram_cell[   40638] = 32'h59ab634a;
    ram_cell[   40639] = 32'hc73449e0;
    ram_cell[   40640] = 32'hc536bccd;
    ram_cell[   40641] = 32'h4cd957ba;
    ram_cell[   40642] = 32'h7bd6cd41;
    ram_cell[   40643] = 32'h36cf3245;
    ram_cell[   40644] = 32'he0582f73;
    ram_cell[   40645] = 32'ha19b5009;
    ram_cell[   40646] = 32'h9aecd896;
    ram_cell[   40647] = 32'hd2097461;
    ram_cell[   40648] = 32'h0d30b0bd;
    ram_cell[   40649] = 32'hce4dc69a;
    ram_cell[   40650] = 32'h1e392524;
    ram_cell[   40651] = 32'h16d26e41;
    ram_cell[   40652] = 32'h0631b8e1;
    ram_cell[   40653] = 32'hd6dd01a2;
    ram_cell[   40654] = 32'h867913c8;
    ram_cell[   40655] = 32'ha764ca18;
    ram_cell[   40656] = 32'ha74bc6cd;
    ram_cell[   40657] = 32'h0e5760e5;
    ram_cell[   40658] = 32'h4e103ec4;
    ram_cell[   40659] = 32'h1dfa9a2b;
    ram_cell[   40660] = 32'h098802df;
    ram_cell[   40661] = 32'h46c151a5;
    ram_cell[   40662] = 32'h80a800cd;
    ram_cell[   40663] = 32'h547630bc;
    ram_cell[   40664] = 32'h473204cb;
    ram_cell[   40665] = 32'h9ef456b2;
    ram_cell[   40666] = 32'h7ee0fc8e;
    ram_cell[   40667] = 32'hf7f9285d;
    ram_cell[   40668] = 32'h5d976365;
    ram_cell[   40669] = 32'hd4304fee;
    ram_cell[   40670] = 32'hb430b0bd;
    ram_cell[   40671] = 32'he639e10c;
    ram_cell[   40672] = 32'h082220a0;
    ram_cell[   40673] = 32'hdef42209;
    ram_cell[   40674] = 32'h87d9750e;
    ram_cell[   40675] = 32'h55067a46;
    ram_cell[   40676] = 32'hec43f621;
    ram_cell[   40677] = 32'ha78da4cf;
    ram_cell[   40678] = 32'hf738c72c;
    ram_cell[   40679] = 32'h7f67a2e5;
    ram_cell[   40680] = 32'ha095c07e;
    ram_cell[   40681] = 32'ha45a205a;
    ram_cell[   40682] = 32'h4277ac1d;
    ram_cell[   40683] = 32'ha7c0213d;
    ram_cell[   40684] = 32'heefdb3d9;
    ram_cell[   40685] = 32'h7ed4bcff;
    ram_cell[   40686] = 32'h49d74982;
    ram_cell[   40687] = 32'h3a1a950b;
    ram_cell[   40688] = 32'h39cad869;
    ram_cell[   40689] = 32'h28ab3729;
    ram_cell[   40690] = 32'h63069dcc;
    ram_cell[   40691] = 32'h2a4bec8d;
    ram_cell[   40692] = 32'h5398481d;
    ram_cell[   40693] = 32'hc969d2bd;
    ram_cell[   40694] = 32'h42147872;
    ram_cell[   40695] = 32'he7e9e32e;
    ram_cell[   40696] = 32'h22f297aa;
    ram_cell[   40697] = 32'hc3c54292;
    ram_cell[   40698] = 32'he2838473;
    ram_cell[   40699] = 32'hebb507da;
    ram_cell[   40700] = 32'h7d3be093;
    ram_cell[   40701] = 32'hb1eafb41;
    ram_cell[   40702] = 32'h618331d0;
    ram_cell[   40703] = 32'h62072be3;
    ram_cell[   40704] = 32'head38549;
    ram_cell[   40705] = 32'h3627a57c;
    ram_cell[   40706] = 32'h24de646d;
    ram_cell[   40707] = 32'haf6d2f03;
    ram_cell[   40708] = 32'h2aa842ba;
    ram_cell[   40709] = 32'h9297b629;
    ram_cell[   40710] = 32'hf0be05fd;
    ram_cell[   40711] = 32'h762f8a3f;
    ram_cell[   40712] = 32'h8e1e860b;
    ram_cell[   40713] = 32'h615cc22e;
    ram_cell[   40714] = 32'h41886061;
    ram_cell[   40715] = 32'h7e0d93fd;
    ram_cell[   40716] = 32'h3c37c5ce;
    ram_cell[   40717] = 32'ha70f26eb;
    ram_cell[   40718] = 32'h1460f9b6;
    ram_cell[   40719] = 32'hb78f66b2;
    ram_cell[   40720] = 32'hc333b948;
    ram_cell[   40721] = 32'hddea2c25;
    ram_cell[   40722] = 32'haa1096f2;
    ram_cell[   40723] = 32'h2f4b53c3;
    ram_cell[   40724] = 32'h6e827f0e;
    ram_cell[   40725] = 32'hac4cadd3;
    ram_cell[   40726] = 32'h0d58bf05;
    ram_cell[   40727] = 32'hdefdbbd4;
    ram_cell[   40728] = 32'h723ebd2c;
    ram_cell[   40729] = 32'hfbcaf8f8;
    ram_cell[   40730] = 32'hc294e479;
    ram_cell[   40731] = 32'ha80e78b8;
    ram_cell[   40732] = 32'h5ee9cab0;
    ram_cell[   40733] = 32'h5841e10a;
    ram_cell[   40734] = 32'h0b703337;
    ram_cell[   40735] = 32'h5d45d208;
    ram_cell[   40736] = 32'hbb3efb81;
    ram_cell[   40737] = 32'h3f3848b5;
    ram_cell[   40738] = 32'hd299f98e;
    ram_cell[   40739] = 32'hbb33ffc9;
    ram_cell[   40740] = 32'h0ff46570;
    ram_cell[   40741] = 32'h654dff7e;
    ram_cell[   40742] = 32'hb5ae2b2a;
    ram_cell[   40743] = 32'h9733a834;
    ram_cell[   40744] = 32'h5145372f;
    ram_cell[   40745] = 32'h05620d9b;
    ram_cell[   40746] = 32'h6ce07716;
    ram_cell[   40747] = 32'h1b36a9f4;
    ram_cell[   40748] = 32'hdfb2787f;
    ram_cell[   40749] = 32'h13d5b516;
    ram_cell[   40750] = 32'hffe00be3;
    ram_cell[   40751] = 32'h27dab426;
    ram_cell[   40752] = 32'h4ef89efa;
    ram_cell[   40753] = 32'ha851e7e3;
    ram_cell[   40754] = 32'heb52ad00;
    ram_cell[   40755] = 32'h4063ff9c;
    ram_cell[   40756] = 32'h90cf1049;
    ram_cell[   40757] = 32'h5dd1eb52;
    ram_cell[   40758] = 32'h8c290530;
    ram_cell[   40759] = 32'h2b3ec1f1;
    ram_cell[   40760] = 32'h26656b78;
    ram_cell[   40761] = 32'hb45835ad;
    ram_cell[   40762] = 32'h219ea74e;
    ram_cell[   40763] = 32'h5204c8ff;
    ram_cell[   40764] = 32'hd1056309;
    ram_cell[   40765] = 32'h240092e0;
    ram_cell[   40766] = 32'h123d38d9;
    ram_cell[   40767] = 32'h73c331b4;
    ram_cell[   40768] = 32'hb05bb3c2;
    ram_cell[   40769] = 32'haa785cf2;
    ram_cell[   40770] = 32'ha25df120;
    ram_cell[   40771] = 32'hde5edec5;
    ram_cell[   40772] = 32'hd08b4d0c;
    ram_cell[   40773] = 32'hc593c1f1;
    ram_cell[   40774] = 32'hb67f43a8;
    ram_cell[   40775] = 32'ha331894a;
    ram_cell[   40776] = 32'h5c671ba0;
    ram_cell[   40777] = 32'h5b0bce05;
    ram_cell[   40778] = 32'h2b1ef455;
    ram_cell[   40779] = 32'h58bbf188;
    ram_cell[   40780] = 32'h05aca1cb;
    ram_cell[   40781] = 32'h4cd83d5f;
    ram_cell[   40782] = 32'h0c68315d;
    ram_cell[   40783] = 32'hb0d40332;
    ram_cell[   40784] = 32'hd348f978;
    ram_cell[   40785] = 32'h16446d7a;
    ram_cell[   40786] = 32'h59b9bf7e;
    ram_cell[   40787] = 32'h7409c43b;
    ram_cell[   40788] = 32'hc2087489;
    ram_cell[   40789] = 32'hd6b46290;
    ram_cell[   40790] = 32'h98b00dc6;
    ram_cell[   40791] = 32'h907c2d05;
    ram_cell[   40792] = 32'h5d27cf75;
    ram_cell[   40793] = 32'hca66f22e;
    ram_cell[   40794] = 32'h20b42af4;
    ram_cell[   40795] = 32'hd36d0e2c;
    ram_cell[   40796] = 32'ha2ed5093;
    ram_cell[   40797] = 32'h6741b0b0;
    ram_cell[   40798] = 32'h99496fba;
    ram_cell[   40799] = 32'h4b6e06de;
    ram_cell[   40800] = 32'h1954ce19;
    ram_cell[   40801] = 32'hb021dcd0;
    ram_cell[   40802] = 32'hffc5b0c2;
    ram_cell[   40803] = 32'h8a4490dd;
    ram_cell[   40804] = 32'hf5e69f63;
    ram_cell[   40805] = 32'h8ca20e4d;
    ram_cell[   40806] = 32'h577c6ffa;
    ram_cell[   40807] = 32'h63844888;
    ram_cell[   40808] = 32'h1263b233;
    ram_cell[   40809] = 32'hed344db9;
    ram_cell[   40810] = 32'hc6ad522b;
    ram_cell[   40811] = 32'h3b9457f3;
    ram_cell[   40812] = 32'h13c6deae;
    ram_cell[   40813] = 32'he28e4ade;
    ram_cell[   40814] = 32'hc42df414;
    ram_cell[   40815] = 32'h4400dcf7;
    ram_cell[   40816] = 32'ha31fd5fd;
    ram_cell[   40817] = 32'hcbe64090;
    ram_cell[   40818] = 32'h18d24b1a;
    ram_cell[   40819] = 32'hac9fdfc1;
    ram_cell[   40820] = 32'hbb911d89;
    ram_cell[   40821] = 32'hd19ab0d4;
    ram_cell[   40822] = 32'he239a584;
    ram_cell[   40823] = 32'h1eb4f1f9;
    ram_cell[   40824] = 32'h2640beeb;
    ram_cell[   40825] = 32'hfe54de6a;
    ram_cell[   40826] = 32'hf1cb7410;
    ram_cell[   40827] = 32'h100128d0;
    ram_cell[   40828] = 32'he92fb605;
    ram_cell[   40829] = 32'ha582ac34;
    ram_cell[   40830] = 32'hc2172e99;
    ram_cell[   40831] = 32'hb296fbf8;
    ram_cell[   40832] = 32'hf5f91963;
    ram_cell[   40833] = 32'h5dca9af4;
    ram_cell[   40834] = 32'heca7b276;
    ram_cell[   40835] = 32'h2f10a124;
    ram_cell[   40836] = 32'hd3e0edae;
    ram_cell[   40837] = 32'hfccb1803;
    ram_cell[   40838] = 32'h9624b1d7;
    ram_cell[   40839] = 32'h07503387;
    ram_cell[   40840] = 32'h4ab9f3bf;
    ram_cell[   40841] = 32'he9c2cb3d;
    ram_cell[   40842] = 32'hdf0fd404;
    ram_cell[   40843] = 32'h53e5246b;
    ram_cell[   40844] = 32'hb90f31f8;
    ram_cell[   40845] = 32'h394e5475;
    ram_cell[   40846] = 32'hf9fa9745;
    ram_cell[   40847] = 32'h4ada4518;
    ram_cell[   40848] = 32'h773952ff;
    ram_cell[   40849] = 32'h32c426fe;
    ram_cell[   40850] = 32'hdc113606;
    ram_cell[   40851] = 32'hf5447406;
    ram_cell[   40852] = 32'h75787c18;
    ram_cell[   40853] = 32'h2f00d1c2;
    ram_cell[   40854] = 32'h2400cee0;
    ram_cell[   40855] = 32'h18fcfa76;
    ram_cell[   40856] = 32'h35cb6f58;
    ram_cell[   40857] = 32'he7df72b1;
    ram_cell[   40858] = 32'h9349c6d6;
    ram_cell[   40859] = 32'h75aab5b5;
    ram_cell[   40860] = 32'h9e64b6c6;
    ram_cell[   40861] = 32'h4a6742c2;
    ram_cell[   40862] = 32'h89362c31;
    ram_cell[   40863] = 32'h1b0ea55c;
    ram_cell[   40864] = 32'h1bb6626f;
    ram_cell[   40865] = 32'h808aa275;
    ram_cell[   40866] = 32'hded8ecbc;
    ram_cell[   40867] = 32'heb1a5ba5;
    ram_cell[   40868] = 32'h0bd7e109;
    ram_cell[   40869] = 32'hf29267e5;
    ram_cell[   40870] = 32'h948db73c;
    ram_cell[   40871] = 32'hc5f152b2;
    ram_cell[   40872] = 32'h7d6907eb;
    ram_cell[   40873] = 32'h7c63665d;
    ram_cell[   40874] = 32'hbea669bf;
    ram_cell[   40875] = 32'he7d2529f;
    ram_cell[   40876] = 32'h34e17223;
    ram_cell[   40877] = 32'h64f5a698;
    ram_cell[   40878] = 32'h2d5bac6a;
    ram_cell[   40879] = 32'h347a1156;
    ram_cell[   40880] = 32'h59ecaeef;
    ram_cell[   40881] = 32'h7731746b;
    ram_cell[   40882] = 32'hd2e12e74;
    ram_cell[   40883] = 32'haa1da220;
    ram_cell[   40884] = 32'hd31d8a62;
    ram_cell[   40885] = 32'h72881a07;
    ram_cell[   40886] = 32'h547a727e;
    ram_cell[   40887] = 32'h2e0380bf;
    ram_cell[   40888] = 32'h225e4209;
    ram_cell[   40889] = 32'hd1f5bcb3;
    ram_cell[   40890] = 32'h25655bbe;
    ram_cell[   40891] = 32'hdcf18feb;
    ram_cell[   40892] = 32'h1cecabd7;
    ram_cell[   40893] = 32'ha46e1ff5;
    ram_cell[   40894] = 32'h896513a5;
    ram_cell[   40895] = 32'h20ec8492;
    ram_cell[   40896] = 32'hfb52ec71;
    ram_cell[   40897] = 32'h02f7e880;
    ram_cell[   40898] = 32'h98051bee;
    ram_cell[   40899] = 32'h671ac1ae;
    ram_cell[   40900] = 32'h6152ca2a;
    ram_cell[   40901] = 32'h634e7dc3;
    ram_cell[   40902] = 32'h21e4347e;
    ram_cell[   40903] = 32'h3747cec8;
    ram_cell[   40904] = 32'h38e6e89e;
    ram_cell[   40905] = 32'h84d36d24;
    ram_cell[   40906] = 32'h17d9502c;
    ram_cell[   40907] = 32'h47ab767f;
    ram_cell[   40908] = 32'h84d067af;
    ram_cell[   40909] = 32'hd4d22d6c;
    ram_cell[   40910] = 32'h7b7f328c;
    ram_cell[   40911] = 32'h34f79278;
    ram_cell[   40912] = 32'h0e505e99;
    ram_cell[   40913] = 32'h25db9b65;
    ram_cell[   40914] = 32'hee1248b7;
    ram_cell[   40915] = 32'hea0068c8;
    ram_cell[   40916] = 32'hf1bf110b;
    ram_cell[   40917] = 32'h5f7aab0b;
    ram_cell[   40918] = 32'h7ead1581;
    ram_cell[   40919] = 32'hc68c5614;
    ram_cell[   40920] = 32'hbf705f8c;
    ram_cell[   40921] = 32'h5b14281d;
    ram_cell[   40922] = 32'h5d7da47c;
    ram_cell[   40923] = 32'h6f70df22;
    ram_cell[   40924] = 32'h44518824;
    ram_cell[   40925] = 32'h551aa5bc;
    ram_cell[   40926] = 32'haa206bac;
    ram_cell[   40927] = 32'hf2920b13;
    ram_cell[   40928] = 32'h01fe51c6;
    ram_cell[   40929] = 32'h26f4c41a;
    ram_cell[   40930] = 32'hae1473d5;
    ram_cell[   40931] = 32'h6d8fe794;
    ram_cell[   40932] = 32'hac9fc6a5;
    ram_cell[   40933] = 32'h2d861260;
    ram_cell[   40934] = 32'h2a3d9f3e;
    ram_cell[   40935] = 32'hc8778f71;
    ram_cell[   40936] = 32'h7cf89408;
    ram_cell[   40937] = 32'h99d414f9;
    ram_cell[   40938] = 32'hcd3f6207;
    ram_cell[   40939] = 32'ha82374c4;
    ram_cell[   40940] = 32'hc983ea97;
    ram_cell[   40941] = 32'h2e3e3a17;
    ram_cell[   40942] = 32'h9f2a75af;
    ram_cell[   40943] = 32'h2664fa53;
    ram_cell[   40944] = 32'h2aa19b23;
    ram_cell[   40945] = 32'h1e3a0edd;
    ram_cell[   40946] = 32'hdab9e17f;
    ram_cell[   40947] = 32'h3751376f;
    ram_cell[   40948] = 32'he216a793;
    ram_cell[   40949] = 32'h650c039e;
    ram_cell[   40950] = 32'hdefbd153;
    ram_cell[   40951] = 32'h0d3072b4;
    ram_cell[   40952] = 32'h62e0ce69;
    ram_cell[   40953] = 32'h70654910;
    ram_cell[   40954] = 32'hf7c0f5ee;
    ram_cell[   40955] = 32'h5e87c5de;
    ram_cell[   40956] = 32'h09fb62ed;
    ram_cell[   40957] = 32'hab921aa0;
    ram_cell[   40958] = 32'h5da5233b;
    ram_cell[   40959] = 32'h980b9d9e;
    ram_cell[   40960] = 32'h17314533;
    ram_cell[   40961] = 32'h3b848893;
    ram_cell[   40962] = 32'hf4e156b5;
    ram_cell[   40963] = 32'hed9ca396;
    ram_cell[   40964] = 32'h8faf23bf;
    ram_cell[   40965] = 32'ha2290daf;
    ram_cell[   40966] = 32'he92bad7a;
    ram_cell[   40967] = 32'h233b55fb;
    ram_cell[   40968] = 32'h72531e23;
    ram_cell[   40969] = 32'hcbe03620;
    ram_cell[   40970] = 32'h76ce43b2;
    ram_cell[   40971] = 32'h78d7247a;
    ram_cell[   40972] = 32'h23a8ad87;
    ram_cell[   40973] = 32'h27ee23cd;
    ram_cell[   40974] = 32'h162515e4;
    ram_cell[   40975] = 32'h935b9990;
    ram_cell[   40976] = 32'he2497801;
    ram_cell[   40977] = 32'ha324127a;
    ram_cell[   40978] = 32'h9153a9e1;
    ram_cell[   40979] = 32'h75143bb2;
    ram_cell[   40980] = 32'h2dbac318;
    ram_cell[   40981] = 32'h0bf4f0eb;
    ram_cell[   40982] = 32'h599bf7dd;
    ram_cell[   40983] = 32'hddf6f61b;
    ram_cell[   40984] = 32'h7f02b656;
    ram_cell[   40985] = 32'h839581d4;
    ram_cell[   40986] = 32'h0cfc751b;
    ram_cell[   40987] = 32'h075f6dc7;
    ram_cell[   40988] = 32'he1a3f69e;
    ram_cell[   40989] = 32'h2713d295;
    ram_cell[   40990] = 32'hef993299;
    ram_cell[   40991] = 32'h5d990e42;
    ram_cell[   40992] = 32'hfd2490bd;
    ram_cell[   40993] = 32'h2aa584aa;
    ram_cell[   40994] = 32'haa8307f6;
    ram_cell[   40995] = 32'h65e5f686;
    ram_cell[   40996] = 32'h2c892c24;
    ram_cell[   40997] = 32'hafdea191;
    ram_cell[   40998] = 32'ha430757b;
    ram_cell[   40999] = 32'h2340cbb1;
    ram_cell[   41000] = 32'h1069d063;
    ram_cell[   41001] = 32'hb34ee607;
    ram_cell[   41002] = 32'h31f20297;
    ram_cell[   41003] = 32'h7c3ea38a;
    ram_cell[   41004] = 32'hb29d9b62;
    ram_cell[   41005] = 32'h68bdb524;
    ram_cell[   41006] = 32'h377e6738;
    ram_cell[   41007] = 32'h1c58f9b3;
    ram_cell[   41008] = 32'h8240d941;
    ram_cell[   41009] = 32'he3088634;
    ram_cell[   41010] = 32'he7f19d8b;
    ram_cell[   41011] = 32'hc0bde897;
    ram_cell[   41012] = 32'h23b70290;
    ram_cell[   41013] = 32'h99d9805c;
    ram_cell[   41014] = 32'h75e52db2;
    ram_cell[   41015] = 32'h13faaa7b;
    ram_cell[   41016] = 32'h521034ca;
    ram_cell[   41017] = 32'h072213da;
    ram_cell[   41018] = 32'h20eb5f1c;
    ram_cell[   41019] = 32'h69979af2;
    ram_cell[   41020] = 32'h23319f64;
    ram_cell[   41021] = 32'h004b4d1a;
    ram_cell[   41022] = 32'h24888d52;
    ram_cell[   41023] = 32'h93fd24fa;
    ram_cell[   41024] = 32'hf0dc6f74;
    ram_cell[   41025] = 32'h12627cc7;
    ram_cell[   41026] = 32'h67ca2ca9;
    ram_cell[   41027] = 32'hc7f81bbf;
    ram_cell[   41028] = 32'hba2cf6f8;
    ram_cell[   41029] = 32'h583e68ae;
    ram_cell[   41030] = 32'h19d3158b;
    ram_cell[   41031] = 32'hc6264ba6;
    ram_cell[   41032] = 32'h8ff4d0be;
    ram_cell[   41033] = 32'hc05ca1b0;
    ram_cell[   41034] = 32'ha7565899;
    ram_cell[   41035] = 32'hd1be7828;
    ram_cell[   41036] = 32'hccfab920;
    ram_cell[   41037] = 32'h794de1f7;
    ram_cell[   41038] = 32'h006e8849;
    ram_cell[   41039] = 32'h054d3859;
    ram_cell[   41040] = 32'he4100b2d;
    ram_cell[   41041] = 32'h39ed60ee;
    ram_cell[   41042] = 32'he8b59d71;
    ram_cell[   41043] = 32'h3ff1e8ae;
    ram_cell[   41044] = 32'hfa617df2;
    ram_cell[   41045] = 32'h3addded3;
    ram_cell[   41046] = 32'h278e3141;
    ram_cell[   41047] = 32'hf79d4c8a;
    ram_cell[   41048] = 32'h65d67ab6;
    ram_cell[   41049] = 32'he72bd284;
    ram_cell[   41050] = 32'h5c7a5898;
    ram_cell[   41051] = 32'h5d168b42;
    ram_cell[   41052] = 32'he800c3ff;
    ram_cell[   41053] = 32'h4f8c52a0;
    ram_cell[   41054] = 32'hc5d0032f;
    ram_cell[   41055] = 32'hf0fe5a77;
    ram_cell[   41056] = 32'h9951c650;
    ram_cell[   41057] = 32'h2e2e91ac;
    ram_cell[   41058] = 32'h0a979f34;
    ram_cell[   41059] = 32'hca3b8771;
    ram_cell[   41060] = 32'hf721882b;
    ram_cell[   41061] = 32'h6be28282;
    ram_cell[   41062] = 32'hb2e3279a;
    ram_cell[   41063] = 32'hbf52cf14;
    ram_cell[   41064] = 32'ha6bb9d2b;
    ram_cell[   41065] = 32'h88173312;
    ram_cell[   41066] = 32'h64f85f9e;
    ram_cell[   41067] = 32'hfc84c815;
    ram_cell[   41068] = 32'h714167cc;
    ram_cell[   41069] = 32'h85cc8a2c;
    ram_cell[   41070] = 32'hf603f4cb;
    ram_cell[   41071] = 32'hd74ae731;
    ram_cell[   41072] = 32'h8b0879fd;
    ram_cell[   41073] = 32'hc553dee3;
    ram_cell[   41074] = 32'hf600db7c;
    ram_cell[   41075] = 32'h56e60924;
    ram_cell[   41076] = 32'hbd6806ef;
    ram_cell[   41077] = 32'h3340e6c7;
    ram_cell[   41078] = 32'h3c55039b;
    ram_cell[   41079] = 32'hbf637021;
    ram_cell[   41080] = 32'h00311bc5;
    ram_cell[   41081] = 32'h69ed6bfc;
    ram_cell[   41082] = 32'h162ce35e;
    ram_cell[   41083] = 32'h2012b355;
    ram_cell[   41084] = 32'h3ae5f179;
    ram_cell[   41085] = 32'h89aa2667;
    ram_cell[   41086] = 32'hd1d3ec19;
    ram_cell[   41087] = 32'ha69244a4;
    ram_cell[   41088] = 32'h89ea4679;
    ram_cell[   41089] = 32'h84517af2;
    ram_cell[   41090] = 32'h59d9a95f;
    ram_cell[   41091] = 32'h8a44a860;
    ram_cell[   41092] = 32'h923898f0;
    ram_cell[   41093] = 32'hcbfddb3f;
    ram_cell[   41094] = 32'h66e5730a;
    ram_cell[   41095] = 32'h8237571c;
    ram_cell[   41096] = 32'hf80afe65;
    ram_cell[   41097] = 32'h9e4fac9c;
    ram_cell[   41098] = 32'ha965f2f7;
    ram_cell[   41099] = 32'hddb2f934;
    ram_cell[   41100] = 32'h25579f00;
    ram_cell[   41101] = 32'h37d02399;
    ram_cell[   41102] = 32'he176a3be;
    ram_cell[   41103] = 32'h5ac1034e;
    ram_cell[   41104] = 32'h70c532fd;
    ram_cell[   41105] = 32'h5b8da755;
    ram_cell[   41106] = 32'ha0b8b13f;
    ram_cell[   41107] = 32'h6e453155;
    ram_cell[   41108] = 32'h41da2b20;
    ram_cell[   41109] = 32'h3653a652;
    ram_cell[   41110] = 32'hb0a04bab;
    ram_cell[   41111] = 32'h007f3238;
    ram_cell[   41112] = 32'hdd7f38c6;
    ram_cell[   41113] = 32'hab3b498b;
    ram_cell[   41114] = 32'h3c4bdd2e;
    ram_cell[   41115] = 32'hf13c402a;
    ram_cell[   41116] = 32'h85fa6387;
    ram_cell[   41117] = 32'heee3d5f1;
    ram_cell[   41118] = 32'h6fa6f6e9;
    ram_cell[   41119] = 32'hd4e1c660;
    ram_cell[   41120] = 32'hbc3a8af1;
    ram_cell[   41121] = 32'h74c064e3;
    ram_cell[   41122] = 32'h302e34d9;
    ram_cell[   41123] = 32'h5c45e65b;
    ram_cell[   41124] = 32'hb3f2d2bb;
    ram_cell[   41125] = 32'hdf0a3fca;
    ram_cell[   41126] = 32'h89b89342;
    ram_cell[   41127] = 32'h8bc900d8;
    ram_cell[   41128] = 32'h06119c4d;
    ram_cell[   41129] = 32'h9e7b71e5;
    ram_cell[   41130] = 32'he66f7aa0;
    ram_cell[   41131] = 32'h0daefdc4;
    ram_cell[   41132] = 32'h5d3081bb;
    ram_cell[   41133] = 32'hb14e0ee2;
    ram_cell[   41134] = 32'h309b7d3a;
    ram_cell[   41135] = 32'h84706189;
    ram_cell[   41136] = 32'h3743cabf;
    ram_cell[   41137] = 32'h64b04902;
    ram_cell[   41138] = 32'hab46e332;
    ram_cell[   41139] = 32'haa507c71;
    ram_cell[   41140] = 32'h9d7e1ce1;
    ram_cell[   41141] = 32'hebf91b32;
    ram_cell[   41142] = 32'h5ab42790;
    ram_cell[   41143] = 32'ha0592ea6;
    ram_cell[   41144] = 32'h585096de;
    ram_cell[   41145] = 32'h6f381206;
    ram_cell[   41146] = 32'hc82e56a0;
    ram_cell[   41147] = 32'hcd490838;
    ram_cell[   41148] = 32'h457943c0;
    ram_cell[   41149] = 32'h0830f6c3;
    ram_cell[   41150] = 32'h406aea2a;
    ram_cell[   41151] = 32'h53eb2b76;
    ram_cell[   41152] = 32'h6f16efe9;
    ram_cell[   41153] = 32'hae397ca3;
    ram_cell[   41154] = 32'h0d44f43b;
    ram_cell[   41155] = 32'h4774d86d;
    ram_cell[   41156] = 32'hb1dcaff8;
    ram_cell[   41157] = 32'h92107158;
    ram_cell[   41158] = 32'hb57860fa;
    ram_cell[   41159] = 32'he0b2857a;
    ram_cell[   41160] = 32'h8b6eb7db;
    ram_cell[   41161] = 32'hbc1362ff;
    ram_cell[   41162] = 32'h64b321a1;
    ram_cell[   41163] = 32'hd2f5678e;
    ram_cell[   41164] = 32'hf6481999;
    ram_cell[   41165] = 32'h047ab06b;
    ram_cell[   41166] = 32'h96b6e315;
    ram_cell[   41167] = 32'hfa030630;
    ram_cell[   41168] = 32'h1bf424ba;
    ram_cell[   41169] = 32'h924adc8a;
    ram_cell[   41170] = 32'h4571831c;
    ram_cell[   41171] = 32'hff221f29;
    ram_cell[   41172] = 32'hb7cf13c8;
    ram_cell[   41173] = 32'h8762104e;
    ram_cell[   41174] = 32'h76e73eff;
    ram_cell[   41175] = 32'h6c5c0053;
    ram_cell[   41176] = 32'hdc0caf5b;
    ram_cell[   41177] = 32'h9f8f2828;
    ram_cell[   41178] = 32'hd72ed034;
    ram_cell[   41179] = 32'hfc690c13;
    ram_cell[   41180] = 32'hae997751;
    ram_cell[   41181] = 32'h8fffe8ef;
    ram_cell[   41182] = 32'hd79cc7dd;
    ram_cell[   41183] = 32'h2a5afe56;
    ram_cell[   41184] = 32'h2683eb54;
    ram_cell[   41185] = 32'he0ba22b7;
    ram_cell[   41186] = 32'hb97a3aa6;
    ram_cell[   41187] = 32'h87335d32;
    ram_cell[   41188] = 32'h31adb7d3;
    ram_cell[   41189] = 32'hf1a45895;
    ram_cell[   41190] = 32'hede98b2f;
    ram_cell[   41191] = 32'hd916b0ee;
    ram_cell[   41192] = 32'h004ab82f;
    ram_cell[   41193] = 32'hd880b65e;
    ram_cell[   41194] = 32'had18f5f9;
    ram_cell[   41195] = 32'h511d7bb9;
    ram_cell[   41196] = 32'hfd683b92;
    ram_cell[   41197] = 32'h85b29998;
    ram_cell[   41198] = 32'h538c9062;
    ram_cell[   41199] = 32'h54478af1;
    ram_cell[   41200] = 32'h1806a75b;
    ram_cell[   41201] = 32'h92217003;
    ram_cell[   41202] = 32'hc7d456b0;
    ram_cell[   41203] = 32'h7e3c8d59;
    ram_cell[   41204] = 32'hf64534c3;
    ram_cell[   41205] = 32'hbd4cf819;
    ram_cell[   41206] = 32'hd50ff129;
    ram_cell[   41207] = 32'h52b3d63e;
    ram_cell[   41208] = 32'hbd1ab27f;
    ram_cell[   41209] = 32'h557c6069;
    ram_cell[   41210] = 32'h88c72120;
    ram_cell[   41211] = 32'h1f70690f;
    ram_cell[   41212] = 32'h9f4d06ad;
    ram_cell[   41213] = 32'h4a25f046;
    ram_cell[   41214] = 32'hed8d6208;
    ram_cell[   41215] = 32'h94f0d466;
    ram_cell[   41216] = 32'h6d147d56;
    ram_cell[   41217] = 32'hf1d20e08;
    ram_cell[   41218] = 32'h1ce0c80b;
    ram_cell[   41219] = 32'hc11b9044;
    ram_cell[   41220] = 32'h7a5eafce;
    ram_cell[   41221] = 32'hb2856a77;
    ram_cell[   41222] = 32'h3799c604;
    ram_cell[   41223] = 32'h08ce94c7;
    ram_cell[   41224] = 32'h4fc8d600;
    ram_cell[   41225] = 32'hb2351d28;
    ram_cell[   41226] = 32'he8fb90c4;
    ram_cell[   41227] = 32'hc329fd94;
    ram_cell[   41228] = 32'h6b4853ed;
    ram_cell[   41229] = 32'hf7cc201c;
    ram_cell[   41230] = 32'ha8350366;
    ram_cell[   41231] = 32'h5303822e;
    ram_cell[   41232] = 32'h451643a3;
    ram_cell[   41233] = 32'he7529f30;
    ram_cell[   41234] = 32'h72adbe28;
    ram_cell[   41235] = 32'h3e0cefba;
    ram_cell[   41236] = 32'h36f3c6f5;
    ram_cell[   41237] = 32'h0aae1a57;
    ram_cell[   41238] = 32'hfba13799;
    ram_cell[   41239] = 32'h070cb018;
    ram_cell[   41240] = 32'hb9c66991;
    ram_cell[   41241] = 32'h13b2c4b2;
    ram_cell[   41242] = 32'h0f815ef1;
    ram_cell[   41243] = 32'h0ff463ce;
    ram_cell[   41244] = 32'h0404d988;
    ram_cell[   41245] = 32'h01f3ff7b;
    ram_cell[   41246] = 32'h70b09032;
    ram_cell[   41247] = 32'h1ee06c38;
    ram_cell[   41248] = 32'h16b3b9a2;
    ram_cell[   41249] = 32'h0d2b5ab5;
    ram_cell[   41250] = 32'h82f03d6c;
    ram_cell[   41251] = 32'h6de779ff;
    ram_cell[   41252] = 32'h2b10d105;
    ram_cell[   41253] = 32'h2d7c5ab4;
    ram_cell[   41254] = 32'h9cc34c47;
    ram_cell[   41255] = 32'h68214033;
    ram_cell[   41256] = 32'h7f46884f;
    ram_cell[   41257] = 32'ha77b6559;
    ram_cell[   41258] = 32'hceafad09;
    ram_cell[   41259] = 32'h21c92f56;
    ram_cell[   41260] = 32'h0e4b3204;
    ram_cell[   41261] = 32'h298e59af;
    ram_cell[   41262] = 32'hbec8095d;
    ram_cell[   41263] = 32'h1cc22941;
    ram_cell[   41264] = 32'h47440030;
    ram_cell[   41265] = 32'h8edec60b;
    ram_cell[   41266] = 32'h888321c3;
    ram_cell[   41267] = 32'hd9254951;
    ram_cell[   41268] = 32'hddbd6a74;
    ram_cell[   41269] = 32'hf37d86a2;
    ram_cell[   41270] = 32'h52a89b0a;
    ram_cell[   41271] = 32'h2fd7f1a3;
    ram_cell[   41272] = 32'h59ba1dd4;
    ram_cell[   41273] = 32'h52bdba37;
    ram_cell[   41274] = 32'h878c4b78;
    ram_cell[   41275] = 32'hd58e381f;
    ram_cell[   41276] = 32'h613273ce;
    ram_cell[   41277] = 32'h7726311e;
    ram_cell[   41278] = 32'h301766f0;
    ram_cell[   41279] = 32'h2b03cd26;
    ram_cell[   41280] = 32'ha31cb9c4;
    ram_cell[   41281] = 32'h87ab0edd;
    ram_cell[   41282] = 32'h1241a18b;
    ram_cell[   41283] = 32'h53a118c1;
    ram_cell[   41284] = 32'hbe2e9437;
    ram_cell[   41285] = 32'h4f661584;
    ram_cell[   41286] = 32'h5ff7ac23;
    ram_cell[   41287] = 32'h515fef8a;
    ram_cell[   41288] = 32'h88e462c9;
    ram_cell[   41289] = 32'hf3b44915;
    ram_cell[   41290] = 32'hbd5c3ebd;
    ram_cell[   41291] = 32'h96d0d208;
    ram_cell[   41292] = 32'h160809fe;
    ram_cell[   41293] = 32'h6dc5ecca;
    ram_cell[   41294] = 32'h22bdc519;
    ram_cell[   41295] = 32'h2bacca7e;
    ram_cell[   41296] = 32'h1c2b8516;
    ram_cell[   41297] = 32'he36f5a07;
    ram_cell[   41298] = 32'he9c214a2;
    ram_cell[   41299] = 32'ha50573ba;
    ram_cell[   41300] = 32'h625c90d8;
    ram_cell[   41301] = 32'ha5da6cba;
    ram_cell[   41302] = 32'hd962eac4;
    ram_cell[   41303] = 32'haa3ead09;
    ram_cell[   41304] = 32'h8b947cef;
    ram_cell[   41305] = 32'hccc8dc86;
    ram_cell[   41306] = 32'h3dcb77f3;
    ram_cell[   41307] = 32'h31e8bea4;
    ram_cell[   41308] = 32'hc99435f9;
    ram_cell[   41309] = 32'h0ecd694b;
    ram_cell[   41310] = 32'hb33aae41;
    ram_cell[   41311] = 32'hf2720a62;
    ram_cell[   41312] = 32'h1fcd27e7;
    ram_cell[   41313] = 32'h0b84a52f;
    ram_cell[   41314] = 32'h1153271a;
    ram_cell[   41315] = 32'ha2934068;
    ram_cell[   41316] = 32'hd864bc5e;
    ram_cell[   41317] = 32'h5c706b2a;
    ram_cell[   41318] = 32'hce71092f;
    ram_cell[   41319] = 32'hd2835628;
    ram_cell[   41320] = 32'h69acc853;
    ram_cell[   41321] = 32'hf3ed37d3;
    ram_cell[   41322] = 32'h7f5fdb38;
    ram_cell[   41323] = 32'hbd97e9eb;
    ram_cell[   41324] = 32'h5bc74471;
    ram_cell[   41325] = 32'h8f89a0f3;
    ram_cell[   41326] = 32'h0cc64f9f;
    ram_cell[   41327] = 32'h5ba6dffd;
    ram_cell[   41328] = 32'ha398acd9;
    ram_cell[   41329] = 32'hbee92ea0;
    ram_cell[   41330] = 32'hde888cfa;
    ram_cell[   41331] = 32'h577de1a9;
    ram_cell[   41332] = 32'h8525d8b1;
    ram_cell[   41333] = 32'hf7670013;
    ram_cell[   41334] = 32'h0ac4ea7c;
    ram_cell[   41335] = 32'h07e2fe44;
    ram_cell[   41336] = 32'h6628644d;
    ram_cell[   41337] = 32'h838631d3;
    ram_cell[   41338] = 32'hb0288605;
    ram_cell[   41339] = 32'h2bea4948;
    ram_cell[   41340] = 32'h394cf07e;
    ram_cell[   41341] = 32'h8a83cd0e;
    ram_cell[   41342] = 32'h5d5fb763;
    ram_cell[   41343] = 32'h8294e7e5;
    ram_cell[   41344] = 32'hd02c0fb4;
    ram_cell[   41345] = 32'h4dc1b256;
    ram_cell[   41346] = 32'ha3225948;
    ram_cell[   41347] = 32'hc6566b58;
    ram_cell[   41348] = 32'hba705e33;
    ram_cell[   41349] = 32'h9a8030a3;
    ram_cell[   41350] = 32'h79cfb4d2;
    ram_cell[   41351] = 32'hb29a247a;
    ram_cell[   41352] = 32'h8253d1a5;
    ram_cell[   41353] = 32'h4e5c519c;
    ram_cell[   41354] = 32'hd670ff6e;
    ram_cell[   41355] = 32'he070c4b2;
    ram_cell[   41356] = 32'ha6e53d54;
    ram_cell[   41357] = 32'he5443cc9;
    ram_cell[   41358] = 32'haf3288cf;
    ram_cell[   41359] = 32'h02ba4129;
    ram_cell[   41360] = 32'ha99b5fa5;
    ram_cell[   41361] = 32'hb9994988;
    ram_cell[   41362] = 32'hab3db0ec;
    ram_cell[   41363] = 32'hcb1764f0;
    ram_cell[   41364] = 32'hf040e392;
    ram_cell[   41365] = 32'hc33a5047;
    ram_cell[   41366] = 32'h9eb1858b;
    ram_cell[   41367] = 32'h486735b9;
    ram_cell[   41368] = 32'hd2772148;
    ram_cell[   41369] = 32'h60ebfbfe;
    ram_cell[   41370] = 32'h5505d1d3;
    ram_cell[   41371] = 32'hbbc0f6b7;
    ram_cell[   41372] = 32'h2b3545c8;
    ram_cell[   41373] = 32'h055d1847;
    ram_cell[   41374] = 32'ha34aebc3;
    ram_cell[   41375] = 32'hac220208;
    ram_cell[   41376] = 32'h235b2bc3;
    ram_cell[   41377] = 32'hc1927a47;
    ram_cell[   41378] = 32'h9294294e;
    ram_cell[   41379] = 32'h1d1e1e4c;
    ram_cell[   41380] = 32'h73b1922c;
    ram_cell[   41381] = 32'h246d075c;
    ram_cell[   41382] = 32'hc805a4a2;
    ram_cell[   41383] = 32'h528b7286;
    ram_cell[   41384] = 32'h94d145ca;
    ram_cell[   41385] = 32'h70232de7;
    ram_cell[   41386] = 32'h69e87541;
    ram_cell[   41387] = 32'h918ff92c;
    ram_cell[   41388] = 32'h557f1420;
    ram_cell[   41389] = 32'ha9d43e21;
    ram_cell[   41390] = 32'hd71221b9;
    ram_cell[   41391] = 32'hfdd1c03c;
    ram_cell[   41392] = 32'h08522836;
    ram_cell[   41393] = 32'h72f75ef5;
    ram_cell[   41394] = 32'hde44664c;
    ram_cell[   41395] = 32'h9ad78dbd;
    ram_cell[   41396] = 32'h39b0d9be;
    ram_cell[   41397] = 32'h8919383a;
    ram_cell[   41398] = 32'h499fe602;
    ram_cell[   41399] = 32'h660ab8a5;
    ram_cell[   41400] = 32'h29298eab;
    ram_cell[   41401] = 32'h025706ea;
    ram_cell[   41402] = 32'hdc4ee9b1;
    ram_cell[   41403] = 32'ha957200e;
    ram_cell[   41404] = 32'h7b8c2dc1;
    ram_cell[   41405] = 32'hc3024d57;
    ram_cell[   41406] = 32'h9dbf49da;
    ram_cell[   41407] = 32'h6a69195b;
    ram_cell[   41408] = 32'h22709b8f;
    ram_cell[   41409] = 32'h9772eb61;
    ram_cell[   41410] = 32'hbb151841;
    ram_cell[   41411] = 32'h783d3cf4;
    ram_cell[   41412] = 32'h15f7a350;
    ram_cell[   41413] = 32'hcce2649f;
    ram_cell[   41414] = 32'ha35170bb;
    ram_cell[   41415] = 32'hbe789b25;
    ram_cell[   41416] = 32'h5d605d2e;
    ram_cell[   41417] = 32'ha4615436;
    ram_cell[   41418] = 32'hf62b9a99;
    ram_cell[   41419] = 32'h6c8f9af3;
    ram_cell[   41420] = 32'h137c3cee;
    ram_cell[   41421] = 32'h391deed3;
    ram_cell[   41422] = 32'h41190f76;
    ram_cell[   41423] = 32'h980538ab;
    ram_cell[   41424] = 32'haa12bfee;
    ram_cell[   41425] = 32'h16760c41;
    ram_cell[   41426] = 32'h6ee346c6;
    ram_cell[   41427] = 32'h51457e57;
    ram_cell[   41428] = 32'h4e97373c;
    ram_cell[   41429] = 32'h50bc592c;
    ram_cell[   41430] = 32'h077b56d2;
    ram_cell[   41431] = 32'hfed075ef;
    ram_cell[   41432] = 32'ha7b44315;
    ram_cell[   41433] = 32'h21cb5997;
    ram_cell[   41434] = 32'hec5f1523;
    ram_cell[   41435] = 32'hfe0ec98b;
    ram_cell[   41436] = 32'hceeada0f;
    ram_cell[   41437] = 32'h14be44c1;
    ram_cell[   41438] = 32'h102d2c97;
    ram_cell[   41439] = 32'h360edecc;
    ram_cell[   41440] = 32'h0c30bae7;
    ram_cell[   41441] = 32'h37fa92c2;
    ram_cell[   41442] = 32'h0724159c;
    ram_cell[   41443] = 32'ha9374fc9;
    ram_cell[   41444] = 32'hb677e86f;
    ram_cell[   41445] = 32'he6372413;
    ram_cell[   41446] = 32'hc2aab94a;
    ram_cell[   41447] = 32'hdf8c95ef;
    ram_cell[   41448] = 32'h868591b3;
    ram_cell[   41449] = 32'hea1043bc;
    ram_cell[   41450] = 32'h3583f4d1;
    ram_cell[   41451] = 32'h6a153c4d;
    ram_cell[   41452] = 32'h1e3fd39b;
    ram_cell[   41453] = 32'h01a24b8e;
    ram_cell[   41454] = 32'hfaf98b99;
    ram_cell[   41455] = 32'h25513c9c;
    ram_cell[   41456] = 32'h22c2c131;
    ram_cell[   41457] = 32'h096427f3;
    ram_cell[   41458] = 32'hbf45ac14;
    ram_cell[   41459] = 32'hd98c5f07;
    ram_cell[   41460] = 32'h3354155d;
    ram_cell[   41461] = 32'hb144431d;
    ram_cell[   41462] = 32'hc750855e;
    ram_cell[   41463] = 32'h512e4558;
    ram_cell[   41464] = 32'h5cb57ec0;
    ram_cell[   41465] = 32'hb9c6a718;
    ram_cell[   41466] = 32'h31fefb58;
    ram_cell[   41467] = 32'hd4922adf;
    ram_cell[   41468] = 32'h4d8fead3;
    ram_cell[   41469] = 32'h78719fe6;
    ram_cell[   41470] = 32'hc312f2f3;
    ram_cell[   41471] = 32'hffb3c67e;
    ram_cell[   41472] = 32'haa518e7f;
    ram_cell[   41473] = 32'h231e7efc;
    ram_cell[   41474] = 32'hb1513875;
    ram_cell[   41475] = 32'h62c3a962;
    ram_cell[   41476] = 32'h5e31bd4d;
    ram_cell[   41477] = 32'h7b019436;
    ram_cell[   41478] = 32'h7e009e99;
    ram_cell[   41479] = 32'h9fecb2d9;
    ram_cell[   41480] = 32'h64233cbd;
    ram_cell[   41481] = 32'h420f8203;
    ram_cell[   41482] = 32'h9539ec0f;
    ram_cell[   41483] = 32'h07f391c4;
    ram_cell[   41484] = 32'h166cd966;
    ram_cell[   41485] = 32'h5865cd6a;
    ram_cell[   41486] = 32'h3b85f9da;
    ram_cell[   41487] = 32'h3be38a9c;
    ram_cell[   41488] = 32'h1543c2a8;
    ram_cell[   41489] = 32'h7f348ccf;
    ram_cell[   41490] = 32'hd3158e37;
    ram_cell[   41491] = 32'h611e7200;
    ram_cell[   41492] = 32'h649095ed;
    ram_cell[   41493] = 32'hcba9977d;
    ram_cell[   41494] = 32'hb4e19d30;
    ram_cell[   41495] = 32'hf7715c6e;
    ram_cell[   41496] = 32'h2e376257;
    ram_cell[   41497] = 32'hb48bba22;
    ram_cell[   41498] = 32'hd618f6d1;
    ram_cell[   41499] = 32'hb32c1241;
    ram_cell[   41500] = 32'h85ea0c7d;
    ram_cell[   41501] = 32'hb1eb79b0;
    ram_cell[   41502] = 32'h3812e25b;
    ram_cell[   41503] = 32'h1353b44a;
    ram_cell[   41504] = 32'hcb72cded;
    ram_cell[   41505] = 32'h245b32a7;
    ram_cell[   41506] = 32'hb437c914;
    ram_cell[   41507] = 32'hc3680a57;
    ram_cell[   41508] = 32'h3c1da4e6;
    ram_cell[   41509] = 32'hdc13aaae;
    ram_cell[   41510] = 32'hee781585;
    ram_cell[   41511] = 32'h836abb6d;
    ram_cell[   41512] = 32'h5841dfda;
    ram_cell[   41513] = 32'h87618cc8;
    ram_cell[   41514] = 32'hed358d89;
    ram_cell[   41515] = 32'hb8859d8e;
    ram_cell[   41516] = 32'h5341d258;
    ram_cell[   41517] = 32'h847e496d;
    ram_cell[   41518] = 32'h1e3bebe7;
    ram_cell[   41519] = 32'h47a5f8a7;
    ram_cell[   41520] = 32'h00fa7d89;
    ram_cell[   41521] = 32'hf9fd0a29;
    ram_cell[   41522] = 32'hc7dc2583;
    ram_cell[   41523] = 32'h6637bc68;
    ram_cell[   41524] = 32'h824a0dbf;
    ram_cell[   41525] = 32'h644941a6;
    ram_cell[   41526] = 32'he28d58ad;
    ram_cell[   41527] = 32'haf424e33;
    ram_cell[   41528] = 32'h85b1c10e;
    ram_cell[   41529] = 32'h24a0721d;
    ram_cell[   41530] = 32'h454cef1b;
    ram_cell[   41531] = 32'he7a9ca3b;
    ram_cell[   41532] = 32'h1ebd4bab;
    ram_cell[   41533] = 32'h2a1f931b;
    ram_cell[   41534] = 32'h68135e21;
    ram_cell[   41535] = 32'h1400d7e8;
    ram_cell[   41536] = 32'hf389af67;
    ram_cell[   41537] = 32'hc7bcb2e2;
    ram_cell[   41538] = 32'h49e107c4;
    ram_cell[   41539] = 32'h4996a294;
    ram_cell[   41540] = 32'h6b9e3eea;
    ram_cell[   41541] = 32'h58ed3130;
    ram_cell[   41542] = 32'h11394844;
    ram_cell[   41543] = 32'h6ad24920;
    ram_cell[   41544] = 32'ha5d6afb0;
    ram_cell[   41545] = 32'h8cfbb7d5;
    ram_cell[   41546] = 32'h14a2713a;
    ram_cell[   41547] = 32'h5c0786d1;
    ram_cell[   41548] = 32'h39160600;
    ram_cell[   41549] = 32'h5b74a16b;
    ram_cell[   41550] = 32'h7a4e9aa6;
    ram_cell[   41551] = 32'h44b20d2d;
    ram_cell[   41552] = 32'h982fb0da;
    ram_cell[   41553] = 32'h52c0bd0f;
    ram_cell[   41554] = 32'hc8ed0fc3;
    ram_cell[   41555] = 32'hb4f7c14b;
    ram_cell[   41556] = 32'h245e0163;
    ram_cell[   41557] = 32'h74a0fa13;
    ram_cell[   41558] = 32'hda38aba4;
    ram_cell[   41559] = 32'he7dd9d91;
    ram_cell[   41560] = 32'hcfe911f4;
    ram_cell[   41561] = 32'hbc6985ba;
    ram_cell[   41562] = 32'hcccedc95;
    ram_cell[   41563] = 32'h5752506f;
    ram_cell[   41564] = 32'hc5f750f7;
    ram_cell[   41565] = 32'h70e40bcc;
    ram_cell[   41566] = 32'hf85faedf;
    ram_cell[   41567] = 32'h41584185;
    ram_cell[   41568] = 32'hd2cfcd07;
    ram_cell[   41569] = 32'hee2f12c8;
    ram_cell[   41570] = 32'hf25abba7;
    ram_cell[   41571] = 32'ha8f3ae95;
    ram_cell[   41572] = 32'h1993978b;
    ram_cell[   41573] = 32'hfc4de255;
    ram_cell[   41574] = 32'hf56f5fa2;
    ram_cell[   41575] = 32'h494f2f24;
    ram_cell[   41576] = 32'h93386fbb;
    ram_cell[   41577] = 32'hb25e6385;
    ram_cell[   41578] = 32'h44de754a;
    ram_cell[   41579] = 32'hb6c702e3;
    ram_cell[   41580] = 32'h679421fc;
    ram_cell[   41581] = 32'hbc489779;
    ram_cell[   41582] = 32'h4a01d796;
    ram_cell[   41583] = 32'hdfdbf758;
    ram_cell[   41584] = 32'hb9cfe58b;
    ram_cell[   41585] = 32'h0bb654c5;
    ram_cell[   41586] = 32'h8ee25096;
    ram_cell[   41587] = 32'hb0745447;
    ram_cell[   41588] = 32'hc8f42fac;
    ram_cell[   41589] = 32'hf124066d;
    ram_cell[   41590] = 32'h19db9cab;
    ram_cell[   41591] = 32'h5781d525;
    ram_cell[   41592] = 32'h5aab7947;
    ram_cell[   41593] = 32'h7466a80e;
    ram_cell[   41594] = 32'h65fdf032;
    ram_cell[   41595] = 32'h9d4c7d8c;
    ram_cell[   41596] = 32'hc464a463;
    ram_cell[   41597] = 32'h383e7da4;
    ram_cell[   41598] = 32'h744947c6;
    ram_cell[   41599] = 32'h6695f77b;
    ram_cell[   41600] = 32'hb00350b8;
    ram_cell[   41601] = 32'h92cb0207;
    ram_cell[   41602] = 32'h9799ae47;
    ram_cell[   41603] = 32'hf468f6b5;
    ram_cell[   41604] = 32'h551f4dc8;
    ram_cell[   41605] = 32'h957d6dd1;
    ram_cell[   41606] = 32'h2d158ff1;
    ram_cell[   41607] = 32'hfcaf298b;
    ram_cell[   41608] = 32'h77eacce9;
    ram_cell[   41609] = 32'hf0d85c6f;
    ram_cell[   41610] = 32'h69cca964;
    ram_cell[   41611] = 32'h95e1e177;
    ram_cell[   41612] = 32'h64a147a8;
    ram_cell[   41613] = 32'hf5f533b4;
    ram_cell[   41614] = 32'h38277adb;
    ram_cell[   41615] = 32'h8018e6b6;
    ram_cell[   41616] = 32'h4f64a055;
    ram_cell[   41617] = 32'he10a5e06;
    ram_cell[   41618] = 32'ha166d816;
    ram_cell[   41619] = 32'ha0ccf0a1;
    ram_cell[   41620] = 32'h514cbd8e;
    ram_cell[   41621] = 32'heae0b92c;
    ram_cell[   41622] = 32'h759c5837;
    ram_cell[   41623] = 32'h67d49f60;
    ram_cell[   41624] = 32'h878d7bd3;
    ram_cell[   41625] = 32'h23957aa6;
    ram_cell[   41626] = 32'h4e8c0b09;
    ram_cell[   41627] = 32'ha022e084;
    ram_cell[   41628] = 32'h4b382855;
    ram_cell[   41629] = 32'h12e8cede;
    ram_cell[   41630] = 32'ha1d2e848;
    ram_cell[   41631] = 32'hf4a694e4;
    ram_cell[   41632] = 32'h11e4f2aa;
    ram_cell[   41633] = 32'h3710f36f;
    ram_cell[   41634] = 32'hb01b80da;
    ram_cell[   41635] = 32'h9f845b76;
    ram_cell[   41636] = 32'h8259c031;
    ram_cell[   41637] = 32'hf9fa835f;
    ram_cell[   41638] = 32'h8dac1121;
    ram_cell[   41639] = 32'hfbf456b5;
    ram_cell[   41640] = 32'h18a4e46a;
    ram_cell[   41641] = 32'h44275418;
    ram_cell[   41642] = 32'hc8495ab7;
    ram_cell[   41643] = 32'h1c70f263;
    ram_cell[   41644] = 32'h7655ff95;
    ram_cell[   41645] = 32'h776dd56c;
    ram_cell[   41646] = 32'h94ae175a;
    ram_cell[   41647] = 32'h4eb7c269;
    ram_cell[   41648] = 32'hc5b0b985;
    ram_cell[   41649] = 32'hf45b7a6c;
    ram_cell[   41650] = 32'he9d2f509;
    ram_cell[   41651] = 32'h62515695;
    ram_cell[   41652] = 32'hb01b077a;
    ram_cell[   41653] = 32'h057eb182;
    ram_cell[   41654] = 32'h7b0199b8;
    ram_cell[   41655] = 32'h6191f6d5;
    ram_cell[   41656] = 32'h16255aa8;
    ram_cell[   41657] = 32'h4c66ed8b;
    ram_cell[   41658] = 32'hcea24626;
    ram_cell[   41659] = 32'h45ae7b16;
    ram_cell[   41660] = 32'ha2694e8f;
    ram_cell[   41661] = 32'hca3b9384;
    ram_cell[   41662] = 32'hf7642b81;
    ram_cell[   41663] = 32'h12e07173;
    ram_cell[   41664] = 32'hede7acd1;
    ram_cell[   41665] = 32'hbbc3490d;
    ram_cell[   41666] = 32'hc530c781;
    ram_cell[   41667] = 32'h58ca8af9;
    ram_cell[   41668] = 32'h42240473;
    ram_cell[   41669] = 32'h9d5ab029;
    ram_cell[   41670] = 32'h4f9cb59a;
    ram_cell[   41671] = 32'h97c0d78e;
    ram_cell[   41672] = 32'h3bd358d7;
    ram_cell[   41673] = 32'h70f1edd0;
    ram_cell[   41674] = 32'h82389b70;
    ram_cell[   41675] = 32'h96c3684e;
    ram_cell[   41676] = 32'hfacbe70d;
    ram_cell[   41677] = 32'h9352ff94;
    ram_cell[   41678] = 32'h4470c2d4;
    ram_cell[   41679] = 32'h9e43b13c;
    ram_cell[   41680] = 32'he9f83985;
    ram_cell[   41681] = 32'h11b35180;
    ram_cell[   41682] = 32'h8135cda6;
    ram_cell[   41683] = 32'h20f68c79;
    ram_cell[   41684] = 32'h44e3e400;
    ram_cell[   41685] = 32'h75f768f4;
    ram_cell[   41686] = 32'h3590b9bc;
    ram_cell[   41687] = 32'h40101ac3;
    ram_cell[   41688] = 32'h10c9fe7b;
    ram_cell[   41689] = 32'he52ee614;
    ram_cell[   41690] = 32'h5d0cd355;
    ram_cell[   41691] = 32'h4b9ed3a2;
    ram_cell[   41692] = 32'he0774b8f;
    ram_cell[   41693] = 32'hc705e728;
    ram_cell[   41694] = 32'h84479b5a;
    ram_cell[   41695] = 32'h5ea1ee2b;
    ram_cell[   41696] = 32'hcd39fe30;
    ram_cell[   41697] = 32'h965f8d99;
    ram_cell[   41698] = 32'h8c6b243a;
    ram_cell[   41699] = 32'h05e8d7d8;
    ram_cell[   41700] = 32'hc5bce1bb;
    ram_cell[   41701] = 32'hc26abfb4;
    ram_cell[   41702] = 32'hd803b466;
    ram_cell[   41703] = 32'h6b17b8ad;
    ram_cell[   41704] = 32'h9dc29074;
    ram_cell[   41705] = 32'h096c8d02;
    ram_cell[   41706] = 32'hbc1195b6;
    ram_cell[   41707] = 32'he09e195b;
    ram_cell[   41708] = 32'h0225f73a;
    ram_cell[   41709] = 32'h18bc6b5a;
    ram_cell[   41710] = 32'h061f3389;
    ram_cell[   41711] = 32'h8fa66df3;
    ram_cell[   41712] = 32'h9602e8ca;
    ram_cell[   41713] = 32'h5c3b3f2f;
    ram_cell[   41714] = 32'hf503308a;
    ram_cell[   41715] = 32'h571fa527;
    ram_cell[   41716] = 32'h077a33ee;
    ram_cell[   41717] = 32'hd1335fde;
    ram_cell[   41718] = 32'hef5e51e9;
    ram_cell[   41719] = 32'hc9d28d31;
    ram_cell[   41720] = 32'h1910cc76;
    ram_cell[   41721] = 32'he823909d;
    ram_cell[   41722] = 32'hea8d3032;
    ram_cell[   41723] = 32'h66214450;
    ram_cell[   41724] = 32'hbfadba26;
    ram_cell[   41725] = 32'h15bfc42b;
    ram_cell[   41726] = 32'h6ead02cb;
    ram_cell[   41727] = 32'heee04452;
    ram_cell[   41728] = 32'hf14b1418;
    ram_cell[   41729] = 32'h315c11da;
    ram_cell[   41730] = 32'hf6b2735f;
    ram_cell[   41731] = 32'hfb57444d;
    ram_cell[   41732] = 32'h194c2cba;
    ram_cell[   41733] = 32'h763f61a3;
    ram_cell[   41734] = 32'he4b2c7fc;
    ram_cell[   41735] = 32'h33df2b65;
    ram_cell[   41736] = 32'h179a7dc3;
    ram_cell[   41737] = 32'h630a9c16;
    ram_cell[   41738] = 32'h24057b50;
    ram_cell[   41739] = 32'h2124be2f;
    ram_cell[   41740] = 32'hfd63c4cc;
    ram_cell[   41741] = 32'h0786b555;
    ram_cell[   41742] = 32'h42892bce;
    ram_cell[   41743] = 32'h319d7d84;
    ram_cell[   41744] = 32'h3688c589;
    ram_cell[   41745] = 32'hacb4d25b;
    ram_cell[   41746] = 32'hbcb720fa;
    ram_cell[   41747] = 32'hb7baa1f6;
    ram_cell[   41748] = 32'h8b5d7d01;
    ram_cell[   41749] = 32'hdbb4dbd1;
    ram_cell[   41750] = 32'he66108a1;
    ram_cell[   41751] = 32'ha3d09094;
    ram_cell[   41752] = 32'hf38ab137;
    ram_cell[   41753] = 32'h4f9b8086;
    ram_cell[   41754] = 32'h9bb16bfb;
    ram_cell[   41755] = 32'hbeffdce5;
    ram_cell[   41756] = 32'h8a15260b;
    ram_cell[   41757] = 32'hdfa65f11;
    ram_cell[   41758] = 32'hf68208fd;
    ram_cell[   41759] = 32'h8b26fa86;
    ram_cell[   41760] = 32'h35864179;
    ram_cell[   41761] = 32'h5bf1c5a4;
    ram_cell[   41762] = 32'h053b7583;
    ram_cell[   41763] = 32'h899fcb3b;
    ram_cell[   41764] = 32'h727d5fe1;
    ram_cell[   41765] = 32'hb8f64522;
    ram_cell[   41766] = 32'hd9095845;
    ram_cell[   41767] = 32'h1ff6f8bc;
    ram_cell[   41768] = 32'h54732587;
    ram_cell[   41769] = 32'h33a6c1c7;
    ram_cell[   41770] = 32'h6e0cc22c;
    ram_cell[   41771] = 32'h2b9526e7;
    ram_cell[   41772] = 32'hf200f7c1;
    ram_cell[   41773] = 32'h26b39380;
    ram_cell[   41774] = 32'hcb03a1cf;
    ram_cell[   41775] = 32'h1342bd96;
    ram_cell[   41776] = 32'h9d71e863;
    ram_cell[   41777] = 32'hfc09d20c;
    ram_cell[   41778] = 32'hdaa124f7;
    ram_cell[   41779] = 32'hc25d25c3;
    ram_cell[   41780] = 32'h4757b577;
    ram_cell[   41781] = 32'h2a963f7b;
    ram_cell[   41782] = 32'hbc7b0ee8;
    ram_cell[   41783] = 32'heaa46854;
    ram_cell[   41784] = 32'he5c25a8f;
    ram_cell[   41785] = 32'h05fbe6f1;
    ram_cell[   41786] = 32'hc6cd3228;
    ram_cell[   41787] = 32'hbbcd2ef3;
    ram_cell[   41788] = 32'h55d31ce5;
    ram_cell[   41789] = 32'ha87748c5;
    ram_cell[   41790] = 32'h827e180f;
    ram_cell[   41791] = 32'ha714814e;
    ram_cell[   41792] = 32'h69f0ab91;
    ram_cell[   41793] = 32'h4d3b002b;
    ram_cell[   41794] = 32'hacfdb3df;
    ram_cell[   41795] = 32'h916c66ce;
    ram_cell[   41796] = 32'h3d804a20;
    ram_cell[   41797] = 32'ha44c9376;
    ram_cell[   41798] = 32'he9c9f11d;
    ram_cell[   41799] = 32'h26fc2b56;
    ram_cell[   41800] = 32'h7634d256;
    ram_cell[   41801] = 32'h47c81c5b;
    ram_cell[   41802] = 32'h28b51568;
    ram_cell[   41803] = 32'h69d7c59a;
    ram_cell[   41804] = 32'h6b8650cb;
    ram_cell[   41805] = 32'hf11a5895;
    ram_cell[   41806] = 32'heaa3049f;
    ram_cell[   41807] = 32'h2a371287;
    ram_cell[   41808] = 32'hb7493b24;
    ram_cell[   41809] = 32'h9871ca42;
    ram_cell[   41810] = 32'hf52e206c;
    ram_cell[   41811] = 32'hd3cb1006;
    ram_cell[   41812] = 32'h1aeba114;
    ram_cell[   41813] = 32'hfe846185;
    ram_cell[   41814] = 32'h10d7e593;
    ram_cell[   41815] = 32'hcef41f16;
    ram_cell[   41816] = 32'h95cdd39d;
    ram_cell[   41817] = 32'h305e7090;
    ram_cell[   41818] = 32'h5f4556a0;
    ram_cell[   41819] = 32'h51b66728;
    ram_cell[   41820] = 32'h45f337e4;
    ram_cell[   41821] = 32'h337e5f6d;
    ram_cell[   41822] = 32'h0fc9aeca;
    ram_cell[   41823] = 32'ha09a9b7a;
    ram_cell[   41824] = 32'hbbc0cce1;
    ram_cell[   41825] = 32'hc235d98f;
    ram_cell[   41826] = 32'he64d5aad;
    ram_cell[   41827] = 32'h5ccd541a;
    ram_cell[   41828] = 32'ha21f72d5;
    ram_cell[   41829] = 32'h0507a4d9;
    ram_cell[   41830] = 32'h38ed7801;
    ram_cell[   41831] = 32'hc7be661f;
    ram_cell[   41832] = 32'haefc80f0;
    ram_cell[   41833] = 32'h3b403029;
    ram_cell[   41834] = 32'ha37d1fb4;
    ram_cell[   41835] = 32'h89d9514e;
    ram_cell[   41836] = 32'h1c36c071;
    ram_cell[   41837] = 32'h7eeb05e4;
    ram_cell[   41838] = 32'h47f2b5dc;
    ram_cell[   41839] = 32'h79640e5a;
    ram_cell[   41840] = 32'hcaaf00b0;
    ram_cell[   41841] = 32'hc6fe5029;
    ram_cell[   41842] = 32'h5b291fe1;
    ram_cell[   41843] = 32'hbc1cf8f0;
    ram_cell[   41844] = 32'haafea9fe;
    ram_cell[   41845] = 32'h29fd1678;
    ram_cell[   41846] = 32'h7475c83d;
    ram_cell[   41847] = 32'hc2170e48;
    ram_cell[   41848] = 32'hbd334499;
    ram_cell[   41849] = 32'h0af2fb4d;
    ram_cell[   41850] = 32'h18937940;
    ram_cell[   41851] = 32'hc3997769;
    ram_cell[   41852] = 32'hb7e78f73;
    ram_cell[   41853] = 32'hb8fb8083;
    ram_cell[   41854] = 32'hf6c2c131;
    ram_cell[   41855] = 32'h2f608d19;
    ram_cell[   41856] = 32'he0f48093;
    ram_cell[   41857] = 32'h4b743ab0;
    ram_cell[   41858] = 32'hf2b9535d;
    ram_cell[   41859] = 32'h863a6f3a;
    ram_cell[   41860] = 32'h329dab5c;
    ram_cell[   41861] = 32'hbe15ea8d;
    ram_cell[   41862] = 32'h528d4020;
    ram_cell[   41863] = 32'h20b2a51c;
    ram_cell[   41864] = 32'h3ad2278e;
    ram_cell[   41865] = 32'hab90dc93;
    ram_cell[   41866] = 32'h52e6fdf4;
    ram_cell[   41867] = 32'h09e1b34a;
    ram_cell[   41868] = 32'h76104d7f;
    ram_cell[   41869] = 32'h03ae1127;
    ram_cell[   41870] = 32'h33be6134;
    ram_cell[   41871] = 32'h7d9b07ff;
    ram_cell[   41872] = 32'hd795aa5f;
    ram_cell[   41873] = 32'h2811d6bb;
    ram_cell[   41874] = 32'hcd3c8de3;
    ram_cell[   41875] = 32'h240b0037;
    ram_cell[   41876] = 32'h1fd69479;
    ram_cell[   41877] = 32'hff6c6772;
    ram_cell[   41878] = 32'h272330cb;
    ram_cell[   41879] = 32'h4ec2a0fc;
    ram_cell[   41880] = 32'hbae09f33;
    ram_cell[   41881] = 32'h2af2b3f3;
    ram_cell[   41882] = 32'h250c9f7a;
    ram_cell[   41883] = 32'h62072978;
    ram_cell[   41884] = 32'hd463f1ae;
    ram_cell[   41885] = 32'h77abfb6b;
    ram_cell[   41886] = 32'h29b207c3;
    ram_cell[   41887] = 32'h37ae5a4b;
    ram_cell[   41888] = 32'h9df9ff6d;
    ram_cell[   41889] = 32'h9a01d2f5;
    ram_cell[   41890] = 32'hbb4e3a65;
    ram_cell[   41891] = 32'h4d5301b8;
    ram_cell[   41892] = 32'h60727729;
    ram_cell[   41893] = 32'hbc63738a;
    ram_cell[   41894] = 32'h48d3b4f2;
    ram_cell[   41895] = 32'hdb50af28;
    ram_cell[   41896] = 32'ha76d9f90;
    ram_cell[   41897] = 32'h78179786;
    ram_cell[   41898] = 32'h79b36f97;
    ram_cell[   41899] = 32'h0916ab96;
    ram_cell[   41900] = 32'hf288e410;
    ram_cell[   41901] = 32'h8f9e9e9d;
    ram_cell[   41902] = 32'hf7688a72;
    ram_cell[   41903] = 32'h92232cc7;
    ram_cell[   41904] = 32'hd47de388;
    ram_cell[   41905] = 32'he84ad379;
    ram_cell[   41906] = 32'ha0d27477;
    ram_cell[   41907] = 32'h51537a37;
    ram_cell[   41908] = 32'h31b332f4;
    ram_cell[   41909] = 32'h7d72e478;
    ram_cell[   41910] = 32'h34d43d72;
    ram_cell[   41911] = 32'hbe7b924e;
    ram_cell[   41912] = 32'h26417ad8;
    ram_cell[   41913] = 32'h8753e020;
    ram_cell[   41914] = 32'hee5b160e;
    ram_cell[   41915] = 32'h3357d1d4;
    ram_cell[   41916] = 32'h25e19918;
    ram_cell[   41917] = 32'hfb1fd280;
    ram_cell[   41918] = 32'h52553f0e;
    ram_cell[   41919] = 32'ha339ff39;
    ram_cell[   41920] = 32'hc7efac22;
    ram_cell[   41921] = 32'hee2fe041;
    ram_cell[   41922] = 32'hf23690ef;
    ram_cell[   41923] = 32'hdda0137a;
    ram_cell[   41924] = 32'hb6399bc4;
    ram_cell[   41925] = 32'h1af1631c;
    ram_cell[   41926] = 32'he6d12d39;
    ram_cell[   41927] = 32'h01dc10d9;
    ram_cell[   41928] = 32'h398bde78;
    ram_cell[   41929] = 32'h09642299;
    ram_cell[   41930] = 32'hd227c4fd;
    ram_cell[   41931] = 32'h77964285;
    ram_cell[   41932] = 32'h887fbab7;
    ram_cell[   41933] = 32'h43db5335;
    ram_cell[   41934] = 32'h6a8ce031;
    ram_cell[   41935] = 32'hf7376a8d;
    ram_cell[   41936] = 32'hc95a1765;
    ram_cell[   41937] = 32'h13435303;
    ram_cell[   41938] = 32'h47a88fb2;
    ram_cell[   41939] = 32'h9a615d2c;
    ram_cell[   41940] = 32'he5f213c0;
    ram_cell[   41941] = 32'heb11ca68;
    ram_cell[   41942] = 32'h49749aad;
    ram_cell[   41943] = 32'h2c1045c0;
    ram_cell[   41944] = 32'h2028dc5f;
    ram_cell[   41945] = 32'hc2e51016;
    ram_cell[   41946] = 32'h6d400267;
    ram_cell[   41947] = 32'h980d1caf;
    ram_cell[   41948] = 32'ha5746c56;
    ram_cell[   41949] = 32'hbca29e7d;
    ram_cell[   41950] = 32'h1026fd8f;
    ram_cell[   41951] = 32'h3e1c2649;
    ram_cell[   41952] = 32'hd2cb2cc5;
    ram_cell[   41953] = 32'h43118ef4;
    ram_cell[   41954] = 32'h42252c69;
    ram_cell[   41955] = 32'h89db9f4e;
    ram_cell[   41956] = 32'he1db0da3;
    ram_cell[   41957] = 32'hec8d6d0e;
    ram_cell[   41958] = 32'hf27def04;
    ram_cell[   41959] = 32'h8689149d;
    ram_cell[   41960] = 32'h50c6d5c2;
    ram_cell[   41961] = 32'had2d4add;
    ram_cell[   41962] = 32'hb484b43b;
    ram_cell[   41963] = 32'h653c99af;
    ram_cell[   41964] = 32'hb640aedf;
    ram_cell[   41965] = 32'ha4f9f90e;
    ram_cell[   41966] = 32'h13df450c;
    ram_cell[   41967] = 32'hf6180342;
    ram_cell[   41968] = 32'h3b124723;
    ram_cell[   41969] = 32'h931f6ea9;
    ram_cell[   41970] = 32'h8b9e76fd;
    ram_cell[   41971] = 32'h4868b1a8;
    ram_cell[   41972] = 32'hfc3563dc;
    ram_cell[   41973] = 32'hefa18c16;
    ram_cell[   41974] = 32'h7936b3a0;
    ram_cell[   41975] = 32'h0b7abd4e;
    ram_cell[   41976] = 32'h580bb414;
    ram_cell[   41977] = 32'hd948c9df;
    ram_cell[   41978] = 32'h7f2997d2;
    ram_cell[   41979] = 32'h2e1077fb;
    ram_cell[   41980] = 32'hfa226ef7;
    ram_cell[   41981] = 32'h73e597ec;
    ram_cell[   41982] = 32'h930d748e;
    ram_cell[   41983] = 32'h9011a905;
    ram_cell[   41984] = 32'ha3c2db21;
    ram_cell[   41985] = 32'h975e76d1;
    ram_cell[   41986] = 32'hf708c1a7;
    ram_cell[   41987] = 32'hf1aa68f9;
    ram_cell[   41988] = 32'hac4e10c3;
    ram_cell[   41989] = 32'ha80ff00f;
    ram_cell[   41990] = 32'hf03ffba2;
    ram_cell[   41991] = 32'hcb29af29;
    ram_cell[   41992] = 32'h7afbcb03;
    ram_cell[   41993] = 32'h24d52fe6;
    ram_cell[   41994] = 32'hc0a52883;
    ram_cell[   41995] = 32'he07bb6b2;
    ram_cell[   41996] = 32'hb46d6e4e;
    ram_cell[   41997] = 32'h84c18934;
    ram_cell[   41998] = 32'h4bf4ae98;
    ram_cell[   41999] = 32'h62775374;
    ram_cell[   42000] = 32'h6fdef2c9;
    ram_cell[   42001] = 32'h6e465137;
    ram_cell[   42002] = 32'hffb2a8cf;
    ram_cell[   42003] = 32'ha94f8b0b;
    ram_cell[   42004] = 32'h72664d25;
    ram_cell[   42005] = 32'h537070aa;
    ram_cell[   42006] = 32'hf4905d3d;
    ram_cell[   42007] = 32'h8534b680;
    ram_cell[   42008] = 32'hc65de3ea;
    ram_cell[   42009] = 32'h75931a0f;
    ram_cell[   42010] = 32'h2065ca4f;
    ram_cell[   42011] = 32'h02b04e99;
    ram_cell[   42012] = 32'hb4630eab;
    ram_cell[   42013] = 32'hb84f7506;
    ram_cell[   42014] = 32'h0683be65;
    ram_cell[   42015] = 32'h8df57aba;
    ram_cell[   42016] = 32'h1eb8dd06;
    ram_cell[   42017] = 32'h9558f6f7;
    ram_cell[   42018] = 32'h30f2e28e;
    ram_cell[   42019] = 32'h8872812c;
    ram_cell[   42020] = 32'hd180127b;
    ram_cell[   42021] = 32'hd2557268;
    ram_cell[   42022] = 32'h1cef06bf;
    ram_cell[   42023] = 32'h4849f92b;
    ram_cell[   42024] = 32'h127a6c92;
    ram_cell[   42025] = 32'h26a84e02;
    ram_cell[   42026] = 32'h7d140c8f;
    ram_cell[   42027] = 32'h3b2d7c1a;
    ram_cell[   42028] = 32'h45faa82c;
    ram_cell[   42029] = 32'h8784f41c;
    ram_cell[   42030] = 32'h1f5d0779;
    ram_cell[   42031] = 32'hd7d6527c;
    ram_cell[   42032] = 32'h882ea390;
    ram_cell[   42033] = 32'h062d8a06;
    ram_cell[   42034] = 32'h6817da85;
    ram_cell[   42035] = 32'h0ff6cece;
    ram_cell[   42036] = 32'h4ab3c631;
    ram_cell[   42037] = 32'h66b703b4;
    ram_cell[   42038] = 32'h0717c692;
    ram_cell[   42039] = 32'h44f45ace;
    ram_cell[   42040] = 32'h1b6b97a1;
    ram_cell[   42041] = 32'h34247d2d;
    ram_cell[   42042] = 32'h543acf0a;
    ram_cell[   42043] = 32'hb50538a4;
    ram_cell[   42044] = 32'h71fa6866;
    ram_cell[   42045] = 32'h115b6f23;
    ram_cell[   42046] = 32'h75306710;
    ram_cell[   42047] = 32'hf35947f2;
    ram_cell[   42048] = 32'h0a29ea56;
    ram_cell[   42049] = 32'h00fe1a64;
    ram_cell[   42050] = 32'h6f717dec;
    ram_cell[   42051] = 32'h37e79643;
    ram_cell[   42052] = 32'ha4b1242f;
    ram_cell[   42053] = 32'h54234f04;
    ram_cell[   42054] = 32'h1a482d59;
    ram_cell[   42055] = 32'h89bca7a0;
    ram_cell[   42056] = 32'h091281bb;
    ram_cell[   42057] = 32'hc5b70dea;
    ram_cell[   42058] = 32'h2252edce;
    ram_cell[   42059] = 32'h5ba214b0;
    ram_cell[   42060] = 32'hede5f07b;
    ram_cell[   42061] = 32'h4796ebe8;
    ram_cell[   42062] = 32'hc570e880;
    ram_cell[   42063] = 32'h2cdb8ce9;
    ram_cell[   42064] = 32'hc5021581;
    ram_cell[   42065] = 32'h7eb5053b;
    ram_cell[   42066] = 32'hae00d71f;
    ram_cell[   42067] = 32'h5856dc0b;
    ram_cell[   42068] = 32'h606a3a4c;
    ram_cell[   42069] = 32'hc3362dfd;
    ram_cell[   42070] = 32'ha41f7ed9;
    ram_cell[   42071] = 32'h3b10c919;
    ram_cell[   42072] = 32'h314c364b;
    ram_cell[   42073] = 32'hb6e54147;
    ram_cell[   42074] = 32'h3d767523;
    ram_cell[   42075] = 32'h81312484;
    ram_cell[   42076] = 32'hae7f52e6;
    ram_cell[   42077] = 32'he3880091;
    ram_cell[   42078] = 32'h5b722309;
    ram_cell[   42079] = 32'he3ceb5c7;
    ram_cell[   42080] = 32'h711acaa0;
    ram_cell[   42081] = 32'h560c4795;
    ram_cell[   42082] = 32'h73de0370;
    ram_cell[   42083] = 32'hf3d1f70b;
    ram_cell[   42084] = 32'hd36597ed;
    ram_cell[   42085] = 32'h9048ebd0;
    ram_cell[   42086] = 32'haf7461df;
    ram_cell[   42087] = 32'h5cb8c392;
    ram_cell[   42088] = 32'hdcf05eeb;
    ram_cell[   42089] = 32'hc3565358;
    ram_cell[   42090] = 32'h45992e5a;
    ram_cell[   42091] = 32'h8718ecf1;
    ram_cell[   42092] = 32'h67e9b5dd;
    ram_cell[   42093] = 32'h3bee8bbf;
    ram_cell[   42094] = 32'h912ebfad;
    ram_cell[   42095] = 32'hc1723428;
    ram_cell[   42096] = 32'hdc112720;
    ram_cell[   42097] = 32'hc4e194dc;
    ram_cell[   42098] = 32'h826b6b17;
    ram_cell[   42099] = 32'hd9f16cbe;
    ram_cell[   42100] = 32'h1c82a186;
    ram_cell[   42101] = 32'hcaf2a368;
    ram_cell[   42102] = 32'h7ba91e91;
    ram_cell[   42103] = 32'hed342688;
    ram_cell[   42104] = 32'h9396cec8;
    ram_cell[   42105] = 32'hf7d04fc0;
    ram_cell[   42106] = 32'hdb25f46d;
    ram_cell[   42107] = 32'h20a5c1ab;
    ram_cell[   42108] = 32'h4ce68c2e;
    ram_cell[   42109] = 32'hae3c7982;
    ram_cell[   42110] = 32'ha48a3741;
    ram_cell[   42111] = 32'hdbfb2677;
    ram_cell[   42112] = 32'hd36438ce;
    ram_cell[   42113] = 32'h9aa56c40;
    ram_cell[   42114] = 32'h2390584f;
    ram_cell[   42115] = 32'h5841c1ef;
    ram_cell[   42116] = 32'hc0d2882a;
    ram_cell[   42117] = 32'h58117e60;
    ram_cell[   42118] = 32'h0272e67c;
    ram_cell[   42119] = 32'h08eb8b7b;
    ram_cell[   42120] = 32'h231078a5;
    ram_cell[   42121] = 32'hebf955e1;
    ram_cell[   42122] = 32'h81ab3729;
    ram_cell[   42123] = 32'hecf5ae6e;
    ram_cell[   42124] = 32'h37868a13;
    ram_cell[   42125] = 32'hff8579d8;
    ram_cell[   42126] = 32'h3b08b1d4;
    ram_cell[   42127] = 32'h140bc072;
    ram_cell[   42128] = 32'h87ab279d;
    ram_cell[   42129] = 32'h19b38348;
    ram_cell[   42130] = 32'hffa0b62a;
    ram_cell[   42131] = 32'hb29cbc83;
    ram_cell[   42132] = 32'hf1656569;
    ram_cell[   42133] = 32'h006c2f44;
    ram_cell[   42134] = 32'h6970301e;
    ram_cell[   42135] = 32'h83f81d31;
    ram_cell[   42136] = 32'h3a99a611;
    ram_cell[   42137] = 32'hd5a77f50;
    ram_cell[   42138] = 32'heea056ff;
    ram_cell[   42139] = 32'h1249a5a9;
    ram_cell[   42140] = 32'hbed6f9f3;
    ram_cell[   42141] = 32'h568cbbce;
    ram_cell[   42142] = 32'he06ed200;
    ram_cell[   42143] = 32'h2306c8c9;
    ram_cell[   42144] = 32'hdc2bf04e;
    ram_cell[   42145] = 32'h97d3ae02;
    ram_cell[   42146] = 32'ha34c2375;
    ram_cell[   42147] = 32'h87893982;
    ram_cell[   42148] = 32'h9d9d5714;
    ram_cell[   42149] = 32'hd1e182b6;
    ram_cell[   42150] = 32'h7fbd17fc;
    ram_cell[   42151] = 32'hb80e8586;
    ram_cell[   42152] = 32'h02085b3f;
    ram_cell[   42153] = 32'h713a3ffd;
    ram_cell[   42154] = 32'h874f2ddd;
    ram_cell[   42155] = 32'h1af7c177;
    ram_cell[   42156] = 32'he0a70211;
    ram_cell[   42157] = 32'h478d1db2;
    ram_cell[   42158] = 32'h0a20c110;
    ram_cell[   42159] = 32'hcbc98d83;
    ram_cell[   42160] = 32'h33ac66ec;
    ram_cell[   42161] = 32'h84b001f2;
    ram_cell[   42162] = 32'heed3092f;
    ram_cell[   42163] = 32'h6068acf3;
    ram_cell[   42164] = 32'hcf5d6f05;
    ram_cell[   42165] = 32'hdd18ccee;
    ram_cell[   42166] = 32'hcc6cf8f3;
    ram_cell[   42167] = 32'h8bf4e220;
    ram_cell[   42168] = 32'h003478f3;
    ram_cell[   42169] = 32'hf015a6d7;
    ram_cell[   42170] = 32'h07fb2baa;
    ram_cell[   42171] = 32'h67ed436b;
    ram_cell[   42172] = 32'h78961d01;
    ram_cell[   42173] = 32'h819dbe2a;
    ram_cell[   42174] = 32'h000bbd20;
    ram_cell[   42175] = 32'hd6fef660;
    ram_cell[   42176] = 32'h2b40f113;
    ram_cell[   42177] = 32'h3c72191a;
    ram_cell[   42178] = 32'h86e1d83f;
    ram_cell[   42179] = 32'h74f8a1b3;
    ram_cell[   42180] = 32'h611f4306;
    ram_cell[   42181] = 32'h54cb8f18;
    ram_cell[   42182] = 32'h3688bfa6;
    ram_cell[   42183] = 32'he6568277;
    ram_cell[   42184] = 32'h427977c8;
    ram_cell[   42185] = 32'haffd563d;
    ram_cell[   42186] = 32'h6f65222d;
    ram_cell[   42187] = 32'h6aa53762;
    ram_cell[   42188] = 32'h3baeb82e;
    ram_cell[   42189] = 32'hd0022d59;
    ram_cell[   42190] = 32'hf13084d6;
    ram_cell[   42191] = 32'hf3f45e7d;
    ram_cell[   42192] = 32'h124aedb9;
    ram_cell[   42193] = 32'hf442a35b;
    ram_cell[   42194] = 32'h79705955;
    ram_cell[   42195] = 32'h681dac35;
    ram_cell[   42196] = 32'h08a5b06b;
    ram_cell[   42197] = 32'h2aff3eed;
    ram_cell[   42198] = 32'hdc537b19;
    ram_cell[   42199] = 32'h22a1ff5c;
    ram_cell[   42200] = 32'h9cb82bec;
    ram_cell[   42201] = 32'h46a6b4bb;
    ram_cell[   42202] = 32'h8c9e7295;
    ram_cell[   42203] = 32'hc3043bdc;
    ram_cell[   42204] = 32'h26589229;
    ram_cell[   42205] = 32'h99e1aa34;
    ram_cell[   42206] = 32'h534381d8;
    ram_cell[   42207] = 32'h4c755e5d;
    ram_cell[   42208] = 32'hf72f40db;
    ram_cell[   42209] = 32'h4a58a6e0;
    ram_cell[   42210] = 32'hba42667d;
    ram_cell[   42211] = 32'hdd131c68;
    ram_cell[   42212] = 32'h4ea537ea;
    ram_cell[   42213] = 32'h48237a2e;
    ram_cell[   42214] = 32'hc2375aff;
    ram_cell[   42215] = 32'he8d79d9e;
    ram_cell[   42216] = 32'h16efdf64;
    ram_cell[   42217] = 32'h0dafcb8e;
    ram_cell[   42218] = 32'h6a5617bb;
    ram_cell[   42219] = 32'hd45b4946;
    ram_cell[   42220] = 32'hc7f05a4d;
    ram_cell[   42221] = 32'hbd238280;
    ram_cell[   42222] = 32'h5b585b0d;
    ram_cell[   42223] = 32'hb7a0187b;
    ram_cell[   42224] = 32'h99bf74bc;
    ram_cell[   42225] = 32'h42bb62f3;
    ram_cell[   42226] = 32'hb4c10cd4;
    ram_cell[   42227] = 32'h0c65f487;
    ram_cell[   42228] = 32'h78962b32;
    ram_cell[   42229] = 32'h27545134;
    ram_cell[   42230] = 32'h6ccdfc0b;
    ram_cell[   42231] = 32'h32049796;
    ram_cell[   42232] = 32'h19106df2;
    ram_cell[   42233] = 32'h47862e70;
    ram_cell[   42234] = 32'h72a9cc8f;
    ram_cell[   42235] = 32'hd93a38cb;
    ram_cell[   42236] = 32'h109ab43c;
    ram_cell[   42237] = 32'h435cdfca;
    ram_cell[   42238] = 32'hdca05bbf;
    ram_cell[   42239] = 32'hac13db74;
    ram_cell[   42240] = 32'h5512b255;
    ram_cell[   42241] = 32'hf67df477;
    ram_cell[   42242] = 32'he30172a7;
    ram_cell[   42243] = 32'hdcb67ccf;
    ram_cell[   42244] = 32'had444742;
    ram_cell[   42245] = 32'h1d13761b;
    ram_cell[   42246] = 32'h06714549;
    ram_cell[   42247] = 32'h41577eab;
    ram_cell[   42248] = 32'h849e57ec;
    ram_cell[   42249] = 32'h8f643c04;
    ram_cell[   42250] = 32'hb9b541da;
    ram_cell[   42251] = 32'hf315a221;
    ram_cell[   42252] = 32'h289fdb2b;
    ram_cell[   42253] = 32'he6115712;
    ram_cell[   42254] = 32'h4a16e791;
    ram_cell[   42255] = 32'h36c2e116;
    ram_cell[   42256] = 32'hd8bff10a;
    ram_cell[   42257] = 32'h3b9d4461;
    ram_cell[   42258] = 32'hf075e789;
    ram_cell[   42259] = 32'h28025add;
    ram_cell[   42260] = 32'h13ef9e7f;
    ram_cell[   42261] = 32'h4ddc75fd;
    ram_cell[   42262] = 32'hbce1a054;
    ram_cell[   42263] = 32'hccb10551;
    ram_cell[   42264] = 32'h5baeab83;
    ram_cell[   42265] = 32'h8d0b4fb7;
    ram_cell[   42266] = 32'h539c1e8b;
    ram_cell[   42267] = 32'hde006fca;
    ram_cell[   42268] = 32'h9ebf7acd;
    ram_cell[   42269] = 32'h45cf6976;
    ram_cell[   42270] = 32'h766036ac;
    ram_cell[   42271] = 32'h4326fc35;
    ram_cell[   42272] = 32'h000ab810;
    ram_cell[   42273] = 32'hd8096b97;
    ram_cell[   42274] = 32'h358746d7;
    ram_cell[   42275] = 32'h28e3e8eb;
    ram_cell[   42276] = 32'h746c9617;
    ram_cell[   42277] = 32'h7c85eab9;
    ram_cell[   42278] = 32'hfe2abce2;
    ram_cell[   42279] = 32'h54aed2df;
    ram_cell[   42280] = 32'h512e0f1e;
    ram_cell[   42281] = 32'hc1ee7faf;
    ram_cell[   42282] = 32'h33ef7f21;
    ram_cell[   42283] = 32'h658e987b;
    ram_cell[   42284] = 32'h63aae56f;
    ram_cell[   42285] = 32'h22d81612;
    ram_cell[   42286] = 32'h87ad8b6a;
    ram_cell[   42287] = 32'h44d575c9;
    ram_cell[   42288] = 32'hded794f5;
    ram_cell[   42289] = 32'h250965c8;
    ram_cell[   42290] = 32'ha992ed5c;
    ram_cell[   42291] = 32'h1be6228c;
    ram_cell[   42292] = 32'h55239a8a;
    ram_cell[   42293] = 32'h8b65ab7a;
    ram_cell[   42294] = 32'h71022481;
    ram_cell[   42295] = 32'h8b4fe5a8;
    ram_cell[   42296] = 32'h2857b8e7;
    ram_cell[   42297] = 32'h3d235edc;
    ram_cell[   42298] = 32'h2a9879d2;
    ram_cell[   42299] = 32'h8d066cf4;
    ram_cell[   42300] = 32'h5fe00b2a;
    ram_cell[   42301] = 32'h0bf5f9af;
    ram_cell[   42302] = 32'hb43bb180;
    ram_cell[   42303] = 32'h05b60522;
    ram_cell[   42304] = 32'h9cd5c386;
    ram_cell[   42305] = 32'hbbfbbd35;
    ram_cell[   42306] = 32'ha2b812d2;
    ram_cell[   42307] = 32'h18c3e6e2;
    ram_cell[   42308] = 32'h5991d3a4;
    ram_cell[   42309] = 32'h16ac26fe;
    ram_cell[   42310] = 32'h4a1f103f;
    ram_cell[   42311] = 32'heeb0bec7;
    ram_cell[   42312] = 32'h84e5b196;
    ram_cell[   42313] = 32'hf70346a5;
    ram_cell[   42314] = 32'h309bdc69;
    ram_cell[   42315] = 32'h32c0eab0;
    ram_cell[   42316] = 32'h2fb97212;
    ram_cell[   42317] = 32'h9e758b62;
    ram_cell[   42318] = 32'h4c796719;
    ram_cell[   42319] = 32'h4b4512f4;
    ram_cell[   42320] = 32'h685ff807;
    ram_cell[   42321] = 32'h7adfb405;
    ram_cell[   42322] = 32'h9818dc79;
    ram_cell[   42323] = 32'h805d7d50;
    ram_cell[   42324] = 32'hf5a5e077;
    ram_cell[   42325] = 32'h4a18610a;
    ram_cell[   42326] = 32'h0628a62c;
    ram_cell[   42327] = 32'h3f6dacdd;
    ram_cell[   42328] = 32'hf4874d52;
    ram_cell[   42329] = 32'h200353e9;
    ram_cell[   42330] = 32'h6e02613c;
    ram_cell[   42331] = 32'hb56bd093;
    ram_cell[   42332] = 32'hccbe7d17;
    ram_cell[   42333] = 32'hceb4d8fe;
    ram_cell[   42334] = 32'h7030c2a4;
    ram_cell[   42335] = 32'h70de2166;
    ram_cell[   42336] = 32'hc73b2284;
    ram_cell[   42337] = 32'h0f462a26;
    ram_cell[   42338] = 32'h72364843;
    ram_cell[   42339] = 32'h1c3cef51;
    ram_cell[   42340] = 32'h38a732e8;
    ram_cell[   42341] = 32'h3f57a70a;
    ram_cell[   42342] = 32'hf270b640;
    ram_cell[   42343] = 32'h4d58e7bb;
    ram_cell[   42344] = 32'he8867502;
    ram_cell[   42345] = 32'hde0d1b42;
    ram_cell[   42346] = 32'he17162ed;
    ram_cell[   42347] = 32'h44eb1e28;
    ram_cell[   42348] = 32'h5cf9d841;
    ram_cell[   42349] = 32'h1c991e69;
    ram_cell[   42350] = 32'hdef55ce5;
    ram_cell[   42351] = 32'h42d0ce88;
    ram_cell[   42352] = 32'hafd10136;
    ram_cell[   42353] = 32'hca8be3be;
    ram_cell[   42354] = 32'he60bd8d1;
    ram_cell[   42355] = 32'hd514f008;
    ram_cell[   42356] = 32'hc6f76909;
    ram_cell[   42357] = 32'h0159e5c5;
    ram_cell[   42358] = 32'hfd565e16;
    ram_cell[   42359] = 32'hf137ac19;
    ram_cell[   42360] = 32'h13ccd4e9;
    ram_cell[   42361] = 32'h0aef00da;
    ram_cell[   42362] = 32'h619b493d;
    ram_cell[   42363] = 32'h94372656;
    ram_cell[   42364] = 32'h3c073829;
    ram_cell[   42365] = 32'h89afb0bc;
    ram_cell[   42366] = 32'hb3ffcda9;
    ram_cell[   42367] = 32'h51cd87f8;
    ram_cell[   42368] = 32'h0535cb23;
    ram_cell[   42369] = 32'h3cacaa9d;
    ram_cell[   42370] = 32'h7ea89e9f;
    ram_cell[   42371] = 32'hcd9531e2;
    ram_cell[   42372] = 32'h89e229de;
    ram_cell[   42373] = 32'h5f174599;
    ram_cell[   42374] = 32'h6349791b;
    ram_cell[   42375] = 32'h9ad77457;
    ram_cell[   42376] = 32'h389514f5;
    ram_cell[   42377] = 32'hbfe9d54e;
    ram_cell[   42378] = 32'h8a420ae4;
    ram_cell[   42379] = 32'h466397c4;
    ram_cell[   42380] = 32'hb54df810;
    ram_cell[   42381] = 32'h53b475ac;
    ram_cell[   42382] = 32'ha4b8d50c;
    ram_cell[   42383] = 32'h2ef95887;
    ram_cell[   42384] = 32'hec9fa6a0;
    ram_cell[   42385] = 32'h901aac97;
    ram_cell[   42386] = 32'h56a831f8;
    ram_cell[   42387] = 32'h92517586;
    ram_cell[   42388] = 32'h6b261257;
    ram_cell[   42389] = 32'hc916df62;
    ram_cell[   42390] = 32'h4d897b8f;
    ram_cell[   42391] = 32'h99618e6f;
    ram_cell[   42392] = 32'hf06772a3;
    ram_cell[   42393] = 32'h15984afa;
    ram_cell[   42394] = 32'h278c8cd0;
    ram_cell[   42395] = 32'h8cf87a0a;
    ram_cell[   42396] = 32'h41df56f9;
    ram_cell[   42397] = 32'hc540e4da;
    ram_cell[   42398] = 32'ha0a51ad9;
    ram_cell[   42399] = 32'ha31d30eb;
    ram_cell[   42400] = 32'hf856a423;
    ram_cell[   42401] = 32'h394d01ca;
    ram_cell[   42402] = 32'hb7e76509;
    ram_cell[   42403] = 32'h0590666d;
    ram_cell[   42404] = 32'hf583da23;
    ram_cell[   42405] = 32'hec50f9cb;
    ram_cell[   42406] = 32'h545fa230;
    ram_cell[   42407] = 32'h5906943b;
    ram_cell[   42408] = 32'hd781b2b1;
    ram_cell[   42409] = 32'h91f553a3;
    ram_cell[   42410] = 32'h87b107c2;
    ram_cell[   42411] = 32'h57647602;
    ram_cell[   42412] = 32'h584040af;
    ram_cell[   42413] = 32'h400be630;
    ram_cell[   42414] = 32'h0ee13165;
    ram_cell[   42415] = 32'hf5e6bf05;
    ram_cell[   42416] = 32'h9df748be;
    ram_cell[   42417] = 32'hc4c6b596;
    ram_cell[   42418] = 32'h1aa5e121;
    ram_cell[   42419] = 32'ha3e3c543;
    ram_cell[   42420] = 32'h5e5c15e3;
    ram_cell[   42421] = 32'h0f3c97c7;
    ram_cell[   42422] = 32'hbc21d46c;
    ram_cell[   42423] = 32'hb59b4aa6;
    ram_cell[   42424] = 32'hd6ac2bff;
    ram_cell[   42425] = 32'h0f801425;
    ram_cell[   42426] = 32'h64a862fb;
    ram_cell[   42427] = 32'h54015394;
    ram_cell[   42428] = 32'h40abb858;
    ram_cell[   42429] = 32'h5a5ed4b2;
    ram_cell[   42430] = 32'h3533f795;
    ram_cell[   42431] = 32'h3e9e4743;
    ram_cell[   42432] = 32'h0b011303;
    ram_cell[   42433] = 32'he1385a90;
    ram_cell[   42434] = 32'h49d4e574;
    ram_cell[   42435] = 32'hb2d24900;
    ram_cell[   42436] = 32'h2436c3a6;
    ram_cell[   42437] = 32'hd32e47bf;
    ram_cell[   42438] = 32'h4087f872;
    ram_cell[   42439] = 32'ha5215906;
    ram_cell[   42440] = 32'h2143f89e;
    ram_cell[   42441] = 32'h42db4d1e;
    ram_cell[   42442] = 32'hd0322174;
    ram_cell[   42443] = 32'h335be932;
    ram_cell[   42444] = 32'hbf4bc936;
    ram_cell[   42445] = 32'hfd9ab189;
    ram_cell[   42446] = 32'hf73c96ff;
    ram_cell[   42447] = 32'hf6d9563c;
    ram_cell[   42448] = 32'h47e097a6;
    ram_cell[   42449] = 32'hfa550e1b;
    ram_cell[   42450] = 32'hed80ebe5;
    ram_cell[   42451] = 32'h46c0ed62;
    ram_cell[   42452] = 32'h8e10fda1;
    ram_cell[   42453] = 32'h851110e5;
    ram_cell[   42454] = 32'h9cf11fb1;
    ram_cell[   42455] = 32'haa06c819;
    ram_cell[   42456] = 32'ha4996e77;
    ram_cell[   42457] = 32'h4a716a79;
    ram_cell[   42458] = 32'h2ad6c678;
    ram_cell[   42459] = 32'h318b992f;
    ram_cell[   42460] = 32'hdc385ef3;
    ram_cell[   42461] = 32'h6c776692;
    ram_cell[   42462] = 32'h082d72bf;
    ram_cell[   42463] = 32'hdd29660e;
    ram_cell[   42464] = 32'ha1583d00;
    ram_cell[   42465] = 32'h681a062e;
    ram_cell[   42466] = 32'h7e1d371c;
    ram_cell[   42467] = 32'hee179f58;
    ram_cell[   42468] = 32'h6777aae9;
    ram_cell[   42469] = 32'h71f71147;
    ram_cell[   42470] = 32'h4335cc88;
    ram_cell[   42471] = 32'he77310e0;
    ram_cell[   42472] = 32'h0bf2b93e;
    ram_cell[   42473] = 32'hfb8413d7;
    ram_cell[   42474] = 32'hc7361edb;
    ram_cell[   42475] = 32'h40738bab;
    ram_cell[   42476] = 32'h8ed76ca0;
    ram_cell[   42477] = 32'hf95a5696;
    ram_cell[   42478] = 32'h64287159;
    ram_cell[   42479] = 32'hf1c98a07;
    ram_cell[   42480] = 32'h15c6357d;
    ram_cell[   42481] = 32'h115907b5;
    ram_cell[   42482] = 32'he6bd232f;
    ram_cell[   42483] = 32'h789478d5;
    ram_cell[   42484] = 32'h9c3daace;
    ram_cell[   42485] = 32'h2e84601d;
    ram_cell[   42486] = 32'h340034b7;
    ram_cell[   42487] = 32'h2369efa8;
    ram_cell[   42488] = 32'h90624e62;
    ram_cell[   42489] = 32'h6137fc6a;
    ram_cell[   42490] = 32'hb51c841f;
    ram_cell[   42491] = 32'h220aa196;
    ram_cell[   42492] = 32'hb0608587;
    ram_cell[   42493] = 32'h3ad867c1;
    ram_cell[   42494] = 32'h761207e7;
    ram_cell[   42495] = 32'h8779917b;
    ram_cell[   42496] = 32'hfd619fa6;
    ram_cell[   42497] = 32'h801253af;
    ram_cell[   42498] = 32'h8f7c6208;
    ram_cell[   42499] = 32'h23d2c1ed;
    ram_cell[   42500] = 32'ha0cabb57;
    ram_cell[   42501] = 32'haf9c87c0;
    ram_cell[   42502] = 32'hfae63c07;
    ram_cell[   42503] = 32'h13ee31a4;
    ram_cell[   42504] = 32'hecbd0051;
    ram_cell[   42505] = 32'he7c80301;
    ram_cell[   42506] = 32'h05744856;
    ram_cell[   42507] = 32'hd6a28252;
    ram_cell[   42508] = 32'h045000fa;
    ram_cell[   42509] = 32'haff59b8e;
    ram_cell[   42510] = 32'h52719e91;
    ram_cell[   42511] = 32'h03706e9e;
    ram_cell[   42512] = 32'h4f73f621;
    ram_cell[   42513] = 32'h1ebe7b2d;
    ram_cell[   42514] = 32'h72c4dd2e;
    ram_cell[   42515] = 32'hc36c304d;
    ram_cell[   42516] = 32'hf50d2d0b;
    ram_cell[   42517] = 32'h398eb53f;
    ram_cell[   42518] = 32'h734c65b3;
    ram_cell[   42519] = 32'h17507b86;
    ram_cell[   42520] = 32'h680ef254;
    ram_cell[   42521] = 32'hc5843028;
    ram_cell[   42522] = 32'ha04e1b15;
    ram_cell[   42523] = 32'hc6e1c8ea;
    ram_cell[   42524] = 32'hcda99f18;
    ram_cell[   42525] = 32'h1720ec51;
    ram_cell[   42526] = 32'ha723efa0;
    ram_cell[   42527] = 32'h01d34f18;
    ram_cell[   42528] = 32'h3594c754;
    ram_cell[   42529] = 32'hbdab6180;
    ram_cell[   42530] = 32'h98ec6f1a;
    ram_cell[   42531] = 32'he5ca62fb;
    ram_cell[   42532] = 32'h8e9e88e8;
    ram_cell[   42533] = 32'hc51373c8;
    ram_cell[   42534] = 32'h92f6b954;
    ram_cell[   42535] = 32'h2a2544f2;
    ram_cell[   42536] = 32'hd570f31e;
    ram_cell[   42537] = 32'h9159468e;
    ram_cell[   42538] = 32'hcf89ed7b;
    ram_cell[   42539] = 32'h4e6e967b;
    ram_cell[   42540] = 32'h480c1305;
    ram_cell[   42541] = 32'h40b244bb;
    ram_cell[   42542] = 32'h61103700;
    ram_cell[   42543] = 32'ha3b4ab70;
    ram_cell[   42544] = 32'hcc9713fb;
    ram_cell[   42545] = 32'hc1bf69e3;
    ram_cell[   42546] = 32'hc7913872;
    ram_cell[   42547] = 32'h042696a1;
    ram_cell[   42548] = 32'h029a11f2;
    ram_cell[   42549] = 32'hd464c155;
    ram_cell[   42550] = 32'h41996ae1;
    ram_cell[   42551] = 32'h6203b1b1;
    ram_cell[   42552] = 32'h78cebd59;
    ram_cell[   42553] = 32'hab1b9460;
    ram_cell[   42554] = 32'h2b231970;
    ram_cell[   42555] = 32'h63ad54cc;
    ram_cell[   42556] = 32'h05b5e3ab;
    ram_cell[   42557] = 32'haf6a5e10;
    ram_cell[   42558] = 32'hed936222;
    ram_cell[   42559] = 32'h0df7ab7c;
    ram_cell[   42560] = 32'h592099e9;
    ram_cell[   42561] = 32'h8e940f9c;
    ram_cell[   42562] = 32'h13f17055;
    ram_cell[   42563] = 32'hdf54899d;
    ram_cell[   42564] = 32'h4de9294c;
    ram_cell[   42565] = 32'h0b1f46f5;
    ram_cell[   42566] = 32'hbf77c520;
    ram_cell[   42567] = 32'he98435c5;
    ram_cell[   42568] = 32'h9efd4032;
    ram_cell[   42569] = 32'hc22f0567;
    ram_cell[   42570] = 32'h6813f510;
    ram_cell[   42571] = 32'hd5e4dfe1;
    ram_cell[   42572] = 32'h1710deb7;
    ram_cell[   42573] = 32'he5989f68;
    ram_cell[   42574] = 32'he3bf4b3e;
    ram_cell[   42575] = 32'hbdc9a6e3;
    ram_cell[   42576] = 32'h5160db08;
    ram_cell[   42577] = 32'h3e72a76f;
    ram_cell[   42578] = 32'h84f8d287;
    ram_cell[   42579] = 32'h481a940e;
    ram_cell[   42580] = 32'h35c792bb;
    ram_cell[   42581] = 32'h536b7bcf;
    ram_cell[   42582] = 32'he68b3371;
    ram_cell[   42583] = 32'h71e38060;
    ram_cell[   42584] = 32'hf8fbabd7;
    ram_cell[   42585] = 32'hff4dae82;
    ram_cell[   42586] = 32'hc476d387;
    ram_cell[   42587] = 32'hce7b0e06;
    ram_cell[   42588] = 32'hd8eeadaf;
    ram_cell[   42589] = 32'h2ea2efe2;
    ram_cell[   42590] = 32'hb85b8d84;
    ram_cell[   42591] = 32'hce5bc3b7;
    ram_cell[   42592] = 32'h754f6a46;
    ram_cell[   42593] = 32'h2c963d08;
    ram_cell[   42594] = 32'h48753bc3;
    ram_cell[   42595] = 32'h21b0644f;
    ram_cell[   42596] = 32'h8d02e2fa;
    ram_cell[   42597] = 32'h4420f807;
    ram_cell[   42598] = 32'h70f06bd7;
    ram_cell[   42599] = 32'hb6c16a0e;
    ram_cell[   42600] = 32'h8fbc5da2;
    ram_cell[   42601] = 32'hb8de4dcf;
    ram_cell[   42602] = 32'h9dae74f9;
    ram_cell[   42603] = 32'h7985c58f;
    ram_cell[   42604] = 32'h488bfccb;
    ram_cell[   42605] = 32'h517ffdcb;
    ram_cell[   42606] = 32'h7e5c78a0;
    ram_cell[   42607] = 32'h430c26f6;
    ram_cell[   42608] = 32'h5dd77d6f;
    ram_cell[   42609] = 32'h9a5e1030;
    ram_cell[   42610] = 32'h8cddec50;
    ram_cell[   42611] = 32'h60a35745;
    ram_cell[   42612] = 32'hd0ed2ecd;
    ram_cell[   42613] = 32'h07d56f99;
    ram_cell[   42614] = 32'h3f27c66b;
    ram_cell[   42615] = 32'haa2a4517;
    ram_cell[   42616] = 32'h6697940a;
    ram_cell[   42617] = 32'ha0264637;
    ram_cell[   42618] = 32'h98b855a5;
    ram_cell[   42619] = 32'ha6cf2329;
    ram_cell[   42620] = 32'h77b1ce1b;
    ram_cell[   42621] = 32'h70bb5d7c;
    ram_cell[   42622] = 32'h3ea6142f;
    ram_cell[   42623] = 32'h5d58d808;
    ram_cell[   42624] = 32'hb73aa6c1;
    ram_cell[   42625] = 32'h1f1e9275;
    ram_cell[   42626] = 32'h0a986278;
    ram_cell[   42627] = 32'h8599dd2d;
    ram_cell[   42628] = 32'h6f3c07ce;
    ram_cell[   42629] = 32'h3f7ed452;
    ram_cell[   42630] = 32'h50d9f32e;
    ram_cell[   42631] = 32'h90dab6ce;
    ram_cell[   42632] = 32'he01e4cd3;
    ram_cell[   42633] = 32'hd8542715;
    ram_cell[   42634] = 32'h4b794971;
    ram_cell[   42635] = 32'h3c9ba692;
    ram_cell[   42636] = 32'hf8ea533b;
    ram_cell[   42637] = 32'h205082b6;
    ram_cell[   42638] = 32'he5bb9845;
    ram_cell[   42639] = 32'h93557662;
    ram_cell[   42640] = 32'hd92546e4;
    ram_cell[   42641] = 32'hde79a0d9;
    ram_cell[   42642] = 32'hf7118042;
    ram_cell[   42643] = 32'ha6a91daa;
    ram_cell[   42644] = 32'h33adfa3b;
    ram_cell[   42645] = 32'hfa9e2429;
    ram_cell[   42646] = 32'h4701d9fe;
    ram_cell[   42647] = 32'h54e5c6da;
    ram_cell[   42648] = 32'hb1ddcb38;
    ram_cell[   42649] = 32'he45e00cf;
    ram_cell[   42650] = 32'h3287ee2a;
    ram_cell[   42651] = 32'h6d5a24bf;
    ram_cell[   42652] = 32'h85481249;
    ram_cell[   42653] = 32'hed314b48;
    ram_cell[   42654] = 32'h395d4691;
    ram_cell[   42655] = 32'h1dd95c1a;
    ram_cell[   42656] = 32'heae65705;
    ram_cell[   42657] = 32'h4ff9f9fa;
    ram_cell[   42658] = 32'h71bef5a1;
    ram_cell[   42659] = 32'hec064704;
    ram_cell[   42660] = 32'h5e4af871;
    ram_cell[   42661] = 32'hc35e43c6;
    ram_cell[   42662] = 32'h8f6ef567;
    ram_cell[   42663] = 32'h41393683;
    ram_cell[   42664] = 32'h122f886c;
    ram_cell[   42665] = 32'hb2244759;
    ram_cell[   42666] = 32'h1f2939d9;
    ram_cell[   42667] = 32'hf4ea6752;
    ram_cell[   42668] = 32'h40f2fe68;
    ram_cell[   42669] = 32'h1d608d76;
    ram_cell[   42670] = 32'h03c5d687;
    ram_cell[   42671] = 32'h10837d63;
    ram_cell[   42672] = 32'h0cb9498c;
    ram_cell[   42673] = 32'h8fecf3e9;
    ram_cell[   42674] = 32'h02f93e5d;
    ram_cell[   42675] = 32'h46b61f49;
    ram_cell[   42676] = 32'h091f5ae4;
    ram_cell[   42677] = 32'hb4ef7734;
    ram_cell[   42678] = 32'h8f4a4dcc;
    ram_cell[   42679] = 32'h7db7a967;
    ram_cell[   42680] = 32'h8ce58fc9;
    ram_cell[   42681] = 32'h5914a41d;
    ram_cell[   42682] = 32'h8406aba5;
    ram_cell[   42683] = 32'h752b67ea;
    ram_cell[   42684] = 32'he8b4916f;
    ram_cell[   42685] = 32'hdd9c6cea;
    ram_cell[   42686] = 32'hfd1a9427;
    ram_cell[   42687] = 32'ha4bc49a5;
    ram_cell[   42688] = 32'hee6d4562;
    ram_cell[   42689] = 32'h97afbc67;
    ram_cell[   42690] = 32'h219b86db;
    ram_cell[   42691] = 32'hd18da630;
    ram_cell[   42692] = 32'h1259dda9;
    ram_cell[   42693] = 32'h6f1ce864;
    ram_cell[   42694] = 32'hae26d8bd;
    ram_cell[   42695] = 32'h8d253be1;
    ram_cell[   42696] = 32'hfc194f47;
    ram_cell[   42697] = 32'hdc073c87;
    ram_cell[   42698] = 32'hc0471ce2;
    ram_cell[   42699] = 32'hd2cfa9f2;
    ram_cell[   42700] = 32'h8732be68;
    ram_cell[   42701] = 32'hf9b6040f;
    ram_cell[   42702] = 32'h66555cff;
    ram_cell[   42703] = 32'hb25de645;
    ram_cell[   42704] = 32'h60e96058;
    ram_cell[   42705] = 32'hd0823b2a;
    ram_cell[   42706] = 32'ha224a359;
    ram_cell[   42707] = 32'hedf87b81;
    ram_cell[   42708] = 32'h9f1d86f6;
    ram_cell[   42709] = 32'h551b2c6e;
    ram_cell[   42710] = 32'h2de26ff2;
    ram_cell[   42711] = 32'h063bbeb9;
    ram_cell[   42712] = 32'hedb04db7;
    ram_cell[   42713] = 32'h0280b0ea;
    ram_cell[   42714] = 32'hf5cf5f94;
    ram_cell[   42715] = 32'h28511807;
    ram_cell[   42716] = 32'hbc6be403;
    ram_cell[   42717] = 32'h379931b9;
    ram_cell[   42718] = 32'h2106ec39;
    ram_cell[   42719] = 32'hc9ab63dc;
    ram_cell[   42720] = 32'hc209252f;
    ram_cell[   42721] = 32'ha0ee641b;
    ram_cell[   42722] = 32'h81e0dc8e;
    ram_cell[   42723] = 32'h8364ddcf;
    ram_cell[   42724] = 32'ha30f6a07;
    ram_cell[   42725] = 32'hc95938bb;
    ram_cell[   42726] = 32'h6e4b2a8d;
    ram_cell[   42727] = 32'h4edfae9f;
    ram_cell[   42728] = 32'hb4da8a6b;
    ram_cell[   42729] = 32'hca2c17ac;
    ram_cell[   42730] = 32'h9181da3f;
    ram_cell[   42731] = 32'hee5205ca;
    ram_cell[   42732] = 32'haff90e48;
    ram_cell[   42733] = 32'h7547de64;
    ram_cell[   42734] = 32'h3c9c5180;
    ram_cell[   42735] = 32'hd8e00306;
    ram_cell[   42736] = 32'haa3a6f21;
    ram_cell[   42737] = 32'haed5c3cb;
    ram_cell[   42738] = 32'hfb8ddfdb;
    ram_cell[   42739] = 32'h60b9d361;
    ram_cell[   42740] = 32'haf431629;
    ram_cell[   42741] = 32'hbf83ccf5;
    ram_cell[   42742] = 32'hd2234ebc;
    ram_cell[   42743] = 32'hf4d1709c;
    ram_cell[   42744] = 32'h1ae735d1;
    ram_cell[   42745] = 32'h608bc1f9;
    ram_cell[   42746] = 32'h95d2e8c2;
    ram_cell[   42747] = 32'h6d39cf07;
    ram_cell[   42748] = 32'hcfe6a5d0;
    ram_cell[   42749] = 32'h98e2761f;
    ram_cell[   42750] = 32'hafa359c9;
    ram_cell[   42751] = 32'hc741fabd;
    ram_cell[   42752] = 32'h78ef402f;
    ram_cell[   42753] = 32'hce6469ac;
    ram_cell[   42754] = 32'h4ae6c52d;
    ram_cell[   42755] = 32'he70a8deb;
    ram_cell[   42756] = 32'haebcdcca;
    ram_cell[   42757] = 32'hc50ecf02;
    ram_cell[   42758] = 32'hbc63aa10;
    ram_cell[   42759] = 32'h0f83f165;
    ram_cell[   42760] = 32'h2cda3014;
    ram_cell[   42761] = 32'h968de5b0;
    ram_cell[   42762] = 32'h2cf3408e;
    ram_cell[   42763] = 32'hc40665c7;
    ram_cell[   42764] = 32'h0bf34b15;
    ram_cell[   42765] = 32'h12117ce6;
    ram_cell[   42766] = 32'ha6253d56;
    ram_cell[   42767] = 32'hd99100d3;
    ram_cell[   42768] = 32'hb3a98765;
    ram_cell[   42769] = 32'hed88fdb8;
    ram_cell[   42770] = 32'h875b29c6;
    ram_cell[   42771] = 32'hfe102b3c;
    ram_cell[   42772] = 32'h6109e20c;
    ram_cell[   42773] = 32'h66e9980e;
    ram_cell[   42774] = 32'ha5c1ad98;
    ram_cell[   42775] = 32'h153763c6;
    ram_cell[   42776] = 32'h30294534;
    ram_cell[   42777] = 32'h0fb47138;
    ram_cell[   42778] = 32'hf65ad4fa;
    ram_cell[   42779] = 32'hd4826766;
    ram_cell[   42780] = 32'h650d7812;
    ram_cell[   42781] = 32'ha87a98c1;
    ram_cell[   42782] = 32'he6718f72;
    ram_cell[   42783] = 32'h3a9f723e;
    ram_cell[   42784] = 32'h4e3bec0f;
    ram_cell[   42785] = 32'haf461401;
    ram_cell[   42786] = 32'h4ca2e985;
    ram_cell[   42787] = 32'hab0c7b74;
    ram_cell[   42788] = 32'ha3a5c7db;
    ram_cell[   42789] = 32'h8f22abd6;
    ram_cell[   42790] = 32'h003ae847;
    ram_cell[   42791] = 32'hb12ba78c;
    ram_cell[   42792] = 32'h8733e252;
    ram_cell[   42793] = 32'ha9a5e124;
    ram_cell[   42794] = 32'h169b1c0f;
    ram_cell[   42795] = 32'h5d7f3616;
    ram_cell[   42796] = 32'h19a38a5c;
    ram_cell[   42797] = 32'h41f79deb;
    ram_cell[   42798] = 32'h736cf982;
    ram_cell[   42799] = 32'hccb25960;
    ram_cell[   42800] = 32'h9615e895;
    ram_cell[   42801] = 32'h55b82511;
    ram_cell[   42802] = 32'h3f76ae30;
    ram_cell[   42803] = 32'h3092f701;
    ram_cell[   42804] = 32'hd88630ed;
    ram_cell[   42805] = 32'h192c1b04;
    ram_cell[   42806] = 32'hc21b0610;
    ram_cell[   42807] = 32'h9fb3a46d;
    ram_cell[   42808] = 32'ha4615655;
    ram_cell[   42809] = 32'h4fd78afe;
    ram_cell[   42810] = 32'h69e6eef5;
    ram_cell[   42811] = 32'h132adbe1;
    ram_cell[   42812] = 32'hb6d48d12;
    ram_cell[   42813] = 32'hb42ffe27;
    ram_cell[   42814] = 32'hb0cb7c6f;
    ram_cell[   42815] = 32'h81fb7b16;
    ram_cell[   42816] = 32'hac3e238f;
    ram_cell[   42817] = 32'hf08f3bbb;
    ram_cell[   42818] = 32'h327d4d28;
    ram_cell[   42819] = 32'h1930f393;
    ram_cell[   42820] = 32'h9e0c9443;
    ram_cell[   42821] = 32'hcac81034;
    ram_cell[   42822] = 32'hfc67402b;
    ram_cell[   42823] = 32'ha730046e;
    ram_cell[   42824] = 32'h49abbe5c;
    ram_cell[   42825] = 32'h235ea463;
    ram_cell[   42826] = 32'h78d05894;
    ram_cell[   42827] = 32'hc966c1d4;
    ram_cell[   42828] = 32'h2fe45bdf;
    ram_cell[   42829] = 32'hfe2bf5e1;
    ram_cell[   42830] = 32'hc529f980;
    ram_cell[   42831] = 32'h4afffb27;
    ram_cell[   42832] = 32'ha540c858;
    ram_cell[   42833] = 32'hb85059d9;
    ram_cell[   42834] = 32'h3e41549b;
    ram_cell[   42835] = 32'hab46c0e3;
    ram_cell[   42836] = 32'hfe0372c5;
    ram_cell[   42837] = 32'h356b3302;
    ram_cell[   42838] = 32'ha5c0b84c;
    ram_cell[   42839] = 32'h1ebb8b6b;
    ram_cell[   42840] = 32'h9929acb1;
    ram_cell[   42841] = 32'h5a96f915;
    ram_cell[   42842] = 32'hc52074e6;
    ram_cell[   42843] = 32'h26fb545a;
    ram_cell[   42844] = 32'h85b3ed25;
    ram_cell[   42845] = 32'h4e8f9e04;
    ram_cell[   42846] = 32'ha4b254ba;
    ram_cell[   42847] = 32'ha99b63f6;
    ram_cell[   42848] = 32'hf8f32b9b;
    ram_cell[   42849] = 32'h7945a7c4;
    ram_cell[   42850] = 32'h6ad62b0b;
    ram_cell[   42851] = 32'h8ffce97f;
    ram_cell[   42852] = 32'hc98ccddc;
    ram_cell[   42853] = 32'h76bd02f7;
    ram_cell[   42854] = 32'h0c47ddaf;
    ram_cell[   42855] = 32'h2ac930cd;
    ram_cell[   42856] = 32'ha6006942;
    ram_cell[   42857] = 32'ha3944253;
    ram_cell[   42858] = 32'h084d985d;
    ram_cell[   42859] = 32'h159b01ac;
    ram_cell[   42860] = 32'hcfbc31ea;
    ram_cell[   42861] = 32'h08533e3f;
    ram_cell[   42862] = 32'h7c4954ad;
    ram_cell[   42863] = 32'h6431cdad;
    ram_cell[   42864] = 32'h2e38a71d;
    ram_cell[   42865] = 32'hb931e26a;
    ram_cell[   42866] = 32'h1ee57a9d;
    ram_cell[   42867] = 32'h4cc98821;
    ram_cell[   42868] = 32'h19f5471a;
    ram_cell[   42869] = 32'h77bd17d5;
    ram_cell[   42870] = 32'h4403bb21;
    ram_cell[   42871] = 32'h21a0e7e3;
    ram_cell[   42872] = 32'hb5c7e281;
    ram_cell[   42873] = 32'h4699f581;
    ram_cell[   42874] = 32'h95b6e42f;
    ram_cell[   42875] = 32'h67c0ef72;
    ram_cell[   42876] = 32'h0a335887;
    ram_cell[   42877] = 32'h82f34590;
    ram_cell[   42878] = 32'h89ff1b5e;
    ram_cell[   42879] = 32'h666d05e7;
    ram_cell[   42880] = 32'hf8d18342;
    ram_cell[   42881] = 32'hdb777f4b;
    ram_cell[   42882] = 32'h723f68fc;
    ram_cell[   42883] = 32'h7bcb6e3e;
    ram_cell[   42884] = 32'h49ddc3b8;
    ram_cell[   42885] = 32'h587d95a7;
    ram_cell[   42886] = 32'he40aa6b7;
    ram_cell[   42887] = 32'h502e354e;
    ram_cell[   42888] = 32'h28ef4b0c;
    ram_cell[   42889] = 32'hd3da6c75;
    ram_cell[   42890] = 32'h35b04fcf;
    ram_cell[   42891] = 32'h86fdc4e3;
    ram_cell[   42892] = 32'h6ebdea3c;
    ram_cell[   42893] = 32'hb65dff92;
    ram_cell[   42894] = 32'hd4d10d78;
    ram_cell[   42895] = 32'ha5588745;
    ram_cell[   42896] = 32'ha8ed82b2;
    ram_cell[   42897] = 32'hdb587d08;
    ram_cell[   42898] = 32'h0aad068d;
    ram_cell[   42899] = 32'h8c06555e;
    ram_cell[   42900] = 32'ha2f6e020;
    ram_cell[   42901] = 32'h4e0404c7;
    ram_cell[   42902] = 32'h8a1593c1;
    ram_cell[   42903] = 32'hebfb0aed;
    ram_cell[   42904] = 32'h5083237a;
    ram_cell[   42905] = 32'hb19b3a4e;
    ram_cell[   42906] = 32'he2cb5bdf;
    ram_cell[   42907] = 32'h966ff056;
    ram_cell[   42908] = 32'h2244e572;
    ram_cell[   42909] = 32'h87d83991;
    ram_cell[   42910] = 32'h6997dfd5;
    ram_cell[   42911] = 32'h362bff91;
    ram_cell[   42912] = 32'hf50a8229;
    ram_cell[   42913] = 32'h96bcb699;
    ram_cell[   42914] = 32'h699e6cb1;
    ram_cell[   42915] = 32'h9b0ceb5a;
    ram_cell[   42916] = 32'h9054a0ec;
    ram_cell[   42917] = 32'hfd2bf781;
    ram_cell[   42918] = 32'h39ce3c3c;
    ram_cell[   42919] = 32'hc1e40ce9;
    ram_cell[   42920] = 32'hdc9cbdaa;
    ram_cell[   42921] = 32'h19b0694b;
    ram_cell[   42922] = 32'hc84e2424;
    ram_cell[   42923] = 32'h8f7de0ac;
    ram_cell[   42924] = 32'hea6203db;
    ram_cell[   42925] = 32'h73a4050f;
    ram_cell[   42926] = 32'hb3840649;
    ram_cell[   42927] = 32'h78e086b6;
    ram_cell[   42928] = 32'h49530c8f;
    ram_cell[   42929] = 32'h6172b770;
    ram_cell[   42930] = 32'h0ea8bd1d;
    ram_cell[   42931] = 32'h50bce512;
    ram_cell[   42932] = 32'h6274df6c;
    ram_cell[   42933] = 32'he065821d;
    ram_cell[   42934] = 32'h2c483926;
    ram_cell[   42935] = 32'hfc74c209;
    ram_cell[   42936] = 32'h52addb92;
    ram_cell[   42937] = 32'h9b9e12cb;
    ram_cell[   42938] = 32'h77879ad6;
    ram_cell[   42939] = 32'h09f78c85;
    ram_cell[   42940] = 32'ha55e9b1d;
    ram_cell[   42941] = 32'hfe61035c;
    ram_cell[   42942] = 32'h2dc2a1f2;
    ram_cell[   42943] = 32'h1ab485a9;
    ram_cell[   42944] = 32'h1790fb01;
    ram_cell[   42945] = 32'h9962a6f9;
    ram_cell[   42946] = 32'hd596c5dd;
    ram_cell[   42947] = 32'ha9a55de7;
    ram_cell[   42948] = 32'h0ff0e4cf;
    ram_cell[   42949] = 32'hf3b77515;
    ram_cell[   42950] = 32'h2a773dcb;
    ram_cell[   42951] = 32'h0c9a7448;
    ram_cell[   42952] = 32'h06a52cff;
    ram_cell[   42953] = 32'hc6134130;
    ram_cell[   42954] = 32'h1e5026cc;
    ram_cell[   42955] = 32'heea6f43f;
    ram_cell[   42956] = 32'h01c8b72c;
    ram_cell[   42957] = 32'hd65a2d7b;
    ram_cell[   42958] = 32'h19688455;
    ram_cell[   42959] = 32'h602c4183;
    ram_cell[   42960] = 32'hb62bed5a;
    ram_cell[   42961] = 32'h7ac01fb9;
    ram_cell[   42962] = 32'hd80ae314;
    ram_cell[   42963] = 32'h0f5ab915;
    ram_cell[   42964] = 32'hb3e188df;
    ram_cell[   42965] = 32'hdc701700;
    ram_cell[   42966] = 32'h75d51d53;
    ram_cell[   42967] = 32'h25915051;
    ram_cell[   42968] = 32'hf8e4ef60;
    ram_cell[   42969] = 32'h82bbad15;
    ram_cell[   42970] = 32'h1ef6121a;
    ram_cell[   42971] = 32'h98f82018;
    ram_cell[   42972] = 32'he6eb8216;
    ram_cell[   42973] = 32'h503adad0;
    ram_cell[   42974] = 32'h514daa48;
    ram_cell[   42975] = 32'hfad06d2c;
    ram_cell[   42976] = 32'ha0dd15a8;
    ram_cell[   42977] = 32'h06df13e9;
    ram_cell[   42978] = 32'hea63fc1e;
    ram_cell[   42979] = 32'h058fbee4;
    ram_cell[   42980] = 32'h0d7a4e72;
    ram_cell[   42981] = 32'h597b41be;
    ram_cell[   42982] = 32'hbf766abe;
    ram_cell[   42983] = 32'h39015020;
    ram_cell[   42984] = 32'h77a5dea0;
    ram_cell[   42985] = 32'h754c3806;
    ram_cell[   42986] = 32'h0f6018d7;
    ram_cell[   42987] = 32'ha74b77e4;
    ram_cell[   42988] = 32'hccf7a16a;
    ram_cell[   42989] = 32'hf27bd6b2;
    ram_cell[   42990] = 32'h6e0fc564;
    ram_cell[   42991] = 32'h1114dde6;
    ram_cell[   42992] = 32'h8b219fee;
    ram_cell[   42993] = 32'hf5bf5ab3;
    ram_cell[   42994] = 32'hbcce4e36;
    ram_cell[   42995] = 32'hc66b7ef8;
    ram_cell[   42996] = 32'he01b0e86;
    ram_cell[   42997] = 32'h3613d0de;
    ram_cell[   42998] = 32'hfa942b62;
    ram_cell[   42999] = 32'h59647dca;
    ram_cell[   43000] = 32'h714ba0f8;
    ram_cell[   43001] = 32'h8e1ad9e8;
    ram_cell[   43002] = 32'h5abb4d1c;
    ram_cell[   43003] = 32'h0d425be6;
    ram_cell[   43004] = 32'h4e4e739f;
    ram_cell[   43005] = 32'h041f2924;
    ram_cell[   43006] = 32'ha9b361cf;
    ram_cell[   43007] = 32'h327cba07;
    ram_cell[   43008] = 32'h10863fd7;
    ram_cell[   43009] = 32'h7fe0d3b9;
    ram_cell[   43010] = 32'h1ad15adc;
    ram_cell[   43011] = 32'h27c1d7b9;
    ram_cell[   43012] = 32'he3427442;
    ram_cell[   43013] = 32'h229ea7ab;
    ram_cell[   43014] = 32'hb16be639;
    ram_cell[   43015] = 32'hb15013d0;
    ram_cell[   43016] = 32'h32e08fa3;
    ram_cell[   43017] = 32'h4dd31bd8;
    ram_cell[   43018] = 32'he271cfbb;
    ram_cell[   43019] = 32'h40ff1ce7;
    ram_cell[   43020] = 32'h69b217af;
    ram_cell[   43021] = 32'h41d47504;
    ram_cell[   43022] = 32'h0aa2c039;
    ram_cell[   43023] = 32'ha20e3857;
    ram_cell[   43024] = 32'h99f384c2;
    ram_cell[   43025] = 32'h371c41c8;
    ram_cell[   43026] = 32'h461b5ba7;
    ram_cell[   43027] = 32'hbac9232d;
    ram_cell[   43028] = 32'hc510c627;
    ram_cell[   43029] = 32'h14823858;
    ram_cell[   43030] = 32'h711c4386;
    ram_cell[   43031] = 32'h33df38b0;
    ram_cell[   43032] = 32'h3e2b781e;
    ram_cell[   43033] = 32'h1e2d9254;
    ram_cell[   43034] = 32'ha6d17b61;
    ram_cell[   43035] = 32'h7470b9cb;
    ram_cell[   43036] = 32'h9255625e;
    ram_cell[   43037] = 32'h4170d224;
    ram_cell[   43038] = 32'h4d32966e;
    ram_cell[   43039] = 32'h82ee3f51;
    ram_cell[   43040] = 32'h3564e942;
    ram_cell[   43041] = 32'he072569b;
    ram_cell[   43042] = 32'h4b53b09b;
    ram_cell[   43043] = 32'h82930f50;
    ram_cell[   43044] = 32'he2161c06;
    ram_cell[   43045] = 32'hce3ca20a;
    ram_cell[   43046] = 32'h3a07260f;
    ram_cell[   43047] = 32'h2a9cd50c;
    ram_cell[   43048] = 32'h1269cd83;
    ram_cell[   43049] = 32'h10b92e16;
    ram_cell[   43050] = 32'h5816f29c;
    ram_cell[   43051] = 32'h94167d71;
    ram_cell[   43052] = 32'h6a49b3f7;
    ram_cell[   43053] = 32'hf8c7b5b5;
    ram_cell[   43054] = 32'h80e287ed;
    ram_cell[   43055] = 32'h35abaa8d;
    ram_cell[   43056] = 32'h9cb792c5;
    ram_cell[   43057] = 32'h7e0efc2b;
    ram_cell[   43058] = 32'h79f6d36e;
    ram_cell[   43059] = 32'hbbc5fc5f;
    ram_cell[   43060] = 32'h980f7c6a;
    ram_cell[   43061] = 32'hd09f6872;
    ram_cell[   43062] = 32'hc7e074a7;
    ram_cell[   43063] = 32'h0ea5ad30;
    ram_cell[   43064] = 32'h3d5240b8;
    ram_cell[   43065] = 32'hdedb322e;
    ram_cell[   43066] = 32'h6b377888;
    ram_cell[   43067] = 32'h3a483a01;
    ram_cell[   43068] = 32'h15d2a01a;
    ram_cell[   43069] = 32'hd2090612;
    ram_cell[   43070] = 32'hf9b2d068;
    ram_cell[   43071] = 32'heba3d86b;
    ram_cell[   43072] = 32'hf55882f2;
    ram_cell[   43073] = 32'h2a846792;
    ram_cell[   43074] = 32'h771947d1;
    ram_cell[   43075] = 32'h219d66bf;
    ram_cell[   43076] = 32'h908da747;
    ram_cell[   43077] = 32'h333acaf7;
    ram_cell[   43078] = 32'hc830842d;
    ram_cell[   43079] = 32'h23b02332;
    ram_cell[   43080] = 32'h5e012254;
    ram_cell[   43081] = 32'h8dd8b033;
    ram_cell[   43082] = 32'h70fc8572;
    ram_cell[   43083] = 32'h55b15a23;
    ram_cell[   43084] = 32'hb187ea2b;
    ram_cell[   43085] = 32'h79210bde;
    ram_cell[   43086] = 32'h35d3e339;
    ram_cell[   43087] = 32'h42921ea2;
    ram_cell[   43088] = 32'h51e81c6b;
    ram_cell[   43089] = 32'h4f94bec9;
    ram_cell[   43090] = 32'h29b1ace8;
    ram_cell[   43091] = 32'h628cc59e;
    ram_cell[   43092] = 32'hab9a1920;
    ram_cell[   43093] = 32'haa5fa046;
    ram_cell[   43094] = 32'hc591411c;
    ram_cell[   43095] = 32'hdf08a314;
    ram_cell[   43096] = 32'hd9c9c105;
    ram_cell[   43097] = 32'h1f318974;
    ram_cell[   43098] = 32'h0f2c34c3;
    ram_cell[   43099] = 32'h4d1bd1b4;
    ram_cell[   43100] = 32'h3c64f544;
    ram_cell[   43101] = 32'ha2b0a782;
    ram_cell[   43102] = 32'h23ec1457;
    ram_cell[   43103] = 32'h2c0afc62;
    ram_cell[   43104] = 32'h61b8a695;
    ram_cell[   43105] = 32'he4eed06b;
    ram_cell[   43106] = 32'h745d10e4;
    ram_cell[   43107] = 32'h7f864732;
    ram_cell[   43108] = 32'he81e7049;
    ram_cell[   43109] = 32'h5f02f5fc;
    ram_cell[   43110] = 32'h8a50079d;
    ram_cell[   43111] = 32'h5120980d;
    ram_cell[   43112] = 32'h054e20e9;
    ram_cell[   43113] = 32'hb2e9d93b;
    ram_cell[   43114] = 32'ha392384c;
    ram_cell[   43115] = 32'h503a6cb5;
    ram_cell[   43116] = 32'hf3de4744;
    ram_cell[   43117] = 32'hf6b5614e;
    ram_cell[   43118] = 32'hc00e86a5;
    ram_cell[   43119] = 32'hcac8f0f0;
    ram_cell[   43120] = 32'hdc865145;
    ram_cell[   43121] = 32'h67e8284f;
    ram_cell[   43122] = 32'h10fb4f4d;
    ram_cell[   43123] = 32'h504e1a13;
    ram_cell[   43124] = 32'hc1da31ad;
    ram_cell[   43125] = 32'hefc9e1f1;
    ram_cell[   43126] = 32'h90325971;
    ram_cell[   43127] = 32'h852550ed;
    ram_cell[   43128] = 32'h06a4ecfd;
    ram_cell[   43129] = 32'h18271138;
    ram_cell[   43130] = 32'hf1aa8a50;
    ram_cell[   43131] = 32'hd7ce6fd4;
    ram_cell[   43132] = 32'h1a2d2764;
    ram_cell[   43133] = 32'h9e05ba3f;
    ram_cell[   43134] = 32'ha040928d;
    ram_cell[   43135] = 32'h642069e2;
    ram_cell[   43136] = 32'h083ff352;
    ram_cell[   43137] = 32'h4e116c0d;
    ram_cell[   43138] = 32'hbaf3901b;
    ram_cell[   43139] = 32'h21ba16ee;
    ram_cell[   43140] = 32'hda4718ec;
    ram_cell[   43141] = 32'hee1bf206;
    ram_cell[   43142] = 32'h782422f9;
    ram_cell[   43143] = 32'h2e288c9e;
    ram_cell[   43144] = 32'h1f237fbf;
    ram_cell[   43145] = 32'h4309cbcf;
    ram_cell[   43146] = 32'ha96b68b1;
    ram_cell[   43147] = 32'hacd41227;
    ram_cell[   43148] = 32'he9d326ae;
    ram_cell[   43149] = 32'h76499b36;
    ram_cell[   43150] = 32'hd887ae93;
    ram_cell[   43151] = 32'hc54ba390;
    ram_cell[   43152] = 32'h17d5b3d5;
    ram_cell[   43153] = 32'h47dba8d0;
    ram_cell[   43154] = 32'hf3bb2628;
    ram_cell[   43155] = 32'h5cbf63e2;
    ram_cell[   43156] = 32'h5582e1a6;
    ram_cell[   43157] = 32'h97961e32;
    ram_cell[   43158] = 32'h88308bac;
    ram_cell[   43159] = 32'hfaac7b33;
    ram_cell[   43160] = 32'h5788f32b;
    ram_cell[   43161] = 32'h6d4e73d5;
    ram_cell[   43162] = 32'h1b40b721;
    ram_cell[   43163] = 32'h822ed57c;
    ram_cell[   43164] = 32'h02a3ced1;
    ram_cell[   43165] = 32'h7a63149d;
    ram_cell[   43166] = 32'h4f3e2e8a;
    ram_cell[   43167] = 32'h3fcf7395;
    ram_cell[   43168] = 32'hb7cd0994;
    ram_cell[   43169] = 32'h76885f2e;
    ram_cell[   43170] = 32'h2682459c;
    ram_cell[   43171] = 32'hda0bf79c;
    ram_cell[   43172] = 32'hf0561587;
    ram_cell[   43173] = 32'hc5d3f363;
    ram_cell[   43174] = 32'h9c49df3f;
    ram_cell[   43175] = 32'h540fdcaf;
    ram_cell[   43176] = 32'hddc8d6c0;
    ram_cell[   43177] = 32'h26882344;
    ram_cell[   43178] = 32'h78e114b1;
    ram_cell[   43179] = 32'h39fd0d75;
    ram_cell[   43180] = 32'h1469ebd6;
    ram_cell[   43181] = 32'h43fc1967;
    ram_cell[   43182] = 32'h72bb3c61;
    ram_cell[   43183] = 32'h50a7148e;
    ram_cell[   43184] = 32'hc62751c9;
    ram_cell[   43185] = 32'hacdb7a53;
    ram_cell[   43186] = 32'h9a0b35ab;
    ram_cell[   43187] = 32'hc9dfd631;
    ram_cell[   43188] = 32'hdad60ee1;
    ram_cell[   43189] = 32'hffb2a531;
    ram_cell[   43190] = 32'had09feb3;
    ram_cell[   43191] = 32'h151c47b3;
    ram_cell[   43192] = 32'h8f2e5d91;
    ram_cell[   43193] = 32'h9c006014;
    ram_cell[   43194] = 32'h47c0545a;
    ram_cell[   43195] = 32'h8799ad59;
    ram_cell[   43196] = 32'h1f828fb6;
    ram_cell[   43197] = 32'h3e76e563;
    ram_cell[   43198] = 32'he02f9932;
    ram_cell[   43199] = 32'hcd3f0138;
    ram_cell[   43200] = 32'h7ab1b28f;
    ram_cell[   43201] = 32'hcf77d386;
    ram_cell[   43202] = 32'hb4b5c30f;
    ram_cell[   43203] = 32'h3773dad3;
    ram_cell[   43204] = 32'h809c063b;
    ram_cell[   43205] = 32'h1271041f;
    ram_cell[   43206] = 32'h26310706;
    ram_cell[   43207] = 32'hf1c977bb;
    ram_cell[   43208] = 32'ha9260156;
    ram_cell[   43209] = 32'h0d98d81e;
    ram_cell[   43210] = 32'hee41a574;
    ram_cell[   43211] = 32'h7e4de8be;
    ram_cell[   43212] = 32'h27ed6089;
    ram_cell[   43213] = 32'h4cb67cb9;
    ram_cell[   43214] = 32'h3779c097;
    ram_cell[   43215] = 32'hbd4c2246;
    ram_cell[   43216] = 32'hbff6a25e;
    ram_cell[   43217] = 32'h9b39c1f3;
    ram_cell[   43218] = 32'h7222d7f8;
    ram_cell[   43219] = 32'h25f05c80;
    ram_cell[   43220] = 32'he9b20017;
    ram_cell[   43221] = 32'hf489744a;
    ram_cell[   43222] = 32'hcabf790d;
    ram_cell[   43223] = 32'he3ce64af;
    ram_cell[   43224] = 32'ha87a7a41;
    ram_cell[   43225] = 32'hfc29c18c;
    ram_cell[   43226] = 32'h1d2d9562;
    ram_cell[   43227] = 32'hcc4d7938;
    ram_cell[   43228] = 32'haa72748b;
    ram_cell[   43229] = 32'h0f80e1f2;
    ram_cell[   43230] = 32'hb34f5644;
    ram_cell[   43231] = 32'h9ee949df;
    ram_cell[   43232] = 32'hab615cd4;
    ram_cell[   43233] = 32'h89e22168;
    ram_cell[   43234] = 32'h11a3c31e;
    ram_cell[   43235] = 32'h120f4296;
    ram_cell[   43236] = 32'h1d7e2051;
    ram_cell[   43237] = 32'h74d5bfa7;
    ram_cell[   43238] = 32'h78eb22df;
    ram_cell[   43239] = 32'hca5446cb;
    ram_cell[   43240] = 32'hbaf954ee;
    ram_cell[   43241] = 32'h9c65c960;
    ram_cell[   43242] = 32'h8f0cf652;
    ram_cell[   43243] = 32'h228729b4;
    ram_cell[   43244] = 32'h89cba649;
    ram_cell[   43245] = 32'hcee7d7ee;
    ram_cell[   43246] = 32'h04541363;
    ram_cell[   43247] = 32'h29078854;
    ram_cell[   43248] = 32'h31dc6797;
    ram_cell[   43249] = 32'he22e19f9;
    ram_cell[   43250] = 32'h9a46245c;
    ram_cell[   43251] = 32'h50724575;
    ram_cell[   43252] = 32'h0b6fc6d4;
    ram_cell[   43253] = 32'h2a57ecb5;
    ram_cell[   43254] = 32'hc19bf27e;
    ram_cell[   43255] = 32'h0f619b44;
    ram_cell[   43256] = 32'hfc4818c4;
    ram_cell[   43257] = 32'h76907272;
    ram_cell[   43258] = 32'h9d1b8c66;
    ram_cell[   43259] = 32'h855d70db;
    ram_cell[   43260] = 32'h1841c118;
    ram_cell[   43261] = 32'h2ee7fcc0;
    ram_cell[   43262] = 32'he61c36a3;
    ram_cell[   43263] = 32'ha8102f2b;
    ram_cell[   43264] = 32'h4347dd17;
    ram_cell[   43265] = 32'h3d491d90;
    ram_cell[   43266] = 32'h984a049b;
    ram_cell[   43267] = 32'hf7b9a93d;
    ram_cell[   43268] = 32'hd3b88c5b;
    ram_cell[   43269] = 32'ha108efc9;
    ram_cell[   43270] = 32'h84fc1c2c;
    ram_cell[   43271] = 32'h13a20148;
    ram_cell[   43272] = 32'h17ba1413;
    ram_cell[   43273] = 32'h7575b2ba;
    ram_cell[   43274] = 32'h33aae21d;
    ram_cell[   43275] = 32'hd5154406;
    ram_cell[   43276] = 32'he2db74d3;
    ram_cell[   43277] = 32'hee46800a;
    ram_cell[   43278] = 32'haf5855ba;
    ram_cell[   43279] = 32'h84dea5d7;
    ram_cell[   43280] = 32'h3a18476b;
    ram_cell[   43281] = 32'h4f40092d;
    ram_cell[   43282] = 32'h862b9b76;
    ram_cell[   43283] = 32'ha2be5265;
    ram_cell[   43284] = 32'ha9d0ec13;
    ram_cell[   43285] = 32'h64d4f976;
    ram_cell[   43286] = 32'hd7a1c4a7;
    ram_cell[   43287] = 32'h87f275e4;
    ram_cell[   43288] = 32'he89d46dd;
    ram_cell[   43289] = 32'h6ad6f3be;
    ram_cell[   43290] = 32'h6214204a;
    ram_cell[   43291] = 32'hf1fe6818;
    ram_cell[   43292] = 32'h1e750d03;
    ram_cell[   43293] = 32'hb1a50e09;
    ram_cell[   43294] = 32'h65144a32;
    ram_cell[   43295] = 32'h0e860f7d;
    ram_cell[   43296] = 32'h62e36a71;
    ram_cell[   43297] = 32'h258f1c48;
    ram_cell[   43298] = 32'h391a3d45;
    ram_cell[   43299] = 32'hf1ea1822;
    ram_cell[   43300] = 32'h222df8cd;
    ram_cell[   43301] = 32'h9b2478f7;
    ram_cell[   43302] = 32'h561e2785;
    ram_cell[   43303] = 32'h3b4f8117;
    ram_cell[   43304] = 32'hd6059ba4;
    ram_cell[   43305] = 32'h17a2a55e;
    ram_cell[   43306] = 32'h7f18b45a;
    ram_cell[   43307] = 32'h6071d043;
    ram_cell[   43308] = 32'h191d029a;
    ram_cell[   43309] = 32'h85a2f662;
    ram_cell[   43310] = 32'hb25b31ba;
    ram_cell[   43311] = 32'hc8d17d87;
    ram_cell[   43312] = 32'hed76b658;
    ram_cell[   43313] = 32'h596e56fd;
    ram_cell[   43314] = 32'hf12136e0;
    ram_cell[   43315] = 32'hd39f1a0f;
    ram_cell[   43316] = 32'h46ac02d0;
    ram_cell[   43317] = 32'h7ca94299;
    ram_cell[   43318] = 32'haa16c15a;
    ram_cell[   43319] = 32'hef818ccc;
    ram_cell[   43320] = 32'h331f694d;
    ram_cell[   43321] = 32'h903837b1;
    ram_cell[   43322] = 32'h9f819b91;
    ram_cell[   43323] = 32'h4254c8bc;
    ram_cell[   43324] = 32'h84647ab3;
    ram_cell[   43325] = 32'h3cf88cd2;
    ram_cell[   43326] = 32'h898f5d5b;
    ram_cell[   43327] = 32'h130f0c18;
    ram_cell[   43328] = 32'hf737a846;
    ram_cell[   43329] = 32'hfa072baa;
    ram_cell[   43330] = 32'h8a3398b6;
    ram_cell[   43331] = 32'h74b81440;
    ram_cell[   43332] = 32'h95abf4e1;
    ram_cell[   43333] = 32'ha1a4aff3;
    ram_cell[   43334] = 32'h346c83bc;
    ram_cell[   43335] = 32'hc8163f23;
    ram_cell[   43336] = 32'h36499dae;
    ram_cell[   43337] = 32'hce8bc409;
    ram_cell[   43338] = 32'hde2e28cc;
    ram_cell[   43339] = 32'h71ebde53;
    ram_cell[   43340] = 32'h817b61b5;
    ram_cell[   43341] = 32'h868da02a;
    ram_cell[   43342] = 32'h4e3a5fb2;
    ram_cell[   43343] = 32'hb97c3a1c;
    ram_cell[   43344] = 32'h02a49bfb;
    ram_cell[   43345] = 32'h0cc7f9c3;
    ram_cell[   43346] = 32'h54f07c20;
    ram_cell[   43347] = 32'h9806a8b6;
    ram_cell[   43348] = 32'hbb5a6f21;
    ram_cell[   43349] = 32'h84f7416c;
    ram_cell[   43350] = 32'hc1ee1faa;
    ram_cell[   43351] = 32'h5cbfd8ab;
    ram_cell[   43352] = 32'hea75a7f6;
    ram_cell[   43353] = 32'he0be7184;
    ram_cell[   43354] = 32'hb86a76a9;
    ram_cell[   43355] = 32'h215a1731;
    ram_cell[   43356] = 32'h0c5ce42f;
    ram_cell[   43357] = 32'h49e886b7;
    ram_cell[   43358] = 32'h019ca560;
    ram_cell[   43359] = 32'h5da2fc0b;
    ram_cell[   43360] = 32'h6c45b240;
    ram_cell[   43361] = 32'ha4026bd0;
    ram_cell[   43362] = 32'h079005ed;
    ram_cell[   43363] = 32'he663afee;
    ram_cell[   43364] = 32'h5e6aa166;
    ram_cell[   43365] = 32'he78e602d;
    ram_cell[   43366] = 32'h481a5c5d;
    ram_cell[   43367] = 32'hf5ba2d81;
    ram_cell[   43368] = 32'h885181f7;
    ram_cell[   43369] = 32'hbac71e89;
    ram_cell[   43370] = 32'h0e9bdaf5;
    ram_cell[   43371] = 32'hcf6c6630;
    ram_cell[   43372] = 32'hb69da1e8;
    ram_cell[   43373] = 32'h550917a8;
    ram_cell[   43374] = 32'h41ac7162;
    ram_cell[   43375] = 32'h67d1e586;
    ram_cell[   43376] = 32'he72ff5d9;
    ram_cell[   43377] = 32'hc7e85eb2;
    ram_cell[   43378] = 32'h3a2344a4;
    ram_cell[   43379] = 32'h738c3de0;
    ram_cell[   43380] = 32'h1b577fdb;
    ram_cell[   43381] = 32'h2f690e66;
    ram_cell[   43382] = 32'hfdb1f5cc;
    ram_cell[   43383] = 32'h918aef12;
    ram_cell[   43384] = 32'hfc793272;
    ram_cell[   43385] = 32'h404d03d1;
    ram_cell[   43386] = 32'h85d85bc5;
    ram_cell[   43387] = 32'hc5609aee;
    ram_cell[   43388] = 32'hb40b71d6;
    ram_cell[   43389] = 32'h2a4cb163;
    ram_cell[   43390] = 32'hf5473110;
    ram_cell[   43391] = 32'h81a812e7;
    ram_cell[   43392] = 32'hc3ecfd78;
    ram_cell[   43393] = 32'hfae691ef;
    ram_cell[   43394] = 32'h523b9d73;
    ram_cell[   43395] = 32'h743944dc;
    ram_cell[   43396] = 32'h4f016167;
    ram_cell[   43397] = 32'hc2535b45;
    ram_cell[   43398] = 32'h9498a2d2;
    ram_cell[   43399] = 32'h08b02cca;
    ram_cell[   43400] = 32'hf8bccae6;
    ram_cell[   43401] = 32'hcbc52f7a;
    ram_cell[   43402] = 32'hdb867905;
    ram_cell[   43403] = 32'hdd7f0a1b;
    ram_cell[   43404] = 32'h1f5a9bbc;
    ram_cell[   43405] = 32'h18a8c4b1;
    ram_cell[   43406] = 32'h1646aa21;
    ram_cell[   43407] = 32'h10109046;
    ram_cell[   43408] = 32'hf570e2e1;
    ram_cell[   43409] = 32'hb62d3d99;
    ram_cell[   43410] = 32'h36db49c7;
    ram_cell[   43411] = 32'hea0adb17;
    ram_cell[   43412] = 32'h8804283b;
    ram_cell[   43413] = 32'hd449bd35;
    ram_cell[   43414] = 32'h10fba324;
    ram_cell[   43415] = 32'hf0e8f278;
    ram_cell[   43416] = 32'h42f9f262;
    ram_cell[   43417] = 32'h50a08144;
    ram_cell[   43418] = 32'h2e26492f;
    ram_cell[   43419] = 32'h7543a82d;
    ram_cell[   43420] = 32'h2e3e83bb;
    ram_cell[   43421] = 32'hd625a15f;
    ram_cell[   43422] = 32'h33019e92;
    ram_cell[   43423] = 32'h251b6673;
    ram_cell[   43424] = 32'hdf54d737;
    ram_cell[   43425] = 32'hf8c73552;
    ram_cell[   43426] = 32'h1c832333;
    ram_cell[   43427] = 32'had204b42;
    ram_cell[   43428] = 32'h63e77368;
    ram_cell[   43429] = 32'hf936f7d8;
    ram_cell[   43430] = 32'h2fa165be;
    ram_cell[   43431] = 32'h99f0be47;
    ram_cell[   43432] = 32'hc6ae9f70;
    ram_cell[   43433] = 32'h46c5d180;
    ram_cell[   43434] = 32'hfb91e92d;
    ram_cell[   43435] = 32'h53864f59;
    ram_cell[   43436] = 32'hdafcc6d0;
    ram_cell[   43437] = 32'hc9bc90db;
    ram_cell[   43438] = 32'hdf265c23;
    ram_cell[   43439] = 32'hcd93cf5f;
    ram_cell[   43440] = 32'h321e0a23;
    ram_cell[   43441] = 32'h170f9402;
    ram_cell[   43442] = 32'ha9ce2f72;
    ram_cell[   43443] = 32'hc9e42921;
    ram_cell[   43444] = 32'h9a2388fa;
    ram_cell[   43445] = 32'h006e5b2e;
    ram_cell[   43446] = 32'hc5d20b9b;
    ram_cell[   43447] = 32'h5d2ccb21;
    ram_cell[   43448] = 32'h49927b50;
    ram_cell[   43449] = 32'hf0cb6b30;
    ram_cell[   43450] = 32'h17ddb2ba;
    ram_cell[   43451] = 32'hcf1da56a;
    ram_cell[   43452] = 32'h73304d7f;
    ram_cell[   43453] = 32'he163669e;
    ram_cell[   43454] = 32'h1f54cfd6;
    ram_cell[   43455] = 32'h473c7ae2;
    ram_cell[   43456] = 32'h9fc27fe3;
    ram_cell[   43457] = 32'h6be4f3b3;
    ram_cell[   43458] = 32'h990c533b;
    ram_cell[   43459] = 32'h21d2d4cd;
    ram_cell[   43460] = 32'h06ef4dda;
    ram_cell[   43461] = 32'hdb8b81cf;
    ram_cell[   43462] = 32'h21b23713;
    ram_cell[   43463] = 32'h24a384e0;
    ram_cell[   43464] = 32'h2d9f20c1;
    ram_cell[   43465] = 32'h9caaf34e;
    ram_cell[   43466] = 32'h5ccc4a99;
    ram_cell[   43467] = 32'h3c6c6548;
    ram_cell[   43468] = 32'hf85d4fae;
    ram_cell[   43469] = 32'h52a655a9;
    ram_cell[   43470] = 32'h3ec03602;
    ram_cell[   43471] = 32'h0661dd41;
    ram_cell[   43472] = 32'h103da72d;
    ram_cell[   43473] = 32'hb785ceef;
    ram_cell[   43474] = 32'h5a46ca05;
    ram_cell[   43475] = 32'hd1866184;
    ram_cell[   43476] = 32'h562fa13f;
    ram_cell[   43477] = 32'h0a513470;
    ram_cell[   43478] = 32'haefd72ea;
    ram_cell[   43479] = 32'h18a5c7e3;
    ram_cell[   43480] = 32'h475a7941;
    ram_cell[   43481] = 32'hec1e5380;
    ram_cell[   43482] = 32'h40ba3b81;
    ram_cell[   43483] = 32'h540d75ec;
    ram_cell[   43484] = 32'h52624910;
    ram_cell[   43485] = 32'hea6e6001;
    ram_cell[   43486] = 32'h2f3e0d6d;
    ram_cell[   43487] = 32'hbecae6a0;
    ram_cell[   43488] = 32'h793adee1;
    ram_cell[   43489] = 32'h3054d505;
    ram_cell[   43490] = 32'h6cf7f11a;
    ram_cell[   43491] = 32'h41c6aad7;
    ram_cell[   43492] = 32'hbfeb4116;
    ram_cell[   43493] = 32'hf4326135;
    ram_cell[   43494] = 32'h5e651c7f;
    ram_cell[   43495] = 32'hcc481346;
    ram_cell[   43496] = 32'hb36865e7;
    ram_cell[   43497] = 32'h84856826;
    ram_cell[   43498] = 32'h528db93e;
    ram_cell[   43499] = 32'h25211b9f;
    ram_cell[   43500] = 32'hdb7cc6d2;
    ram_cell[   43501] = 32'hc5589770;
    ram_cell[   43502] = 32'hd5f6cb0a;
    ram_cell[   43503] = 32'h606566a8;
    ram_cell[   43504] = 32'h947d3f39;
    ram_cell[   43505] = 32'h5360a779;
    ram_cell[   43506] = 32'he759d022;
    ram_cell[   43507] = 32'h95ca3aef;
    ram_cell[   43508] = 32'h2b3eb0f2;
    ram_cell[   43509] = 32'hc4307aa8;
    ram_cell[   43510] = 32'h16d820fc;
    ram_cell[   43511] = 32'h262becc6;
    ram_cell[   43512] = 32'hda2a236e;
    ram_cell[   43513] = 32'h171cdadb;
    ram_cell[   43514] = 32'hf4aa3297;
    ram_cell[   43515] = 32'h6e403ca8;
    ram_cell[   43516] = 32'h6655fb85;
    ram_cell[   43517] = 32'he599439b;
    ram_cell[   43518] = 32'hfa6ae7ac;
    ram_cell[   43519] = 32'hbb9bc909;
    ram_cell[   43520] = 32'hc7a68c31;
    ram_cell[   43521] = 32'h0d8c2190;
    ram_cell[   43522] = 32'hd50834e5;
    ram_cell[   43523] = 32'hc6085ed4;
    ram_cell[   43524] = 32'h7ea1214f;
    ram_cell[   43525] = 32'ha4f85178;
    ram_cell[   43526] = 32'h494e51c3;
    ram_cell[   43527] = 32'h9f706914;
    ram_cell[   43528] = 32'hc6d6a231;
    ram_cell[   43529] = 32'haa5e72a8;
    ram_cell[   43530] = 32'h2fcef2e3;
    ram_cell[   43531] = 32'h55bc0e6b;
    ram_cell[   43532] = 32'h1218c5a1;
    ram_cell[   43533] = 32'h75e6b753;
    ram_cell[   43534] = 32'h8225dde5;
    ram_cell[   43535] = 32'h93b719c9;
    ram_cell[   43536] = 32'h43fd766a;
    ram_cell[   43537] = 32'h6448f89c;
    ram_cell[   43538] = 32'h41564212;
    ram_cell[   43539] = 32'h94b2083c;
    ram_cell[   43540] = 32'h542288c3;
    ram_cell[   43541] = 32'h0cc2109f;
    ram_cell[   43542] = 32'h9f619f08;
    ram_cell[   43543] = 32'h8415445c;
    ram_cell[   43544] = 32'hcdfb8b27;
    ram_cell[   43545] = 32'hcbd69066;
    ram_cell[   43546] = 32'hafbc4e0d;
    ram_cell[   43547] = 32'h53fd555a;
    ram_cell[   43548] = 32'heccb0849;
    ram_cell[   43549] = 32'h1f32ba2c;
    ram_cell[   43550] = 32'h5d3c760e;
    ram_cell[   43551] = 32'heab8e3b3;
    ram_cell[   43552] = 32'h8f68605f;
    ram_cell[   43553] = 32'hccfc1e3e;
    ram_cell[   43554] = 32'h52fcbe96;
    ram_cell[   43555] = 32'h9f9962b6;
    ram_cell[   43556] = 32'hafb44806;
    ram_cell[   43557] = 32'hdb3aabe6;
    ram_cell[   43558] = 32'h251d69d1;
    ram_cell[   43559] = 32'had36c4f2;
    ram_cell[   43560] = 32'hffc85652;
    ram_cell[   43561] = 32'h3f575116;
    ram_cell[   43562] = 32'h03ba07a7;
    ram_cell[   43563] = 32'hdd5d341a;
    ram_cell[   43564] = 32'h25cabe3a;
    ram_cell[   43565] = 32'he81645f6;
    ram_cell[   43566] = 32'h9c33ddf4;
    ram_cell[   43567] = 32'h42822f94;
    ram_cell[   43568] = 32'h14961819;
    ram_cell[   43569] = 32'ha12556c3;
    ram_cell[   43570] = 32'hbe99cde6;
    ram_cell[   43571] = 32'h3019f6fb;
    ram_cell[   43572] = 32'h1516cc89;
    ram_cell[   43573] = 32'hea16b8ff;
    ram_cell[   43574] = 32'hb489573f;
    ram_cell[   43575] = 32'hfabc55b5;
    ram_cell[   43576] = 32'h1f75718f;
    ram_cell[   43577] = 32'hd90e58d0;
    ram_cell[   43578] = 32'h2a65aa1f;
    ram_cell[   43579] = 32'hbd08a673;
    ram_cell[   43580] = 32'h95132274;
    ram_cell[   43581] = 32'hb7e18176;
    ram_cell[   43582] = 32'h2210635d;
    ram_cell[   43583] = 32'h1e4e851c;
    ram_cell[   43584] = 32'ha1daf14b;
    ram_cell[   43585] = 32'h3ccbb3fe;
    ram_cell[   43586] = 32'h9f75c3b1;
    ram_cell[   43587] = 32'h1e0c8faa;
    ram_cell[   43588] = 32'h37a7fe5b;
    ram_cell[   43589] = 32'h69cae6bd;
    ram_cell[   43590] = 32'h6783803b;
    ram_cell[   43591] = 32'h03adb402;
    ram_cell[   43592] = 32'h8ef82eab;
    ram_cell[   43593] = 32'hdd09731b;
    ram_cell[   43594] = 32'h7c45aa16;
    ram_cell[   43595] = 32'hc0cfe757;
    ram_cell[   43596] = 32'h9ea1208e;
    ram_cell[   43597] = 32'h47cb4137;
    ram_cell[   43598] = 32'ha96b9012;
    ram_cell[   43599] = 32'h607d6210;
    ram_cell[   43600] = 32'h3e0acc40;
    ram_cell[   43601] = 32'h2bdd7da4;
    ram_cell[   43602] = 32'ha6050f82;
    ram_cell[   43603] = 32'hc670048a;
    ram_cell[   43604] = 32'haf948e72;
    ram_cell[   43605] = 32'hd3d9ea1c;
    ram_cell[   43606] = 32'hcb14cff8;
    ram_cell[   43607] = 32'hdedbfd40;
    ram_cell[   43608] = 32'he4bc86a0;
    ram_cell[   43609] = 32'hf7f33e34;
    ram_cell[   43610] = 32'hca63cb26;
    ram_cell[   43611] = 32'h6095074b;
    ram_cell[   43612] = 32'h5d5ef3df;
    ram_cell[   43613] = 32'h28ca1f75;
    ram_cell[   43614] = 32'hd59321b9;
    ram_cell[   43615] = 32'hcd4e30b6;
    ram_cell[   43616] = 32'h9d161036;
    ram_cell[   43617] = 32'h9b527108;
    ram_cell[   43618] = 32'hee0fc7ec;
    ram_cell[   43619] = 32'h4d04916b;
    ram_cell[   43620] = 32'hd31d9126;
    ram_cell[   43621] = 32'hf3a16fef;
    ram_cell[   43622] = 32'h80a10499;
    ram_cell[   43623] = 32'hf83fbf90;
    ram_cell[   43624] = 32'h8326d30c;
    ram_cell[   43625] = 32'hee980e44;
    ram_cell[   43626] = 32'h080f531e;
    ram_cell[   43627] = 32'h4aa3ebec;
    ram_cell[   43628] = 32'h10ee1dbf;
    ram_cell[   43629] = 32'hc90f95cb;
    ram_cell[   43630] = 32'hcf9aec33;
    ram_cell[   43631] = 32'h13739204;
    ram_cell[   43632] = 32'h06790e2d;
    ram_cell[   43633] = 32'haf7f9f2e;
    ram_cell[   43634] = 32'h811e69a2;
    ram_cell[   43635] = 32'hb05c1e59;
    ram_cell[   43636] = 32'h6327a2ef;
    ram_cell[   43637] = 32'h63647e9c;
    ram_cell[   43638] = 32'ha1c5dfe6;
    ram_cell[   43639] = 32'hbd986aa6;
    ram_cell[   43640] = 32'h22922702;
    ram_cell[   43641] = 32'h333d0fd6;
    ram_cell[   43642] = 32'h6e30a496;
    ram_cell[   43643] = 32'h2c327725;
    ram_cell[   43644] = 32'h7be3ad3d;
    ram_cell[   43645] = 32'h4d444be0;
    ram_cell[   43646] = 32'h444ecbeb;
    ram_cell[   43647] = 32'h2f3362d1;
    ram_cell[   43648] = 32'h26f4b8c9;
    ram_cell[   43649] = 32'h6e1c4c9b;
    ram_cell[   43650] = 32'h9028852d;
    ram_cell[   43651] = 32'hb9b52523;
    ram_cell[   43652] = 32'h3775f1f9;
    ram_cell[   43653] = 32'h418a3ad0;
    ram_cell[   43654] = 32'h34392c97;
    ram_cell[   43655] = 32'ha59bc0f7;
    ram_cell[   43656] = 32'hec84e6b2;
    ram_cell[   43657] = 32'he6051173;
    ram_cell[   43658] = 32'h621fe0fa;
    ram_cell[   43659] = 32'h9c0265f1;
    ram_cell[   43660] = 32'h3f4b0e4b;
    ram_cell[   43661] = 32'he090e669;
    ram_cell[   43662] = 32'hf39ebb17;
    ram_cell[   43663] = 32'h2a739c8a;
    ram_cell[   43664] = 32'h3b6d1cc3;
    ram_cell[   43665] = 32'hea661731;
    ram_cell[   43666] = 32'h51297fdd;
    ram_cell[   43667] = 32'h6780f8b1;
    ram_cell[   43668] = 32'h58f83883;
    ram_cell[   43669] = 32'hd0a7fd1b;
    ram_cell[   43670] = 32'h039bca3c;
    ram_cell[   43671] = 32'h4a349a2d;
    ram_cell[   43672] = 32'h5c3b8ec0;
    ram_cell[   43673] = 32'h3ad1729f;
    ram_cell[   43674] = 32'h5de1bfca;
    ram_cell[   43675] = 32'hc107b0ee;
    ram_cell[   43676] = 32'h741d3166;
    ram_cell[   43677] = 32'hd12dd886;
    ram_cell[   43678] = 32'h3efcc6ba;
    ram_cell[   43679] = 32'h9062c682;
    ram_cell[   43680] = 32'h8970439f;
    ram_cell[   43681] = 32'h4ca4c835;
    ram_cell[   43682] = 32'ha8a6504f;
    ram_cell[   43683] = 32'h7e6195dd;
    ram_cell[   43684] = 32'h8d7cc284;
    ram_cell[   43685] = 32'h097ea73c;
    ram_cell[   43686] = 32'hf3257029;
    ram_cell[   43687] = 32'h989f4464;
    ram_cell[   43688] = 32'hb5163515;
    ram_cell[   43689] = 32'h1d62de13;
    ram_cell[   43690] = 32'h659a4777;
    ram_cell[   43691] = 32'h03e197d3;
    ram_cell[   43692] = 32'h3a61fcdd;
    ram_cell[   43693] = 32'h7cae8c62;
    ram_cell[   43694] = 32'h650a1d0f;
    ram_cell[   43695] = 32'h7098e53b;
    ram_cell[   43696] = 32'h183eb200;
    ram_cell[   43697] = 32'h1af77e3f;
    ram_cell[   43698] = 32'hf487d2fb;
    ram_cell[   43699] = 32'hc8016e80;
    ram_cell[   43700] = 32'h04809d6e;
    ram_cell[   43701] = 32'h70985a0f;
    ram_cell[   43702] = 32'hb6930a02;
    ram_cell[   43703] = 32'hb7a0d216;
    ram_cell[   43704] = 32'h1a6fae61;
    ram_cell[   43705] = 32'hb985dcc5;
    ram_cell[   43706] = 32'h6a9a3752;
    ram_cell[   43707] = 32'hb2d01b82;
    ram_cell[   43708] = 32'hd8f465c2;
    ram_cell[   43709] = 32'h918b7bb5;
    ram_cell[   43710] = 32'h9c699c57;
    ram_cell[   43711] = 32'headdbe53;
    ram_cell[   43712] = 32'h197d91d1;
    ram_cell[   43713] = 32'hd3c6374d;
    ram_cell[   43714] = 32'h4ad96309;
    ram_cell[   43715] = 32'hba4fa986;
    ram_cell[   43716] = 32'h3ccb3c64;
    ram_cell[   43717] = 32'h47ac935f;
    ram_cell[   43718] = 32'h93ef0c44;
    ram_cell[   43719] = 32'he7e6cd78;
    ram_cell[   43720] = 32'h60b2e834;
    ram_cell[   43721] = 32'hee04844a;
    ram_cell[   43722] = 32'h5b489b56;
    ram_cell[   43723] = 32'h2739f380;
    ram_cell[   43724] = 32'hb958357d;
    ram_cell[   43725] = 32'h640fcecf;
    ram_cell[   43726] = 32'h4a401134;
    ram_cell[   43727] = 32'ha4b0200a;
    ram_cell[   43728] = 32'h7b0921a5;
    ram_cell[   43729] = 32'he2c9d930;
    ram_cell[   43730] = 32'h68dbba5f;
    ram_cell[   43731] = 32'h442e0dd5;
    ram_cell[   43732] = 32'h2f3bb2eb;
    ram_cell[   43733] = 32'hdcf549b9;
    ram_cell[   43734] = 32'h9e188bdb;
    ram_cell[   43735] = 32'h34e4a306;
    ram_cell[   43736] = 32'hc0ea765d;
    ram_cell[   43737] = 32'hf89b4622;
    ram_cell[   43738] = 32'h87aade13;
    ram_cell[   43739] = 32'h17de961e;
    ram_cell[   43740] = 32'h425e66c9;
    ram_cell[   43741] = 32'h1bb42184;
    ram_cell[   43742] = 32'h925fbceb;
    ram_cell[   43743] = 32'h6bd6a4f0;
    ram_cell[   43744] = 32'h222dd4e2;
    ram_cell[   43745] = 32'hebc4debb;
    ram_cell[   43746] = 32'h7fab79bb;
    ram_cell[   43747] = 32'h61b36891;
    ram_cell[   43748] = 32'h6aa3b28b;
    ram_cell[   43749] = 32'h6c800a94;
    ram_cell[   43750] = 32'hac3ed64c;
    ram_cell[   43751] = 32'h4404906f;
    ram_cell[   43752] = 32'hedf6118d;
    ram_cell[   43753] = 32'hf1c731d2;
    ram_cell[   43754] = 32'h53ba3706;
    ram_cell[   43755] = 32'hea405263;
    ram_cell[   43756] = 32'hacb005da;
    ram_cell[   43757] = 32'h6d22fc69;
    ram_cell[   43758] = 32'h7dd7b443;
    ram_cell[   43759] = 32'h137e7ca3;
    ram_cell[   43760] = 32'h37b63aec;
    ram_cell[   43761] = 32'hf73f9204;
    ram_cell[   43762] = 32'h3ec492cc;
    ram_cell[   43763] = 32'hf54c7863;
    ram_cell[   43764] = 32'h639dee0b;
    ram_cell[   43765] = 32'hb150756b;
    ram_cell[   43766] = 32'h36f8604d;
    ram_cell[   43767] = 32'h0b036a2d;
    ram_cell[   43768] = 32'h6848070e;
    ram_cell[   43769] = 32'hb55fef0d;
    ram_cell[   43770] = 32'hde0ba834;
    ram_cell[   43771] = 32'h6169b598;
    ram_cell[   43772] = 32'h459373fd;
    ram_cell[   43773] = 32'h65636a7b;
    ram_cell[   43774] = 32'h6f519fb6;
    ram_cell[   43775] = 32'h7abbd213;
    ram_cell[   43776] = 32'h57840f44;
    ram_cell[   43777] = 32'h19eac9f0;
    ram_cell[   43778] = 32'h17c851ce;
    ram_cell[   43779] = 32'h771b80d0;
    ram_cell[   43780] = 32'hcdb8c4cc;
    ram_cell[   43781] = 32'ha7c49175;
    ram_cell[   43782] = 32'h675a416b;
    ram_cell[   43783] = 32'hdd0f6b50;
    ram_cell[   43784] = 32'he98b0a94;
    ram_cell[   43785] = 32'h74f71a1f;
    ram_cell[   43786] = 32'hb8fd7f8a;
    ram_cell[   43787] = 32'h3c122fcf;
    ram_cell[   43788] = 32'hcc1d7136;
    ram_cell[   43789] = 32'h09029043;
    ram_cell[   43790] = 32'hbf63c8d1;
    ram_cell[   43791] = 32'h3a344d45;
    ram_cell[   43792] = 32'hb2d9b098;
    ram_cell[   43793] = 32'h40b9ac86;
    ram_cell[   43794] = 32'h13052baf;
    ram_cell[   43795] = 32'h7957bd48;
    ram_cell[   43796] = 32'h254d6b72;
    ram_cell[   43797] = 32'h67462f45;
    ram_cell[   43798] = 32'h61a647a2;
    ram_cell[   43799] = 32'h44734e54;
    ram_cell[   43800] = 32'h006234df;
    ram_cell[   43801] = 32'h540389ad;
    ram_cell[   43802] = 32'hc214b7e3;
    ram_cell[   43803] = 32'hc540837c;
    ram_cell[   43804] = 32'h93576eda;
    ram_cell[   43805] = 32'h721454de;
    ram_cell[   43806] = 32'h00930649;
    ram_cell[   43807] = 32'h2a073908;
    ram_cell[   43808] = 32'h01aa5e7c;
    ram_cell[   43809] = 32'h0b4138dd;
    ram_cell[   43810] = 32'h5ec61209;
    ram_cell[   43811] = 32'h650c2d32;
    ram_cell[   43812] = 32'h4507dffe;
    ram_cell[   43813] = 32'h0079ab1b;
    ram_cell[   43814] = 32'h3c881141;
    ram_cell[   43815] = 32'h7dc4a6bd;
    ram_cell[   43816] = 32'hdee05762;
    ram_cell[   43817] = 32'hb6c16916;
    ram_cell[   43818] = 32'h2ac08cb9;
    ram_cell[   43819] = 32'hb2bf2c23;
    ram_cell[   43820] = 32'h45f02f4b;
    ram_cell[   43821] = 32'h138d2e77;
    ram_cell[   43822] = 32'h20fb8575;
    ram_cell[   43823] = 32'h09031802;
    ram_cell[   43824] = 32'h20eada2e;
    ram_cell[   43825] = 32'h65ce40f6;
    ram_cell[   43826] = 32'he2dac10d;
    ram_cell[   43827] = 32'hb1e4c570;
    ram_cell[   43828] = 32'h9f257cef;
    ram_cell[   43829] = 32'h01aaf199;
    ram_cell[   43830] = 32'he7f6d7bc;
    ram_cell[   43831] = 32'h7075df3d;
    ram_cell[   43832] = 32'h8cd678e0;
    ram_cell[   43833] = 32'h28266c21;
    ram_cell[   43834] = 32'h1dc01182;
    ram_cell[   43835] = 32'h0a17ae0a;
    ram_cell[   43836] = 32'h7121d5e1;
    ram_cell[   43837] = 32'h9db5f7c3;
    ram_cell[   43838] = 32'h5fb9172d;
    ram_cell[   43839] = 32'hb46f83f1;
    ram_cell[   43840] = 32'h17df990b;
    ram_cell[   43841] = 32'h446429c8;
    ram_cell[   43842] = 32'hfe227d99;
    ram_cell[   43843] = 32'h67d23da8;
    ram_cell[   43844] = 32'h7253f0ed;
    ram_cell[   43845] = 32'h79f60ca2;
    ram_cell[   43846] = 32'h8e7d1b89;
    ram_cell[   43847] = 32'hba8643a8;
    ram_cell[   43848] = 32'h094d1156;
    ram_cell[   43849] = 32'h5b2ee73f;
    ram_cell[   43850] = 32'h301ed2c2;
    ram_cell[   43851] = 32'hfce8f4c2;
    ram_cell[   43852] = 32'h208f2901;
    ram_cell[   43853] = 32'h76b4a040;
    ram_cell[   43854] = 32'hd4113add;
    ram_cell[   43855] = 32'h0b9fea77;
    ram_cell[   43856] = 32'h2e1ee9ab;
    ram_cell[   43857] = 32'h1e78c42f;
    ram_cell[   43858] = 32'h19f589cf;
    ram_cell[   43859] = 32'hbfa13674;
    ram_cell[   43860] = 32'hc531e923;
    ram_cell[   43861] = 32'h39ff93ca;
    ram_cell[   43862] = 32'h3dd6fdab;
    ram_cell[   43863] = 32'h212fc00c;
    ram_cell[   43864] = 32'h5e682f4a;
    ram_cell[   43865] = 32'h12f608f4;
    ram_cell[   43866] = 32'h0214959f;
    ram_cell[   43867] = 32'hd3eafd36;
    ram_cell[   43868] = 32'hfebf4363;
    ram_cell[   43869] = 32'h583d90e5;
    ram_cell[   43870] = 32'h5511f659;
    ram_cell[   43871] = 32'h29252748;
    ram_cell[   43872] = 32'h2c28b537;
    ram_cell[   43873] = 32'h25eff54f;
    ram_cell[   43874] = 32'h51851a77;
    ram_cell[   43875] = 32'h01d8462f;
    ram_cell[   43876] = 32'he48e79ff;
    ram_cell[   43877] = 32'hb632f220;
    ram_cell[   43878] = 32'h24369ada;
    ram_cell[   43879] = 32'hafe67856;
    ram_cell[   43880] = 32'h788e598e;
    ram_cell[   43881] = 32'h9913f228;
    ram_cell[   43882] = 32'h57aab07d;
    ram_cell[   43883] = 32'h770e29e1;
    ram_cell[   43884] = 32'h6081064d;
    ram_cell[   43885] = 32'h7881076f;
    ram_cell[   43886] = 32'h31a4c380;
    ram_cell[   43887] = 32'h4fd4f750;
    ram_cell[   43888] = 32'hc180bf5d;
    ram_cell[   43889] = 32'h82eaaac1;
    ram_cell[   43890] = 32'h5c762f3d;
    ram_cell[   43891] = 32'h7993babf;
    ram_cell[   43892] = 32'h294fee06;
    ram_cell[   43893] = 32'hccf261b7;
    ram_cell[   43894] = 32'h41200fb2;
    ram_cell[   43895] = 32'hed32ea19;
    ram_cell[   43896] = 32'h427f7b02;
    ram_cell[   43897] = 32'h4e29d155;
    ram_cell[   43898] = 32'h8b8037f1;
    ram_cell[   43899] = 32'h3a23cbef;
    ram_cell[   43900] = 32'haacbed1b;
    ram_cell[   43901] = 32'h731175b9;
    ram_cell[   43902] = 32'h41e18d19;
    ram_cell[   43903] = 32'h6dada7fe;
    ram_cell[   43904] = 32'ha6040302;
    ram_cell[   43905] = 32'h6fde1a0b;
    ram_cell[   43906] = 32'h9fa05f37;
    ram_cell[   43907] = 32'hb3ba90a1;
    ram_cell[   43908] = 32'heb6b55ae;
    ram_cell[   43909] = 32'h60e4f13b;
    ram_cell[   43910] = 32'hce78c490;
    ram_cell[   43911] = 32'h2f2e38e1;
    ram_cell[   43912] = 32'ha1300560;
    ram_cell[   43913] = 32'h4d034c4a;
    ram_cell[   43914] = 32'h71864bc0;
    ram_cell[   43915] = 32'hd25c053b;
    ram_cell[   43916] = 32'hd029e2aa;
    ram_cell[   43917] = 32'hebe905d6;
    ram_cell[   43918] = 32'ha835182e;
    ram_cell[   43919] = 32'h20f1cae5;
    ram_cell[   43920] = 32'hef362846;
    ram_cell[   43921] = 32'h92e27805;
    ram_cell[   43922] = 32'heb67512a;
    ram_cell[   43923] = 32'hc9857432;
    ram_cell[   43924] = 32'ha6019084;
    ram_cell[   43925] = 32'ha1b00841;
    ram_cell[   43926] = 32'h060c804e;
    ram_cell[   43927] = 32'h2ecd7108;
    ram_cell[   43928] = 32'h37e9ea77;
    ram_cell[   43929] = 32'h689a4f88;
    ram_cell[   43930] = 32'h6ae613eb;
    ram_cell[   43931] = 32'h15d524ee;
    ram_cell[   43932] = 32'h6226b5c4;
    ram_cell[   43933] = 32'hcd75e055;
    ram_cell[   43934] = 32'hc4c0eb81;
    ram_cell[   43935] = 32'hfa0850eb;
    ram_cell[   43936] = 32'h7ce646f7;
    ram_cell[   43937] = 32'h63a2d628;
    ram_cell[   43938] = 32'h4557a6ff;
    ram_cell[   43939] = 32'h4131d2df;
    ram_cell[   43940] = 32'h74c9a244;
    ram_cell[   43941] = 32'h07d24c8c;
    ram_cell[   43942] = 32'h31a23f08;
    ram_cell[   43943] = 32'h391ae122;
    ram_cell[   43944] = 32'h02514471;
    ram_cell[   43945] = 32'h6782032d;
    ram_cell[   43946] = 32'hc7e8afb5;
    ram_cell[   43947] = 32'h8d221cc9;
    ram_cell[   43948] = 32'hd4c069a5;
    ram_cell[   43949] = 32'h41a2fce2;
    ram_cell[   43950] = 32'h8b4bc134;
    ram_cell[   43951] = 32'h01bd0491;
    ram_cell[   43952] = 32'hf07c62fe;
    ram_cell[   43953] = 32'hd6ebb1ae;
    ram_cell[   43954] = 32'h5b69fe18;
    ram_cell[   43955] = 32'h8e5afb9b;
    ram_cell[   43956] = 32'h7d4b861b;
    ram_cell[   43957] = 32'h4216bf78;
    ram_cell[   43958] = 32'h3712c6db;
    ram_cell[   43959] = 32'h3a0df547;
    ram_cell[   43960] = 32'h8d7dbe8f;
    ram_cell[   43961] = 32'h14226423;
    ram_cell[   43962] = 32'h2630cb42;
    ram_cell[   43963] = 32'h0d686213;
    ram_cell[   43964] = 32'hf8b0bc05;
    ram_cell[   43965] = 32'h500f2023;
    ram_cell[   43966] = 32'h551aa47b;
    ram_cell[   43967] = 32'h3d82052b;
    ram_cell[   43968] = 32'h71806b48;
    ram_cell[   43969] = 32'hb06c4a78;
    ram_cell[   43970] = 32'h61adba22;
    ram_cell[   43971] = 32'h79105edf;
    ram_cell[   43972] = 32'hd2d7f290;
    ram_cell[   43973] = 32'hcf0ea2db;
    ram_cell[   43974] = 32'h1840ec65;
    ram_cell[   43975] = 32'hea9c790b;
    ram_cell[   43976] = 32'h1fc0978c;
    ram_cell[   43977] = 32'hd38665b0;
    ram_cell[   43978] = 32'hd03527f6;
    ram_cell[   43979] = 32'hf892ce10;
    ram_cell[   43980] = 32'h64057819;
    ram_cell[   43981] = 32'h0106a4a9;
    ram_cell[   43982] = 32'hb5465eef;
    ram_cell[   43983] = 32'h533585e4;
    ram_cell[   43984] = 32'hc232bf06;
    ram_cell[   43985] = 32'hd9b12870;
    ram_cell[   43986] = 32'h2e427a69;
    ram_cell[   43987] = 32'h3a7c5bcb;
    ram_cell[   43988] = 32'hd4a9643b;
    ram_cell[   43989] = 32'hc1817a0c;
    ram_cell[   43990] = 32'hb06334c7;
    ram_cell[   43991] = 32'h1697be40;
    ram_cell[   43992] = 32'h155722d3;
    ram_cell[   43993] = 32'h480c89df;
    ram_cell[   43994] = 32'h622ddf3a;
    ram_cell[   43995] = 32'hfeb2993f;
    ram_cell[   43996] = 32'he95158a6;
    ram_cell[   43997] = 32'hf1466a26;
    ram_cell[   43998] = 32'h8ab79b2b;
    ram_cell[   43999] = 32'h092a1f0d;
    ram_cell[   44000] = 32'h81ac0cde;
    ram_cell[   44001] = 32'h6b3e45db;
    ram_cell[   44002] = 32'h85936c90;
    ram_cell[   44003] = 32'h66131dbd;
    ram_cell[   44004] = 32'h9d510d0f;
    ram_cell[   44005] = 32'h019b896b;
    ram_cell[   44006] = 32'h05aa34bd;
    ram_cell[   44007] = 32'hf078b89d;
    ram_cell[   44008] = 32'h43ca3daf;
    ram_cell[   44009] = 32'h7ed097ef;
    ram_cell[   44010] = 32'h1e245ecf;
    ram_cell[   44011] = 32'hbbf01ca9;
    ram_cell[   44012] = 32'h0a5ac6ea;
    ram_cell[   44013] = 32'h1dd15b97;
    ram_cell[   44014] = 32'h98857203;
    ram_cell[   44015] = 32'h81169e08;
    ram_cell[   44016] = 32'hf1e25247;
    ram_cell[   44017] = 32'h98cf399a;
    ram_cell[   44018] = 32'hfbc63a53;
    ram_cell[   44019] = 32'h49419350;
    ram_cell[   44020] = 32'hd62878f2;
    ram_cell[   44021] = 32'h95695200;
    ram_cell[   44022] = 32'h931a369b;
    ram_cell[   44023] = 32'h371d9eac;
    ram_cell[   44024] = 32'h2b8fadfe;
    ram_cell[   44025] = 32'h7d395b55;
    ram_cell[   44026] = 32'hb296b137;
    ram_cell[   44027] = 32'h2e829090;
    ram_cell[   44028] = 32'h11c639c6;
    ram_cell[   44029] = 32'h0ae9f0c0;
    ram_cell[   44030] = 32'h6157fa31;
    ram_cell[   44031] = 32'ha930f265;
    ram_cell[   44032] = 32'h4a77c099;
    ram_cell[   44033] = 32'h6e822e4b;
    ram_cell[   44034] = 32'hc905532b;
    ram_cell[   44035] = 32'h19634d55;
    ram_cell[   44036] = 32'h1b6a94b1;
    ram_cell[   44037] = 32'h6d0dde93;
    ram_cell[   44038] = 32'h079dc5bc;
    ram_cell[   44039] = 32'h40a96441;
    ram_cell[   44040] = 32'h519215e6;
    ram_cell[   44041] = 32'h717480cc;
    ram_cell[   44042] = 32'he8b6bea8;
    ram_cell[   44043] = 32'h68ec6afd;
    ram_cell[   44044] = 32'h05fcf3b6;
    ram_cell[   44045] = 32'h33fd446f;
    ram_cell[   44046] = 32'h869a01b9;
    ram_cell[   44047] = 32'hebd7b9ba;
    ram_cell[   44048] = 32'h16f48d7b;
    ram_cell[   44049] = 32'h4ed6f19b;
    ram_cell[   44050] = 32'h088bad8a;
    ram_cell[   44051] = 32'hb79a6d37;
    ram_cell[   44052] = 32'h23377a41;
    ram_cell[   44053] = 32'hb2b26435;
    ram_cell[   44054] = 32'h96d8b96c;
    ram_cell[   44055] = 32'h0f33f78a;
    ram_cell[   44056] = 32'hb0fa630e;
    ram_cell[   44057] = 32'h6a45d070;
    ram_cell[   44058] = 32'h92f1780f;
    ram_cell[   44059] = 32'hb159f79e;
    ram_cell[   44060] = 32'ha5c16649;
    ram_cell[   44061] = 32'h25ff17ca;
    ram_cell[   44062] = 32'h5d88ecf2;
    ram_cell[   44063] = 32'h54d37ed0;
    ram_cell[   44064] = 32'hae7cf7b2;
    ram_cell[   44065] = 32'h4115007c;
    ram_cell[   44066] = 32'h9ef3a3e2;
    ram_cell[   44067] = 32'he729bd83;
    ram_cell[   44068] = 32'h99100d39;
    ram_cell[   44069] = 32'hfc523e4c;
    ram_cell[   44070] = 32'h2c070e7b;
    ram_cell[   44071] = 32'h72d2e826;
    ram_cell[   44072] = 32'had19ae6b;
    ram_cell[   44073] = 32'h0d25c981;
    ram_cell[   44074] = 32'h2cd64106;
    ram_cell[   44075] = 32'h6a850b9b;
    ram_cell[   44076] = 32'h32002c35;
    ram_cell[   44077] = 32'h522d276c;
    ram_cell[   44078] = 32'h53fbe7ac;
    ram_cell[   44079] = 32'h7e3d1f56;
    ram_cell[   44080] = 32'hd7ae70fd;
    ram_cell[   44081] = 32'h59703f7f;
    ram_cell[   44082] = 32'h084653bd;
    ram_cell[   44083] = 32'h49da978a;
    ram_cell[   44084] = 32'hb72519dc;
    ram_cell[   44085] = 32'h43acb78c;
    ram_cell[   44086] = 32'h42177185;
    ram_cell[   44087] = 32'h2ca23e6d;
    ram_cell[   44088] = 32'h0f066ccd;
    ram_cell[   44089] = 32'h28c40564;
    ram_cell[   44090] = 32'hdee3bff6;
    ram_cell[   44091] = 32'h92b19bd0;
    ram_cell[   44092] = 32'h1c8b8d4a;
    ram_cell[   44093] = 32'hcb9977c5;
    ram_cell[   44094] = 32'h1026ad7b;
    ram_cell[   44095] = 32'ha0ed8fcf;
    ram_cell[   44096] = 32'h4e08ddaf;
    ram_cell[   44097] = 32'hecd3bd7b;
    ram_cell[   44098] = 32'hb0931382;
    ram_cell[   44099] = 32'ha6634721;
    ram_cell[   44100] = 32'h3322f7b6;
    ram_cell[   44101] = 32'hd0c6bebb;
    ram_cell[   44102] = 32'h441bb111;
    ram_cell[   44103] = 32'h269b1bfc;
    ram_cell[   44104] = 32'haf05f129;
    ram_cell[   44105] = 32'ha53402de;
    ram_cell[   44106] = 32'h622f8295;
    ram_cell[   44107] = 32'h98e87e9f;
    ram_cell[   44108] = 32'h0c745144;
    ram_cell[   44109] = 32'h27218a10;
    ram_cell[   44110] = 32'hee8b12c1;
    ram_cell[   44111] = 32'h432c5b45;
    ram_cell[   44112] = 32'hd8d16297;
    ram_cell[   44113] = 32'h15488ab6;
    ram_cell[   44114] = 32'hc354a3ed;
    ram_cell[   44115] = 32'ha65cb5cd;
    ram_cell[   44116] = 32'h77fe701c;
    ram_cell[   44117] = 32'h222a9dbb;
    ram_cell[   44118] = 32'he4dfb4de;
    ram_cell[   44119] = 32'hc3a03840;
    ram_cell[   44120] = 32'h46542b57;
    ram_cell[   44121] = 32'ha1148e9c;
    ram_cell[   44122] = 32'h0b1516ed;
    ram_cell[   44123] = 32'h553944e2;
    ram_cell[   44124] = 32'hea547a9c;
    ram_cell[   44125] = 32'h4cf30a46;
    ram_cell[   44126] = 32'h7f979fbf;
    ram_cell[   44127] = 32'hcf47d8d1;
    ram_cell[   44128] = 32'hfcd0ccf4;
    ram_cell[   44129] = 32'hc42bb23b;
    ram_cell[   44130] = 32'h45476672;
    ram_cell[   44131] = 32'ha7338e1d;
    ram_cell[   44132] = 32'h03d0828f;
    ram_cell[   44133] = 32'hf6df1c55;
    ram_cell[   44134] = 32'h25c4d1b5;
    ram_cell[   44135] = 32'hb2a143e1;
    ram_cell[   44136] = 32'hfbe285c3;
    ram_cell[   44137] = 32'h781c61dd;
    ram_cell[   44138] = 32'h06a35250;
    ram_cell[   44139] = 32'h6428fa0c;
    ram_cell[   44140] = 32'h4ab7b814;
    ram_cell[   44141] = 32'h632d4a5f;
    ram_cell[   44142] = 32'h8ba9f502;
    ram_cell[   44143] = 32'hbc345031;
    ram_cell[   44144] = 32'h21edaeed;
    ram_cell[   44145] = 32'hee2dc5e9;
    ram_cell[   44146] = 32'h5e45ca2d;
    ram_cell[   44147] = 32'hd1dab4ba;
    ram_cell[   44148] = 32'h0bc64c89;
    ram_cell[   44149] = 32'h98de5688;
    ram_cell[   44150] = 32'h10de683c;
    ram_cell[   44151] = 32'h3c9f1e70;
    ram_cell[   44152] = 32'h78a1c7d0;
    ram_cell[   44153] = 32'hb453f99a;
    ram_cell[   44154] = 32'h07d2b6de;
    ram_cell[   44155] = 32'hc96f69f5;
    ram_cell[   44156] = 32'h3a629566;
    ram_cell[   44157] = 32'h8caf5df8;
    ram_cell[   44158] = 32'h1c98ba87;
    ram_cell[   44159] = 32'hda4415be;
    ram_cell[   44160] = 32'h32357303;
    ram_cell[   44161] = 32'h709d3bd0;
    ram_cell[   44162] = 32'h2846329a;
    ram_cell[   44163] = 32'hb246c80c;
    ram_cell[   44164] = 32'h8530532d;
    ram_cell[   44165] = 32'hd56045f6;
    ram_cell[   44166] = 32'h5d734d34;
    ram_cell[   44167] = 32'h21116e95;
    ram_cell[   44168] = 32'hbe6817d3;
    ram_cell[   44169] = 32'h960b53dc;
    ram_cell[   44170] = 32'hc4db332b;
    ram_cell[   44171] = 32'h1c26ae29;
    ram_cell[   44172] = 32'h398f0333;
    ram_cell[   44173] = 32'h629257f4;
    ram_cell[   44174] = 32'h86120be4;
    ram_cell[   44175] = 32'h4f819215;
    ram_cell[   44176] = 32'hcbaccbff;
    ram_cell[   44177] = 32'h2e321f1a;
    ram_cell[   44178] = 32'h3dc727b7;
    ram_cell[   44179] = 32'hbd9156ef;
    ram_cell[   44180] = 32'h0a15f7c6;
    ram_cell[   44181] = 32'hd6a699e1;
    ram_cell[   44182] = 32'h53dc15ed;
    ram_cell[   44183] = 32'h52ecfc8b;
    ram_cell[   44184] = 32'h801332de;
    ram_cell[   44185] = 32'hb625bd93;
    ram_cell[   44186] = 32'h1c72c323;
    ram_cell[   44187] = 32'h1a18b853;
    ram_cell[   44188] = 32'h7a84f572;
    ram_cell[   44189] = 32'hf5ded012;
    ram_cell[   44190] = 32'h6158100d;
    ram_cell[   44191] = 32'hd49e4623;
    ram_cell[   44192] = 32'h0141bd3f;
    ram_cell[   44193] = 32'h8926b75f;
    ram_cell[   44194] = 32'h846e794c;
    ram_cell[   44195] = 32'h064ac71c;
    ram_cell[   44196] = 32'hff5250ee;
    ram_cell[   44197] = 32'hb23c8086;
    ram_cell[   44198] = 32'hfd04846e;
    ram_cell[   44199] = 32'h8468132a;
    ram_cell[   44200] = 32'h1aca42f7;
    ram_cell[   44201] = 32'h00b21dae;
    ram_cell[   44202] = 32'h1efb4427;
    ram_cell[   44203] = 32'h2ba8dda0;
    ram_cell[   44204] = 32'h259309be;
    ram_cell[   44205] = 32'hf98daeb9;
    ram_cell[   44206] = 32'h0a276b03;
    ram_cell[   44207] = 32'h86cda852;
    ram_cell[   44208] = 32'h51dfca01;
    ram_cell[   44209] = 32'hb2823a35;
    ram_cell[   44210] = 32'h731a02ed;
    ram_cell[   44211] = 32'h8a01a99b;
    ram_cell[   44212] = 32'hfdc90778;
    ram_cell[   44213] = 32'h5f40b470;
    ram_cell[   44214] = 32'haa610d98;
    ram_cell[   44215] = 32'h75364a5f;
    ram_cell[   44216] = 32'hc51f2f00;
    ram_cell[   44217] = 32'hcc7aa864;
    ram_cell[   44218] = 32'h5e4971cc;
    ram_cell[   44219] = 32'had028afc;
    ram_cell[   44220] = 32'h438eb0a5;
    ram_cell[   44221] = 32'hdbc223f7;
    ram_cell[   44222] = 32'h60b0db00;
    ram_cell[   44223] = 32'h55c9fa4c;
    ram_cell[   44224] = 32'h74c4b60e;
    ram_cell[   44225] = 32'h81d31128;
    ram_cell[   44226] = 32'h6a39f8af;
    ram_cell[   44227] = 32'h53b31488;
    ram_cell[   44228] = 32'had5aadc5;
    ram_cell[   44229] = 32'h9f83a5cd;
    ram_cell[   44230] = 32'h1524112a;
    ram_cell[   44231] = 32'hf2388245;
    ram_cell[   44232] = 32'h6b45de4b;
    ram_cell[   44233] = 32'hfee8aef0;
    ram_cell[   44234] = 32'ha4759816;
    ram_cell[   44235] = 32'hc1b914bf;
    ram_cell[   44236] = 32'h8ffee6ab;
    ram_cell[   44237] = 32'hc1d6918e;
    ram_cell[   44238] = 32'h23cf102f;
    ram_cell[   44239] = 32'h6a56e32a;
    ram_cell[   44240] = 32'h499d6332;
    ram_cell[   44241] = 32'hb4e6e301;
    ram_cell[   44242] = 32'hf41e9c0f;
    ram_cell[   44243] = 32'h28c14722;
    ram_cell[   44244] = 32'hb33dc968;
    ram_cell[   44245] = 32'h455da74e;
    ram_cell[   44246] = 32'h17262cfc;
    ram_cell[   44247] = 32'hdb913684;
    ram_cell[   44248] = 32'h9c425af9;
    ram_cell[   44249] = 32'h571787cd;
    ram_cell[   44250] = 32'h38ba42b3;
    ram_cell[   44251] = 32'hf57ca540;
    ram_cell[   44252] = 32'h165c49f5;
    ram_cell[   44253] = 32'h87128c36;
    ram_cell[   44254] = 32'hfe142fcd;
    ram_cell[   44255] = 32'h41220d3e;
    ram_cell[   44256] = 32'hce81c060;
    ram_cell[   44257] = 32'hca5e7454;
    ram_cell[   44258] = 32'ha6982afe;
    ram_cell[   44259] = 32'had8c1ee7;
    ram_cell[   44260] = 32'h1957f9f4;
    ram_cell[   44261] = 32'h8b23c73a;
    ram_cell[   44262] = 32'h203aa4a9;
    ram_cell[   44263] = 32'h5d0e2947;
    ram_cell[   44264] = 32'hfd4bac72;
    ram_cell[   44265] = 32'h4a819441;
    ram_cell[   44266] = 32'h7886c00e;
    ram_cell[   44267] = 32'h80dbd2ef;
    ram_cell[   44268] = 32'hdc027449;
    ram_cell[   44269] = 32'h1a6e7880;
    ram_cell[   44270] = 32'h0225030a;
    ram_cell[   44271] = 32'hae6e2018;
    ram_cell[   44272] = 32'hc812e922;
    ram_cell[   44273] = 32'hd565da7c;
    ram_cell[   44274] = 32'hc5d90c96;
    ram_cell[   44275] = 32'h00ec5b42;
    ram_cell[   44276] = 32'hd1686d68;
    ram_cell[   44277] = 32'hf908edf1;
    ram_cell[   44278] = 32'hb42ecbbe;
    ram_cell[   44279] = 32'h00a5e4fe;
    ram_cell[   44280] = 32'hc2f4a781;
    ram_cell[   44281] = 32'h4f161966;
    ram_cell[   44282] = 32'h2ddd3a66;
    ram_cell[   44283] = 32'hba83b364;
    ram_cell[   44284] = 32'hdd348514;
    ram_cell[   44285] = 32'hca520828;
    ram_cell[   44286] = 32'h05d2879f;
    ram_cell[   44287] = 32'h6ce2e406;
    ram_cell[   44288] = 32'h6d5a8dfa;
    ram_cell[   44289] = 32'h93f97ca3;
    ram_cell[   44290] = 32'h975a7dd3;
    ram_cell[   44291] = 32'h31fad9fe;
    ram_cell[   44292] = 32'he62dd01b;
    ram_cell[   44293] = 32'hba3d9d0b;
    ram_cell[   44294] = 32'h28c01609;
    ram_cell[   44295] = 32'ha5873c89;
    ram_cell[   44296] = 32'h158b8bf8;
    ram_cell[   44297] = 32'h6c9d85bb;
    ram_cell[   44298] = 32'h417acedc;
    ram_cell[   44299] = 32'h3c43304b;
    ram_cell[   44300] = 32'h11a09d67;
    ram_cell[   44301] = 32'hc2e76ead;
    ram_cell[   44302] = 32'ha92dcbd3;
    ram_cell[   44303] = 32'h4067676a;
    ram_cell[   44304] = 32'h92725472;
    ram_cell[   44305] = 32'h4e7e9dc8;
    ram_cell[   44306] = 32'h3d5eaa86;
    ram_cell[   44307] = 32'h76eb017b;
    ram_cell[   44308] = 32'hf2f3b740;
    ram_cell[   44309] = 32'h65b3ed76;
    ram_cell[   44310] = 32'hd895bbf1;
    ram_cell[   44311] = 32'h656be9f6;
    ram_cell[   44312] = 32'hf9ee9b1a;
    ram_cell[   44313] = 32'haf8617ce;
    ram_cell[   44314] = 32'hdf070851;
    ram_cell[   44315] = 32'h4458ed82;
    ram_cell[   44316] = 32'ha63f356c;
    ram_cell[   44317] = 32'h16212ba2;
    ram_cell[   44318] = 32'h86e55f64;
    ram_cell[   44319] = 32'h042a616a;
    ram_cell[   44320] = 32'h594364c4;
    ram_cell[   44321] = 32'h1918283a;
    ram_cell[   44322] = 32'h6c7b38b0;
    ram_cell[   44323] = 32'h2cb022af;
    ram_cell[   44324] = 32'h13d75da2;
    ram_cell[   44325] = 32'h11e883bb;
    ram_cell[   44326] = 32'h9ca56525;
    ram_cell[   44327] = 32'h2add5663;
    ram_cell[   44328] = 32'he9aef5e9;
    ram_cell[   44329] = 32'h664d94d8;
    ram_cell[   44330] = 32'hba6c7eda;
    ram_cell[   44331] = 32'h8826d2c0;
    ram_cell[   44332] = 32'h8a96a471;
    ram_cell[   44333] = 32'h1bfd31b0;
    ram_cell[   44334] = 32'h4b44e72e;
    ram_cell[   44335] = 32'h7ab240e6;
    ram_cell[   44336] = 32'h731e8bbf;
    ram_cell[   44337] = 32'he2cf34ee;
    ram_cell[   44338] = 32'ha17eebf8;
    ram_cell[   44339] = 32'he2d88267;
    ram_cell[   44340] = 32'h580e41ee;
    ram_cell[   44341] = 32'hec5d99e9;
    ram_cell[   44342] = 32'h8a1d126a;
    ram_cell[   44343] = 32'h5cdbc658;
    ram_cell[   44344] = 32'he328da54;
    ram_cell[   44345] = 32'h4986dcbe;
    ram_cell[   44346] = 32'he743ea21;
    ram_cell[   44347] = 32'hf7606968;
    ram_cell[   44348] = 32'h803da93a;
    ram_cell[   44349] = 32'hde8a750b;
    ram_cell[   44350] = 32'h314cb825;
    ram_cell[   44351] = 32'h64744572;
    ram_cell[   44352] = 32'h26159180;
    ram_cell[   44353] = 32'h8e91a21c;
    ram_cell[   44354] = 32'hc3b330f0;
    ram_cell[   44355] = 32'hcea5a119;
    ram_cell[   44356] = 32'hc7a4e90b;
    ram_cell[   44357] = 32'h0feb5d80;
    ram_cell[   44358] = 32'h096aa71d;
    ram_cell[   44359] = 32'h4fc4372b;
    ram_cell[   44360] = 32'ha330f1c5;
    ram_cell[   44361] = 32'h81ba31e4;
    ram_cell[   44362] = 32'h5fe63881;
    ram_cell[   44363] = 32'h692e89a4;
    ram_cell[   44364] = 32'h48d70100;
    ram_cell[   44365] = 32'he7d35ca7;
    ram_cell[   44366] = 32'h421e1495;
    ram_cell[   44367] = 32'h3be34b57;
    ram_cell[   44368] = 32'haabf4715;
    ram_cell[   44369] = 32'h69867791;
    ram_cell[   44370] = 32'h259d3c11;
    ram_cell[   44371] = 32'h2987e7f5;
    ram_cell[   44372] = 32'hc2bed72d;
    ram_cell[   44373] = 32'hf4f34d8d;
    ram_cell[   44374] = 32'h2b3f75a3;
    ram_cell[   44375] = 32'h08f21a72;
    ram_cell[   44376] = 32'h4af398ab;
    ram_cell[   44377] = 32'h6ab0fc9c;
    ram_cell[   44378] = 32'h35c22225;
    ram_cell[   44379] = 32'hbefa9723;
    ram_cell[   44380] = 32'h020c4bd8;
    ram_cell[   44381] = 32'hcf12e662;
    ram_cell[   44382] = 32'h2e343f4e;
    ram_cell[   44383] = 32'he0943023;
    ram_cell[   44384] = 32'h141ee030;
    ram_cell[   44385] = 32'hd459b3e8;
    ram_cell[   44386] = 32'hbe210645;
    ram_cell[   44387] = 32'h2e9e5625;
    ram_cell[   44388] = 32'h1ddcc653;
    ram_cell[   44389] = 32'h1a11ea3b;
    ram_cell[   44390] = 32'h9220f048;
    ram_cell[   44391] = 32'h9f59787d;
    ram_cell[   44392] = 32'h5d9d7891;
    ram_cell[   44393] = 32'hfc5a0dd1;
    ram_cell[   44394] = 32'h2becb5e1;
    ram_cell[   44395] = 32'hd5b1c4b8;
    ram_cell[   44396] = 32'h98e08221;
    ram_cell[   44397] = 32'h9c13f90b;
    ram_cell[   44398] = 32'ha144e0a2;
    ram_cell[   44399] = 32'hab66836a;
    ram_cell[   44400] = 32'h7d26d1cb;
    ram_cell[   44401] = 32'h3b93f12e;
    ram_cell[   44402] = 32'h4cba1b81;
    ram_cell[   44403] = 32'ha75f0d96;
    ram_cell[   44404] = 32'h6b3b57db;
    ram_cell[   44405] = 32'hfad3dbd1;
    ram_cell[   44406] = 32'h00872f32;
    ram_cell[   44407] = 32'h45fa53f2;
    ram_cell[   44408] = 32'hde5f8d8f;
    ram_cell[   44409] = 32'hb67f4222;
    ram_cell[   44410] = 32'h4931d306;
    ram_cell[   44411] = 32'h636827ea;
    ram_cell[   44412] = 32'h7f7126cb;
    ram_cell[   44413] = 32'h7ffabd80;
    ram_cell[   44414] = 32'he9d58d22;
    ram_cell[   44415] = 32'h11367207;
    ram_cell[   44416] = 32'h23426a25;
    ram_cell[   44417] = 32'h61bdefaa;
    ram_cell[   44418] = 32'h692fdc80;
    ram_cell[   44419] = 32'hfba14485;
    ram_cell[   44420] = 32'hbbd78336;
    ram_cell[   44421] = 32'hd2cba590;
    ram_cell[   44422] = 32'h086f2678;
    ram_cell[   44423] = 32'h2b69989b;
    ram_cell[   44424] = 32'hc61dea5e;
    ram_cell[   44425] = 32'haeaf7482;
    ram_cell[   44426] = 32'h8c3f26b4;
    ram_cell[   44427] = 32'he7c98f01;
    ram_cell[   44428] = 32'ha67aa4f1;
    ram_cell[   44429] = 32'he9e90574;
    ram_cell[   44430] = 32'h77ac5d15;
    ram_cell[   44431] = 32'h1d432429;
    ram_cell[   44432] = 32'he3e765dc;
    ram_cell[   44433] = 32'ha8dbf35e;
    ram_cell[   44434] = 32'h9e25c248;
    ram_cell[   44435] = 32'h6e369728;
    ram_cell[   44436] = 32'h1fadc51b;
    ram_cell[   44437] = 32'h8f5864a4;
    ram_cell[   44438] = 32'h4e47385a;
    ram_cell[   44439] = 32'hf9538061;
    ram_cell[   44440] = 32'h6d42b104;
    ram_cell[   44441] = 32'hc593d64c;
    ram_cell[   44442] = 32'hb810af26;
    ram_cell[   44443] = 32'h3357f4ad;
    ram_cell[   44444] = 32'h399120ea;
    ram_cell[   44445] = 32'he7d4e57c;
    ram_cell[   44446] = 32'hb835bd3d;
    ram_cell[   44447] = 32'h636e2389;
    ram_cell[   44448] = 32'hf93c94d3;
    ram_cell[   44449] = 32'h7cec2660;
    ram_cell[   44450] = 32'h5e3f0ca4;
    ram_cell[   44451] = 32'hcc2f85f8;
    ram_cell[   44452] = 32'h02bf67a5;
    ram_cell[   44453] = 32'h8710304a;
    ram_cell[   44454] = 32'h840e2452;
    ram_cell[   44455] = 32'h03b480aa;
    ram_cell[   44456] = 32'h55c316f4;
    ram_cell[   44457] = 32'h7a50455f;
    ram_cell[   44458] = 32'h45629c36;
    ram_cell[   44459] = 32'h421d62a6;
    ram_cell[   44460] = 32'hf7d6b39b;
    ram_cell[   44461] = 32'h5c5523b9;
    ram_cell[   44462] = 32'ha5bbcf9a;
    ram_cell[   44463] = 32'h8be0f635;
    ram_cell[   44464] = 32'h9f21a977;
    ram_cell[   44465] = 32'h8a429a70;
    ram_cell[   44466] = 32'hae7bde27;
    ram_cell[   44467] = 32'h58f89289;
    ram_cell[   44468] = 32'ha0093dea;
    ram_cell[   44469] = 32'h00a2746e;
    ram_cell[   44470] = 32'h722d07b0;
    ram_cell[   44471] = 32'hca10c3a3;
    ram_cell[   44472] = 32'h030b9553;
    ram_cell[   44473] = 32'ha80351f3;
    ram_cell[   44474] = 32'h4b4537be;
    ram_cell[   44475] = 32'h075e8abd;
    ram_cell[   44476] = 32'h7cde0eff;
    ram_cell[   44477] = 32'h1469e000;
    ram_cell[   44478] = 32'h62d60386;
    ram_cell[   44479] = 32'hf0371969;
    ram_cell[   44480] = 32'h2daa9fcb;
    ram_cell[   44481] = 32'h4816dccc;
    ram_cell[   44482] = 32'hd81d3b68;
    ram_cell[   44483] = 32'h48fed684;
    ram_cell[   44484] = 32'ha10be64b;
    ram_cell[   44485] = 32'h42c4e3ff;
    ram_cell[   44486] = 32'ha65c4725;
    ram_cell[   44487] = 32'hfb3b2201;
    ram_cell[   44488] = 32'he31cca3b;
    ram_cell[   44489] = 32'h7710108c;
    ram_cell[   44490] = 32'h36847c57;
    ram_cell[   44491] = 32'h4eba2b71;
    ram_cell[   44492] = 32'h6c96988d;
    ram_cell[   44493] = 32'h4e5cfbfa;
    ram_cell[   44494] = 32'h504c294c;
    ram_cell[   44495] = 32'h6452be21;
    ram_cell[   44496] = 32'h71292f64;
    ram_cell[   44497] = 32'hd61b4f13;
    ram_cell[   44498] = 32'hbc93d13c;
    ram_cell[   44499] = 32'hd8ccce9d;
    ram_cell[   44500] = 32'h96481a10;
    ram_cell[   44501] = 32'hbfd7a905;
    ram_cell[   44502] = 32'hb92c0cca;
    ram_cell[   44503] = 32'h58c3d67c;
    ram_cell[   44504] = 32'h76aa6f6c;
    ram_cell[   44505] = 32'hb846bc71;
    ram_cell[   44506] = 32'h7d48ee5e;
    ram_cell[   44507] = 32'h6385ac53;
    ram_cell[   44508] = 32'h7617d22e;
    ram_cell[   44509] = 32'h29d87499;
    ram_cell[   44510] = 32'hd82f1bb8;
    ram_cell[   44511] = 32'hef5ceeba;
    ram_cell[   44512] = 32'h907113c6;
    ram_cell[   44513] = 32'h0c95454f;
    ram_cell[   44514] = 32'hce34e22d;
    ram_cell[   44515] = 32'h70b39e5d;
    ram_cell[   44516] = 32'h6600006e;
    ram_cell[   44517] = 32'hdea40fd1;
    ram_cell[   44518] = 32'h0e236d4b;
    ram_cell[   44519] = 32'h00b5a14f;
    ram_cell[   44520] = 32'heee9cd62;
    ram_cell[   44521] = 32'h631cf66a;
    ram_cell[   44522] = 32'h44ca932f;
    ram_cell[   44523] = 32'h0fabe8ad;
    ram_cell[   44524] = 32'he8b56b5e;
    ram_cell[   44525] = 32'haa5dc1c3;
    ram_cell[   44526] = 32'h6fab0cfe;
    ram_cell[   44527] = 32'h1fe61bf3;
    ram_cell[   44528] = 32'hf0ea6b16;
    ram_cell[   44529] = 32'h113f5779;
    ram_cell[   44530] = 32'h920fffd4;
    ram_cell[   44531] = 32'h667ec1f6;
    ram_cell[   44532] = 32'h4b7cf4b2;
    ram_cell[   44533] = 32'h4e6e4cd5;
    ram_cell[   44534] = 32'hc51acbfc;
    ram_cell[   44535] = 32'hf2d8fb6d;
    ram_cell[   44536] = 32'hc94b4855;
    ram_cell[   44537] = 32'hb26d53aa;
    ram_cell[   44538] = 32'h5f60e097;
    ram_cell[   44539] = 32'h25e14a85;
    ram_cell[   44540] = 32'h483c2d3f;
    ram_cell[   44541] = 32'h9acfaa9b;
    ram_cell[   44542] = 32'h440e136c;
    ram_cell[   44543] = 32'h1cc51a25;
    ram_cell[   44544] = 32'h93adf2bc;
    ram_cell[   44545] = 32'h25bb5c8b;
    ram_cell[   44546] = 32'h6a8d8ce9;
    ram_cell[   44547] = 32'hf1cb8923;
    ram_cell[   44548] = 32'he1ff7eb9;
    ram_cell[   44549] = 32'h6168da6a;
    ram_cell[   44550] = 32'hfd932384;
    ram_cell[   44551] = 32'h055531fc;
    ram_cell[   44552] = 32'hfa0098d9;
    ram_cell[   44553] = 32'h6e53aa88;
    ram_cell[   44554] = 32'h98230bae;
    ram_cell[   44555] = 32'h0fb239f3;
    ram_cell[   44556] = 32'hba92bb3a;
    ram_cell[   44557] = 32'hc12af34f;
    ram_cell[   44558] = 32'hfcd37a0a;
    ram_cell[   44559] = 32'h6f781b8a;
    ram_cell[   44560] = 32'h6d5b353d;
    ram_cell[   44561] = 32'h43586ec3;
    ram_cell[   44562] = 32'h59e74c35;
    ram_cell[   44563] = 32'h258ad792;
    ram_cell[   44564] = 32'h2acfef68;
    ram_cell[   44565] = 32'h25c323cc;
    ram_cell[   44566] = 32'h09c592ee;
    ram_cell[   44567] = 32'ha21167b7;
    ram_cell[   44568] = 32'h66a9bd2e;
    ram_cell[   44569] = 32'hcbf2937e;
    ram_cell[   44570] = 32'h260ce739;
    ram_cell[   44571] = 32'h5b6ece1a;
    ram_cell[   44572] = 32'h7fb6143c;
    ram_cell[   44573] = 32'h818abc43;
    ram_cell[   44574] = 32'hb9ce3e75;
    ram_cell[   44575] = 32'h7c0a76ec;
    ram_cell[   44576] = 32'h870598ce;
    ram_cell[   44577] = 32'h1f87288c;
    ram_cell[   44578] = 32'hc9c6933f;
    ram_cell[   44579] = 32'hd4c45840;
    ram_cell[   44580] = 32'h8fe8c645;
    ram_cell[   44581] = 32'h633dd921;
    ram_cell[   44582] = 32'h25d7f8c8;
    ram_cell[   44583] = 32'hab37478d;
    ram_cell[   44584] = 32'h04fc80aa;
    ram_cell[   44585] = 32'h58245e7a;
    ram_cell[   44586] = 32'hcb14688d;
    ram_cell[   44587] = 32'h5bc9d803;
    ram_cell[   44588] = 32'h2be08910;
    ram_cell[   44589] = 32'h6f0d0443;
    ram_cell[   44590] = 32'h1e179a9f;
    ram_cell[   44591] = 32'h7c85bd78;
    ram_cell[   44592] = 32'h7a60b0e6;
    ram_cell[   44593] = 32'h1bbe3e1b;
    ram_cell[   44594] = 32'hf4972857;
    ram_cell[   44595] = 32'h4117fb1b;
    ram_cell[   44596] = 32'h90c0a583;
    ram_cell[   44597] = 32'hac7342fc;
    ram_cell[   44598] = 32'h51f7a47d;
    ram_cell[   44599] = 32'h7f8d8f97;
    ram_cell[   44600] = 32'h44ebe497;
    ram_cell[   44601] = 32'h86dc48a4;
    ram_cell[   44602] = 32'h5b07116c;
    ram_cell[   44603] = 32'h098fff17;
    ram_cell[   44604] = 32'h9c586fa1;
    ram_cell[   44605] = 32'he6166ade;
    ram_cell[   44606] = 32'h09b49290;
    ram_cell[   44607] = 32'hc0a59cf7;
    ram_cell[   44608] = 32'h4f6bb22d;
    ram_cell[   44609] = 32'h83b69865;
    ram_cell[   44610] = 32'habaf9bac;
    ram_cell[   44611] = 32'hbdbb604a;
    ram_cell[   44612] = 32'h68db973b;
    ram_cell[   44613] = 32'h97c2c4ed;
    ram_cell[   44614] = 32'haee286b7;
    ram_cell[   44615] = 32'h55cc9405;
    ram_cell[   44616] = 32'hed79b65d;
    ram_cell[   44617] = 32'h1173845e;
    ram_cell[   44618] = 32'h7cf8afee;
    ram_cell[   44619] = 32'h3051e0a3;
    ram_cell[   44620] = 32'h1849aa19;
    ram_cell[   44621] = 32'hff0ec087;
    ram_cell[   44622] = 32'h79aa7dd5;
    ram_cell[   44623] = 32'h428ec264;
    ram_cell[   44624] = 32'hc040e575;
    ram_cell[   44625] = 32'h6603b013;
    ram_cell[   44626] = 32'h6bce5e72;
    ram_cell[   44627] = 32'hec163852;
    ram_cell[   44628] = 32'h36925357;
    ram_cell[   44629] = 32'h8b0b494d;
    ram_cell[   44630] = 32'h8ffbe621;
    ram_cell[   44631] = 32'h73b7629d;
    ram_cell[   44632] = 32'h3425f386;
    ram_cell[   44633] = 32'heac5f2c7;
    ram_cell[   44634] = 32'hfe363213;
    ram_cell[   44635] = 32'hc11c5877;
    ram_cell[   44636] = 32'he0b6cf4f;
    ram_cell[   44637] = 32'h5c99c923;
    ram_cell[   44638] = 32'h84ce9123;
    ram_cell[   44639] = 32'h39581e6d;
    ram_cell[   44640] = 32'hcf0f920c;
    ram_cell[   44641] = 32'h102d458e;
    ram_cell[   44642] = 32'h524f49fb;
    ram_cell[   44643] = 32'h0a2bfd9a;
    ram_cell[   44644] = 32'hce76a5df;
    ram_cell[   44645] = 32'h6fdb6a72;
    ram_cell[   44646] = 32'ha8d9d0b4;
    ram_cell[   44647] = 32'h9fd75f51;
    ram_cell[   44648] = 32'hc82a0afa;
    ram_cell[   44649] = 32'h49b5e87f;
    ram_cell[   44650] = 32'h1a680610;
    ram_cell[   44651] = 32'h9ddcc823;
    ram_cell[   44652] = 32'he22244bb;
    ram_cell[   44653] = 32'h4fa831e2;
    ram_cell[   44654] = 32'hda65c7fc;
    ram_cell[   44655] = 32'hc188eed8;
    ram_cell[   44656] = 32'h0f1bef31;
    ram_cell[   44657] = 32'h897c6774;
    ram_cell[   44658] = 32'h5f6b795a;
    ram_cell[   44659] = 32'h08740cea;
    ram_cell[   44660] = 32'hbb1b1ffc;
    ram_cell[   44661] = 32'ha9771d6f;
    ram_cell[   44662] = 32'hf67302b7;
    ram_cell[   44663] = 32'he09503ed;
    ram_cell[   44664] = 32'h2f0145ca;
    ram_cell[   44665] = 32'h5d7f0105;
    ram_cell[   44666] = 32'hfb730db7;
    ram_cell[   44667] = 32'h81bc0d44;
    ram_cell[   44668] = 32'ha8e74a25;
    ram_cell[   44669] = 32'h515cbf7b;
    ram_cell[   44670] = 32'h9fbb0cc9;
    ram_cell[   44671] = 32'h209d8625;
    ram_cell[   44672] = 32'hd6df125d;
    ram_cell[   44673] = 32'h627ce596;
    ram_cell[   44674] = 32'h97a7e931;
    ram_cell[   44675] = 32'he64de851;
    ram_cell[   44676] = 32'h7cd17830;
    ram_cell[   44677] = 32'h5200634c;
    ram_cell[   44678] = 32'haf48fc09;
    ram_cell[   44679] = 32'h2cca3c0f;
    ram_cell[   44680] = 32'h9b44850b;
    ram_cell[   44681] = 32'hb87f019f;
    ram_cell[   44682] = 32'h770ab9d2;
    ram_cell[   44683] = 32'h843a386c;
    ram_cell[   44684] = 32'h03c9836a;
    ram_cell[   44685] = 32'h797bea6c;
    ram_cell[   44686] = 32'h1c42a294;
    ram_cell[   44687] = 32'h142963c9;
    ram_cell[   44688] = 32'h970bfbf1;
    ram_cell[   44689] = 32'h8ead6468;
    ram_cell[   44690] = 32'h7b69b8b0;
    ram_cell[   44691] = 32'h58e33097;
    ram_cell[   44692] = 32'hb7d8faff;
    ram_cell[   44693] = 32'ha51410fd;
    ram_cell[   44694] = 32'h78cd2551;
    ram_cell[   44695] = 32'h868030fe;
    ram_cell[   44696] = 32'h0ae52999;
    ram_cell[   44697] = 32'h6a63597a;
    ram_cell[   44698] = 32'h541c90d9;
    ram_cell[   44699] = 32'he4589af0;
    ram_cell[   44700] = 32'hb34e8227;
    ram_cell[   44701] = 32'h6412737d;
    ram_cell[   44702] = 32'ha4f592a3;
    ram_cell[   44703] = 32'h6ded7e87;
    ram_cell[   44704] = 32'hbda9fc96;
    ram_cell[   44705] = 32'hbe7a061e;
    ram_cell[   44706] = 32'he2ba6981;
    ram_cell[   44707] = 32'h4d16f84f;
    ram_cell[   44708] = 32'h250c9b9d;
    ram_cell[   44709] = 32'had08b632;
    ram_cell[   44710] = 32'hfcc14112;
    ram_cell[   44711] = 32'h19724e81;
    ram_cell[   44712] = 32'h3d6260c1;
    ram_cell[   44713] = 32'h3f6904fa;
    ram_cell[   44714] = 32'h2e0598d0;
    ram_cell[   44715] = 32'hbe5df025;
    ram_cell[   44716] = 32'he96325c1;
    ram_cell[   44717] = 32'h4f54eb62;
    ram_cell[   44718] = 32'h0bade0e9;
    ram_cell[   44719] = 32'hfbcfb5b2;
    ram_cell[   44720] = 32'h1b72b383;
    ram_cell[   44721] = 32'h957bbb30;
    ram_cell[   44722] = 32'h19038f17;
    ram_cell[   44723] = 32'h34ebd9ef;
    ram_cell[   44724] = 32'h3110562b;
    ram_cell[   44725] = 32'h355e08ed;
    ram_cell[   44726] = 32'he30dc30d;
    ram_cell[   44727] = 32'h62026a06;
    ram_cell[   44728] = 32'hb03f9bc4;
    ram_cell[   44729] = 32'h2095a29d;
    ram_cell[   44730] = 32'h0da4e504;
    ram_cell[   44731] = 32'hc4fcaf06;
    ram_cell[   44732] = 32'h95deb6ef;
    ram_cell[   44733] = 32'hdf885499;
    ram_cell[   44734] = 32'hc0885ab3;
    ram_cell[   44735] = 32'h2312daec;
    ram_cell[   44736] = 32'hcc95b651;
    ram_cell[   44737] = 32'h917fde55;
    ram_cell[   44738] = 32'hc2eb80ff;
    ram_cell[   44739] = 32'h78b62714;
    ram_cell[   44740] = 32'h9278557b;
    ram_cell[   44741] = 32'h5e99e8ec;
    ram_cell[   44742] = 32'h6bd6bf68;
    ram_cell[   44743] = 32'hfd0eadd2;
    ram_cell[   44744] = 32'h1c002807;
    ram_cell[   44745] = 32'hba4bbf5b;
    ram_cell[   44746] = 32'h8160a896;
    ram_cell[   44747] = 32'h6d5661e8;
    ram_cell[   44748] = 32'h17490429;
    ram_cell[   44749] = 32'h72b689d6;
    ram_cell[   44750] = 32'h32784bc6;
    ram_cell[   44751] = 32'h00b4a884;
    ram_cell[   44752] = 32'h21870a6d;
    ram_cell[   44753] = 32'h3410ba24;
    ram_cell[   44754] = 32'h1c434f0d;
    ram_cell[   44755] = 32'hc8f32595;
    ram_cell[   44756] = 32'hee953d66;
    ram_cell[   44757] = 32'hb21a384e;
    ram_cell[   44758] = 32'hf9413ba1;
    ram_cell[   44759] = 32'hc17a5d8d;
    ram_cell[   44760] = 32'hb2f75126;
    ram_cell[   44761] = 32'h3ab8d69e;
    ram_cell[   44762] = 32'h2a17ee89;
    ram_cell[   44763] = 32'h2a729c1c;
    ram_cell[   44764] = 32'h9e5a1651;
    ram_cell[   44765] = 32'h5d12cd0d;
    ram_cell[   44766] = 32'h0653bd15;
    ram_cell[   44767] = 32'h6910d221;
    ram_cell[   44768] = 32'h2889570f;
    ram_cell[   44769] = 32'h3d314728;
    ram_cell[   44770] = 32'h99caab5e;
    ram_cell[   44771] = 32'hfa2eea99;
    ram_cell[   44772] = 32'he2cca876;
    ram_cell[   44773] = 32'h850f0ed8;
    ram_cell[   44774] = 32'ha8657c37;
    ram_cell[   44775] = 32'h5c1a8fdb;
    ram_cell[   44776] = 32'h41404183;
    ram_cell[   44777] = 32'h75b55e47;
    ram_cell[   44778] = 32'h99a0f376;
    ram_cell[   44779] = 32'h427b2955;
    ram_cell[   44780] = 32'h3fb72085;
    ram_cell[   44781] = 32'h4f0bae58;
    ram_cell[   44782] = 32'h0da65fc1;
    ram_cell[   44783] = 32'h1f84b324;
    ram_cell[   44784] = 32'h60e844e5;
    ram_cell[   44785] = 32'h22122d43;
    ram_cell[   44786] = 32'h2d01762c;
    ram_cell[   44787] = 32'h3e458485;
    ram_cell[   44788] = 32'h3bf0c0e4;
    ram_cell[   44789] = 32'h50cc05d5;
    ram_cell[   44790] = 32'h6d60b018;
    ram_cell[   44791] = 32'hf2542290;
    ram_cell[   44792] = 32'h7676e6f2;
    ram_cell[   44793] = 32'h63c4767b;
    ram_cell[   44794] = 32'h4048f318;
    ram_cell[   44795] = 32'h5f9ec246;
    ram_cell[   44796] = 32'hbd1ef96f;
    ram_cell[   44797] = 32'haf8aa846;
    ram_cell[   44798] = 32'h7c612184;
    ram_cell[   44799] = 32'he8d75fbd;
    ram_cell[   44800] = 32'h230168d4;
    ram_cell[   44801] = 32'ha8448311;
    ram_cell[   44802] = 32'h798cad9b;
    ram_cell[   44803] = 32'hb66337d4;
    ram_cell[   44804] = 32'h76912994;
    ram_cell[   44805] = 32'heed841be;
    ram_cell[   44806] = 32'h173cc30a;
    ram_cell[   44807] = 32'h19243ec6;
    ram_cell[   44808] = 32'hb0d5573a;
    ram_cell[   44809] = 32'h1a0a5e20;
    ram_cell[   44810] = 32'h82cdebee;
    ram_cell[   44811] = 32'h344fc324;
    ram_cell[   44812] = 32'h3c95938b;
    ram_cell[   44813] = 32'h304baf1a;
    ram_cell[   44814] = 32'h4909b8ea;
    ram_cell[   44815] = 32'hd6c7cda9;
    ram_cell[   44816] = 32'hf2edfc70;
    ram_cell[   44817] = 32'h9ead7261;
    ram_cell[   44818] = 32'hc8cb58bf;
    ram_cell[   44819] = 32'hd6ecfb2d;
    ram_cell[   44820] = 32'h17c12931;
    ram_cell[   44821] = 32'h5b45b719;
    ram_cell[   44822] = 32'hb2c8d6d1;
    ram_cell[   44823] = 32'h6279354c;
    ram_cell[   44824] = 32'had7df580;
    ram_cell[   44825] = 32'h85cc1c4e;
    ram_cell[   44826] = 32'ha022fcc2;
    ram_cell[   44827] = 32'h2de6b97a;
    ram_cell[   44828] = 32'h0367a15c;
    ram_cell[   44829] = 32'haa2c442f;
    ram_cell[   44830] = 32'h7a42fea0;
    ram_cell[   44831] = 32'h2a07bad6;
    ram_cell[   44832] = 32'h5ab5151e;
    ram_cell[   44833] = 32'h2f8415d7;
    ram_cell[   44834] = 32'h147048c1;
    ram_cell[   44835] = 32'h31b01c9a;
    ram_cell[   44836] = 32'hfdab4b2d;
    ram_cell[   44837] = 32'hf1003b52;
    ram_cell[   44838] = 32'ha9eb29d1;
    ram_cell[   44839] = 32'h53a8f277;
    ram_cell[   44840] = 32'h50eac415;
    ram_cell[   44841] = 32'h97d7da9a;
    ram_cell[   44842] = 32'hd8b20016;
    ram_cell[   44843] = 32'hc41df3c1;
    ram_cell[   44844] = 32'h4b7d4f2e;
    ram_cell[   44845] = 32'hdfb5675a;
    ram_cell[   44846] = 32'h70998769;
    ram_cell[   44847] = 32'h263d11d4;
    ram_cell[   44848] = 32'h37c42b59;
    ram_cell[   44849] = 32'h31a15504;
    ram_cell[   44850] = 32'h03f6f87d;
    ram_cell[   44851] = 32'h29c5a765;
    ram_cell[   44852] = 32'h6648dac2;
    ram_cell[   44853] = 32'h6c7a8456;
    ram_cell[   44854] = 32'hc42060a4;
    ram_cell[   44855] = 32'h09518ecc;
    ram_cell[   44856] = 32'h1619f1ae;
    ram_cell[   44857] = 32'hb3a71c14;
    ram_cell[   44858] = 32'ha70ece6f;
    ram_cell[   44859] = 32'hc02f81a9;
    ram_cell[   44860] = 32'he602e73d;
    ram_cell[   44861] = 32'hf6deaab0;
    ram_cell[   44862] = 32'hbc40af4f;
    ram_cell[   44863] = 32'h4152d5e4;
    ram_cell[   44864] = 32'h00975c60;
    ram_cell[   44865] = 32'h459f1c05;
    ram_cell[   44866] = 32'h4e1dbb07;
    ram_cell[   44867] = 32'h348e1993;
    ram_cell[   44868] = 32'h19fa8ffb;
    ram_cell[   44869] = 32'h0a4eee4c;
    ram_cell[   44870] = 32'hddd00762;
    ram_cell[   44871] = 32'h24a115dd;
    ram_cell[   44872] = 32'h3fcf283d;
    ram_cell[   44873] = 32'hf46c3a20;
    ram_cell[   44874] = 32'h6e535678;
    ram_cell[   44875] = 32'hc65f5890;
    ram_cell[   44876] = 32'hfdfe6816;
    ram_cell[   44877] = 32'ha55fa12b;
    ram_cell[   44878] = 32'hdb4a82c1;
    ram_cell[   44879] = 32'h334e65ed;
    ram_cell[   44880] = 32'h8a6d2027;
    ram_cell[   44881] = 32'h4a7ee488;
    ram_cell[   44882] = 32'h47547af3;
    ram_cell[   44883] = 32'h3602f64e;
    ram_cell[   44884] = 32'h07289872;
    ram_cell[   44885] = 32'hb8b70b26;
    ram_cell[   44886] = 32'h0b59e9c1;
    ram_cell[   44887] = 32'h6b51a2c4;
    ram_cell[   44888] = 32'h2491c147;
    ram_cell[   44889] = 32'h1807bb11;
    ram_cell[   44890] = 32'h76b0e7d9;
    ram_cell[   44891] = 32'hc664aeb0;
    ram_cell[   44892] = 32'h8ed697d5;
    ram_cell[   44893] = 32'h20b78c08;
    ram_cell[   44894] = 32'hd6b9ed4b;
    ram_cell[   44895] = 32'h1076864d;
    ram_cell[   44896] = 32'h628b299f;
    ram_cell[   44897] = 32'h0675d048;
    ram_cell[   44898] = 32'hb31ef755;
    ram_cell[   44899] = 32'h0835181b;
    ram_cell[   44900] = 32'hfc1e234d;
    ram_cell[   44901] = 32'h22ef98f7;
    ram_cell[   44902] = 32'h1dedffa1;
    ram_cell[   44903] = 32'hc2b0d82d;
    ram_cell[   44904] = 32'hd261ec3f;
    ram_cell[   44905] = 32'h99b187fe;
    ram_cell[   44906] = 32'hb5b58cc7;
    ram_cell[   44907] = 32'h9129a7e0;
    ram_cell[   44908] = 32'hfad82f3e;
    ram_cell[   44909] = 32'h72cb72c9;
    ram_cell[   44910] = 32'h09cc94af;
    ram_cell[   44911] = 32'h7dc58892;
    ram_cell[   44912] = 32'h5881bf39;
    ram_cell[   44913] = 32'hae32eacb;
    ram_cell[   44914] = 32'h35a007ee;
    ram_cell[   44915] = 32'h3a34ff71;
    ram_cell[   44916] = 32'h460e6cdb;
    ram_cell[   44917] = 32'hf9f95d0b;
    ram_cell[   44918] = 32'hf38c4c61;
    ram_cell[   44919] = 32'hf7599275;
    ram_cell[   44920] = 32'h14837f37;
    ram_cell[   44921] = 32'h2f76e08a;
    ram_cell[   44922] = 32'hb831ba03;
    ram_cell[   44923] = 32'hc5664c68;
    ram_cell[   44924] = 32'hc0f08f6e;
    ram_cell[   44925] = 32'h144e2e70;
    ram_cell[   44926] = 32'hea2ab151;
    ram_cell[   44927] = 32'h135d23e1;
    ram_cell[   44928] = 32'h4224b601;
    ram_cell[   44929] = 32'hc3308785;
    ram_cell[   44930] = 32'h1a098a0f;
    ram_cell[   44931] = 32'h5483bdba;
    ram_cell[   44932] = 32'h074a7f70;
    ram_cell[   44933] = 32'he3339359;
    ram_cell[   44934] = 32'h92582668;
    ram_cell[   44935] = 32'hb01f63d6;
    ram_cell[   44936] = 32'h014fdf9e;
    ram_cell[   44937] = 32'hed6224c2;
    ram_cell[   44938] = 32'h09e398f0;
    ram_cell[   44939] = 32'h969cfc2e;
    ram_cell[   44940] = 32'h5ea163bb;
    ram_cell[   44941] = 32'h16a1dc5f;
    ram_cell[   44942] = 32'h0d5d5ced;
    ram_cell[   44943] = 32'h463ae784;
    ram_cell[   44944] = 32'hcbd6b85d;
    ram_cell[   44945] = 32'hcd4e72ec;
    ram_cell[   44946] = 32'h8d323a2e;
    ram_cell[   44947] = 32'h812697b4;
    ram_cell[   44948] = 32'h62fb875b;
    ram_cell[   44949] = 32'h232abb38;
    ram_cell[   44950] = 32'h6c48419e;
    ram_cell[   44951] = 32'h240509fe;
    ram_cell[   44952] = 32'h7c74e1dc;
    ram_cell[   44953] = 32'h019f8074;
    ram_cell[   44954] = 32'h505708be;
    ram_cell[   44955] = 32'h54d6f245;
    ram_cell[   44956] = 32'h134dcdb5;
    ram_cell[   44957] = 32'h33427425;
    ram_cell[   44958] = 32'hdc03f0d7;
    ram_cell[   44959] = 32'h3e2a5f19;
    ram_cell[   44960] = 32'h9ce3c58f;
    ram_cell[   44961] = 32'hd16f14cf;
    ram_cell[   44962] = 32'hd7b331f3;
    ram_cell[   44963] = 32'hdd7ad6ce;
    ram_cell[   44964] = 32'he9d4b049;
    ram_cell[   44965] = 32'h352be15f;
    ram_cell[   44966] = 32'hab5aefe8;
    ram_cell[   44967] = 32'h579b4d03;
    ram_cell[   44968] = 32'he89616b2;
    ram_cell[   44969] = 32'ha17c6bb8;
    ram_cell[   44970] = 32'ha551fb56;
    ram_cell[   44971] = 32'hfa2f8dfa;
    ram_cell[   44972] = 32'hf04ec484;
    ram_cell[   44973] = 32'he4844da7;
    ram_cell[   44974] = 32'h9d69aa90;
    ram_cell[   44975] = 32'he4f276fd;
    ram_cell[   44976] = 32'he7ac8c03;
    ram_cell[   44977] = 32'h93a29c5c;
    ram_cell[   44978] = 32'hb04b67fd;
    ram_cell[   44979] = 32'hb670d996;
    ram_cell[   44980] = 32'h54221b59;
    ram_cell[   44981] = 32'h7b5936cc;
    ram_cell[   44982] = 32'h26737f01;
    ram_cell[   44983] = 32'h039967c9;
    ram_cell[   44984] = 32'h86a87c78;
    ram_cell[   44985] = 32'h45c290c6;
    ram_cell[   44986] = 32'h1b62d217;
    ram_cell[   44987] = 32'he962d9e7;
    ram_cell[   44988] = 32'h6b4266f9;
    ram_cell[   44989] = 32'h7628d852;
    ram_cell[   44990] = 32'h6ba123bf;
    ram_cell[   44991] = 32'h06daa083;
    ram_cell[   44992] = 32'hf24cc0a4;
    ram_cell[   44993] = 32'haf592076;
    ram_cell[   44994] = 32'hc9fe6b9d;
    ram_cell[   44995] = 32'habf9e92d;
    ram_cell[   44996] = 32'h124a47b0;
    ram_cell[   44997] = 32'h05f1cee2;
    ram_cell[   44998] = 32'h18545b8b;
    ram_cell[   44999] = 32'ha0c9e430;
    ram_cell[   45000] = 32'habcaaa5e;
    ram_cell[   45001] = 32'h050325b2;
    ram_cell[   45002] = 32'h827ca918;
    ram_cell[   45003] = 32'h972deeaa;
    ram_cell[   45004] = 32'h89e8edcd;
    ram_cell[   45005] = 32'h89e50e44;
    ram_cell[   45006] = 32'hab1e3eae;
    ram_cell[   45007] = 32'hb8ca846d;
    ram_cell[   45008] = 32'h4f343530;
    ram_cell[   45009] = 32'hc8ab0e26;
    ram_cell[   45010] = 32'hab54d2f7;
    ram_cell[   45011] = 32'ha3d83939;
    ram_cell[   45012] = 32'h22fe9caa;
    ram_cell[   45013] = 32'h2d42ac7e;
    ram_cell[   45014] = 32'he321a7f8;
    ram_cell[   45015] = 32'h336ebd10;
    ram_cell[   45016] = 32'h8ec88273;
    ram_cell[   45017] = 32'h38e3b276;
    ram_cell[   45018] = 32'hbae6f47e;
    ram_cell[   45019] = 32'h9d9370ab;
    ram_cell[   45020] = 32'h92bb9f9e;
    ram_cell[   45021] = 32'h5ddeda37;
    ram_cell[   45022] = 32'h35b38aa2;
    ram_cell[   45023] = 32'heccdd7b9;
    ram_cell[   45024] = 32'h78e2dd6d;
    ram_cell[   45025] = 32'h062b2ab8;
    ram_cell[   45026] = 32'h54cba837;
    ram_cell[   45027] = 32'h773687bd;
    ram_cell[   45028] = 32'h36eecc74;
    ram_cell[   45029] = 32'ha0ddeee9;
    ram_cell[   45030] = 32'hae174064;
    ram_cell[   45031] = 32'h24d725e5;
    ram_cell[   45032] = 32'hd9994abd;
    ram_cell[   45033] = 32'hf749bb5e;
    ram_cell[   45034] = 32'h6de8201b;
    ram_cell[   45035] = 32'h6de5e86a;
    ram_cell[   45036] = 32'h5924521e;
    ram_cell[   45037] = 32'hb808a81e;
    ram_cell[   45038] = 32'h2ea066c3;
    ram_cell[   45039] = 32'hbb31ffb7;
    ram_cell[   45040] = 32'h5a5bdba8;
    ram_cell[   45041] = 32'h6fdfc4e2;
    ram_cell[   45042] = 32'h294c0ede;
    ram_cell[   45043] = 32'h0c53d4e8;
    ram_cell[   45044] = 32'h17042543;
    ram_cell[   45045] = 32'h76dd733b;
    ram_cell[   45046] = 32'h2f9a23f1;
    ram_cell[   45047] = 32'h61e12bba;
    ram_cell[   45048] = 32'h3060f193;
    ram_cell[   45049] = 32'h849ad8ae;
    ram_cell[   45050] = 32'he2526978;
    ram_cell[   45051] = 32'hdd680844;
    ram_cell[   45052] = 32'h7046adc9;
    ram_cell[   45053] = 32'hf8cbe81a;
    ram_cell[   45054] = 32'h2b6a41a4;
    ram_cell[   45055] = 32'h82c96676;
    ram_cell[   45056] = 32'h909d1421;
    ram_cell[   45057] = 32'h76e4930b;
    ram_cell[   45058] = 32'hbb1b2dfa;
    ram_cell[   45059] = 32'h091d2c7a;
    ram_cell[   45060] = 32'he38a1fbc;
    ram_cell[   45061] = 32'h065694d4;
    ram_cell[   45062] = 32'h96531970;
    ram_cell[   45063] = 32'hcbd2e6c3;
    ram_cell[   45064] = 32'hbdbd3dbf;
    ram_cell[   45065] = 32'h2a5cfeba;
    ram_cell[   45066] = 32'h38318a4d;
    ram_cell[   45067] = 32'hab34fd4f;
    ram_cell[   45068] = 32'h0a52eded;
    ram_cell[   45069] = 32'h6238fddb;
    ram_cell[   45070] = 32'h5110959b;
    ram_cell[   45071] = 32'h69611991;
    ram_cell[   45072] = 32'h40e83e71;
    ram_cell[   45073] = 32'hb5279d19;
    ram_cell[   45074] = 32'hb3fdd567;
    ram_cell[   45075] = 32'h1462a003;
    ram_cell[   45076] = 32'h5a6c2968;
    ram_cell[   45077] = 32'had19a9fe;
    ram_cell[   45078] = 32'haf4fbfb3;
    ram_cell[   45079] = 32'he256745f;
    ram_cell[   45080] = 32'h65d24e36;
    ram_cell[   45081] = 32'h34be0892;
    ram_cell[   45082] = 32'h59dab7ae;
    ram_cell[   45083] = 32'hfd5598fc;
    ram_cell[   45084] = 32'heef9bc5b;
    ram_cell[   45085] = 32'h9beee2c5;
    ram_cell[   45086] = 32'hba6d6f11;
    ram_cell[   45087] = 32'haa1b2d40;
    ram_cell[   45088] = 32'ha4263b70;
    ram_cell[   45089] = 32'hd1a32465;
    ram_cell[   45090] = 32'hfbea6baa;
    ram_cell[   45091] = 32'h2bdc887a;
    ram_cell[   45092] = 32'h6be33afe;
    ram_cell[   45093] = 32'h200c466c;
    ram_cell[   45094] = 32'h5e193e52;
    ram_cell[   45095] = 32'h28975cf8;
    ram_cell[   45096] = 32'h1317b0a4;
    ram_cell[   45097] = 32'h82b524dc;
    ram_cell[   45098] = 32'hc0e10da5;
    ram_cell[   45099] = 32'h4a75f543;
    ram_cell[   45100] = 32'h68d0b193;
    ram_cell[   45101] = 32'he8e48c31;
    ram_cell[   45102] = 32'h65d68895;
    ram_cell[   45103] = 32'h4d62a996;
    ram_cell[   45104] = 32'h65081b29;
    ram_cell[   45105] = 32'h35098b3b;
    ram_cell[   45106] = 32'h3d8de2a6;
    ram_cell[   45107] = 32'h3f18d145;
    ram_cell[   45108] = 32'hb941e619;
    ram_cell[   45109] = 32'ha91d9bac;
    ram_cell[   45110] = 32'h221d1c57;
    ram_cell[   45111] = 32'hb822b30a;
    ram_cell[   45112] = 32'haa56e4a6;
    ram_cell[   45113] = 32'hf9ca14c3;
    ram_cell[   45114] = 32'hb7d0ec38;
    ram_cell[   45115] = 32'h93f8f2c5;
    ram_cell[   45116] = 32'h3f83fcfa;
    ram_cell[   45117] = 32'h2f204dfd;
    ram_cell[   45118] = 32'hfc770f4c;
    ram_cell[   45119] = 32'h63c8d0db;
    ram_cell[   45120] = 32'h85a7a23c;
    ram_cell[   45121] = 32'hc55572a1;
    ram_cell[   45122] = 32'h16ae97b6;
    ram_cell[   45123] = 32'h58b19c4d;
    ram_cell[   45124] = 32'h93b6ee0e;
    ram_cell[   45125] = 32'hc1f6eef0;
    ram_cell[   45126] = 32'h2517817e;
    ram_cell[   45127] = 32'hc02fd465;
    ram_cell[   45128] = 32'h1048e478;
    ram_cell[   45129] = 32'h4e7d4959;
    ram_cell[   45130] = 32'h1a3f7055;
    ram_cell[   45131] = 32'hfb0dabd6;
    ram_cell[   45132] = 32'hfc593650;
    ram_cell[   45133] = 32'h757838b1;
    ram_cell[   45134] = 32'h9183d153;
    ram_cell[   45135] = 32'h9c93c785;
    ram_cell[   45136] = 32'h95f939d9;
    ram_cell[   45137] = 32'h6040b90b;
    ram_cell[   45138] = 32'hf387451e;
    ram_cell[   45139] = 32'h551dd14d;
    ram_cell[   45140] = 32'hfaf1974f;
    ram_cell[   45141] = 32'h62f4df33;
    ram_cell[   45142] = 32'he0242fa6;
    ram_cell[   45143] = 32'h974a8774;
    ram_cell[   45144] = 32'hbe6fe279;
    ram_cell[   45145] = 32'h36d525fb;
    ram_cell[   45146] = 32'h85471431;
    ram_cell[   45147] = 32'h7e80956c;
    ram_cell[   45148] = 32'hd94fadb5;
    ram_cell[   45149] = 32'h63598135;
    ram_cell[   45150] = 32'ha58def8d;
    ram_cell[   45151] = 32'h409be8a9;
    ram_cell[   45152] = 32'h9249f165;
    ram_cell[   45153] = 32'he5b9bbfa;
    ram_cell[   45154] = 32'h3688e030;
    ram_cell[   45155] = 32'hbbeb293f;
    ram_cell[   45156] = 32'hb2a076df;
    ram_cell[   45157] = 32'hc14b8dc4;
    ram_cell[   45158] = 32'h00a593d5;
    ram_cell[   45159] = 32'haa380321;
    ram_cell[   45160] = 32'hac7461be;
    ram_cell[   45161] = 32'h26c62d99;
    ram_cell[   45162] = 32'h0431688c;
    ram_cell[   45163] = 32'hf1136bba;
    ram_cell[   45164] = 32'h6434199e;
    ram_cell[   45165] = 32'hd0c295e5;
    ram_cell[   45166] = 32'h4ff99cbd;
    ram_cell[   45167] = 32'hd752c0c1;
    ram_cell[   45168] = 32'hb7a719d4;
    ram_cell[   45169] = 32'hea88cf63;
    ram_cell[   45170] = 32'hb0977705;
    ram_cell[   45171] = 32'h1e1b56c7;
    ram_cell[   45172] = 32'he09e5e0b;
    ram_cell[   45173] = 32'h417a53a9;
    ram_cell[   45174] = 32'he3b321d9;
    ram_cell[   45175] = 32'hdbbca4ff;
    ram_cell[   45176] = 32'h4e9d1039;
    ram_cell[   45177] = 32'hd4db48b4;
    ram_cell[   45178] = 32'h4e8122bb;
    ram_cell[   45179] = 32'hb8ade5c3;
    ram_cell[   45180] = 32'hdcb70b8a;
    ram_cell[   45181] = 32'h520ea4ab;
    ram_cell[   45182] = 32'hbeb7750e;
    ram_cell[   45183] = 32'h518ce4aa;
    ram_cell[   45184] = 32'h57d6bf52;
    ram_cell[   45185] = 32'h5895c023;
    ram_cell[   45186] = 32'hec093b92;
    ram_cell[   45187] = 32'h4e3d0721;
    ram_cell[   45188] = 32'h511df62b;
    ram_cell[   45189] = 32'h167fc944;
    ram_cell[   45190] = 32'h099ce47f;
    ram_cell[   45191] = 32'h4aef0a43;
    ram_cell[   45192] = 32'ha0ef639f;
    ram_cell[   45193] = 32'h9eb6afad;
    ram_cell[   45194] = 32'h3854a0e8;
    ram_cell[   45195] = 32'h1a3a39f2;
    ram_cell[   45196] = 32'h3ac1f176;
    ram_cell[   45197] = 32'h0ebd85be;
    ram_cell[   45198] = 32'h8107474d;
    ram_cell[   45199] = 32'h8f93c904;
    ram_cell[   45200] = 32'h79320c87;
    ram_cell[   45201] = 32'hf0edbe7f;
    ram_cell[   45202] = 32'hcf68144d;
    ram_cell[   45203] = 32'hfb05b2cc;
    ram_cell[   45204] = 32'h11d22a37;
    ram_cell[   45205] = 32'h27b6ee55;
    ram_cell[   45206] = 32'h9a82ee0d;
    ram_cell[   45207] = 32'h2843ece5;
    ram_cell[   45208] = 32'hf2d22a87;
    ram_cell[   45209] = 32'h35382bbe;
    ram_cell[   45210] = 32'h4be841c4;
    ram_cell[   45211] = 32'h1a8ec0fb;
    ram_cell[   45212] = 32'h7ed3c3b2;
    ram_cell[   45213] = 32'h8d9d1c89;
    ram_cell[   45214] = 32'h72a54b9f;
    ram_cell[   45215] = 32'hf973555e;
    ram_cell[   45216] = 32'h4b31acf2;
    ram_cell[   45217] = 32'hb042ff16;
    ram_cell[   45218] = 32'h8df69138;
    ram_cell[   45219] = 32'hef37329e;
    ram_cell[   45220] = 32'h1c6854cd;
    ram_cell[   45221] = 32'h27119e38;
    ram_cell[   45222] = 32'h8121cce7;
    ram_cell[   45223] = 32'h5ce3c5be;
    ram_cell[   45224] = 32'h9bf9b655;
    ram_cell[   45225] = 32'h2aad166f;
    ram_cell[   45226] = 32'h7c339550;
    ram_cell[   45227] = 32'hdd8b043f;
    ram_cell[   45228] = 32'h9949f433;
    ram_cell[   45229] = 32'h9b5ee46d;
    ram_cell[   45230] = 32'hb49770d5;
    ram_cell[   45231] = 32'h0cfa27eb;
    ram_cell[   45232] = 32'h82a2722e;
    ram_cell[   45233] = 32'h1e171c36;
    ram_cell[   45234] = 32'ha2b13d37;
    ram_cell[   45235] = 32'hccaebb1e;
    ram_cell[   45236] = 32'h6552e4b1;
    ram_cell[   45237] = 32'hc6100879;
    ram_cell[   45238] = 32'h8baf3218;
    ram_cell[   45239] = 32'hd8551029;
    ram_cell[   45240] = 32'hcdce8364;
    ram_cell[   45241] = 32'h3d599576;
    ram_cell[   45242] = 32'ha15fcb82;
    ram_cell[   45243] = 32'hbf0df100;
    ram_cell[   45244] = 32'h5abd1051;
    ram_cell[   45245] = 32'h2799fc42;
    ram_cell[   45246] = 32'h3186991b;
    ram_cell[   45247] = 32'h8e5f77e9;
    ram_cell[   45248] = 32'h3194d593;
    ram_cell[   45249] = 32'h74df5006;
    ram_cell[   45250] = 32'h5a37512d;
    ram_cell[   45251] = 32'h2fa47d10;
    ram_cell[   45252] = 32'hf4a0a592;
    ram_cell[   45253] = 32'haaf5c621;
    ram_cell[   45254] = 32'he5f24098;
    ram_cell[   45255] = 32'hce744d99;
    ram_cell[   45256] = 32'h4f54f8ae;
    ram_cell[   45257] = 32'h8922c6bf;
    ram_cell[   45258] = 32'hea9723f6;
    ram_cell[   45259] = 32'he66e4cbf;
    ram_cell[   45260] = 32'hfabc4832;
    ram_cell[   45261] = 32'h2df8325c;
    ram_cell[   45262] = 32'h1f01c5f0;
    ram_cell[   45263] = 32'hb44053e9;
    ram_cell[   45264] = 32'hfe4fc97c;
    ram_cell[   45265] = 32'h7b988617;
    ram_cell[   45266] = 32'hfa558938;
    ram_cell[   45267] = 32'h6f11e4d1;
    ram_cell[   45268] = 32'h01c680ea;
    ram_cell[   45269] = 32'h0f1c9cc5;
    ram_cell[   45270] = 32'hcd8fd4c6;
    ram_cell[   45271] = 32'hb3320fad;
    ram_cell[   45272] = 32'h757e9d8d;
    ram_cell[   45273] = 32'hd7a580fe;
    ram_cell[   45274] = 32'h3c508cfe;
    ram_cell[   45275] = 32'h86977580;
    ram_cell[   45276] = 32'h001b1554;
    ram_cell[   45277] = 32'h0d87a732;
    ram_cell[   45278] = 32'h493ac9e0;
    ram_cell[   45279] = 32'h672adb8b;
    ram_cell[   45280] = 32'hd6d61475;
    ram_cell[   45281] = 32'h247763c6;
    ram_cell[   45282] = 32'h13023489;
    ram_cell[   45283] = 32'heff42f04;
    ram_cell[   45284] = 32'h6795e7a4;
    ram_cell[   45285] = 32'hc69c383a;
    ram_cell[   45286] = 32'h0a3c2365;
    ram_cell[   45287] = 32'h31b91ac2;
    ram_cell[   45288] = 32'h7ec720dc;
    ram_cell[   45289] = 32'hc30d297c;
    ram_cell[   45290] = 32'had4616ee;
    ram_cell[   45291] = 32'h994b1288;
    ram_cell[   45292] = 32'h715d58fd;
    ram_cell[   45293] = 32'hfe3e4f2e;
    ram_cell[   45294] = 32'hd7a22e6f;
    ram_cell[   45295] = 32'hfa11e6ee;
    ram_cell[   45296] = 32'h28e74635;
    ram_cell[   45297] = 32'hdef351bc;
    ram_cell[   45298] = 32'h84d0f4f8;
    ram_cell[   45299] = 32'hf1bbae22;
    ram_cell[   45300] = 32'h94fa2272;
    ram_cell[   45301] = 32'h39519277;
    ram_cell[   45302] = 32'h8e58c948;
    ram_cell[   45303] = 32'h949d604d;
    ram_cell[   45304] = 32'he4f0ecfe;
    ram_cell[   45305] = 32'h4a542edc;
    ram_cell[   45306] = 32'hbd3fde8a;
    ram_cell[   45307] = 32'h1708cc22;
    ram_cell[   45308] = 32'he985f51f;
    ram_cell[   45309] = 32'hf14eb48c;
    ram_cell[   45310] = 32'h1559518a;
    ram_cell[   45311] = 32'h5c134eee;
    ram_cell[   45312] = 32'hf77127f0;
    ram_cell[   45313] = 32'h36fbff41;
    ram_cell[   45314] = 32'hda1f21d7;
    ram_cell[   45315] = 32'hab5b0ddb;
    ram_cell[   45316] = 32'h5753684c;
    ram_cell[   45317] = 32'he5ceb6f3;
    ram_cell[   45318] = 32'h7c38f69b;
    ram_cell[   45319] = 32'h0fcf4a29;
    ram_cell[   45320] = 32'h9dc0abe5;
    ram_cell[   45321] = 32'h2c40dee3;
    ram_cell[   45322] = 32'h9b69b13c;
    ram_cell[   45323] = 32'h5d12f0b0;
    ram_cell[   45324] = 32'h8c50f4a5;
    ram_cell[   45325] = 32'h48cc488a;
    ram_cell[   45326] = 32'h9f8a29d2;
    ram_cell[   45327] = 32'h7a01f54b;
    ram_cell[   45328] = 32'he58803fc;
    ram_cell[   45329] = 32'h78a5f7df;
    ram_cell[   45330] = 32'h01f6f18e;
    ram_cell[   45331] = 32'h6eb7b8ca;
    ram_cell[   45332] = 32'h599c3892;
    ram_cell[   45333] = 32'h317e66be;
    ram_cell[   45334] = 32'h1daa7a7e;
    ram_cell[   45335] = 32'he36dcdf1;
    ram_cell[   45336] = 32'h31cb96ce;
    ram_cell[   45337] = 32'hf919f079;
    ram_cell[   45338] = 32'h19150d40;
    ram_cell[   45339] = 32'hf7f97541;
    ram_cell[   45340] = 32'h54d03f3e;
    ram_cell[   45341] = 32'he7982ccc;
    ram_cell[   45342] = 32'hcd1388d0;
    ram_cell[   45343] = 32'h60977b5a;
    ram_cell[   45344] = 32'hbf74c239;
    ram_cell[   45345] = 32'h487b9d0d;
    ram_cell[   45346] = 32'hb2448fc8;
    ram_cell[   45347] = 32'h204e0918;
    ram_cell[   45348] = 32'h2e548c5d;
    ram_cell[   45349] = 32'h2498f1e9;
    ram_cell[   45350] = 32'hcb005fb9;
    ram_cell[   45351] = 32'hd7000eb7;
    ram_cell[   45352] = 32'h486c44b9;
    ram_cell[   45353] = 32'h2968a090;
    ram_cell[   45354] = 32'haf12f5ef;
    ram_cell[   45355] = 32'h1f7d20be;
    ram_cell[   45356] = 32'h146bc711;
    ram_cell[   45357] = 32'h553ca3cb;
    ram_cell[   45358] = 32'h934db17e;
    ram_cell[   45359] = 32'h9340cd25;
    ram_cell[   45360] = 32'h838688fb;
    ram_cell[   45361] = 32'h5219692a;
    ram_cell[   45362] = 32'hb30de0e5;
    ram_cell[   45363] = 32'h817af2a7;
    ram_cell[   45364] = 32'h2596ee3e;
    ram_cell[   45365] = 32'h17dbd8c1;
    ram_cell[   45366] = 32'h9bc340db;
    ram_cell[   45367] = 32'hc253d8f4;
    ram_cell[   45368] = 32'hddd67f1e;
    ram_cell[   45369] = 32'hcdbac83b;
    ram_cell[   45370] = 32'hcea46505;
    ram_cell[   45371] = 32'hec1164c7;
    ram_cell[   45372] = 32'hd99a45ed;
    ram_cell[   45373] = 32'h06baa619;
    ram_cell[   45374] = 32'hb9aa3559;
    ram_cell[   45375] = 32'h11044624;
    ram_cell[   45376] = 32'h941bd73c;
    ram_cell[   45377] = 32'h5502110c;
    ram_cell[   45378] = 32'h2925598d;
    ram_cell[   45379] = 32'h4d0da92a;
    ram_cell[   45380] = 32'h3919c029;
    ram_cell[   45381] = 32'h07192081;
    ram_cell[   45382] = 32'hb1f76e03;
    ram_cell[   45383] = 32'h04489d2e;
    ram_cell[   45384] = 32'hd5254cde;
    ram_cell[   45385] = 32'hd6c40cf3;
    ram_cell[   45386] = 32'ha0be63c3;
    ram_cell[   45387] = 32'h083afa70;
    ram_cell[   45388] = 32'ha432c7dc;
    ram_cell[   45389] = 32'h8f180934;
    ram_cell[   45390] = 32'h85b04e15;
    ram_cell[   45391] = 32'h1f7becec;
    ram_cell[   45392] = 32'hb8ffd309;
    ram_cell[   45393] = 32'h47705af5;
    ram_cell[   45394] = 32'hab917ec3;
    ram_cell[   45395] = 32'hdbed639c;
    ram_cell[   45396] = 32'h1fceb285;
    ram_cell[   45397] = 32'h43acd162;
    ram_cell[   45398] = 32'hf35bcaab;
    ram_cell[   45399] = 32'h30ef93da;
    ram_cell[   45400] = 32'h5f02b2a3;
    ram_cell[   45401] = 32'hcc86a922;
    ram_cell[   45402] = 32'h69d47d38;
    ram_cell[   45403] = 32'h5d9f51e7;
    ram_cell[   45404] = 32'h15d6758a;
    ram_cell[   45405] = 32'h3a0f7d23;
    ram_cell[   45406] = 32'hf42e1ccf;
    ram_cell[   45407] = 32'h122d1864;
    ram_cell[   45408] = 32'h2a452de2;
    ram_cell[   45409] = 32'hc30d39e6;
    ram_cell[   45410] = 32'h0e493646;
    ram_cell[   45411] = 32'hd497719b;
    ram_cell[   45412] = 32'hc1b7d88a;
    ram_cell[   45413] = 32'h94e7e01d;
    ram_cell[   45414] = 32'h18882d4e;
    ram_cell[   45415] = 32'h661db11a;
    ram_cell[   45416] = 32'hacbb75eb;
    ram_cell[   45417] = 32'hd2efa2a1;
    ram_cell[   45418] = 32'h9f2a560c;
    ram_cell[   45419] = 32'h5539b427;
    ram_cell[   45420] = 32'h627f72ce;
    ram_cell[   45421] = 32'h452175dd;
    ram_cell[   45422] = 32'h4fc3c433;
    ram_cell[   45423] = 32'h47af1475;
    ram_cell[   45424] = 32'ha0e502fb;
    ram_cell[   45425] = 32'hd26d0c63;
    ram_cell[   45426] = 32'h06b65c65;
    ram_cell[   45427] = 32'h77033d43;
    ram_cell[   45428] = 32'hb4c05274;
    ram_cell[   45429] = 32'h59adf07c;
    ram_cell[   45430] = 32'hbf3afacd;
    ram_cell[   45431] = 32'hc4e39edf;
    ram_cell[   45432] = 32'hbc76b08d;
    ram_cell[   45433] = 32'h2989ebb3;
    ram_cell[   45434] = 32'hcc1c01c5;
    ram_cell[   45435] = 32'h1e2385f2;
    ram_cell[   45436] = 32'h96b9bc0e;
    ram_cell[   45437] = 32'h8ee667c5;
    ram_cell[   45438] = 32'h875cb1e2;
    ram_cell[   45439] = 32'hed493942;
    ram_cell[   45440] = 32'hd342e644;
    ram_cell[   45441] = 32'hf688adc4;
    ram_cell[   45442] = 32'h74d20876;
    ram_cell[   45443] = 32'h4b615520;
    ram_cell[   45444] = 32'hab445235;
    ram_cell[   45445] = 32'h586feafc;
    ram_cell[   45446] = 32'h2d48d095;
    ram_cell[   45447] = 32'h3ebab869;
    ram_cell[   45448] = 32'h11b9c002;
    ram_cell[   45449] = 32'h52788a61;
    ram_cell[   45450] = 32'he18e850f;
    ram_cell[   45451] = 32'h4522f414;
    ram_cell[   45452] = 32'h8ae87433;
    ram_cell[   45453] = 32'h5e7e313c;
    ram_cell[   45454] = 32'hfcaa1c11;
    ram_cell[   45455] = 32'h048f9312;
    ram_cell[   45456] = 32'hbce40b8c;
    ram_cell[   45457] = 32'hb3de32e9;
    ram_cell[   45458] = 32'h6e0c9e5e;
    ram_cell[   45459] = 32'hf41ce227;
    ram_cell[   45460] = 32'hd37d3edc;
    ram_cell[   45461] = 32'hde3872f5;
    ram_cell[   45462] = 32'h2a4ac4de;
    ram_cell[   45463] = 32'h4e6a760f;
    ram_cell[   45464] = 32'h07a22a7f;
    ram_cell[   45465] = 32'h4fae8fa2;
    ram_cell[   45466] = 32'h81b44458;
    ram_cell[   45467] = 32'hfbf0f751;
    ram_cell[   45468] = 32'hc45c8d0f;
    ram_cell[   45469] = 32'hbfb6728a;
    ram_cell[   45470] = 32'h3eb3350f;
    ram_cell[   45471] = 32'h33b275f0;
    ram_cell[   45472] = 32'h4344bb39;
    ram_cell[   45473] = 32'he053fc68;
    ram_cell[   45474] = 32'hcae1647a;
    ram_cell[   45475] = 32'h0e37da28;
    ram_cell[   45476] = 32'h614af60a;
    ram_cell[   45477] = 32'h0003bb14;
    ram_cell[   45478] = 32'ha9402e89;
    ram_cell[   45479] = 32'h1797fdeb;
    ram_cell[   45480] = 32'h15bc01c5;
    ram_cell[   45481] = 32'hbe8845a9;
    ram_cell[   45482] = 32'hd7688d3f;
    ram_cell[   45483] = 32'h7bec9163;
    ram_cell[   45484] = 32'hc9e2ec9c;
    ram_cell[   45485] = 32'heefa30a2;
    ram_cell[   45486] = 32'hb38840fd;
    ram_cell[   45487] = 32'h6f152fc0;
    ram_cell[   45488] = 32'h28d2b540;
    ram_cell[   45489] = 32'h9fd67226;
    ram_cell[   45490] = 32'h0847236d;
    ram_cell[   45491] = 32'h69416ba8;
    ram_cell[   45492] = 32'h34bf9a17;
    ram_cell[   45493] = 32'hd6b9e3e2;
    ram_cell[   45494] = 32'h1422d187;
    ram_cell[   45495] = 32'hdcd38f4a;
    ram_cell[   45496] = 32'h8c19659c;
    ram_cell[   45497] = 32'ha826a044;
    ram_cell[   45498] = 32'hdaf0b1cc;
    ram_cell[   45499] = 32'hdbdf291a;
    ram_cell[   45500] = 32'h8b2fe797;
    ram_cell[   45501] = 32'h239e1781;
    ram_cell[   45502] = 32'hc9595dff;
    ram_cell[   45503] = 32'hb89e2c1c;
    ram_cell[   45504] = 32'hf792c43a;
    ram_cell[   45505] = 32'h505e7584;
    ram_cell[   45506] = 32'he5b3d36c;
    ram_cell[   45507] = 32'h6e835e6b;
    ram_cell[   45508] = 32'h35ccaab7;
    ram_cell[   45509] = 32'h762d9bbf;
    ram_cell[   45510] = 32'h1e4a4275;
    ram_cell[   45511] = 32'h82e3ea4f;
    ram_cell[   45512] = 32'h03ed77ba;
    ram_cell[   45513] = 32'h81c7738b;
    ram_cell[   45514] = 32'hf45241ea;
    ram_cell[   45515] = 32'hfd5ca76b;
    ram_cell[   45516] = 32'h33f7ef30;
    ram_cell[   45517] = 32'h3c820da3;
    ram_cell[   45518] = 32'h7f902920;
    ram_cell[   45519] = 32'he72a5fbe;
    ram_cell[   45520] = 32'h7c9b5c4f;
    ram_cell[   45521] = 32'h124c71de;
    ram_cell[   45522] = 32'heea0e372;
    ram_cell[   45523] = 32'hf870f6f2;
    ram_cell[   45524] = 32'h3b1a6c96;
    ram_cell[   45525] = 32'hc3a047f3;
    ram_cell[   45526] = 32'h84d7fef1;
    ram_cell[   45527] = 32'hd2f32e8d;
    ram_cell[   45528] = 32'h680012ab;
    ram_cell[   45529] = 32'hfd4c257a;
    ram_cell[   45530] = 32'h7157c8e0;
    ram_cell[   45531] = 32'hc2405573;
    ram_cell[   45532] = 32'h67453e56;
    ram_cell[   45533] = 32'hc022c5f7;
    ram_cell[   45534] = 32'h28212e47;
    ram_cell[   45535] = 32'hab30a5f7;
    ram_cell[   45536] = 32'h22cd16ca;
    ram_cell[   45537] = 32'h9427b590;
    ram_cell[   45538] = 32'h2d4593cb;
    ram_cell[   45539] = 32'h95ff88c1;
    ram_cell[   45540] = 32'h2d877351;
    ram_cell[   45541] = 32'h7d3a0d97;
    ram_cell[   45542] = 32'h325f2e20;
    ram_cell[   45543] = 32'h32e4300f;
    ram_cell[   45544] = 32'h03b82f73;
    ram_cell[   45545] = 32'h14367cfc;
    ram_cell[   45546] = 32'h0151e34c;
    ram_cell[   45547] = 32'hb986ce2c;
    ram_cell[   45548] = 32'hc7300240;
    ram_cell[   45549] = 32'hc0f1fd72;
    ram_cell[   45550] = 32'hc2bb6203;
    ram_cell[   45551] = 32'h19bc076b;
    ram_cell[   45552] = 32'hd884a0b9;
    ram_cell[   45553] = 32'h0ce9808e;
    ram_cell[   45554] = 32'he7139e39;
    ram_cell[   45555] = 32'hd8050461;
    ram_cell[   45556] = 32'h8fa272c5;
    ram_cell[   45557] = 32'h45df64ad;
    ram_cell[   45558] = 32'h1a71ec0b;
    ram_cell[   45559] = 32'h55ea385c;
    ram_cell[   45560] = 32'h9c1a20e6;
    ram_cell[   45561] = 32'he4e174e6;
    ram_cell[   45562] = 32'h1f6b4c55;
    ram_cell[   45563] = 32'hfd24e621;
    ram_cell[   45564] = 32'hc54d5bfd;
    ram_cell[   45565] = 32'h70a321f4;
    ram_cell[   45566] = 32'h9f46d11f;
    ram_cell[   45567] = 32'h95007159;
    ram_cell[   45568] = 32'hefba446d;
    ram_cell[   45569] = 32'h3f6dbaaf;
    ram_cell[   45570] = 32'h0d765de2;
    ram_cell[   45571] = 32'h57e52af2;
    ram_cell[   45572] = 32'h537c6704;
    ram_cell[   45573] = 32'h8710cc4d;
    ram_cell[   45574] = 32'h051cbd29;
    ram_cell[   45575] = 32'hee112a53;
    ram_cell[   45576] = 32'he4837cf0;
    ram_cell[   45577] = 32'hf4ec7d36;
    ram_cell[   45578] = 32'hf1f37ac2;
    ram_cell[   45579] = 32'h3b246f69;
    ram_cell[   45580] = 32'h6a427ca2;
    ram_cell[   45581] = 32'hc7b76cb8;
    ram_cell[   45582] = 32'h0f7adddf;
    ram_cell[   45583] = 32'h39eb2564;
    ram_cell[   45584] = 32'h49367ad6;
    ram_cell[   45585] = 32'h2520ddbf;
    ram_cell[   45586] = 32'h9fe1faa3;
    ram_cell[   45587] = 32'hfc27ebd2;
    ram_cell[   45588] = 32'h2bd72861;
    ram_cell[   45589] = 32'hd54cb6bd;
    ram_cell[   45590] = 32'hdf3ab7fc;
    ram_cell[   45591] = 32'hc1f8c77b;
    ram_cell[   45592] = 32'h267f789b;
    ram_cell[   45593] = 32'h38b17d2f;
    ram_cell[   45594] = 32'h2186d093;
    ram_cell[   45595] = 32'he345de23;
    ram_cell[   45596] = 32'h95e06d70;
    ram_cell[   45597] = 32'h9d58e94b;
    ram_cell[   45598] = 32'hacd5b6d7;
    ram_cell[   45599] = 32'h7a7df6d5;
    ram_cell[   45600] = 32'hd11b64f5;
    ram_cell[   45601] = 32'hf51cdebb;
    ram_cell[   45602] = 32'h616ee2b5;
    ram_cell[   45603] = 32'hdbaac58e;
    ram_cell[   45604] = 32'h1ae344e2;
    ram_cell[   45605] = 32'h1cf45320;
    ram_cell[   45606] = 32'hc1a26db5;
    ram_cell[   45607] = 32'h4ecb8b65;
    ram_cell[   45608] = 32'hf32b2d91;
    ram_cell[   45609] = 32'hd9131245;
    ram_cell[   45610] = 32'hfa5dc56d;
    ram_cell[   45611] = 32'h90003716;
    ram_cell[   45612] = 32'he2ba3c45;
    ram_cell[   45613] = 32'h213a8840;
    ram_cell[   45614] = 32'h80ab4822;
    ram_cell[   45615] = 32'h2181532f;
    ram_cell[   45616] = 32'h42039b04;
    ram_cell[   45617] = 32'h644521a2;
    ram_cell[   45618] = 32'hb8fe1aec;
    ram_cell[   45619] = 32'hf7bb1dc3;
    ram_cell[   45620] = 32'h290395c8;
    ram_cell[   45621] = 32'h36dfca37;
    ram_cell[   45622] = 32'he77e4592;
    ram_cell[   45623] = 32'h07e1c7bc;
    ram_cell[   45624] = 32'he6ae11d0;
    ram_cell[   45625] = 32'h2db527c1;
    ram_cell[   45626] = 32'h8ae0f18c;
    ram_cell[   45627] = 32'h44880a99;
    ram_cell[   45628] = 32'h4b68eefc;
    ram_cell[   45629] = 32'hd62bd31c;
    ram_cell[   45630] = 32'h5ddf323d;
    ram_cell[   45631] = 32'h07b5cb28;
    ram_cell[   45632] = 32'h77bf039b;
    ram_cell[   45633] = 32'h4676e8da;
    ram_cell[   45634] = 32'he635f312;
    ram_cell[   45635] = 32'h22ffa7d3;
    ram_cell[   45636] = 32'ha93c0a5e;
    ram_cell[   45637] = 32'h3e2489ad;
    ram_cell[   45638] = 32'h44157b79;
    ram_cell[   45639] = 32'h85f0f12c;
    ram_cell[   45640] = 32'h80f09053;
    ram_cell[   45641] = 32'h5d416fec;
    ram_cell[   45642] = 32'h95ad1236;
    ram_cell[   45643] = 32'h8b0b6253;
    ram_cell[   45644] = 32'h144e2ce9;
    ram_cell[   45645] = 32'h895c6b12;
    ram_cell[   45646] = 32'h754ecd55;
    ram_cell[   45647] = 32'h71df586a;
    ram_cell[   45648] = 32'hfb6dc7bf;
    ram_cell[   45649] = 32'h9ffb3ed9;
    ram_cell[   45650] = 32'ha7d40db6;
    ram_cell[   45651] = 32'h666646e2;
    ram_cell[   45652] = 32'h7a52db74;
    ram_cell[   45653] = 32'h1fde7471;
    ram_cell[   45654] = 32'hb8b19c3a;
    ram_cell[   45655] = 32'h9bbdd612;
    ram_cell[   45656] = 32'h8fe9094a;
    ram_cell[   45657] = 32'h2a149961;
    ram_cell[   45658] = 32'h5d2bb19e;
    ram_cell[   45659] = 32'hcc00b284;
    ram_cell[   45660] = 32'h29456188;
    ram_cell[   45661] = 32'hd1447aba;
    ram_cell[   45662] = 32'ha56bb098;
    ram_cell[   45663] = 32'h1f110844;
    ram_cell[   45664] = 32'h657d7cc8;
    ram_cell[   45665] = 32'hbe237718;
    ram_cell[   45666] = 32'hd53947da;
    ram_cell[   45667] = 32'h56d6588b;
    ram_cell[   45668] = 32'h30f92d24;
    ram_cell[   45669] = 32'h0ed67b97;
    ram_cell[   45670] = 32'h7cc96494;
    ram_cell[   45671] = 32'h108c54bb;
    ram_cell[   45672] = 32'hb6cd8d02;
    ram_cell[   45673] = 32'h5d26390b;
    ram_cell[   45674] = 32'h4348d8a6;
    ram_cell[   45675] = 32'h36be175e;
    ram_cell[   45676] = 32'hca8e2763;
    ram_cell[   45677] = 32'h4c23b795;
    ram_cell[   45678] = 32'he83e6412;
    ram_cell[   45679] = 32'h2e64a70a;
    ram_cell[   45680] = 32'h30c867aa;
    ram_cell[   45681] = 32'he79a2452;
    ram_cell[   45682] = 32'h687843b3;
    ram_cell[   45683] = 32'h3ca6a74c;
    ram_cell[   45684] = 32'hb88611c4;
    ram_cell[   45685] = 32'h9e1b5385;
    ram_cell[   45686] = 32'h29d533b7;
    ram_cell[   45687] = 32'h445f711c;
    ram_cell[   45688] = 32'hc55532be;
    ram_cell[   45689] = 32'hf873520c;
    ram_cell[   45690] = 32'h862c7016;
    ram_cell[   45691] = 32'h37cbe02a;
    ram_cell[   45692] = 32'h2e9975c2;
    ram_cell[   45693] = 32'h1855afe5;
    ram_cell[   45694] = 32'haca921b0;
    ram_cell[   45695] = 32'h8f9840d4;
    ram_cell[   45696] = 32'hfd62e39a;
    ram_cell[   45697] = 32'h0d1f2f00;
    ram_cell[   45698] = 32'hb971303f;
    ram_cell[   45699] = 32'h442567de;
    ram_cell[   45700] = 32'h3fdc4a46;
    ram_cell[   45701] = 32'h40ddd720;
    ram_cell[   45702] = 32'hbd3ca160;
    ram_cell[   45703] = 32'h54e63c72;
    ram_cell[   45704] = 32'h78ae904c;
    ram_cell[   45705] = 32'h62b022c0;
    ram_cell[   45706] = 32'h77c08ae0;
    ram_cell[   45707] = 32'hed832239;
    ram_cell[   45708] = 32'h5b50e233;
    ram_cell[   45709] = 32'h641c18fd;
    ram_cell[   45710] = 32'hd0bd71d2;
    ram_cell[   45711] = 32'hf08100d7;
    ram_cell[   45712] = 32'hfb271648;
    ram_cell[   45713] = 32'hcfa12ae1;
    ram_cell[   45714] = 32'h6636d014;
    ram_cell[   45715] = 32'h220a5718;
    ram_cell[   45716] = 32'hbfb825a2;
    ram_cell[   45717] = 32'hebd6b8ad;
    ram_cell[   45718] = 32'h4257d8aa;
    ram_cell[   45719] = 32'h175825e2;
    ram_cell[   45720] = 32'h01479e55;
    ram_cell[   45721] = 32'h2baf5be6;
    ram_cell[   45722] = 32'h1e24e7f1;
    ram_cell[   45723] = 32'ha431c511;
    ram_cell[   45724] = 32'h1ea9bb6d;
    ram_cell[   45725] = 32'h76190c82;
    ram_cell[   45726] = 32'h861f59c6;
    ram_cell[   45727] = 32'h839a64e5;
    ram_cell[   45728] = 32'h1987a0d0;
    ram_cell[   45729] = 32'h5c4a1d03;
    ram_cell[   45730] = 32'h943c7407;
    ram_cell[   45731] = 32'h35d00205;
    ram_cell[   45732] = 32'h7d455566;
    ram_cell[   45733] = 32'h744a9199;
    ram_cell[   45734] = 32'h7818cbd1;
    ram_cell[   45735] = 32'h3c3db0a7;
    ram_cell[   45736] = 32'h4496db19;
    ram_cell[   45737] = 32'h8e1d1a4c;
    ram_cell[   45738] = 32'hd809d027;
    ram_cell[   45739] = 32'h5027520f;
    ram_cell[   45740] = 32'haeeb8e1a;
    ram_cell[   45741] = 32'hd2457bc2;
    ram_cell[   45742] = 32'h7ac2b8c7;
    ram_cell[   45743] = 32'h65708568;
    ram_cell[   45744] = 32'h6f2dd41f;
    ram_cell[   45745] = 32'h492b47bb;
    ram_cell[   45746] = 32'hb09c1f97;
    ram_cell[   45747] = 32'h9859378e;
    ram_cell[   45748] = 32'hfbfc2ce5;
    ram_cell[   45749] = 32'hfbeae8ce;
    ram_cell[   45750] = 32'h2982c0fc;
    ram_cell[   45751] = 32'h3ad94aa0;
    ram_cell[   45752] = 32'h603ee619;
    ram_cell[   45753] = 32'hcfb57c11;
    ram_cell[   45754] = 32'he5117f45;
    ram_cell[   45755] = 32'h69d576d8;
    ram_cell[   45756] = 32'h12403a9f;
    ram_cell[   45757] = 32'hb2769a8c;
    ram_cell[   45758] = 32'hee4aac8f;
    ram_cell[   45759] = 32'h4170fbb6;
    ram_cell[   45760] = 32'h69738c05;
    ram_cell[   45761] = 32'head64c0e;
    ram_cell[   45762] = 32'hae28f492;
    ram_cell[   45763] = 32'hb065521b;
    ram_cell[   45764] = 32'h825b4105;
    ram_cell[   45765] = 32'h7d01bd3f;
    ram_cell[   45766] = 32'h4c8a26cb;
    ram_cell[   45767] = 32'hd4da5854;
    ram_cell[   45768] = 32'hb53b4777;
    ram_cell[   45769] = 32'h570ba2a5;
    ram_cell[   45770] = 32'h0d187972;
    ram_cell[   45771] = 32'h42df029a;
    ram_cell[   45772] = 32'h3a2881b1;
    ram_cell[   45773] = 32'hca2746f9;
    ram_cell[   45774] = 32'hc7639edc;
    ram_cell[   45775] = 32'hf0d296dd;
    ram_cell[   45776] = 32'h469a77bb;
    ram_cell[   45777] = 32'h48075a82;
    ram_cell[   45778] = 32'h7fc5d280;
    ram_cell[   45779] = 32'h506826e3;
    ram_cell[   45780] = 32'hc484a2ce;
    ram_cell[   45781] = 32'h77e74cee;
    ram_cell[   45782] = 32'h7b71476b;
    ram_cell[   45783] = 32'he60d6244;
    ram_cell[   45784] = 32'h539da1ce;
    ram_cell[   45785] = 32'h8fe41b2c;
    ram_cell[   45786] = 32'hba2f3d52;
    ram_cell[   45787] = 32'h2c543d6c;
    ram_cell[   45788] = 32'he45cba24;
    ram_cell[   45789] = 32'hc98d6fa4;
    ram_cell[   45790] = 32'h9a2649bd;
    ram_cell[   45791] = 32'hd2739e28;
    ram_cell[   45792] = 32'hf68e3f1f;
    ram_cell[   45793] = 32'h0306a19e;
    ram_cell[   45794] = 32'h000bbcbb;
    ram_cell[   45795] = 32'hda1fb4d0;
    ram_cell[   45796] = 32'h406d0d37;
    ram_cell[   45797] = 32'hf36348fc;
    ram_cell[   45798] = 32'h8a3df634;
    ram_cell[   45799] = 32'h9bf4850a;
    ram_cell[   45800] = 32'h0beb3673;
    ram_cell[   45801] = 32'h57da1cef;
    ram_cell[   45802] = 32'h9a74eea6;
    ram_cell[   45803] = 32'h2eded2c9;
    ram_cell[   45804] = 32'hda1c4861;
    ram_cell[   45805] = 32'h1886bf8a;
    ram_cell[   45806] = 32'h795a2bea;
    ram_cell[   45807] = 32'ha614f97a;
    ram_cell[   45808] = 32'h68c859c4;
    ram_cell[   45809] = 32'ha08905e5;
    ram_cell[   45810] = 32'hadd39401;
    ram_cell[   45811] = 32'h18e807c3;
    ram_cell[   45812] = 32'h38b36562;
    ram_cell[   45813] = 32'h8719e2f3;
    ram_cell[   45814] = 32'h9b1129a2;
    ram_cell[   45815] = 32'hc15510d5;
    ram_cell[   45816] = 32'h633859e5;
    ram_cell[   45817] = 32'h65e9909b;
    ram_cell[   45818] = 32'hd8018fad;
    ram_cell[   45819] = 32'h86c2823c;
    ram_cell[   45820] = 32'hd56524b3;
    ram_cell[   45821] = 32'hdd8a12b0;
    ram_cell[   45822] = 32'h01d1d78a;
    ram_cell[   45823] = 32'h6f0a2c59;
    ram_cell[   45824] = 32'hea17b332;
    ram_cell[   45825] = 32'hca3f6199;
    ram_cell[   45826] = 32'h3302fa47;
    ram_cell[   45827] = 32'h15d0ffbc;
    ram_cell[   45828] = 32'hca11fd6b;
    ram_cell[   45829] = 32'h8c80fb91;
    ram_cell[   45830] = 32'h6d725f8d;
    ram_cell[   45831] = 32'hb9119c3c;
    ram_cell[   45832] = 32'h97de366e;
    ram_cell[   45833] = 32'hb4d7be94;
    ram_cell[   45834] = 32'h22f7f4bc;
    ram_cell[   45835] = 32'h718986aa;
    ram_cell[   45836] = 32'h6b70cdc4;
    ram_cell[   45837] = 32'h4d9986c2;
    ram_cell[   45838] = 32'h70cb7b53;
    ram_cell[   45839] = 32'h53e79f3b;
    ram_cell[   45840] = 32'h6ff69104;
    ram_cell[   45841] = 32'h6eed6dc5;
    ram_cell[   45842] = 32'hcd9f860e;
    ram_cell[   45843] = 32'h623c4ba6;
    ram_cell[   45844] = 32'h3103c8fe;
    ram_cell[   45845] = 32'h75f3cde5;
    ram_cell[   45846] = 32'he49c58f3;
    ram_cell[   45847] = 32'h5e3005c8;
    ram_cell[   45848] = 32'h10d0fdf7;
    ram_cell[   45849] = 32'hdfb5aaab;
    ram_cell[   45850] = 32'h86ae0fc8;
    ram_cell[   45851] = 32'h22fa150e;
    ram_cell[   45852] = 32'h0cc138e2;
    ram_cell[   45853] = 32'h5364c310;
    ram_cell[   45854] = 32'hee6c4151;
    ram_cell[   45855] = 32'h9f1b6bfc;
    ram_cell[   45856] = 32'h1c54db24;
    ram_cell[   45857] = 32'h0e22182b;
    ram_cell[   45858] = 32'hce47996c;
    ram_cell[   45859] = 32'h108fe4ed;
    ram_cell[   45860] = 32'h575a95e0;
    ram_cell[   45861] = 32'h1fab67ca;
    ram_cell[   45862] = 32'h92ed0560;
    ram_cell[   45863] = 32'hefea6916;
    ram_cell[   45864] = 32'heb879379;
    ram_cell[   45865] = 32'h09aa9cdb;
    ram_cell[   45866] = 32'hb225b99b;
    ram_cell[   45867] = 32'h0b73f13b;
    ram_cell[   45868] = 32'hf9acc5d9;
    ram_cell[   45869] = 32'h6de7075e;
    ram_cell[   45870] = 32'hc526eb9c;
    ram_cell[   45871] = 32'h43769746;
    ram_cell[   45872] = 32'hd408d77a;
    ram_cell[   45873] = 32'ha90825a0;
    ram_cell[   45874] = 32'h9418bb19;
    ram_cell[   45875] = 32'h24164113;
    ram_cell[   45876] = 32'hf760baf4;
    ram_cell[   45877] = 32'h61298419;
    ram_cell[   45878] = 32'h86025884;
    ram_cell[   45879] = 32'hae72f8e7;
    ram_cell[   45880] = 32'h4d280e44;
    ram_cell[   45881] = 32'h0aa085bf;
    ram_cell[   45882] = 32'hbfab0c1b;
    ram_cell[   45883] = 32'hae0068cc;
    ram_cell[   45884] = 32'ha7421bfe;
    ram_cell[   45885] = 32'h8a1d133f;
    ram_cell[   45886] = 32'h99ba74ef;
    ram_cell[   45887] = 32'h9a3cab30;
    ram_cell[   45888] = 32'hdef8d4cb;
    ram_cell[   45889] = 32'h2a874fa2;
    ram_cell[   45890] = 32'hbd8d1750;
    ram_cell[   45891] = 32'h5f142d5c;
    ram_cell[   45892] = 32'h26e15f05;
    ram_cell[   45893] = 32'h7d2d7eaf;
    ram_cell[   45894] = 32'hbd32c57f;
    ram_cell[   45895] = 32'hc6701341;
    ram_cell[   45896] = 32'h743e2318;
    ram_cell[   45897] = 32'h5c1ab760;
    ram_cell[   45898] = 32'h68ba980d;
    ram_cell[   45899] = 32'hedc5f777;
    ram_cell[   45900] = 32'hfe196b82;
    ram_cell[   45901] = 32'h53b60669;
    ram_cell[   45902] = 32'h4eea539e;
    ram_cell[   45903] = 32'h39c087b4;
    ram_cell[   45904] = 32'ha55e6051;
    ram_cell[   45905] = 32'h13bf55d3;
    ram_cell[   45906] = 32'hdbffc98c;
    ram_cell[   45907] = 32'hb8d34cf8;
    ram_cell[   45908] = 32'hd73be734;
    ram_cell[   45909] = 32'hca85c4b9;
    ram_cell[   45910] = 32'h5a103c6f;
    ram_cell[   45911] = 32'h7aaac7e8;
    ram_cell[   45912] = 32'h5e450fee;
    ram_cell[   45913] = 32'h803d6bb0;
    ram_cell[   45914] = 32'h31d82ed5;
    ram_cell[   45915] = 32'h83680194;
    ram_cell[   45916] = 32'h089ff905;
    ram_cell[   45917] = 32'h0c295457;
    ram_cell[   45918] = 32'hf426839f;
    ram_cell[   45919] = 32'he8588d09;
    ram_cell[   45920] = 32'ha4f1770b;
    ram_cell[   45921] = 32'hf835811f;
    ram_cell[   45922] = 32'h09534d09;
    ram_cell[   45923] = 32'h3e7e8bad;
    ram_cell[   45924] = 32'hc4f38736;
    ram_cell[   45925] = 32'h7febb95a;
    ram_cell[   45926] = 32'hddd65ae0;
    ram_cell[   45927] = 32'ha8cf77c8;
    ram_cell[   45928] = 32'h5511dd45;
    ram_cell[   45929] = 32'he9c4ec74;
    ram_cell[   45930] = 32'hd263d7aa;
    ram_cell[   45931] = 32'hf4334483;
    ram_cell[   45932] = 32'hc6e0cc25;
    ram_cell[   45933] = 32'hdffaff1f;
    ram_cell[   45934] = 32'h513591e5;
    ram_cell[   45935] = 32'heaa08481;
    ram_cell[   45936] = 32'hcc737037;
    ram_cell[   45937] = 32'h91560797;
    ram_cell[   45938] = 32'h263bbb6c;
    ram_cell[   45939] = 32'h5aec3166;
    ram_cell[   45940] = 32'h8f651012;
    ram_cell[   45941] = 32'he32a67c8;
    ram_cell[   45942] = 32'h9151440c;
    ram_cell[   45943] = 32'h0f72932c;
    ram_cell[   45944] = 32'h13638453;
    ram_cell[   45945] = 32'h10c7b9ce;
    ram_cell[   45946] = 32'h2f4727ea;
    ram_cell[   45947] = 32'h5b72abb6;
    ram_cell[   45948] = 32'h43f207c1;
    ram_cell[   45949] = 32'h2bc6377b;
    ram_cell[   45950] = 32'h1f069e29;
    ram_cell[   45951] = 32'h94656e62;
    ram_cell[   45952] = 32'h16bd405f;
    ram_cell[   45953] = 32'h35ad35a8;
    ram_cell[   45954] = 32'h575f70c9;
    ram_cell[   45955] = 32'h71087024;
    ram_cell[   45956] = 32'hbd2a8842;
    ram_cell[   45957] = 32'hf08c4766;
    ram_cell[   45958] = 32'h1708e57e;
    ram_cell[   45959] = 32'h33037f2f;
    ram_cell[   45960] = 32'h83e9a925;
    ram_cell[   45961] = 32'h958ab721;
    ram_cell[   45962] = 32'hbd483128;
    ram_cell[   45963] = 32'h7c4aebf9;
    ram_cell[   45964] = 32'ha45953b5;
    ram_cell[   45965] = 32'h7f543869;
    ram_cell[   45966] = 32'h8a495e60;
    ram_cell[   45967] = 32'hc7b08ca3;
    ram_cell[   45968] = 32'h85cca863;
    ram_cell[   45969] = 32'h716cc973;
    ram_cell[   45970] = 32'ha4f542f9;
    ram_cell[   45971] = 32'h6a35bd85;
    ram_cell[   45972] = 32'hed1be0e0;
    ram_cell[   45973] = 32'hfecdf93d;
    ram_cell[   45974] = 32'h79c6bb92;
    ram_cell[   45975] = 32'he9e71ffd;
    ram_cell[   45976] = 32'hdd3c6bb6;
    ram_cell[   45977] = 32'h77456b3d;
    ram_cell[   45978] = 32'h1aa9ba97;
    ram_cell[   45979] = 32'he6c6d7a8;
    ram_cell[   45980] = 32'h1406f822;
    ram_cell[   45981] = 32'hb5a378f4;
    ram_cell[   45982] = 32'ha7ed2659;
    ram_cell[   45983] = 32'h1a23c908;
    ram_cell[   45984] = 32'h17eb93e6;
    ram_cell[   45985] = 32'h298e1bd3;
    ram_cell[   45986] = 32'he048a9fb;
    ram_cell[   45987] = 32'hdc5cf8e6;
    ram_cell[   45988] = 32'hfdf766b6;
    ram_cell[   45989] = 32'h3a168cca;
    ram_cell[   45990] = 32'h17739b0a;
    ram_cell[   45991] = 32'h66734c8d;
    ram_cell[   45992] = 32'h22d163ee;
    ram_cell[   45993] = 32'h79bf48b6;
    ram_cell[   45994] = 32'h637c30e9;
    ram_cell[   45995] = 32'h16eb95d3;
    ram_cell[   45996] = 32'h74e1038e;
    ram_cell[   45997] = 32'h7a1001b7;
    ram_cell[   45998] = 32'h62f90d30;
    ram_cell[   45999] = 32'hf1d7237d;
    ram_cell[   46000] = 32'h53c7d6c9;
    ram_cell[   46001] = 32'h3e5328b4;
    ram_cell[   46002] = 32'h929190a3;
    ram_cell[   46003] = 32'hc656fa08;
    ram_cell[   46004] = 32'h3a35315c;
    ram_cell[   46005] = 32'h46aec7b5;
    ram_cell[   46006] = 32'h24206db3;
    ram_cell[   46007] = 32'hf07fa47e;
    ram_cell[   46008] = 32'h2b7c2597;
    ram_cell[   46009] = 32'ha9db63ab;
    ram_cell[   46010] = 32'h5055b6cc;
    ram_cell[   46011] = 32'h8fb370c5;
    ram_cell[   46012] = 32'hf783014a;
    ram_cell[   46013] = 32'h45f07458;
    ram_cell[   46014] = 32'h474a1c9f;
    ram_cell[   46015] = 32'h76d07216;
    ram_cell[   46016] = 32'h76b4b84e;
    ram_cell[   46017] = 32'h03620d03;
    ram_cell[   46018] = 32'hd9260f75;
    ram_cell[   46019] = 32'h8e05df81;
    ram_cell[   46020] = 32'hb7e07cd9;
    ram_cell[   46021] = 32'he1da2ed3;
    ram_cell[   46022] = 32'hd4dd339e;
    ram_cell[   46023] = 32'h12415b77;
    ram_cell[   46024] = 32'he533e536;
    ram_cell[   46025] = 32'h6083afff;
    ram_cell[   46026] = 32'h9954289b;
    ram_cell[   46027] = 32'h84a1d02f;
    ram_cell[   46028] = 32'hd719ec12;
    ram_cell[   46029] = 32'h69763c8a;
    ram_cell[   46030] = 32'hb7020077;
    ram_cell[   46031] = 32'h584dbafc;
    ram_cell[   46032] = 32'ha79ce82b;
    ram_cell[   46033] = 32'h3c312531;
    ram_cell[   46034] = 32'h30938106;
    ram_cell[   46035] = 32'h8bb69040;
    ram_cell[   46036] = 32'he44552be;
    ram_cell[   46037] = 32'h7bce0276;
    ram_cell[   46038] = 32'h572c695f;
    ram_cell[   46039] = 32'h53b1142c;
    ram_cell[   46040] = 32'h8fe76cd6;
    ram_cell[   46041] = 32'hb57b413f;
    ram_cell[   46042] = 32'h674650f2;
    ram_cell[   46043] = 32'hd5c32cac;
    ram_cell[   46044] = 32'h64d5e545;
    ram_cell[   46045] = 32'h6a159545;
    ram_cell[   46046] = 32'h78e1c3a0;
    ram_cell[   46047] = 32'hc38ca2b6;
    ram_cell[   46048] = 32'h04ca0053;
    ram_cell[   46049] = 32'heb9ac911;
    ram_cell[   46050] = 32'h0a4e751a;
    ram_cell[   46051] = 32'he84c16e6;
    ram_cell[   46052] = 32'h95054cc0;
    ram_cell[   46053] = 32'h3b86245d;
    ram_cell[   46054] = 32'h4c56971f;
    ram_cell[   46055] = 32'hcc7774a5;
    ram_cell[   46056] = 32'h0fe2ac98;
    ram_cell[   46057] = 32'hf50aeaaa;
    ram_cell[   46058] = 32'h5ed98023;
    ram_cell[   46059] = 32'ha995d898;
    ram_cell[   46060] = 32'h2b24b987;
    ram_cell[   46061] = 32'h079e1bb8;
    ram_cell[   46062] = 32'h1ad90e4e;
    ram_cell[   46063] = 32'h67c659ee;
    ram_cell[   46064] = 32'hdca07c36;
    ram_cell[   46065] = 32'hfca2ba5a;
    ram_cell[   46066] = 32'hee534241;
    ram_cell[   46067] = 32'h4d6970a7;
    ram_cell[   46068] = 32'h2a0874ce;
    ram_cell[   46069] = 32'h74085fbb;
    ram_cell[   46070] = 32'hc7055810;
    ram_cell[   46071] = 32'he54451f6;
    ram_cell[   46072] = 32'h2b60eefa;
    ram_cell[   46073] = 32'h8023158d;
    ram_cell[   46074] = 32'hf38dc0cf;
    ram_cell[   46075] = 32'hfae0e350;
    ram_cell[   46076] = 32'h1f217720;
    ram_cell[   46077] = 32'h65179063;
    ram_cell[   46078] = 32'haf5a24c3;
    ram_cell[   46079] = 32'h934f50e1;
    ram_cell[   46080] = 32'h890c5082;
    ram_cell[   46081] = 32'h59488ea3;
    ram_cell[   46082] = 32'h0cf18f99;
    ram_cell[   46083] = 32'hbd9c6158;
    ram_cell[   46084] = 32'h131a220d;
    ram_cell[   46085] = 32'h49c2fdc1;
    ram_cell[   46086] = 32'hbad24fc8;
    ram_cell[   46087] = 32'h08671594;
    ram_cell[   46088] = 32'hc4036e75;
    ram_cell[   46089] = 32'h845c042e;
    ram_cell[   46090] = 32'h4ff8a927;
    ram_cell[   46091] = 32'hef02afc6;
    ram_cell[   46092] = 32'h09dc94ad;
    ram_cell[   46093] = 32'hcd9383c9;
    ram_cell[   46094] = 32'h283350ac;
    ram_cell[   46095] = 32'h1a5c40f1;
    ram_cell[   46096] = 32'ha19ed16a;
    ram_cell[   46097] = 32'h28a5528d;
    ram_cell[   46098] = 32'h7ff53b16;
    ram_cell[   46099] = 32'h872a6fe0;
    ram_cell[   46100] = 32'h59ebe775;
    ram_cell[   46101] = 32'h9200adee;
    ram_cell[   46102] = 32'ha720f4bd;
    ram_cell[   46103] = 32'h7401a8e9;
    ram_cell[   46104] = 32'h5e670531;
    ram_cell[   46105] = 32'h64fc2ff4;
    ram_cell[   46106] = 32'hcfc3f7c9;
    ram_cell[   46107] = 32'hdc06eeb6;
    ram_cell[   46108] = 32'h3b1e5683;
    ram_cell[   46109] = 32'h1cb3b101;
    ram_cell[   46110] = 32'hc655fc6c;
    ram_cell[   46111] = 32'h32d6d0b4;
    ram_cell[   46112] = 32'h533f6660;
    ram_cell[   46113] = 32'h31ec35a5;
    ram_cell[   46114] = 32'h7e0a171f;
    ram_cell[   46115] = 32'h48729ba0;
    ram_cell[   46116] = 32'h28f4a0d7;
    ram_cell[   46117] = 32'hfabf70f6;
    ram_cell[   46118] = 32'h556860e7;
    ram_cell[   46119] = 32'hb9f426ac;
    ram_cell[   46120] = 32'h6116b390;
    ram_cell[   46121] = 32'hefb7d12b;
    ram_cell[   46122] = 32'hc72a488f;
    ram_cell[   46123] = 32'h7dc8bd29;
    ram_cell[   46124] = 32'h9fbf1148;
    ram_cell[   46125] = 32'h5d3849af;
    ram_cell[   46126] = 32'h2b21b60a;
    ram_cell[   46127] = 32'hb2c07bb7;
    ram_cell[   46128] = 32'hc9bdfd8b;
    ram_cell[   46129] = 32'h34860adf;
    ram_cell[   46130] = 32'h1091196f;
    ram_cell[   46131] = 32'h595f0b7e;
    ram_cell[   46132] = 32'he483753b;
    ram_cell[   46133] = 32'h78552997;
    ram_cell[   46134] = 32'h91771b04;
    ram_cell[   46135] = 32'h26ce1e04;
    ram_cell[   46136] = 32'h366d9f39;
    ram_cell[   46137] = 32'h66379735;
    ram_cell[   46138] = 32'h5df193a4;
    ram_cell[   46139] = 32'h0a985891;
    ram_cell[   46140] = 32'hd5204af9;
    ram_cell[   46141] = 32'hbf8f085a;
    ram_cell[   46142] = 32'hd587c330;
    ram_cell[   46143] = 32'hd629e5ec;
    ram_cell[   46144] = 32'h086cf13d;
    ram_cell[   46145] = 32'h73023bd1;
    ram_cell[   46146] = 32'h78e8d3d1;
    ram_cell[   46147] = 32'h50a1662c;
    ram_cell[   46148] = 32'h4b3df7a2;
    ram_cell[   46149] = 32'h726f3fff;
    ram_cell[   46150] = 32'hacc15a5d;
    ram_cell[   46151] = 32'h0327eca4;
    ram_cell[   46152] = 32'h66af043f;
    ram_cell[   46153] = 32'h26be89b1;
    ram_cell[   46154] = 32'hdafe6dc4;
    ram_cell[   46155] = 32'h66c8d04d;
    ram_cell[   46156] = 32'h76ae40a1;
    ram_cell[   46157] = 32'hb4e65360;
    ram_cell[   46158] = 32'h8ad459ba;
    ram_cell[   46159] = 32'h07603aa3;
    ram_cell[   46160] = 32'h7d4d4645;
    ram_cell[   46161] = 32'hdf1f1982;
    ram_cell[   46162] = 32'hc33a2701;
    ram_cell[   46163] = 32'h2b940543;
    ram_cell[   46164] = 32'hd2a7ec07;
    ram_cell[   46165] = 32'hc12bb60a;
    ram_cell[   46166] = 32'h707fe70c;
    ram_cell[   46167] = 32'h22d80d82;
    ram_cell[   46168] = 32'h3cf87f62;
    ram_cell[   46169] = 32'hc9b8f471;
    ram_cell[   46170] = 32'h5678df52;
    ram_cell[   46171] = 32'h2057dacf;
    ram_cell[   46172] = 32'h6585f616;
    ram_cell[   46173] = 32'hc9f25832;
    ram_cell[   46174] = 32'hcb710293;
    ram_cell[   46175] = 32'h6045adfe;
    ram_cell[   46176] = 32'h1ce92e98;
    ram_cell[   46177] = 32'h733025e7;
    ram_cell[   46178] = 32'hfe754e08;
    ram_cell[   46179] = 32'h32b62936;
    ram_cell[   46180] = 32'h5d2f21c1;
    ram_cell[   46181] = 32'h9ffabec7;
    ram_cell[   46182] = 32'hcf51bdb4;
    ram_cell[   46183] = 32'hac88ba06;
    ram_cell[   46184] = 32'h4020597b;
    ram_cell[   46185] = 32'hcc456bef;
    ram_cell[   46186] = 32'h8aef5780;
    ram_cell[   46187] = 32'hce9cf94f;
    ram_cell[   46188] = 32'h57b802bb;
    ram_cell[   46189] = 32'h63a6e7c3;
    ram_cell[   46190] = 32'he6120638;
    ram_cell[   46191] = 32'h1a3c5b51;
    ram_cell[   46192] = 32'h8b3262ba;
    ram_cell[   46193] = 32'hc1f498b2;
    ram_cell[   46194] = 32'h27b3fc86;
    ram_cell[   46195] = 32'h3a768624;
    ram_cell[   46196] = 32'he35ff3ae;
    ram_cell[   46197] = 32'ha239eebe;
    ram_cell[   46198] = 32'h22e1129f;
    ram_cell[   46199] = 32'hce4648af;
    ram_cell[   46200] = 32'hdbca076a;
    ram_cell[   46201] = 32'hd0d0424e;
    ram_cell[   46202] = 32'hcea5b9f3;
    ram_cell[   46203] = 32'hc95b99b3;
    ram_cell[   46204] = 32'haa2d356a;
    ram_cell[   46205] = 32'h55033539;
    ram_cell[   46206] = 32'h77ba3973;
    ram_cell[   46207] = 32'hb3992a2c;
    ram_cell[   46208] = 32'h83db8330;
    ram_cell[   46209] = 32'hf233187f;
    ram_cell[   46210] = 32'h65f9449c;
    ram_cell[   46211] = 32'h2e4a9a2e;
    ram_cell[   46212] = 32'hc5d5d377;
    ram_cell[   46213] = 32'h69d8963d;
    ram_cell[   46214] = 32'hc08eafce;
    ram_cell[   46215] = 32'h241d5464;
    ram_cell[   46216] = 32'h6131b1b5;
    ram_cell[   46217] = 32'hc3e350bd;
    ram_cell[   46218] = 32'h0afda989;
    ram_cell[   46219] = 32'hc4efc82f;
    ram_cell[   46220] = 32'h11d155ad;
    ram_cell[   46221] = 32'h4f3e7d15;
    ram_cell[   46222] = 32'h5e5926fd;
    ram_cell[   46223] = 32'h64120a20;
    ram_cell[   46224] = 32'h61575708;
    ram_cell[   46225] = 32'h49480b0e;
    ram_cell[   46226] = 32'h51e09449;
    ram_cell[   46227] = 32'h64d1e1a9;
    ram_cell[   46228] = 32'h943cc582;
    ram_cell[   46229] = 32'h94fc8244;
    ram_cell[   46230] = 32'h2f4ca449;
    ram_cell[   46231] = 32'h8633e954;
    ram_cell[   46232] = 32'h19e3fc7a;
    ram_cell[   46233] = 32'hde81d34d;
    ram_cell[   46234] = 32'h2fa5e7b6;
    ram_cell[   46235] = 32'hba0bb1ae;
    ram_cell[   46236] = 32'hf51a5b0f;
    ram_cell[   46237] = 32'h9cbb5c60;
    ram_cell[   46238] = 32'h626712aa;
    ram_cell[   46239] = 32'hc4220ab0;
    ram_cell[   46240] = 32'he62a9ba0;
    ram_cell[   46241] = 32'h322b38f7;
    ram_cell[   46242] = 32'h6a499dbd;
    ram_cell[   46243] = 32'h1220f128;
    ram_cell[   46244] = 32'h41211eb6;
    ram_cell[   46245] = 32'h2afdc17e;
    ram_cell[   46246] = 32'h69f6dc01;
    ram_cell[   46247] = 32'h5308f1bd;
    ram_cell[   46248] = 32'hc1adea7a;
    ram_cell[   46249] = 32'h3e811490;
    ram_cell[   46250] = 32'he8df00b7;
    ram_cell[   46251] = 32'h9d3857b5;
    ram_cell[   46252] = 32'hab25b8d8;
    ram_cell[   46253] = 32'h6e967aef;
    ram_cell[   46254] = 32'hbc7369b0;
    ram_cell[   46255] = 32'h6f4c824f;
    ram_cell[   46256] = 32'h748ac172;
    ram_cell[   46257] = 32'h012e193f;
    ram_cell[   46258] = 32'h705d644a;
    ram_cell[   46259] = 32'hd9b3c92e;
    ram_cell[   46260] = 32'h2ab4fe92;
    ram_cell[   46261] = 32'h8fd7c05f;
    ram_cell[   46262] = 32'h4e4701b3;
    ram_cell[   46263] = 32'h66df872a;
    ram_cell[   46264] = 32'hf870cc99;
    ram_cell[   46265] = 32'h41c17eea;
    ram_cell[   46266] = 32'hcf21760d;
    ram_cell[   46267] = 32'h5a22c960;
    ram_cell[   46268] = 32'hb919b96b;
    ram_cell[   46269] = 32'h3df95acd;
    ram_cell[   46270] = 32'heb755451;
    ram_cell[   46271] = 32'hb32bbf13;
    ram_cell[   46272] = 32'h81baa697;
    ram_cell[   46273] = 32'h5e44465d;
    ram_cell[   46274] = 32'h8813718b;
    ram_cell[   46275] = 32'h311f2d54;
    ram_cell[   46276] = 32'h56aae02b;
    ram_cell[   46277] = 32'ha7710f7c;
    ram_cell[   46278] = 32'h15b18c04;
    ram_cell[   46279] = 32'h368e6ef2;
    ram_cell[   46280] = 32'h1e617409;
    ram_cell[   46281] = 32'h3eca985a;
    ram_cell[   46282] = 32'h564c5f3f;
    ram_cell[   46283] = 32'h138c5ffb;
    ram_cell[   46284] = 32'h87877db3;
    ram_cell[   46285] = 32'h5b740bce;
    ram_cell[   46286] = 32'hc9d51bd6;
    ram_cell[   46287] = 32'h7fc0fdc7;
    ram_cell[   46288] = 32'h995aa539;
    ram_cell[   46289] = 32'h99eba867;
    ram_cell[   46290] = 32'h312da251;
    ram_cell[   46291] = 32'h88969bb2;
    ram_cell[   46292] = 32'h001a8cf9;
    ram_cell[   46293] = 32'hf37af24e;
    ram_cell[   46294] = 32'hf695cf1f;
    ram_cell[   46295] = 32'h04d2de48;
    ram_cell[   46296] = 32'h218e011c;
    ram_cell[   46297] = 32'h08bdb718;
    ram_cell[   46298] = 32'hb9332807;
    ram_cell[   46299] = 32'hc428f4e0;
    ram_cell[   46300] = 32'h859b4085;
    ram_cell[   46301] = 32'h80ac1ddc;
    ram_cell[   46302] = 32'h91a77142;
    ram_cell[   46303] = 32'h58656a0f;
    ram_cell[   46304] = 32'h7589a4dd;
    ram_cell[   46305] = 32'h3b493bf0;
    ram_cell[   46306] = 32'he875be32;
    ram_cell[   46307] = 32'h0c62e3bf;
    ram_cell[   46308] = 32'h3e265542;
    ram_cell[   46309] = 32'h2636fd01;
    ram_cell[   46310] = 32'h15ddefd6;
    ram_cell[   46311] = 32'h2e3fa291;
    ram_cell[   46312] = 32'hcdc203af;
    ram_cell[   46313] = 32'ha2211550;
    ram_cell[   46314] = 32'h0e9ab78c;
    ram_cell[   46315] = 32'h54913ae3;
    ram_cell[   46316] = 32'hc9e11c2f;
    ram_cell[   46317] = 32'h5f86314c;
    ram_cell[   46318] = 32'h8a75f8d8;
    ram_cell[   46319] = 32'h870af77b;
    ram_cell[   46320] = 32'h91614d11;
    ram_cell[   46321] = 32'he5e03dd2;
    ram_cell[   46322] = 32'hefe498ff;
    ram_cell[   46323] = 32'hceebf463;
    ram_cell[   46324] = 32'h5578d5c1;
    ram_cell[   46325] = 32'h707dde1d;
    ram_cell[   46326] = 32'h7c42f04c;
    ram_cell[   46327] = 32'h94b85480;
    ram_cell[   46328] = 32'hacb1ff32;
    ram_cell[   46329] = 32'h6b51c85a;
    ram_cell[   46330] = 32'h15c1992a;
    ram_cell[   46331] = 32'h5304f568;
    ram_cell[   46332] = 32'h8daed6ef;
    ram_cell[   46333] = 32'hdc21d2a7;
    ram_cell[   46334] = 32'h3d73a725;
    ram_cell[   46335] = 32'hf0aaa4a8;
    ram_cell[   46336] = 32'hb5fd29da;
    ram_cell[   46337] = 32'hdf073fce;
    ram_cell[   46338] = 32'h7cffe586;
    ram_cell[   46339] = 32'hec47dc66;
    ram_cell[   46340] = 32'h7294c4f0;
    ram_cell[   46341] = 32'hb7965d76;
    ram_cell[   46342] = 32'hff958b25;
    ram_cell[   46343] = 32'h52b02413;
    ram_cell[   46344] = 32'h4ca8c4d9;
    ram_cell[   46345] = 32'hae960d76;
    ram_cell[   46346] = 32'heed93eb5;
    ram_cell[   46347] = 32'hefcbb32f;
    ram_cell[   46348] = 32'h3f599c61;
    ram_cell[   46349] = 32'h63446d69;
    ram_cell[   46350] = 32'h888abad1;
    ram_cell[   46351] = 32'hcf87ecec;
    ram_cell[   46352] = 32'h198c6b9b;
    ram_cell[   46353] = 32'h1ac0bfef;
    ram_cell[   46354] = 32'h4ff0940a;
    ram_cell[   46355] = 32'h182b3e1a;
    ram_cell[   46356] = 32'h25c0da16;
    ram_cell[   46357] = 32'h56ca73d8;
    ram_cell[   46358] = 32'h72587e38;
    ram_cell[   46359] = 32'h571e4896;
    ram_cell[   46360] = 32'h68c6a63b;
    ram_cell[   46361] = 32'ha2f84284;
    ram_cell[   46362] = 32'h2ad31170;
    ram_cell[   46363] = 32'hcc46be05;
    ram_cell[   46364] = 32'hb4320c38;
    ram_cell[   46365] = 32'h566bedba;
    ram_cell[   46366] = 32'hf7ba2432;
    ram_cell[   46367] = 32'h92dbeb28;
    ram_cell[   46368] = 32'hba0cede7;
    ram_cell[   46369] = 32'h8e5c67ed;
    ram_cell[   46370] = 32'h207edc9d;
    ram_cell[   46371] = 32'hc1674e47;
    ram_cell[   46372] = 32'he01c6433;
    ram_cell[   46373] = 32'hb95e7506;
    ram_cell[   46374] = 32'h743eb4c0;
    ram_cell[   46375] = 32'h635d27f4;
    ram_cell[   46376] = 32'h4b6e7516;
    ram_cell[   46377] = 32'h4b831d3c;
    ram_cell[   46378] = 32'h4f285a9a;
    ram_cell[   46379] = 32'h2f2591bd;
    ram_cell[   46380] = 32'hf06746e3;
    ram_cell[   46381] = 32'h28c8edae;
    ram_cell[   46382] = 32'h0d93277d;
    ram_cell[   46383] = 32'h4926c7a3;
    ram_cell[   46384] = 32'h98005fda;
    ram_cell[   46385] = 32'hf1323709;
    ram_cell[   46386] = 32'h7c3bffd9;
    ram_cell[   46387] = 32'haf43fc7e;
    ram_cell[   46388] = 32'h948713f7;
    ram_cell[   46389] = 32'h8a22eebe;
    ram_cell[   46390] = 32'hf75d4888;
    ram_cell[   46391] = 32'h01825514;
    ram_cell[   46392] = 32'h31f3edd1;
    ram_cell[   46393] = 32'h2146c4ba;
    ram_cell[   46394] = 32'h2b498cdb;
    ram_cell[   46395] = 32'h52c8c623;
    ram_cell[   46396] = 32'hfe8913b9;
    ram_cell[   46397] = 32'h1fb33a40;
    ram_cell[   46398] = 32'h93900bcd;
    ram_cell[   46399] = 32'h2aed1f7f;
    ram_cell[   46400] = 32'he73bbfde;
    ram_cell[   46401] = 32'h28e77e1f;
    ram_cell[   46402] = 32'h2930a17f;
    ram_cell[   46403] = 32'h9207acdb;
    ram_cell[   46404] = 32'ha6ca8345;
    ram_cell[   46405] = 32'h4e2b8263;
    ram_cell[   46406] = 32'hb68f5c23;
    ram_cell[   46407] = 32'hee8b2e3d;
    ram_cell[   46408] = 32'hd36b10d9;
    ram_cell[   46409] = 32'hc7097d68;
    ram_cell[   46410] = 32'haaa80b54;
    ram_cell[   46411] = 32'hbef4c237;
    ram_cell[   46412] = 32'h47e0562d;
    ram_cell[   46413] = 32'hd45a80a2;
    ram_cell[   46414] = 32'h863699e5;
    ram_cell[   46415] = 32'h1dd9a684;
    ram_cell[   46416] = 32'h02a56af1;
    ram_cell[   46417] = 32'h766bb04a;
    ram_cell[   46418] = 32'hb40ddd04;
    ram_cell[   46419] = 32'he722ee45;
    ram_cell[   46420] = 32'hab450a2c;
    ram_cell[   46421] = 32'h4f762022;
    ram_cell[   46422] = 32'he7265ad2;
    ram_cell[   46423] = 32'hb35a7c35;
    ram_cell[   46424] = 32'h619c0276;
    ram_cell[   46425] = 32'h5fe63953;
    ram_cell[   46426] = 32'haa2675b0;
    ram_cell[   46427] = 32'h80f28a5a;
    ram_cell[   46428] = 32'h87f8d36d;
    ram_cell[   46429] = 32'h7e450136;
    ram_cell[   46430] = 32'h17e99d58;
    ram_cell[   46431] = 32'hc0fe3b0f;
    ram_cell[   46432] = 32'hb7840327;
    ram_cell[   46433] = 32'hb78adc6b;
    ram_cell[   46434] = 32'h0fdef21e;
    ram_cell[   46435] = 32'ha56f87f8;
    ram_cell[   46436] = 32'hed5f4fec;
    ram_cell[   46437] = 32'h6f476757;
    ram_cell[   46438] = 32'hea06cc3f;
    ram_cell[   46439] = 32'h944ec507;
    ram_cell[   46440] = 32'h74e76ff5;
    ram_cell[   46441] = 32'hb6ae4145;
    ram_cell[   46442] = 32'h306f5a23;
    ram_cell[   46443] = 32'h7c0ea6fc;
    ram_cell[   46444] = 32'ha060d869;
    ram_cell[   46445] = 32'h87ab70ac;
    ram_cell[   46446] = 32'hc92fc60d;
    ram_cell[   46447] = 32'haab4dbec;
    ram_cell[   46448] = 32'h250a19ce;
    ram_cell[   46449] = 32'h72002f0e;
    ram_cell[   46450] = 32'hc6e08f18;
    ram_cell[   46451] = 32'h87278882;
    ram_cell[   46452] = 32'h52ce4fa6;
    ram_cell[   46453] = 32'h8fd76a7d;
    ram_cell[   46454] = 32'h3750e6f8;
    ram_cell[   46455] = 32'he3bed8db;
    ram_cell[   46456] = 32'hd5fccd12;
    ram_cell[   46457] = 32'h87241b40;
    ram_cell[   46458] = 32'h71a30a97;
    ram_cell[   46459] = 32'h6e3fa765;
    ram_cell[   46460] = 32'h7dffc8aa;
    ram_cell[   46461] = 32'he113eb84;
    ram_cell[   46462] = 32'h4c9104d5;
    ram_cell[   46463] = 32'hbfd87cde;
    ram_cell[   46464] = 32'h26ad4387;
    ram_cell[   46465] = 32'hf81e2a23;
    ram_cell[   46466] = 32'h95c1a581;
    ram_cell[   46467] = 32'h3f496bf9;
    ram_cell[   46468] = 32'hf3dc113f;
    ram_cell[   46469] = 32'h8b139fc9;
    ram_cell[   46470] = 32'h75406586;
    ram_cell[   46471] = 32'hb3ef9acd;
    ram_cell[   46472] = 32'h70062274;
    ram_cell[   46473] = 32'h194d637d;
    ram_cell[   46474] = 32'hb8035e6d;
    ram_cell[   46475] = 32'h6e776aca;
    ram_cell[   46476] = 32'h6df1f8fa;
    ram_cell[   46477] = 32'h76cd7fc0;
    ram_cell[   46478] = 32'h94ed73dd;
    ram_cell[   46479] = 32'h38953a64;
    ram_cell[   46480] = 32'h7a19124f;
    ram_cell[   46481] = 32'had730876;
    ram_cell[   46482] = 32'hecf51b47;
    ram_cell[   46483] = 32'h3ee6dc17;
    ram_cell[   46484] = 32'hda3b7c3a;
    ram_cell[   46485] = 32'hfc7d11fe;
    ram_cell[   46486] = 32'h1fd94ed0;
    ram_cell[   46487] = 32'hc8172bbc;
    ram_cell[   46488] = 32'hf2946909;
    ram_cell[   46489] = 32'h13b8a702;
    ram_cell[   46490] = 32'h9c805c6b;
    ram_cell[   46491] = 32'hf226fdd6;
    ram_cell[   46492] = 32'h8c32058f;
    ram_cell[   46493] = 32'hd27fe15c;
    ram_cell[   46494] = 32'h6325c258;
    ram_cell[   46495] = 32'hf0b4240d;
    ram_cell[   46496] = 32'hb8f16b4e;
    ram_cell[   46497] = 32'h6afbd536;
    ram_cell[   46498] = 32'h8330765d;
    ram_cell[   46499] = 32'h6aa04513;
    ram_cell[   46500] = 32'hb7017653;
    ram_cell[   46501] = 32'h1115fd26;
    ram_cell[   46502] = 32'h812ba1b0;
    ram_cell[   46503] = 32'h2452a3b3;
    ram_cell[   46504] = 32'h20932923;
    ram_cell[   46505] = 32'h62b60213;
    ram_cell[   46506] = 32'h7f14162d;
    ram_cell[   46507] = 32'h2dd5acc2;
    ram_cell[   46508] = 32'h0807c222;
    ram_cell[   46509] = 32'hff9caa86;
    ram_cell[   46510] = 32'h0081d855;
    ram_cell[   46511] = 32'ha03999e3;
    ram_cell[   46512] = 32'h5680878a;
    ram_cell[   46513] = 32'h8745605f;
    ram_cell[   46514] = 32'h5eae028c;
    ram_cell[   46515] = 32'h7cd0706c;
    ram_cell[   46516] = 32'h44a7230a;
    ram_cell[   46517] = 32'h7ad81851;
    ram_cell[   46518] = 32'ha8e28aaf;
    ram_cell[   46519] = 32'ha7c0e8a1;
    ram_cell[   46520] = 32'hf02a37bb;
    ram_cell[   46521] = 32'hb413e88e;
    ram_cell[   46522] = 32'hd657457e;
    ram_cell[   46523] = 32'h59861931;
    ram_cell[   46524] = 32'hd674b1c0;
    ram_cell[   46525] = 32'h86751999;
    ram_cell[   46526] = 32'h26ff2264;
    ram_cell[   46527] = 32'h221d7756;
    ram_cell[   46528] = 32'hfb6e5f38;
    ram_cell[   46529] = 32'h1cdf323c;
    ram_cell[   46530] = 32'h8d206607;
    ram_cell[   46531] = 32'h145041c4;
    ram_cell[   46532] = 32'h1aad9f1b;
    ram_cell[   46533] = 32'h5d34033b;
    ram_cell[   46534] = 32'hd10e5960;
    ram_cell[   46535] = 32'hdf6cfb0f;
    ram_cell[   46536] = 32'h742f3d0e;
    ram_cell[   46537] = 32'h1214949b;
    ram_cell[   46538] = 32'h0941e00c;
    ram_cell[   46539] = 32'h71b49b74;
    ram_cell[   46540] = 32'h9e9185df;
    ram_cell[   46541] = 32'hb2f06227;
    ram_cell[   46542] = 32'h819e5797;
    ram_cell[   46543] = 32'h2232c263;
    ram_cell[   46544] = 32'hf0a1f264;
    ram_cell[   46545] = 32'hdf788f84;
    ram_cell[   46546] = 32'h1d9841ce;
    ram_cell[   46547] = 32'hc456f2d2;
    ram_cell[   46548] = 32'h82a26ba9;
    ram_cell[   46549] = 32'h881c8856;
    ram_cell[   46550] = 32'h89decd30;
    ram_cell[   46551] = 32'h845dc0ea;
    ram_cell[   46552] = 32'h2129ba69;
    ram_cell[   46553] = 32'h619e0a7d;
    ram_cell[   46554] = 32'h95f29bf6;
    ram_cell[   46555] = 32'h2b3460af;
    ram_cell[   46556] = 32'hd5407c7a;
    ram_cell[   46557] = 32'h2ca61423;
    ram_cell[   46558] = 32'h6c01840e;
    ram_cell[   46559] = 32'h6487de9a;
    ram_cell[   46560] = 32'hb5f45254;
    ram_cell[   46561] = 32'h55435a20;
    ram_cell[   46562] = 32'hb570dd15;
    ram_cell[   46563] = 32'h2ecac6b9;
    ram_cell[   46564] = 32'h7e3ae7d7;
    ram_cell[   46565] = 32'ha4c94467;
    ram_cell[   46566] = 32'h0d9b13c0;
    ram_cell[   46567] = 32'h5e6d7236;
    ram_cell[   46568] = 32'hd4875073;
    ram_cell[   46569] = 32'ha0e5cf89;
    ram_cell[   46570] = 32'h23555a8d;
    ram_cell[   46571] = 32'hd561608c;
    ram_cell[   46572] = 32'h1b88d2e7;
    ram_cell[   46573] = 32'h1f7586f3;
    ram_cell[   46574] = 32'hb12de59c;
    ram_cell[   46575] = 32'h1c54b845;
    ram_cell[   46576] = 32'h59867e0f;
    ram_cell[   46577] = 32'hfc8be8a8;
    ram_cell[   46578] = 32'h6d14b281;
    ram_cell[   46579] = 32'hd0ca4780;
    ram_cell[   46580] = 32'hbc64c110;
    ram_cell[   46581] = 32'hdd84cec7;
    ram_cell[   46582] = 32'he5510dae;
    ram_cell[   46583] = 32'hb09bde6b;
    ram_cell[   46584] = 32'he4a7425b;
    ram_cell[   46585] = 32'h1ce7ec10;
    ram_cell[   46586] = 32'ha0df4d20;
    ram_cell[   46587] = 32'he62ab793;
    ram_cell[   46588] = 32'h09a7d5de;
    ram_cell[   46589] = 32'he56ffd9b;
    ram_cell[   46590] = 32'h31b98b72;
    ram_cell[   46591] = 32'hf6d18f05;
    ram_cell[   46592] = 32'hcd502fbb;
    ram_cell[   46593] = 32'h7acb97e0;
    ram_cell[   46594] = 32'h97c0faab;
    ram_cell[   46595] = 32'h012e8bf1;
    ram_cell[   46596] = 32'h86a76bb6;
    ram_cell[   46597] = 32'h29523fa4;
    ram_cell[   46598] = 32'hc7bbc501;
    ram_cell[   46599] = 32'h71557b4e;
    ram_cell[   46600] = 32'h1082b662;
    ram_cell[   46601] = 32'h6d6296a9;
    ram_cell[   46602] = 32'h7771fd65;
    ram_cell[   46603] = 32'hb220243d;
    ram_cell[   46604] = 32'h616b5215;
    ram_cell[   46605] = 32'h70b017b5;
    ram_cell[   46606] = 32'h3a22331f;
    ram_cell[   46607] = 32'h761a2d03;
    ram_cell[   46608] = 32'h98a5c5c6;
    ram_cell[   46609] = 32'h6aacb37c;
    ram_cell[   46610] = 32'h60818d34;
    ram_cell[   46611] = 32'h580568e5;
    ram_cell[   46612] = 32'h9b32c7f9;
    ram_cell[   46613] = 32'hd6a199e1;
    ram_cell[   46614] = 32'hcb9f3d3e;
    ram_cell[   46615] = 32'h46f81d7d;
    ram_cell[   46616] = 32'h9f51ecf4;
    ram_cell[   46617] = 32'h1c286884;
    ram_cell[   46618] = 32'he927ac12;
    ram_cell[   46619] = 32'h66ca9dbc;
    ram_cell[   46620] = 32'h1365f2f4;
    ram_cell[   46621] = 32'h25683bf3;
    ram_cell[   46622] = 32'h91575d8b;
    ram_cell[   46623] = 32'hc3b99550;
    ram_cell[   46624] = 32'h0be8cabe;
    ram_cell[   46625] = 32'h70c1dec7;
    ram_cell[   46626] = 32'h09896a8d;
    ram_cell[   46627] = 32'ha0ab4a80;
    ram_cell[   46628] = 32'h9aaa3f98;
    ram_cell[   46629] = 32'hc01b4474;
    ram_cell[   46630] = 32'hf91a9ee3;
    ram_cell[   46631] = 32'hb2f73a71;
    ram_cell[   46632] = 32'hd967f3f1;
    ram_cell[   46633] = 32'h2f8596d6;
    ram_cell[   46634] = 32'he42cda94;
    ram_cell[   46635] = 32'hbd37fce9;
    ram_cell[   46636] = 32'h6d1c5687;
    ram_cell[   46637] = 32'h431f3af9;
    ram_cell[   46638] = 32'h99f09edb;
    ram_cell[   46639] = 32'h96e58ec8;
    ram_cell[   46640] = 32'h15bd6a4d;
    ram_cell[   46641] = 32'h51cd4def;
    ram_cell[   46642] = 32'haf8d1a5e;
    ram_cell[   46643] = 32'h8becfcc4;
    ram_cell[   46644] = 32'he067c967;
    ram_cell[   46645] = 32'hb2dfa9d4;
    ram_cell[   46646] = 32'hb72e6096;
    ram_cell[   46647] = 32'hab48e1d4;
    ram_cell[   46648] = 32'hc4e681d6;
    ram_cell[   46649] = 32'h4772703d;
    ram_cell[   46650] = 32'h3f0754fd;
    ram_cell[   46651] = 32'hd704dee1;
    ram_cell[   46652] = 32'hc5377596;
    ram_cell[   46653] = 32'hb5c55491;
    ram_cell[   46654] = 32'hfae0c960;
    ram_cell[   46655] = 32'hede39ab3;
    ram_cell[   46656] = 32'h3d998672;
    ram_cell[   46657] = 32'h13630a7a;
    ram_cell[   46658] = 32'hea3f1bfa;
    ram_cell[   46659] = 32'h5eb39734;
    ram_cell[   46660] = 32'haeacf361;
    ram_cell[   46661] = 32'h265111f2;
    ram_cell[   46662] = 32'hf9172ff8;
    ram_cell[   46663] = 32'h75c71592;
    ram_cell[   46664] = 32'hcbcb314d;
    ram_cell[   46665] = 32'hedbca561;
    ram_cell[   46666] = 32'h7c2d4aa9;
    ram_cell[   46667] = 32'h4c1be739;
    ram_cell[   46668] = 32'ha88c5e16;
    ram_cell[   46669] = 32'ha5f2b1c5;
    ram_cell[   46670] = 32'hb01c955b;
    ram_cell[   46671] = 32'hf47d3f37;
    ram_cell[   46672] = 32'h64499b0d;
    ram_cell[   46673] = 32'ha37a7048;
    ram_cell[   46674] = 32'h279477ef;
    ram_cell[   46675] = 32'h979522a8;
    ram_cell[   46676] = 32'h2350e236;
    ram_cell[   46677] = 32'h3ecc409f;
    ram_cell[   46678] = 32'he7ed578a;
    ram_cell[   46679] = 32'h72876bbb;
    ram_cell[   46680] = 32'h3b2b3677;
    ram_cell[   46681] = 32'h1698b8fa;
    ram_cell[   46682] = 32'h2b711ca8;
    ram_cell[   46683] = 32'h95dbe950;
    ram_cell[   46684] = 32'h14b1f1b3;
    ram_cell[   46685] = 32'hda9e0a6b;
    ram_cell[   46686] = 32'h6e41724c;
    ram_cell[   46687] = 32'h55e42c7f;
    ram_cell[   46688] = 32'h36a3b1c2;
    ram_cell[   46689] = 32'hc9d8655a;
    ram_cell[   46690] = 32'h958633ca;
    ram_cell[   46691] = 32'h50473a1e;
    ram_cell[   46692] = 32'hb295e2d9;
    ram_cell[   46693] = 32'ha7e6d0f7;
    ram_cell[   46694] = 32'h0a4f22a5;
    ram_cell[   46695] = 32'h30426b91;
    ram_cell[   46696] = 32'hfe7c0ed0;
    ram_cell[   46697] = 32'he1b163ff;
    ram_cell[   46698] = 32'h03449e4d;
    ram_cell[   46699] = 32'h214e6885;
    ram_cell[   46700] = 32'h8b5a89dc;
    ram_cell[   46701] = 32'h06a43b4e;
    ram_cell[   46702] = 32'h6b15daa2;
    ram_cell[   46703] = 32'h77707d68;
    ram_cell[   46704] = 32'h2dc3e261;
    ram_cell[   46705] = 32'h43ffe159;
    ram_cell[   46706] = 32'h282d79eb;
    ram_cell[   46707] = 32'hede12986;
    ram_cell[   46708] = 32'hea5175a0;
    ram_cell[   46709] = 32'h70110c27;
    ram_cell[   46710] = 32'h8e652d60;
    ram_cell[   46711] = 32'hc9d302ec;
    ram_cell[   46712] = 32'h2fced230;
    ram_cell[   46713] = 32'h88d39a61;
    ram_cell[   46714] = 32'h8253f739;
    ram_cell[   46715] = 32'h2e07dc78;
    ram_cell[   46716] = 32'h9a9b7c1f;
    ram_cell[   46717] = 32'h753a0ac9;
    ram_cell[   46718] = 32'h276d60f4;
    ram_cell[   46719] = 32'h7135c5ca;
    ram_cell[   46720] = 32'h431e793b;
    ram_cell[   46721] = 32'ha990e643;
    ram_cell[   46722] = 32'h890bce79;
    ram_cell[   46723] = 32'h0f9e6495;
    ram_cell[   46724] = 32'habf812a3;
    ram_cell[   46725] = 32'h677239b9;
    ram_cell[   46726] = 32'hdbed30f6;
    ram_cell[   46727] = 32'h2b7d83bf;
    ram_cell[   46728] = 32'hb3577b9e;
    ram_cell[   46729] = 32'h02eb7a19;
    ram_cell[   46730] = 32'hb824069c;
    ram_cell[   46731] = 32'h038fbde2;
    ram_cell[   46732] = 32'hd313a901;
    ram_cell[   46733] = 32'hdb3a2e15;
    ram_cell[   46734] = 32'h4682d940;
    ram_cell[   46735] = 32'hf6ca272c;
    ram_cell[   46736] = 32'h37672372;
    ram_cell[   46737] = 32'hb03858ed;
    ram_cell[   46738] = 32'h4c37a08b;
    ram_cell[   46739] = 32'he1faa273;
    ram_cell[   46740] = 32'h72a79e59;
    ram_cell[   46741] = 32'h0cadede0;
    ram_cell[   46742] = 32'h00883a07;
    ram_cell[   46743] = 32'h54295cce;
    ram_cell[   46744] = 32'h0edbc943;
    ram_cell[   46745] = 32'h5dcc225d;
    ram_cell[   46746] = 32'ha59e9ba5;
    ram_cell[   46747] = 32'h3f03e681;
    ram_cell[   46748] = 32'h95e3844d;
    ram_cell[   46749] = 32'h924fb1d3;
    ram_cell[   46750] = 32'ha51f4931;
    ram_cell[   46751] = 32'ha96bb6b3;
    ram_cell[   46752] = 32'hfb32376c;
    ram_cell[   46753] = 32'h3b27d3a7;
    ram_cell[   46754] = 32'h14788557;
    ram_cell[   46755] = 32'h395672e0;
    ram_cell[   46756] = 32'h274d2168;
    ram_cell[   46757] = 32'h03f91f6e;
    ram_cell[   46758] = 32'hd329f0f9;
    ram_cell[   46759] = 32'h806ea030;
    ram_cell[   46760] = 32'h7caec5a3;
    ram_cell[   46761] = 32'h9cf33974;
    ram_cell[   46762] = 32'h514b6ddb;
    ram_cell[   46763] = 32'h84f28dd5;
    ram_cell[   46764] = 32'hc33c53a4;
    ram_cell[   46765] = 32'h605e0ff3;
    ram_cell[   46766] = 32'h95939409;
    ram_cell[   46767] = 32'h157b51d2;
    ram_cell[   46768] = 32'h77fa6a94;
    ram_cell[   46769] = 32'he58f470d;
    ram_cell[   46770] = 32'hedf20ca6;
    ram_cell[   46771] = 32'h21bb8ae0;
    ram_cell[   46772] = 32'hfc90f2b6;
    ram_cell[   46773] = 32'hd3784557;
    ram_cell[   46774] = 32'hb0f414d1;
    ram_cell[   46775] = 32'hc379e3e3;
    ram_cell[   46776] = 32'hd7b58d49;
    ram_cell[   46777] = 32'he1d8a7e3;
    ram_cell[   46778] = 32'h3af007c0;
    ram_cell[   46779] = 32'h5f9d10c2;
    ram_cell[   46780] = 32'hf871de65;
    ram_cell[   46781] = 32'h6dcd7ab5;
    ram_cell[   46782] = 32'hc809bc61;
    ram_cell[   46783] = 32'h5dd27653;
    ram_cell[   46784] = 32'h34be8ae8;
    ram_cell[   46785] = 32'h12fd53cb;
    ram_cell[   46786] = 32'h4cd1f1ff;
    ram_cell[   46787] = 32'h301d93c2;
    ram_cell[   46788] = 32'h61354dd2;
    ram_cell[   46789] = 32'hb4208b77;
    ram_cell[   46790] = 32'h6f6f7d11;
    ram_cell[   46791] = 32'hf92b04c6;
    ram_cell[   46792] = 32'h4e2b73be;
    ram_cell[   46793] = 32'h4bfffa42;
    ram_cell[   46794] = 32'h2d0c7485;
    ram_cell[   46795] = 32'h2a27f13e;
    ram_cell[   46796] = 32'h261e8c50;
    ram_cell[   46797] = 32'hd28c21ff;
    ram_cell[   46798] = 32'he1de6f45;
    ram_cell[   46799] = 32'h40c0f4d8;
    ram_cell[   46800] = 32'h9a93cd1d;
    ram_cell[   46801] = 32'he2d2f0cf;
    ram_cell[   46802] = 32'h04c67b7f;
    ram_cell[   46803] = 32'h86471489;
    ram_cell[   46804] = 32'hc6d70b20;
    ram_cell[   46805] = 32'h43125089;
    ram_cell[   46806] = 32'hca63dfdd;
    ram_cell[   46807] = 32'h3597b9dc;
    ram_cell[   46808] = 32'h3221e3c7;
    ram_cell[   46809] = 32'h656053a2;
    ram_cell[   46810] = 32'h18278742;
    ram_cell[   46811] = 32'h17970c8f;
    ram_cell[   46812] = 32'hd5cff268;
    ram_cell[   46813] = 32'h09baefbc;
    ram_cell[   46814] = 32'h6ff36f19;
    ram_cell[   46815] = 32'h994296a4;
    ram_cell[   46816] = 32'h0a99bf57;
    ram_cell[   46817] = 32'h4d48c5c7;
    ram_cell[   46818] = 32'hf391a6d2;
    ram_cell[   46819] = 32'h046a4078;
    ram_cell[   46820] = 32'h23167cc6;
    ram_cell[   46821] = 32'ha16bd77b;
    ram_cell[   46822] = 32'h9bf2bec5;
    ram_cell[   46823] = 32'h330d1fef;
    ram_cell[   46824] = 32'h9e966bca;
    ram_cell[   46825] = 32'h8cccda14;
    ram_cell[   46826] = 32'hd4e62986;
    ram_cell[   46827] = 32'hf4a582df;
    ram_cell[   46828] = 32'hc7947c24;
    ram_cell[   46829] = 32'he4008e9b;
    ram_cell[   46830] = 32'h6868d910;
    ram_cell[   46831] = 32'hc8d215ac;
    ram_cell[   46832] = 32'ha84e31df;
    ram_cell[   46833] = 32'hfb8b329a;
    ram_cell[   46834] = 32'hfa0f67fb;
    ram_cell[   46835] = 32'h55d14818;
    ram_cell[   46836] = 32'hab42223a;
    ram_cell[   46837] = 32'h9d9f46ba;
    ram_cell[   46838] = 32'h91a7cd38;
    ram_cell[   46839] = 32'h4cc0bdfb;
    ram_cell[   46840] = 32'h0c177c41;
    ram_cell[   46841] = 32'h4bbd26b6;
    ram_cell[   46842] = 32'h17fd50c0;
    ram_cell[   46843] = 32'h3202d7f0;
    ram_cell[   46844] = 32'h9009acce;
    ram_cell[   46845] = 32'h7784d91e;
    ram_cell[   46846] = 32'hf2683bf3;
    ram_cell[   46847] = 32'h2022d3d1;
    ram_cell[   46848] = 32'h0ac6dfed;
    ram_cell[   46849] = 32'h1b58070d;
    ram_cell[   46850] = 32'hec251a20;
    ram_cell[   46851] = 32'hb53579d9;
    ram_cell[   46852] = 32'h8e9e2e2b;
    ram_cell[   46853] = 32'hc109f539;
    ram_cell[   46854] = 32'h538bfe0b;
    ram_cell[   46855] = 32'hb78dd1a4;
    ram_cell[   46856] = 32'h95fe243f;
    ram_cell[   46857] = 32'h760f4df3;
    ram_cell[   46858] = 32'h99c8253f;
    ram_cell[   46859] = 32'hb1b62188;
    ram_cell[   46860] = 32'h49d0eaff;
    ram_cell[   46861] = 32'h649db199;
    ram_cell[   46862] = 32'ha40df7cb;
    ram_cell[   46863] = 32'hc26efea7;
    ram_cell[   46864] = 32'h0a70db7e;
    ram_cell[   46865] = 32'h8995168a;
    ram_cell[   46866] = 32'he790273a;
    ram_cell[   46867] = 32'h1c5631cb;
    ram_cell[   46868] = 32'h1f30a0e8;
    ram_cell[   46869] = 32'hb2fb0478;
    ram_cell[   46870] = 32'h29cb073b;
    ram_cell[   46871] = 32'h85d6e7a1;
    ram_cell[   46872] = 32'h08fe6aa0;
    ram_cell[   46873] = 32'haeba3f74;
    ram_cell[   46874] = 32'h1b694870;
    ram_cell[   46875] = 32'he19fbb48;
    ram_cell[   46876] = 32'h5e2cd070;
    ram_cell[   46877] = 32'hdd9e543b;
    ram_cell[   46878] = 32'h437cc093;
    ram_cell[   46879] = 32'h1c8cc683;
    ram_cell[   46880] = 32'h30a5f51c;
    ram_cell[   46881] = 32'h214d3a39;
    ram_cell[   46882] = 32'hd0b1c08c;
    ram_cell[   46883] = 32'hf51c3684;
    ram_cell[   46884] = 32'h53cfd164;
    ram_cell[   46885] = 32'he7851b8f;
    ram_cell[   46886] = 32'hcefe2195;
    ram_cell[   46887] = 32'h6f948bd3;
    ram_cell[   46888] = 32'h8e39b027;
    ram_cell[   46889] = 32'he28ea98a;
    ram_cell[   46890] = 32'h12a7635c;
    ram_cell[   46891] = 32'hda90e2c4;
    ram_cell[   46892] = 32'ha5aff921;
    ram_cell[   46893] = 32'h663cf42a;
    ram_cell[   46894] = 32'h61d41727;
    ram_cell[   46895] = 32'hedbdc729;
    ram_cell[   46896] = 32'h6ff6347d;
    ram_cell[   46897] = 32'h17454131;
    ram_cell[   46898] = 32'h82692578;
    ram_cell[   46899] = 32'h6e548fbd;
    ram_cell[   46900] = 32'h47fec973;
    ram_cell[   46901] = 32'h581755f8;
    ram_cell[   46902] = 32'h7b50c2d0;
    ram_cell[   46903] = 32'hbbf1c2af;
    ram_cell[   46904] = 32'h593f54c2;
    ram_cell[   46905] = 32'hbf8cd2bd;
    ram_cell[   46906] = 32'h97583abf;
    ram_cell[   46907] = 32'h844ee38d;
    ram_cell[   46908] = 32'h58c180e7;
    ram_cell[   46909] = 32'h1760caf5;
    ram_cell[   46910] = 32'h399eda7d;
    ram_cell[   46911] = 32'hdb823804;
    ram_cell[   46912] = 32'h63fd3242;
    ram_cell[   46913] = 32'hc02d9291;
    ram_cell[   46914] = 32'h4edc4b8b;
    ram_cell[   46915] = 32'ha7807461;
    ram_cell[   46916] = 32'h590ef7e3;
    ram_cell[   46917] = 32'he673995a;
    ram_cell[   46918] = 32'h50abca3d;
    ram_cell[   46919] = 32'hc8281edd;
    ram_cell[   46920] = 32'h72be94c9;
    ram_cell[   46921] = 32'h9fe391e9;
    ram_cell[   46922] = 32'ha949cb26;
    ram_cell[   46923] = 32'h458b9871;
    ram_cell[   46924] = 32'h5c2abfe7;
    ram_cell[   46925] = 32'h715c7452;
    ram_cell[   46926] = 32'h4ecdbec6;
    ram_cell[   46927] = 32'h029f898d;
    ram_cell[   46928] = 32'hbe818d0e;
    ram_cell[   46929] = 32'h7a42ecca;
    ram_cell[   46930] = 32'h1733baef;
    ram_cell[   46931] = 32'hb09e2981;
    ram_cell[   46932] = 32'hb6cfedf6;
    ram_cell[   46933] = 32'ha728c6c3;
    ram_cell[   46934] = 32'h1668b0ea;
    ram_cell[   46935] = 32'he4ae6397;
    ram_cell[   46936] = 32'h55ddcd55;
    ram_cell[   46937] = 32'h14394951;
    ram_cell[   46938] = 32'he5df8a14;
    ram_cell[   46939] = 32'h5b7cb659;
    ram_cell[   46940] = 32'h028f3dbe;
    ram_cell[   46941] = 32'h18131dc1;
    ram_cell[   46942] = 32'h79a94e12;
    ram_cell[   46943] = 32'ha46065f7;
    ram_cell[   46944] = 32'hcdbcadbc;
    ram_cell[   46945] = 32'he83140e7;
    ram_cell[   46946] = 32'h8c3b28c0;
    ram_cell[   46947] = 32'h7255b09b;
    ram_cell[   46948] = 32'hfdf6b8d5;
    ram_cell[   46949] = 32'hf52afb7c;
    ram_cell[   46950] = 32'h0337cf52;
    ram_cell[   46951] = 32'h2c12e2f9;
    ram_cell[   46952] = 32'h991c4eb2;
    ram_cell[   46953] = 32'h4f11cb93;
    ram_cell[   46954] = 32'hede9c5c1;
    ram_cell[   46955] = 32'ha4a4f040;
    ram_cell[   46956] = 32'h96f15811;
    ram_cell[   46957] = 32'ha965d0cb;
    ram_cell[   46958] = 32'h85b9d119;
    ram_cell[   46959] = 32'h9c615e9b;
    ram_cell[   46960] = 32'ha21a813a;
    ram_cell[   46961] = 32'h24074dc7;
    ram_cell[   46962] = 32'h3e6ee7cc;
    ram_cell[   46963] = 32'h77e6cd85;
    ram_cell[   46964] = 32'h2f12cf68;
    ram_cell[   46965] = 32'h96026627;
    ram_cell[   46966] = 32'h4b0a2725;
    ram_cell[   46967] = 32'h64cad1c1;
    ram_cell[   46968] = 32'h72fb42c3;
    ram_cell[   46969] = 32'h1b5139f9;
    ram_cell[   46970] = 32'hc14f98d1;
    ram_cell[   46971] = 32'hcb16894a;
    ram_cell[   46972] = 32'h69ecd5d0;
    ram_cell[   46973] = 32'h6fac07d7;
    ram_cell[   46974] = 32'hd12ed328;
    ram_cell[   46975] = 32'hd265b5b8;
    ram_cell[   46976] = 32'h86842a47;
    ram_cell[   46977] = 32'hd1a8c7af;
    ram_cell[   46978] = 32'h6aa9b310;
    ram_cell[   46979] = 32'h0802fb96;
    ram_cell[   46980] = 32'h4e439359;
    ram_cell[   46981] = 32'h8c8ec1cb;
    ram_cell[   46982] = 32'h0b494f46;
    ram_cell[   46983] = 32'h66cc08f7;
    ram_cell[   46984] = 32'h262320d5;
    ram_cell[   46985] = 32'hd92f24c5;
    ram_cell[   46986] = 32'hc1a6c965;
    ram_cell[   46987] = 32'h44c4eaae;
    ram_cell[   46988] = 32'h85bec43a;
    ram_cell[   46989] = 32'hbd52bc30;
    ram_cell[   46990] = 32'h49fa73e6;
    ram_cell[   46991] = 32'h937d34d1;
    ram_cell[   46992] = 32'h21b01c8d;
    ram_cell[   46993] = 32'h2f90bae6;
    ram_cell[   46994] = 32'h9aa75346;
    ram_cell[   46995] = 32'h20689f09;
    ram_cell[   46996] = 32'h104220c2;
    ram_cell[   46997] = 32'h62ac6944;
    ram_cell[   46998] = 32'h3bf82b9d;
    ram_cell[   46999] = 32'h4e5ff497;
    ram_cell[   47000] = 32'hb2264497;
    ram_cell[   47001] = 32'he9d9cf52;
    ram_cell[   47002] = 32'h06acc991;
    ram_cell[   47003] = 32'h885223c8;
    ram_cell[   47004] = 32'h4a0c140c;
    ram_cell[   47005] = 32'h4c4ded6f;
    ram_cell[   47006] = 32'h01c5dbb2;
    ram_cell[   47007] = 32'h537b957b;
    ram_cell[   47008] = 32'h0fb4ef15;
    ram_cell[   47009] = 32'h87bf85c8;
    ram_cell[   47010] = 32'h0b3412cd;
    ram_cell[   47011] = 32'h23b8af71;
    ram_cell[   47012] = 32'h55d22afe;
    ram_cell[   47013] = 32'h6084b7be;
    ram_cell[   47014] = 32'h80aa1db7;
    ram_cell[   47015] = 32'h34e91355;
    ram_cell[   47016] = 32'hca2603bb;
    ram_cell[   47017] = 32'he5ca1e86;
    ram_cell[   47018] = 32'h97f7cd33;
    ram_cell[   47019] = 32'h05f641c6;
    ram_cell[   47020] = 32'hbd931553;
    ram_cell[   47021] = 32'h31134138;
    ram_cell[   47022] = 32'h75898ab5;
    ram_cell[   47023] = 32'h6778b794;
    ram_cell[   47024] = 32'hf1d19c0a;
    ram_cell[   47025] = 32'h753e7b37;
    ram_cell[   47026] = 32'h7400a7e0;
    ram_cell[   47027] = 32'h21b89e4c;
    ram_cell[   47028] = 32'hcf4ac681;
    ram_cell[   47029] = 32'h2f1e5847;
    ram_cell[   47030] = 32'h7afb20cd;
    ram_cell[   47031] = 32'h8d8ed0e1;
    ram_cell[   47032] = 32'h74d1bfcb;
    ram_cell[   47033] = 32'h73e2b38e;
    ram_cell[   47034] = 32'h76bcf03c;
    ram_cell[   47035] = 32'hc0c09836;
    ram_cell[   47036] = 32'h799ac9b6;
    ram_cell[   47037] = 32'h22140a48;
    ram_cell[   47038] = 32'h78fe5201;
    ram_cell[   47039] = 32'h2c7f547b;
    ram_cell[   47040] = 32'hd223c571;
    ram_cell[   47041] = 32'h683d9e52;
    ram_cell[   47042] = 32'h4e151dfc;
    ram_cell[   47043] = 32'h1d5ba973;
    ram_cell[   47044] = 32'hdb4fefd7;
    ram_cell[   47045] = 32'hb4b712f5;
    ram_cell[   47046] = 32'h9b082516;
    ram_cell[   47047] = 32'h8e8e5431;
    ram_cell[   47048] = 32'h75da9036;
    ram_cell[   47049] = 32'h557e373b;
    ram_cell[   47050] = 32'hd6418813;
    ram_cell[   47051] = 32'h5a4c4222;
    ram_cell[   47052] = 32'h7c3ec9d1;
    ram_cell[   47053] = 32'h555d53f7;
    ram_cell[   47054] = 32'h27800976;
    ram_cell[   47055] = 32'hed20e443;
    ram_cell[   47056] = 32'hfce21360;
    ram_cell[   47057] = 32'h464a05da;
    ram_cell[   47058] = 32'h5306e26b;
    ram_cell[   47059] = 32'hf83f0bfe;
    ram_cell[   47060] = 32'h5661ed46;
    ram_cell[   47061] = 32'h9a53af55;
    ram_cell[   47062] = 32'h747b67b4;
    ram_cell[   47063] = 32'h29183d8d;
    ram_cell[   47064] = 32'h130a151a;
    ram_cell[   47065] = 32'h77845555;
    ram_cell[   47066] = 32'h3b789fb8;
    ram_cell[   47067] = 32'hbbb46bf9;
    ram_cell[   47068] = 32'hf6cd652c;
    ram_cell[   47069] = 32'h34cd3ded;
    ram_cell[   47070] = 32'hc2446c6b;
    ram_cell[   47071] = 32'h98625fd5;
    ram_cell[   47072] = 32'h408c2957;
    ram_cell[   47073] = 32'hed9f5276;
    ram_cell[   47074] = 32'h88837beb;
    ram_cell[   47075] = 32'h7d52ae93;
    ram_cell[   47076] = 32'hecd344d8;
    ram_cell[   47077] = 32'ha595d326;
    ram_cell[   47078] = 32'hb52e597e;
    ram_cell[   47079] = 32'hf3f99102;
    ram_cell[   47080] = 32'h1b242fc6;
    ram_cell[   47081] = 32'h9ca9e3d7;
    ram_cell[   47082] = 32'h88748764;
    ram_cell[   47083] = 32'h16279149;
    ram_cell[   47084] = 32'h448da2c7;
    ram_cell[   47085] = 32'h44e940e2;
    ram_cell[   47086] = 32'h456ede85;
    ram_cell[   47087] = 32'h57b1be56;
    ram_cell[   47088] = 32'ha75b20c6;
    ram_cell[   47089] = 32'hacbcb681;
    ram_cell[   47090] = 32'h9fcea49a;
    ram_cell[   47091] = 32'hb3392b63;
    ram_cell[   47092] = 32'hec59bdcb;
    ram_cell[   47093] = 32'h2346195a;
    ram_cell[   47094] = 32'hff211806;
    ram_cell[   47095] = 32'hf349e938;
    ram_cell[   47096] = 32'h6bf71688;
    ram_cell[   47097] = 32'hc878ad0b;
    ram_cell[   47098] = 32'hf49efb8f;
    ram_cell[   47099] = 32'h915e725b;
    ram_cell[   47100] = 32'h2dea4824;
    ram_cell[   47101] = 32'h12850fbe;
    ram_cell[   47102] = 32'hf2cab645;
    ram_cell[   47103] = 32'h5e1428e2;
    ram_cell[   47104] = 32'hc7ac7eb0;
    ram_cell[   47105] = 32'h099476d6;
    ram_cell[   47106] = 32'h3290295c;
    ram_cell[   47107] = 32'h80d0aa40;
    ram_cell[   47108] = 32'h94742b4f;
    ram_cell[   47109] = 32'hdfaaa729;
    ram_cell[   47110] = 32'hbc1e8121;
    ram_cell[   47111] = 32'h3d17fbb3;
    ram_cell[   47112] = 32'hcf1bd539;
    ram_cell[   47113] = 32'h0bda1746;
    ram_cell[   47114] = 32'h29c9ad62;
    ram_cell[   47115] = 32'hf9416ff1;
    ram_cell[   47116] = 32'hb8dc244e;
    ram_cell[   47117] = 32'h9414d772;
    ram_cell[   47118] = 32'h9d58f472;
    ram_cell[   47119] = 32'h4fd71b56;
    ram_cell[   47120] = 32'h961f5812;
    ram_cell[   47121] = 32'h430685f4;
    ram_cell[   47122] = 32'h833a5320;
    ram_cell[   47123] = 32'h6b7fde7a;
    ram_cell[   47124] = 32'hacabe0f2;
    ram_cell[   47125] = 32'h725b54b9;
    ram_cell[   47126] = 32'h0e1693ae;
    ram_cell[   47127] = 32'h3454f7ae;
    ram_cell[   47128] = 32'h2ad88801;
    ram_cell[   47129] = 32'h83c4ee4d;
    ram_cell[   47130] = 32'h18aaa7a4;
    ram_cell[   47131] = 32'h192f5e3e;
    ram_cell[   47132] = 32'hb9c02297;
    ram_cell[   47133] = 32'h46a38285;
    ram_cell[   47134] = 32'h73d12d27;
    ram_cell[   47135] = 32'hfe090926;
    ram_cell[   47136] = 32'h22a57613;
    ram_cell[   47137] = 32'hd6c022ad;
    ram_cell[   47138] = 32'hd5ccec4f;
    ram_cell[   47139] = 32'hb6ecf7d2;
    ram_cell[   47140] = 32'hb2eb139d;
    ram_cell[   47141] = 32'hc7c9a2da;
    ram_cell[   47142] = 32'hc50bb23d;
    ram_cell[   47143] = 32'h942fd79f;
    ram_cell[   47144] = 32'ha7969d32;
    ram_cell[   47145] = 32'h1136ffe8;
    ram_cell[   47146] = 32'hb523e584;
    ram_cell[   47147] = 32'h59d71849;
    ram_cell[   47148] = 32'h5f8847ba;
    ram_cell[   47149] = 32'h1c7dab33;
    ram_cell[   47150] = 32'ha6636f49;
    ram_cell[   47151] = 32'hd05a8c03;
    ram_cell[   47152] = 32'h4103ec13;
    ram_cell[   47153] = 32'hb0a9edd4;
    ram_cell[   47154] = 32'hff20f5b8;
    ram_cell[   47155] = 32'hb5c566bd;
    ram_cell[   47156] = 32'h5c44141c;
    ram_cell[   47157] = 32'h936dcaed;
    ram_cell[   47158] = 32'h02e3e6d3;
    ram_cell[   47159] = 32'h14cde3be;
    ram_cell[   47160] = 32'h735c92c5;
    ram_cell[   47161] = 32'haf1fb5ec;
    ram_cell[   47162] = 32'he92b5e3d;
    ram_cell[   47163] = 32'h4b105757;
    ram_cell[   47164] = 32'h17878b15;
    ram_cell[   47165] = 32'h32378de9;
    ram_cell[   47166] = 32'hc84026f4;
    ram_cell[   47167] = 32'hd318937a;
    ram_cell[   47168] = 32'hf8a361ef;
    ram_cell[   47169] = 32'hf186d624;
    ram_cell[   47170] = 32'h3d26dddf;
    ram_cell[   47171] = 32'h57b2b9f3;
    ram_cell[   47172] = 32'h32de3a18;
    ram_cell[   47173] = 32'hce19b2cc;
    ram_cell[   47174] = 32'h37f371c7;
    ram_cell[   47175] = 32'h536b6a88;
    ram_cell[   47176] = 32'h470b905c;
    ram_cell[   47177] = 32'h0ea42a07;
    ram_cell[   47178] = 32'h34a9e04f;
    ram_cell[   47179] = 32'hf64877e3;
    ram_cell[   47180] = 32'h05862278;
    ram_cell[   47181] = 32'hcfd7302a;
    ram_cell[   47182] = 32'hb231488c;
    ram_cell[   47183] = 32'hacf132be;
    ram_cell[   47184] = 32'h4dc04ecb;
    ram_cell[   47185] = 32'h57f8b28d;
    ram_cell[   47186] = 32'h53be0635;
    ram_cell[   47187] = 32'hbfaf06b5;
    ram_cell[   47188] = 32'h3ca42095;
    ram_cell[   47189] = 32'h3ae9aaac;
    ram_cell[   47190] = 32'h41b61b15;
    ram_cell[   47191] = 32'h15a36e2a;
    ram_cell[   47192] = 32'h8b67e267;
    ram_cell[   47193] = 32'he61287a4;
    ram_cell[   47194] = 32'h7ab03785;
    ram_cell[   47195] = 32'hf1958891;
    ram_cell[   47196] = 32'hdb25718e;
    ram_cell[   47197] = 32'hb7fc4c46;
    ram_cell[   47198] = 32'h5b8b1f72;
    ram_cell[   47199] = 32'h6ce440d9;
    ram_cell[   47200] = 32'h3a9b6ea1;
    ram_cell[   47201] = 32'hfcd1a706;
    ram_cell[   47202] = 32'hbb7e82c8;
    ram_cell[   47203] = 32'haee1f49d;
    ram_cell[   47204] = 32'h1598a65d;
    ram_cell[   47205] = 32'h2453f317;
    ram_cell[   47206] = 32'hc7365e59;
    ram_cell[   47207] = 32'h76c39554;
    ram_cell[   47208] = 32'he41a62d3;
    ram_cell[   47209] = 32'hab188233;
    ram_cell[   47210] = 32'hea154713;
    ram_cell[   47211] = 32'h3a473104;
    ram_cell[   47212] = 32'h34b01c03;
    ram_cell[   47213] = 32'h80441950;
    ram_cell[   47214] = 32'hc2e28f8a;
    ram_cell[   47215] = 32'hbb2d75f6;
    ram_cell[   47216] = 32'h62f25c0f;
    ram_cell[   47217] = 32'h32a34c33;
    ram_cell[   47218] = 32'h6d9e770d;
    ram_cell[   47219] = 32'ha1712fec;
    ram_cell[   47220] = 32'h1d46063d;
    ram_cell[   47221] = 32'h7ffcdcc5;
    ram_cell[   47222] = 32'hccc4cac2;
    ram_cell[   47223] = 32'h13eecb21;
    ram_cell[   47224] = 32'h352c81c9;
    ram_cell[   47225] = 32'h4006b740;
    ram_cell[   47226] = 32'h7f5e134d;
    ram_cell[   47227] = 32'h89ca7e3e;
    ram_cell[   47228] = 32'he48389be;
    ram_cell[   47229] = 32'hb1ec5dcf;
    ram_cell[   47230] = 32'h57638734;
    ram_cell[   47231] = 32'h786c53c7;
    ram_cell[   47232] = 32'h41714aad;
    ram_cell[   47233] = 32'hb4b2b3f2;
    ram_cell[   47234] = 32'h7cb06af6;
    ram_cell[   47235] = 32'heacbe12c;
    ram_cell[   47236] = 32'hcbb15102;
    ram_cell[   47237] = 32'h13e2701a;
    ram_cell[   47238] = 32'h92c408d2;
    ram_cell[   47239] = 32'h43054ac4;
    ram_cell[   47240] = 32'heef7ee7a;
    ram_cell[   47241] = 32'h4972e490;
    ram_cell[   47242] = 32'hb9776dcc;
    ram_cell[   47243] = 32'h6c190ebe;
    ram_cell[   47244] = 32'hd46970b4;
    ram_cell[   47245] = 32'h36eabba7;
    ram_cell[   47246] = 32'h776504c2;
    ram_cell[   47247] = 32'he315c092;
    ram_cell[   47248] = 32'h82596b87;
    ram_cell[   47249] = 32'h8fc7c686;
    ram_cell[   47250] = 32'h7d8e2d0b;
    ram_cell[   47251] = 32'hb26f6d6b;
    ram_cell[   47252] = 32'h93186b88;
    ram_cell[   47253] = 32'h3b1213e9;
    ram_cell[   47254] = 32'h762ffe89;
    ram_cell[   47255] = 32'hbd353886;
    ram_cell[   47256] = 32'ha71cce97;
    ram_cell[   47257] = 32'hcce373cf;
    ram_cell[   47258] = 32'h820d3654;
    ram_cell[   47259] = 32'hf278cc7e;
    ram_cell[   47260] = 32'hb5ff58b1;
    ram_cell[   47261] = 32'hc97860b6;
    ram_cell[   47262] = 32'h15996d4e;
    ram_cell[   47263] = 32'h3d06ec2e;
    ram_cell[   47264] = 32'h23663087;
    ram_cell[   47265] = 32'h4c6f6f13;
    ram_cell[   47266] = 32'h17b61feb;
    ram_cell[   47267] = 32'h70bfd580;
    ram_cell[   47268] = 32'hc5243430;
    ram_cell[   47269] = 32'h728f6788;
    ram_cell[   47270] = 32'h2ddd6d3d;
    ram_cell[   47271] = 32'hdb23e156;
    ram_cell[   47272] = 32'h7ef78ed1;
    ram_cell[   47273] = 32'h4bcb3dd8;
    ram_cell[   47274] = 32'h7dde129e;
    ram_cell[   47275] = 32'h9e68ae8c;
    ram_cell[   47276] = 32'h3cb76446;
    ram_cell[   47277] = 32'h6e47d1a9;
    ram_cell[   47278] = 32'hbd316ac0;
    ram_cell[   47279] = 32'h3f2df89c;
    ram_cell[   47280] = 32'hd7de61cf;
    ram_cell[   47281] = 32'h2eeb743f;
    ram_cell[   47282] = 32'ha88c1d8b;
    ram_cell[   47283] = 32'h20776680;
    ram_cell[   47284] = 32'h1b1ab9ff;
    ram_cell[   47285] = 32'h332ef9c6;
    ram_cell[   47286] = 32'ha2d0ad91;
    ram_cell[   47287] = 32'h875e5e83;
    ram_cell[   47288] = 32'h9868ffd6;
    ram_cell[   47289] = 32'hcb007c45;
    ram_cell[   47290] = 32'h1694e9a4;
    ram_cell[   47291] = 32'hd7164a46;
    ram_cell[   47292] = 32'hf2c6d3bc;
    ram_cell[   47293] = 32'h733be0ac;
    ram_cell[   47294] = 32'h781f28e8;
    ram_cell[   47295] = 32'hb6aac007;
    ram_cell[   47296] = 32'hb40b3efa;
    ram_cell[   47297] = 32'h4bc2ad7f;
    ram_cell[   47298] = 32'h46a59672;
    ram_cell[   47299] = 32'hbb0af618;
    ram_cell[   47300] = 32'h436d3da2;
    ram_cell[   47301] = 32'h6d64e0b2;
    ram_cell[   47302] = 32'h7a6671a4;
    ram_cell[   47303] = 32'hd0165cb3;
    ram_cell[   47304] = 32'hc13f041c;
    ram_cell[   47305] = 32'h89f2e067;
    ram_cell[   47306] = 32'he0eed64a;
    ram_cell[   47307] = 32'hbebc45e5;
    ram_cell[   47308] = 32'h6e5baccf;
    ram_cell[   47309] = 32'h888acc35;
    ram_cell[   47310] = 32'h904194bc;
    ram_cell[   47311] = 32'hd7034575;
    ram_cell[   47312] = 32'h9f00b4a2;
    ram_cell[   47313] = 32'h433595fa;
    ram_cell[   47314] = 32'hf42ae0b8;
    ram_cell[   47315] = 32'ha01bdf8e;
    ram_cell[   47316] = 32'hdd2a1ae0;
    ram_cell[   47317] = 32'h593c3b46;
    ram_cell[   47318] = 32'h83b3901b;
    ram_cell[   47319] = 32'h70b01776;
    ram_cell[   47320] = 32'h097338fc;
    ram_cell[   47321] = 32'h891815f6;
    ram_cell[   47322] = 32'h7f82db65;
    ram_cell[   47323] = 32'h052ea266;
    ram_cell[   47324] = 32'h8b7c659f;
    ram_cell[   47325] = 32'hb339c19f;
    ram_cell[   47326] = 32'hc8f5d176;
    ram_cell[   47327] = 32'h0738d401;
    ram_cell[   47328] = 32'h839b2bf7;
    ram_cell[   47329] = 32'h582e1c24;
    ram_cell[   47330] = 32'hbccb5b50;
    ram_cell[   47331] = 32'h74512283;
    ram_cell[   47332] = 32'haddd6f63;
    ram_cell[   47333] = 32'h98305b09;
    ram_cell[   47334] = 32'hab20cb32;
    ram_cell[   47335] = 32'he49d98e3;
    ram_cell[   47336] = 32'h77e40527;
    ram_cell[   47337] = 32'h426d2a67;
    ram_cell[   47338] = 32'h442cd170;
    ram_cell[   47339] = 32'h5cc55455;
    ram_cell[   47340] = 32'h66ae0456;
    ram_cell[   47341] = 32'h574bc98f;
    ram_cell[   47342] = 32'h0d23e4a9;
    ram_cell[   47343] = 32'h24f5248b;
    ram_cell[   47344] = 32'ha7937ccc;
    ram_cell[   47345] = 32'hd6063bf8;
    ram_cell[   47346] = 32'h58350bd6;
    ram_cell[   47347] = 32'h9745a57d;
    ram_cell[   47348] = 32'h7b9d87a7;
    ram_cell[   47349] = 32'h996f48fc;
    ram_cell[   47350] = 32'hd1605d3f;
    ram_cell[   47351] = 32'hda4fdb03;
    ram_cell[   47352] = 32'h33fd488b;
    ram_cell[   47353] = 32'h94d7d0f8;
    ram_cell[   47354] = 32'hfb1bc056;
    ram_cell[   47355] = 32'h8bcbc1ec;
    ram_cell[   47356] = 32'hc46d84da;
    ram_cell[   47357] = 32'h65a49b9e;
    ram_cell[   47358] = 32'haf5a057f;
    ram_cell[   47359] = 32'h5a4157f0;
    ram_cell[   47360] = 32'h06b80916;
    ram_cell[   47361] = 32'hbf1aa562;
    ram_cell[   47362] = 32'hb1ac913b;
    ram_cell[   47363] = 32'hd5af27ef;
    ram_cell[   47364] = 32'h87d378ac;
    ram_cell[   47365] = 32'hbd65c217;
    ram_cell[   47366] = 32'h4823c958;
    ram_cell[   47367] = 32'hb85aaa21;
    ram_cell[   47368] = 32'h2ee8e85b;
    ram_cell[   47369] = 32'h17ee5dd5;
    ram_cell[   47370] = 32'hb912d5c8;
    ram_cell[   47371] = 32'h14885b66;
    ram_cell[   47372] = 32'he657218d;
    ram_cell[   47373] = 32'h42296066;
    ram_cell[   47374] = 32'hde4a95cd;
    ram_cell[   47375] = 32'hbdcc2695;
    ram_cell[   47376] = 32'h9da705a3;
    ram_cell[   47377] = 32'h7b6f3891;
    ram_cell[   47378] = 32'hfd88117c;
    ram_cell[   47379] = 32'h31109198;
    ram_cell[   47380] = 32'hd321796e;
    ram_cell[   47381] = 32'hca890a2a;
    ram_cell[   47382] = 32'h1d849864;
    ram_cell[   47383] = 32'h6998497f;
    ram_cell[   47384] = 32'h7074535f;
    ram_cell[   47385] = 32'h9ac95622;
    ram_cell[   47386] = 32'hd5c6a452;
    ram_cell[   47387] = 32'hf7befdda;
    ram_cell[   47388] = 32'h85c67103;
    ram_cell[   47389] = 32'h5e22b746;
    ram_cell[   47390] = 32'ha0419af3;
    ram_cell[   47391] = 32'hfec65a1e;
    ram_cell[   47392] = 32'hd8076413;
    ram_cell[   47393] = 32'hdb7fa8f2;
    ram_cell[   47394] = 32'hce9632cb;
    ram_cell[   47395] = 32'ha2464193;
    ram_cell[   47396] = 32'h1fafd31c;
    ram_cell[   47397] = 32'he52ce1de;
    ram_cell[   47398] = 32'h89b24ccf;
    ram_cell[   47399] = 32'h9250adba;
    ram_cell[   47400] = 32'h8ebdae16;
    ram_cell[   47401] = 32'hc9b9ca15;
    ram_cell[   47402] = 32'h8e051d56;
    ram_cell[   47403] = 32'hf58d8050;
    ram_cell[   47404] = 32'h2c4614b9;
    ram_cell[   47405] = 32'h9e4c4d18;
    ram_cell[   47406] = 32'hcf3d2abd;
    ram_cell[   47407] = 32'h0a07f711;
    ram_cell[   47408] = 32'h17992280;
    ram_cell[   47409] = 32'ha334dd7d;
    ram_cell[   47410] = 32'hc2aa1318;
    ram_cell[   47411] = 32'h3252a06b;
    ram_cell[   47412] = 32'hfc6ec97d;
    ram_cell[   47413] = 32'h9dd2d5a2;
    ram_cell[   47414] = 32'h60f4a0c4;
    ram_cell[   47415] = 32'h9ec4f389;
    ram_cell[   47416] = 32'h2f5d6d1e;
    ram_cell[   47417] = 32'h25783699;
    ram_cell[   47418] = 32'h379c5aac;
    ram_cell[   47419] = 32'hce2f52bc;
    ram_cell[   47420] = 32'h2c4a18e2;
    ram_cell[   47421] = 32'hf88255c3;
    ram_cell[   47422] = 32'h4d6f1388;
    ram_cell[   47423] = 32'h1b166d17;
    ram_cell[   47424] = 32'ha9109622;
    ram_cell[   47425] = 32'h7775d39c;
    ram_cell[   47426] = 32'h8961b2e4;
    ram_cell[   47427] = 32'h90b59f6c;
    ram_cell[   47428] = 32'h3e2a48bf;
    ram_cell[   47429] = 32'h6c034f40;
    ram_cell[   47430] = 32'haa2880a8;
    ram_cell[   47431] = 32'h454d9ebc;
    ram_cell[   47432] = 32'hec1f7583;
    ram_cell[   47433] = 32'h58e750c4;
    ram_cell[   47434] = 32'heedb4327;
    ram_cell[   47435] = 32'h4e9de0f5;
    ram_cell[   47436] = 32'h8538d41a;
    ram_cell[   47437] = 32'h0492bac3;
    ram_cell[   47438] = 32'h1ca1aa30;
    ram_cell[   47439] = 32'h3b04b6d0;
    ram_cell[   47440] = 32'h02f45cb4;
    ram_cell[   47441] = 32'hb8a95538;
    ram_cell[   47442] = 32'haa573263;
    ram_cell[   47443] = 32'hef7c1827;
    ram_cell[   47444] = 32'hb8cdbbc6;
    ram_cell[   47445] = 32'ha7ff848d;
    ram_cell[   47446] = 32'h65a6b85e;
    ram_cell[   47447] = 32'h4fd29887;
    ram_cell[   47448] = 32'hf1a17463;
    ram_cell[   47449] = 32'h35758cf7;
    ram_cell[   47450] = 32'h0b4d9bd7;
    ram_cell[   47451] = 32'h8bb3e22e;
    ram_cell[   47452] = 32'h8c9c4a2d;
    ram_cell[   47453] = 32'h3119b340;
    ram_cell[   47454] = 32'hdafe12cc;
    ram_cell[   47455] = 32'h06b9ae01;
    ram_cell[   47456] = 32'he947c94c;
    ram_cell[   47457] = 32'hccb516e3;
    ram_cell[   47458] = 32'hcf1793b3;
    ram_cell[   47459] = 32'h8f461b6a;
    ram_cell[   47460] = 32'hb74db346;
    ram_cell[   47461] = 32'he1364c81;
    ram_cell[   47462] = 32'h9eaacb72;
    ram_cell[   47463] = 32'ha2551026;
    ram_cell[   47464] = 32'h964af696;
    ram_cell[   47465] = 32'h52e7964f;
    ram_cell[   47466] = 32'h6854fbba;
    ram_cell[   47467] = 32'h6f6ef3b3;
    ram_cell[   47468] = 32'h143fde62;
    ram_cell[   47469] = 32'hb6cb8c61;
    ram_cell[   47470] = 32'h7040ac15;
    ram_cell[   47471] = 32'h4b3b23a4;
    ram_cell[   47472] = 32'h814c8d2d;
    ram_cell[   47473] = 32'hbea5cb1a;
    ram_cell[   47474] = 32'h8dd5ae3f;
    ram_cell[   47475] = 32'haeef4891;
    ram_cell[   47476] = 32'h0a6d3a0c;
    ram_cell[   47477] = 32'h387b7b7d;
    ram_cell[   47478] = 32'h1871b575;
    ram_cell[   47479] = 32'hb789af3e;
    ram_cell[   47480] = 32'hfbe20dc9;
    ram_cell[   47481] = 32'h49697b6b;
    ram_cell[   47482] = 32'h1ca1b6f5;
    ram_cell[   47483] = 32'hafd34b0d;
    ram_cell[   47484] = 32'h5a6289ff;
    ram_cell[   47485] = 32'h08f9301c;
    ram_cell[   47486] = 32'hb6ba8c51;
    ram_cell[   47487] = 32'h93a5d16a;
    ram_cell[   47488] = 32'hd1101809;
    ram_cell[   47489] = 32'hbe55b500;
    ram_cell[   47490] = 32'hfa96738a;
    ram_cell[   47491] = 32'h9e34117b;
    ram_cell[   47492] = 32'h5598af63;
    ram_cell[   47493] = 32'ha138dc9e;
    ram_cell[   47494] = 32'h433b29a4;
    ram_cell[   47495] = 32'h80202388;
    ram_cell[   47496] = 32'hba49a432;
    ram_cell[   47497] = 32'h7c9b7fba;
    ram_cell[   47498] = 32'h3b84b944;
    ram_cell[   47499] = 32'hea7b045e;
    ram_cell[   47500] = 32'hfa4bd06f;
    ram_cell[   47501] = 32'hacf6e6a8;
    ram_cell[   47502] = 32'h4486eaf3;
    ram_cell[   47503] = 32'hde88abe3;
    ram_cell[   47504] = 32'h8aba9b93;
    ram_cell[   47505] = 32'hcf419cc4;
    ram_cell[   47506] = 32'h80f8cd58;
    ram_cell[   47507] = 32'hca01f823;
    ram_cell[   47508] = 32'h2fa4257a;
    ram_cell[   47509] = 32'h003b713b;
    ram_cell[   47510] = 32'h809fb97d;
    ram_cell[   47511] = 32'hb0f1baa6;
    ram_cell[   47512] = 32'h8eaf4422;
    ram_cell[   47513] = 32'h8a5e5188;
    ram_cell[   47514] = 32'hb3155a65;
    ram_cell[   47515] = 32'h52960a0f;
    ram_cell[   47516] = 32'hdd416613;
    ram_cell[   47517] = 32'h0779fb54;
    ram_cell[   47518] = 32'he3a13ed3;
    ram_cell[   47519] = 32'h3939569e;
    ram_cell[   47520] = 32'h1897ca3e;
    ram_cell[   47521] = 32'hde005526;
    ram_cell[   47522] = 32'h8b9e826b;
    ram_cell[   47523] = 32'h38cdfd91;
    ram_cell[   47524] = 32'hee71cdf8;
    ram_cell[   47525] = 32'h06c2c75a;
    ram_cell[   47526] = 32'hf6571431;
    ram_cell[   47527] = 32'hdc127109;
    ram_cell[   47528] = 32'h60d3aa17;
    ram_cell[   47529] = 32'h583a95b1;
    ram_cell[   47530] = 32'hf646bb71;
    ram_cell[   47531] = 32'h69cff25c;
    ram_cell[   47532] = 32'h7c5e5696;
    ram_cell[   47533] = 32'h7b9c4aa7;
    ram_cell[   47534] = 32'h3e3a2946;
    ram_cell[   47535] = 32'h539789b0;
    ram_cell[   47536] = 32'h2cc59526;
    ram_cell[   47537] = 32'h55e5d7f3;
    ram_cell[   47538] = 32'ha50d76cf;
    ram_cell[   47539] = 32'h84a265c0;
    ram_cell[   47540] = 32'he1142a44;
    ram_cell[   47541] = 32'heb8a910a;
    ram_cell[   47542] = 32'hfc88493f;
    ram_cell[   47543] = 32'h4a2d5b76;
    ram_cell[   47544] = 32'h49c95f29;
    ram_cell[   47545] = 32'h62afd22d;
    ram_cell[   47546] = 32'h51d1412a;
    ram_cell[   47547] = 32'hefef4b30;
    ram_cell[   47548] = 32'h913579ac;
    ram_cell[   47549] = 32'h5814873c;
    ram_cell[   47550] = 32'h6f22591b;
    ram_cell[   47551] = 32'h901a752d;
    ram_cell[   47552] = 32'h5a9aff88;
    ram_cell[   47553] = 32'hf424ef59;
    ram_cell[   47554] = 32'h414731a1;
    ram_cell[   47555] = 32'h800a4dd2;
    ram_cell[   47556] = 32'hea8bea51;
    ram_cell[   47557] = 32'hcb6be107;
    ram_cell[   47558] = 32'h3f9a86cc;
    ram_cell[   47559] = 32'h2f0c15ba;
    ram_cell[   47560] = 32'h71e28682;
    ram_cell[   47561] = 32'ha39e9acd;
    ram_cell[   47562] = 32'hdf02a034;
    ram_cell[   47563] = 32'hc46b77c1;
    ram_cell[   47564] = 32'h3b0d9099;
    ram_cell[   47565] = 32'h7edea3d0;
    ram_cell[   47566] = 32'h828b1c70;
    ram_cell[   47567] = 32'h17eedc2a;
    ram_cell[   47568] = 32'hdcfe0caa;
    ram_cell[   47569] = 32'hafc6108f;
    ram_cell[   47570] = 32'h8883102e;
    ram_cell[   47571] = 32'h5c58b5eb;
    ram_cell[   47572] = 32'hb7084bb9;
    ram_cell[   47573] = 32'h1851932e;
    ram_cell[   47574] = 32'h83c2b809;
    ram_cell[   47575] = 32'h5c64051c;
    ram_cell[   47576] = 32'h7b35bd25;
    ram_cell[   47577] = 32'h1d6de82b;
    ram_cell[   47578] = 32'hcd1deeb8;
    ram_cell[   47579] = 32'he7b92635;
    ram_cell[   47580] = 32'hf43862eb;
    ram_cell[   47581] = 32'hbe1570d4;
    ram_cell[   47582] = 32'h6024785e;
    ram_cell[   47583] = 32'hbf4ace2c;
    ram_cell[   47584] = 32'h6badf30d;
    ram_cell[   47585] = 32'h4fc59640;
    ram_cell[   47586] = 32'h01eb7170;
    ram_cell[   47587] = 32'h99eca5ee;
    ram_cell[   47588] = 32'h7092d267;
    ram_cell[   47589] = 32'hce7a7f32;
    ram_cell[   47590] = 32'h7d57b509;
    ram_cell[   47591] = 32'h01899666;
    ram_cell[   47592] = 32'hf8a74018;
    ram_cell[   47593] = 32'h24c09bc5;
    ram_cell[   47594] = 32'hacdd7875;
    ram_cell[   47595] = 32'h173e0747;
    ram_cell[   47596] = 32'hb1b76982;
    ram_cell[   47597] = 32'hf83abd63;
    ram_cell[   47598] = 32'hc91e0a50;
    ram_cell[   47599] = 32'h94a73451;
    ram_cell[   47600] = 32'ha80ceb1e;
    ram_cell[   47601] = 32'ha0e302d7;
    ram_cell[   47602] = 32'he8f40b59;
    ram_cell[   47603] = 32'h9d7e9ac9;
    ram_cell[   47604] = 32'h60183c98;
    ram_cell[   47605] = 32'he7a60762;
    ram_cell[   47606] = 32'h9aa94af0;
    ram_cell[   47607] = 32'hb4fd0ea5;
    ram_cell[   47608] = 32'h7c485a5e;
    ram_cell[   47609] = 32'h2afd8a1b;
    ram_cell[   47610] = 32'h4c666b78;
    ram_cell[   47611] = 32'h9fbcfc53;
    ram_cell[   47612] = 32'h05e1cb1f;
    ram_cell[   47613] = 32'h4c8a54f8;
    ram_cell[   47614] = 32'hf69363b3;
    ram_cell[   47615] = 32'h6f42c044;
    ram_cell[   47616] = 32'hd71f27af;
    ram_cell[   47617] = 32'hfe9322c4;
    ram_cell[   47618] = 32'h870fd97f;
    ram_cell[   47619] = 32'h8c2b5850;
    ram_cell[   47620] = 32'h9fc3c257;
    ram_cell[   47621] = 32'h7c445908;
    ram_cell[   47622] = 32'hacaa474d;
    ram_cell[   47623] = 32'h4b643b98;
    ram_cell[   47624] = 32'h81abb0a4;
    ram_cell[   47625] = 32'haf8816f7;
    ram_cell[   47626] = 32'h7d2c8775;
    ram_cell[   47627] = 32'h0e85a824;
    ram_cell[   47628] = 32'h58d124e3;
    ram_cell[   47629] = 32'h24d5765d;
    ram_cell[   47630] = 32'hb9cfaf7f;
    ram_cell[   47631] = 32'h4d23f3f1;
    ram_cell[   47632] = 32'h24443d86;
    ram_cell[   47633] = 32'h9bf8b716;
    ram_cell[   47634] = 32'h70f24d02;
    ram_cell[   47635] = 32'hc2d972e5;
    ram_cell[   47636] = 32'hbce7dc83;
    ram_cell[   47637] = 32'h3e9ec28a;
    ram_cell[   47638] = 32'h4ca77e2d;
    ram_cell[   47639] = 32'hda3b394c;
    ram_cell[   47640] = 32'hf06fa178;
    ram_cell[   47641] = 32'he92dbf02;
    ram_cell[   47642] = 32'h0b60053d;
    ram_cell[   47643] = 32'hc3b9ac50;
    ram_cell[   47644] = 32'he5e30a4c;
    ram_cell[   47645] = 32'h2de24921;
    ram_cell[   47646] = 32'hc2d1a2e1;
    ram_cell[   47647] = 32'hab3693e7;
    ram_cell[   47648] = 32'h62313e1f;
    ram_cell[   47649] = 32'hae722f61;
    ram_cell[   47650] = 32'h136a3f25;
    ram_cell[   47651] = 32'h310a8504;
    ram_cell[   47652] = 32'h743b2b9b;
    ram_cell[   47653] = 32'ha292de31;
    ram_cell[   47654] = 32'h88689bce;
    ram_cell[   47655] = 32'h4193a23d;
    ram_cell[   47656] = 32'h282a0429;
    ram_cell[   47657] = 32'h4b82b1df;
    ram_cell[   47658] = 32'h9cf90eaa;
    ram_cell[   47659] = 32'h760416c5;
    ram_cell[   47660] = 32'hbbed53f3;
    ram_cell[   47661] = 32'he7a23bef;
    ram_cell[   47662] = 32'h954318c2;
    ram_cell[   47663] = 32'he9c39911;
    ram_cell[   47664] = 32'h31ca4f17;
    ram_cell[   47665] = 32'h0184266f;
    ram_cell[   47666] = 32'h2c927183;
    ram_cell[   47667] = 32'h76c0f167;
    ram_cell[   47668] = 32'hfb53ba3f;
    ram_cell[   47669] = 32'h0542e1a2;
    ram_cell[   47670] = 32'h21371573;
    ram_cell[   47671] = 32'h3262bb3e;
    ram_cell[   47672] = 32'hb4237a36;
    ram_cell[   47673] = 32'h9e79389a;
    ram_cell[   47674] = 32'hfdfa49a4;
    ram_cell[   47675] = 32'hbed7a71d;
    ram_cell[   47676] = 32'h53daa301;
    ram_cell[   47677] = 32'h892672ee;
    ram_cell[   47678] = 32'h3e46f18a;
    ram_cell[   47679] = 32'h677c8d4b;
    ram_cell[   47680] = 32'hc8724c2c;
    ram_cell[   47681] = 32'h5d7b7ff3;
    ram_cell[   47682] = 32'hd78cca84;
    ram_cell[   47683] = 32'he7270215;
    ram_cell[   47684] = 32'h1a43267a;
    ram_cell[   47685] = 32'h6b24f05d;
    ram_cell[   47686] = 32'h253d3a62;
    ram_cell[   47687] = 32'haa48da05;
    ram_cell[   47688] = 32'hf47ae197;
    ram_cell[   47689] = 32'haf169f76;
    ram_cell[   47690] = 32'hd8362ff5;
    ram_cell[   47691] = 32'h25184813;
    ram_cell[   47692] = 32'h3f33cf47;
    ram_cell[   47693] = 32'hc21052ff;
    ram_cell[   47694] = 32'h8c823321;
    ram_cell[   47695] = 32'h3a310715;
    ram_cell[   47696] = 32'h3d5be7c4;
    ram_cell[   47697] = 32'h8226fa48;
    ram_cell[   47698] = 32'h2830ded3;
    ram_cell[   47699] = 32'h4bf2d9b7;
    ram_cell[   47700] = 32'h936fbb43;
    ram_cell[   47701] = 32'hba4876db;
    ram_cell[   47702] = 32'hf2b34d67;
    ram_cell[   47703] = 32'h38b10f16;
    ram_cell[   47704] = 32'he05ff7ba;
    ram_cell[   47705] = 32'h0a83204d;
    ram_cell[   47706] = 32'h1d0789da;
    ram_cell[   47707] = 32'h276acca2;
    ram_cell[   47708] = 32'h8f1ed69a;
    ram_cell[   47709] = 32'h09387566;
    ram_cell[   47710] = 32'h7050a5f2;
    ram_cell[   47711] = 32'hda5a045a;
    ram_cell[   47712] = 32'hbd7b9be5;
    ram_cell[   47713] = 32'hd7beea7b;
    ram_cell[   47714] = 32'h4c2ee27d;
    ram_cell[   47715] = 32'h1a5f9ba2;
    ram_cell[   47716] = 32'hcb4e3449;
    ram_cell[   47717] = 32'h8c0b1663;
    ram_cell[   47718] = 32'hd6f0c677;
    ram_cell[   47719] = 32'h7c3229b0;
    ram_cell[   47720] = 32'hc385ab4a;
    ram_cell[   47721] = 32'h18216647;
    ram_cell[   47722] = 32'hc441cc23;
    ram_cell[   47723] = 32'h5a279816;
    ram_cell[   47724] = 32'h91fd152e;
    ram_cell[   47725] = 32'he0e3a62e;
    ram_cell[   47726] = 32'h6a58bc52;
    ram_cell[   47727] = 32'hb8077b12;
    ram_cell[   47728] = 32'h05fd6ac5;
    ram_cell[   47729] = 32'h7a43e9ce;
    ram_cell[   47730] = 32'hbba1cb1a;
    ram_cell[   47731] = 32'h67be55a5;
    ram_cell[   47732] = 32'h47974d8c;
    ram_cell[   47733] = 32'h591ba9d9;
    ram_cell[   47734] = 32'h0299b93e;
    ram_cell[   47735] = 32'hec7fef03;
    ram_cell[   47736] = 32'hed93844c;
    ram_cell[   47737] = 32'hfe570dfe;
    ram_cell[   47738] = 32'h3b8904e0;
    ram_cell[   47739] = 32'hb5bf08ee;
    ram_cell[   47740] = 32'h7ed8e40b;
    ram_cell[   47741] = 32'h4d55248d;
    ram_cell[   47742] = 32'h69ce5eb9;
    ram_cell[   47743] = 32'h33e90566;
    ram_cell[   47744] = 32'h93ac8c62;
    ram_cell[   47745] = 32'h4121ba88;
    ram_cell[   47746] = 32'h892f96fb;
    ram_cell[   47747] = 32'h3c970aeb;
    ram_cell[   47748] = 32'h9d09097d;
    ram_cell[   47749] = 32'hcdceae01;
    ram_cell[   47750] = 32'hafb2a089;
    ram_cell[   47751] = 32'h13517075;
    ram_cell[   47752] = 32'h332d015f;
    ram_cell[   47753] = 32'hafc07fa9;
    ram_cell[   47754] = 32'hb2a1b1b0;
    ram_cell[   47755] = 32'h446be6fa;
    ram_cell[   47756] = 32'hf2b3565f;
    ram_cell[   47757] = 32'he194237e;
    ram_cell[   47758] = 32'h3a23c39b;
    ram_cell[   47759] = 32'hcad49b30;
    ram_cell[   47760] = 32'hda1d2a4e;
    ram_cell[   47761] = 32'h5c84c7ba;
    ram_cell[   47762] = 32'h963e249c;
    ram_cell[   47763] = 32'hc6304b2a;
    ram_cell[   47764] = 32'hb11098ac;
    ram_cell[   47765] = 32'h4f7755f6;
    ram_cell[   47766] = 32'hb250adf3;
    ram_cell[   47767] = 32'h98a56929;
    ram_cell[   47768] = 32'h8ebaff71;
    ram_cell[   47769] = 32'h4e79a196;
    ram_cell[   47770] = 32'h8efa796b;
    ram_cell[   47771] = 32'h65e960d8;
    ram_cell[   47772] = 32'hc62c73bf;
    ram_cell[   47773] = 32'hbb22c50c;
    ram_cell[   47774] = 32'h98b05188;
    ram_cell[   47775] = 32'hfc92ce5a;
    ram_cell[   47776] = 32'h9e7907ba;
    ram_cell[   47777] = 32'hcdac94da;
    ram_cell[   47778] = 32'hcaadb7ab;
    ram_cell[   47779] = 32'h0e211a47;
    ram_cell[   47780] = 32'he3599673;
    ram_cell[   47781] = 32'hc8d66320;
    ram_cell[   47782] = 32'h58f097a8;
    ram_cell[   47783] = 32'hce9c3249;
    ram_cell[   47784] = 32'hf8dbcf62;
    ram_cell[   47785] = 32'h4e0c1c88;
    ram_cell[   47786] = 32'h08b63d10;
    ram_cell[   47787] = 32'hbbc0af7a;
    ram_cell[   47788] = 32'h0fd31525;
    ram_cell[   47789] = 32'hcb82028d;
    ram_cell[   47790] = 32'haacc68b4;
    ram_cell[   47791] = 32'hc16a7d7d;
    ram_cell[   47792] = 32'h6fa891e2;
    ram_cell[   47793] = 32'hb5524751;
    ram_cell[   47794] = 32'hcdcf777c;
    ram_cell[   47795] = 32'h0aa4b2bc;
    ram_cell[   47796] = 32'h1b20cf3a;
    ram_cell[   47797] = 32'hee554267;
    ram_cell[   47798] = 32'h2c852b33;
    ram_cell[   47799] = 32'h48f93433;
    ram_cell[   47800] = 32'h416fce5d;
    ram_cell[   47801] = 32'h945d130e;
    ram_cell[   47802] = 32'h8afbefd2;
    ram_cell[   47803] = 32'h9dd1700f;
    ram_cell[   47804] = 32'hade42289;
    ram_cell[   47805] = 32'hed844e47;
    ram_cell[   47806] = 32'h7cf314aa;
    ram_cell[   47807] = 32'ha783773a;
    ram_cell[   47808] = 32'h89a27b04;
    ram_cell[   47809] = 32'ha6933bdd;
    ram_cell[   47810] = 32'h1297084e;
    ram_cell[   47811] = 32'h571faef3;
    ram_cell[   47812] = 32'h78805e8a;
    ram_cell[   47813] = 32'h6a67a79f;
    ram_cell[   47814] = 32'h04f9b74e;
    ram_cell[   47815] = 32'h115725d7;
    ram_cell[   47816] = 32'hc844264c;
    ram_cell[   47817] = 32'h7674db76;
    ram_cell[   47818] = 32'h1250212e;
    ram_cell[   47819] = 32'h9778e3ec;
    ram_cell[   47820] = 32'h08e2d993;
    ram_cell[   47821] = 32'hde8e07bf;
    ram_cell[   47822] = 32'hfaae3a95;
    ram_cell[   47823] = 32'h7e16c81a;
    ram_cell[   47824] = 32'h3e7beb94;
    ram_cell[   47825] = 32'h02250462;
    ram_cell[   47826] = 32'h474765d9;
    ram_cell[   47827] = 32'hba6937c4;
    ram_cell[   47828] = 32'hb2c2c74e;
    ram_cell[   47829] = 32'h3a7cc4ac;
    ram_cell[   47830] = 32'h1dcd25b8;
    ram_cell[   47831] = 32'he6b0a16c;
    ram_cell[   47832] = 32'haf3147ed;
    ram_cell[   47833] = 32'h89009cbc;
    ram_cell[   47834] = 32'he9f1d03a;
    ram_cell[   47835] = 32'h0b337d5e;
    ram_cell[   47836] = 32'hf2271383;
    ram_cell[   47837] = 32'hd552bb0b;
    ram_cell[   47838] = 32'h8f288b05;
    ram_cell[   47839] = 32'hc158d43c;
    ram_cell[   47840] = 32'h67b798a9;
    ram_cell[   47841] = 32'h8abc6a47;
    ram_cell[   47842] = 32'he2679cb4;
    ram_cell[   47843] = 32'h467d0a87;
    ram_cell[   47844] = 32'h56f0102a;
    ram_cell[   47845] = 32'h46a7fd60;
    ram_cell[   47846] = 32'ha570f70b;
    ram_cell[   47847] = 32'h4a45b6c4;
    ram_cell[   47848] = 32'h087c2da4;
    ram_cell[   47849] = 32'h1ed2a8a8;
    ram_cell[   47850] = 32'h727fbba9;
    ram_cell[   47851] = 32'h155bfcec;
    ram_cell[   47852] = 32'h3eb40e79;
    ram_cell[   47853] = 32'he03350e5;
    ram_cell[   47854] = 32'h55b867ca;
    ram_cell[   47855] = 32'hc8ab69e9;
    ram_cell[   47856] = 32'he085b370;
    ram_cell[   47857] = 32'h4d215808;
    ram_cell[   47858] = 32'hd96eadeb;
    ram_cell[   47859] = 32'hb67f2b99;
    ram_cell[   47860] = 32'h502c993f;
    ram_cell[   47861] = 32'h7ef060e4;
    ram_cell[   47862] = 32'h2d0b0f87;
    ram_cell[   47863] = 32'hbc90c738;
    ram_cell[   47864] = 32'h922691cb;
    ram_cell[   47865] = 32'hd46c7081;
    ram_cell[   47866] = 32'h33f356f6;
    ram_cell[   47867] = 32'h509a91a8;
    ram_cell[   47868] = 32'hf29786e0;
    ram_cell[   47869] = 32'h911d2f1a;
    ram_cell[   47870] = 32'h258e5b2a;
    ram_cell[   47871] = 32'haf71758f;
    ram_cell[   47872] = 32'hacc45a89;
    ram_cell[   47873] = 32'h779efa2d;
    ram_cell[   47874] = 32'hb1eeffae;
    ram_cell[   47875] = 32'h64bf6cdc;
    ram_cell[   47876] = 32'h2c303535;
    ram_cell[   47877] = 32'hfcc9e9fa;
    ram_cell[   47878] = 32'hdc0ff7c3;
    ram_cell[   47879] = 32'h56978d64;
    ram_cell[   47880] = 32'h2c0346ed;
    ram_cell[   47881] = 32'ha1e4dfa0;
    ram_cell[   47882] = 32'h316abd56;
    ram_cell[   47883] = 32'h953b280a;
    ram_cell[   47884] = 32'hfd298f98;
    ram_cell[   47885] = 32'h30dcffe8;
    ram_cell[   47886] = 32'h5dff523f;
    ram_cell[   47887] = 32'h03964659;
    ram_cell[   47888] = 32'h2d9ef413;
    ram_cell[   47889] = 32'hc160a187;
    ram_cell[   47890] = 32'h9a0dcdf7;
    ram_cell[   47891] = 32'h378c4db0;
    ram_cell[   47892] = 32'h4a8b9cda;
    ram_cell[   47893] = 32'ha280f926;
    ram_cell[   47894] = 32'haa43cf3d;
    ram_cell[   47895] = 32'h42b74b14;
    ram_cell[   47896] = 32'h209efa07;
    ram_cell[   47897] = 32'hd0f349ee;
    ram_cell[   47898] = 32'haf8a880a;
    ram_cell[   47899] = 32'h16f0566b;
    ram_cell[   47900] = 32'h101aa98a;
    ram_cell[   47901] = 32'hba2c16c9;
    ram_cell[   47902] = 32'h175d5d21;
    ram_cell[   47903] = 32'h7e643a7a;
    ram_cell[   47904] = 32'h0c398c34;
    ram_cell[   47905] = 32'heeba10bc;
    ram_cell[   47906] = 32'h7c7478ae;
    ram_cell[   47907] = 32'hffce07b0;
    ram_cell[   47908] = 32'h3a821a02;
    ram_cell[   47909] = 32'h31402b45;
    ram_cell[   47910] = 32'h5a1575af;
    ram_cell[   47911] = 32'haf8c4765;
    ram_cell[   47912] = 32'h0f54e035;
    ram_cell[   47913] = 32'h6f1b52fe;
    ram_cell[   47914] = 32'hf9ff5e51;
    ram_cell[   47915] = 32'hb861a9bc;
    ram_cell[   47916] = 32'hc110deef;
    ram_cell[   47917] = 32'h8e43be63;
    ram_cell[   47918] = 32'hfe6cbd5b;
    ram_cell[   47919] = 32'he4f79e40;
    ram_cell[   47920] = 32'h32a8dc86;
    ram_cell[   47921] = 32'h063a2511;
    ram_cell[   47922] = 32'h25269655;
    ram_cell[   47923] = 32'h7f32c61e;
    ram_cell[   47924] = 32'h5b82a6ca;
    ram_cell[   47925] = 32'h87eb69c1;
    ram_cell[   47926] = 32'ha0c4dc7f;
    ram_cell[   47927] = 32'hef1a1880;
    ram_cell[   47928] = 32'h8c82f57d;
    ram_cell[   47929] = 32'h83fdc57c;
    ram_cell[   47930] = 32'h38ec9b6b;
    ram_cell[   47931] = 32'hb2b636e6;
    ram_cell[   47932] = 32'h13a16a48;
    ram_cell[   47933] = 32'h17f11d8b;
    ram_cell[   47934] = 32'hfb60d37a;
    ram_cell[   47935] = 32'h3c095949;
    ram_cell[   47936] = 32'hdfdb0e8f;
    ram_cell[   47937] = 32'ha94c3c22;
    ram_cell[   47938] = 32'h8f647845;
    ram_cell[   47939] = 32'habd24430;
    ram_cell[   47940] = 32'hc30fbcd8;
    ram_cell[   47941] = 32'hb683041d;
    ram_cell[   47942] = 32'hb9f45045;
    ram_cell[   47943] = 32'h5d1736f3;
    ram_cell[   47944] = 32'h6df76b42;
    ram_cell[   47945] = 32'h575ef78f;
    ram_cell[   47946] = 32'h24d0dc3d;
    ram_cell[   47947] = 32'h94f937c6;
    ram_cell[   47948] = 32'head608ac;
    ram_cell[   47949] = 32'h0dd51ae7;
    ram_cell[   47950] = 32'h188c5fcc;
    ram_cell[   47951] = 32'h87094fc1;
    ram_cell[   47952] = 32'h6f943293;
    ram_cell[   47953] = 32'h1b2594f2;
    ram_cell[   47954] = 32'hd433ffee;
    ram_cell[   47955] = 32'h99f6f9cc;
    ram_cell[   47956] = 32'hfafe796b;
    ram_cell[   47957] = 32'h4ad25096;
    ram_cell[   47958] = 32'h46124e67;
    ram_cell[   47959] = 32'h826e9856;
    ram_cell[   47960] = 32'hb2d68db2;
    ram_cell[   47961] = 32'hea8d266d;
    ram_cell[   47962] = 32'h4d21c0fb;
    ram_cell[   47963] = 32'hf091d374;
    ram_cell[   47964] = 32'h68c99d85;
    ram_cell[   47965] = 32'hed3fdb0c;
    ram_cell[   47966] = 32'h5306dcc4;
    ram_cell[   47967] = 32'h838e8ca2;
    ram_cell[   47968] = 32'h862cd796;
    ram_cell[   47969] = 32'hb3ac6927;
    ram_cell[   47970] = 32'h89be9d8e;
    ram_cell[   47971] = 32'h50590be9;
    ram_cell[   47972] = 32'he8b72e7b;
    ram_cell[   47973] = 32'ha616fee7;
    ram_cell[   47974] = 32'h41e78bfa;
    ram_cell[   47975] = 32'hc69f43eb;
    ram_cell[   47976] = 32'h69fdf17d;
    ram_cell[   47977] = 32'h17f10728;
    ram_cell[   47978] = 32'hd135e556;
    ram_cell[   47979] = 32'h355f546a;
    ram_cell[   47980] = 32'h98dca923;
    ram_cell[   47981] = 32'he9e3297c;
    ram_cell[   47982] = 32'hafe8ee3e;
    ram_cell[   47983] = 32'hd5ad52c3;
    ram_cell[   47984] = 32'hf9740d71;
    ram_cell[   47985] = 32'hf388f4a1;
    ram_cell[   47986] = 32'ha865c9dc;
    ram_cell[   47987] = 32'hd457e018;
    ram_cell[   47988] = 32'hee1f7bb0;
    ram_cell[   47989] = 32'h23574f96;
    ram_cell[   47990] = 32'h662dbf64;
    ram_cell[   47991] = 32'h16de76c6;
    ram_cell[   47992] = 32'h38f32322;
    ram_cell[   47993] = 32'h87c687fc;
    ram_cell[   47994] = 32'h46d22f84;
    ram_cell[   47995] = 32'h13af14a5;
    ram_cell[   47996] = 32'he2d06229;
    ram_cell[   47997] = 32'h902bd687;
    ram_cell[   47998] = 32'hd1bada10;
    ram_cell[   47999] = 32'h4c1c097c;
    ram_cell[   48000] = 32'hba23166b;
    ram_cell[   48001] = 32'h6d5ad57d;
    ram_cell[   48002] = 32'h95635551;
    ram_cell[   48003] = 32'h8a74e79e;
    ram_cell[   48004] = 32'h38d5dc08;
    ram_cell[   48005] = 32'hebb80fde;
    ram_cell[   48006] = 32'h3282d772;
    ram_cell[   48007] = 32'h350336a0;
    ram_cell[   48008] = 32'h4000dd51;
    ram_cell[   48009] = 32'hc1dbfd8b;
    ram_cell[   48010] = 32'h31a7efcf;
    ram_cell[   48011] = 32'hc669da7d;
    ram_cell[   48012] = 32'hd86e11e1;
    ram_cell[   48013] = 32'hfbf7b695;
    ram_cell[   48014] = 32'h85a10d71;
    ram_cell[   48015] = 32'h65e90f22;
    ram_cell[   48016] = 32'h8656aa7d;
    ram_cell[   48017] = 32'h95e59b96;
    ram_cell[   48018] = 32'h5a8b4b96;
    ram_cell[   48019] = 32'h20bb6458;
    ram_cell[   48020] = 32'h795aff51;
    ram_cell[   48021] = 32'hcd634402;
    ram_cell[   48022] = 32'hc4e122c6;
    ram_cell[   48023] = 32'he7dbde0c;
    ram_cell[   48024] = 32'h797bf5cd;
    ram_cell[   48025] = 32'hb4c586a9;
    ram_cell[   48026] = 32'he5588ca2;
    ram_cell[   48027] = 32'h91443c67;
    ram_cell[   48028] = 32'h5887bf01;
    ram_cell[   48029] = 32'h12f9a28d;
    ram_cell[   48030] = 32'hd507581a;
    ram_cell[   48031] = 32'h690eb0f9;
    ram_cell[   48032] = 32'h17b82fbb;
    ram_cell[   48033] = 32'hec666171;
    ram_cell[   48034] = 32'h9a4ab75b;
    ram_cell[   48035] = 32'h6d813853;
    ram_cell[   48036] = 32'h018aa0b0;
    ram_cell[   48037] = 32'hf78abe81;
    ram_cell[   48038] = 32'ha8f5ff0d;
    ram_cell[   48039] = 32'h0f5c31ba;
    ram_cell[   48040] = 32'hdbf90561;
    ram_cell[   48041] = 32'h48d0a580;
    ram_cell[   48042] = 32'hf1a2f889;
    ram_cell[   48043] = 32'ha43ebb69;
    ram_cell[   48044] = 32'he04514bb;
    ram_cell[   48045] = 32'h9d8699c3;
    ram_cell[   48046] = 32'h2d4172d5;
    ram_cell[   48047] = 32'h49d99e7b;
    ram_cell[   48048] = 32'h8132884e;
    ram_cell[   48049] = 32'h43a755a8;
    ram_cell[   48050] = 32'hfe81ab68;
    ram_cell[   48051] = 32'hc001ea9b;
    ram_cell[   48052] = 32'h740016fb;
    ram_cell[   48053] = 32'h1d8a7733;
    ram_cell[   48054] = 32'ha0b25008;
    ram_cell[   48055] = 32'hccf3934f;
    ram_cell[   48056] = 32'h56e48cf9;
    ram_cell[   48057] = 32'h82769c49;
    ram_cell[   48058] = 32'h32a2360b;
    ram_cell[   48059] = 32'hef03645a;
    ram_cell[   48060] = 32'hbc07c46c;
    ram_cell[   48061] = 32'h01fc454e;
    ram_cell[   48062] = 32'hf4388501;
    ram_cell[   48063] = 32'h6bc9cd0d;
    ram_cell[   48064] = 32'h5ea5d0d5;
    ram_cell[   48065] = 32'hc6851790;
    ram_cell[   48066] = 32'h08504365;
    ram_cell[   48067] = 32'ha37a5428;
    ram_cell[   48068] = 32'hd0a3d86f;
    ram_cell[   48069] = 32'hdd870b33;
    ram_cell[   48070] = 32'hd5b421f2;
    ram_cell[   48071] = 32'h79b6aa65;
    ram_cell[   48072] = 32'ha780f234;
    ram_cell[   48073] = 32'h8a2c3caa;
    ram_cell[   48074] = 32'hc7b489e0;
    ram_cell[   48075] = 32'hffbe432d;
    ram_cell[   48076] = 32'he3119853;
    ram_cell[   48077] = 32'hd0cf7f20;
    ram_cell[   48078] = 32'hf69e7eb6;
    ram_cell[   48079] = 32'h663b9713;
    ram_cell[   48080] = 32'h6d1cc9c5;
    ram_cell[   48081] = 32'h3148d243;
    ram_cell[   48082] = 32'h125452c5;
    ram_cell[   48083] = 32'hfd43bd73;
    ram_cell[   48084] = 32'h2e00398c;
    ram_cell[   48085] = 32'hfd67ce72;
    ram_cell[   48086] = 32'h4d0ef2b6;
    ram_cell[   48087] = 32'h17ea555e;
    ram_cell[   48088] = 32'hd8df9c44;
    ram_cell[   48089] = 32'hb0eca561;
    ram_cell[   48090] = 32'hc0939cd6;
    ram_cell[   48091] = 32'h5f187dab;
    ram_cell[   48092] = 32'h6c4a3521;
    ram_cell[   48093] = 32'hdec85309;
    ram_cell[   48094] = 32'hc6fe9011;
    ram_cell[   48095] = 32'h2a2bb824;
    ram_cell[   48096] = 32'h9f1788eb;
    ram_cell[   48097] = 32'hca944817;
    ram_cell[   48098] = 32'heb9fdd60;
    ram_cell[   48099] = 32'hbf7133c1;
    ram_cell[   48100] = 32'he8e230a1;
    ram_cell[   48101] = 32'h6650e824;
    ram_cell[   48102] = 32'h44dec543;
    ram_cell[   48103] = 32'hda3f30fe;
    ram_cell[   48104] = 32'he9b08f85;
    ram_cell[   48105] = 32'hcd0ed0a3;
    ram_cell[   48106] = 32'h74cf2c65;
    ram_cell[   48107] = 32'h3678fbd0;
    ram_cell[   48108] = 32'h57dcdf29;
    ram_cell[   48109] = 32'h6c003282;
    ram_cell[   48110] = 32'hecfd26e3;
    ram_cell[   48111] = 32'h3ca33b38;
    ram_cell[   48112] = 32'h48b383f0;
    ram_cell[   48113] = 32'hcec61856;
    ram_cell[   48114] = 32'hbdf62ae2;
    ram_cell[   48115] = 32'heefbc7ad;
    ram_cell[   48116] = 32'h6e5ec059;
    ram_cell[   48117] = 32'h2e519f51;
    ram_cell[   48118] = 32'hdf2d7942;
    ram_cell[   48119] = 32'hdf8d22a0;
    ram_cell[   48120] = 32'h994d05fd;
    ram_cell[   48121] = 32'h87c31cbe;
    ram_cell[   48122] = 32'hc8831460;
    ram_cell[   48123] = 32'h9236989e;
    ram_cell[   48124] = 32'h67c6c2d1;
    ram_cell[   48125] = 32'he5c765bc;
    ram_cell[   48126] = 32'h3e3eda47;
    ram_cell[   48127] = 32'h699b3889;
    ram_cell[   48128] = 32'h2dfe5fb5;
    ram_cell[   48129] = 32'h1a04d801;
    ram_cell[   48130] = 32'h52d1447f;
    ram_cell[   48131] = 32'h3500c26e;
    ram_cell[   48132] = 32'h717d7266;
    ram_cell[   48133] = 32'h3c945fbd;
    ram_cell[   48134] = 32'h65dc7d99;
    ram_cell[   48135] = 32'hbc8990b8;
    ram_cell[   48136] = 32'hafb57f05;
    ram_cell[   48137] = 32'hfa8f42a4;
    ram_cell[   48138] = 32'hdd7ea38c;
    ram_cell[   48139] = 32'haec8c712;
    ram_cell[   48140] = 32'ha19b645f;
    ram_cell[   48141] = 32'h028ef75e;
    ram_cell[   48142] = 32'h41e2c239;
    ram_cell[   48143] = 32'hfb32a55e;
    ram_cell[   48144] = 32'hc45cc320;
    ram_cell[   48145] = 32'h666658ca;
    ram_cell[   48146] = 32'ha32e4bf4;
    ram_cell[   48147] = 32'he9d30146;
    ram_cell[   48148] = 32'hee2dbf82;
    ram_cell[   48149] = 32'h7475ce9a;
    ram_cell[   48150] = 32'hdae887b3;
    ram_cell[   48151] = 32'h22fbde23;
    ram_cell[   48152] = 32'h16394309;
    ram_cell[   48153] = 32'hc0f452c9;
    ram_cell[   48154] = 32'h9badd306;
    ram_cell[   48155] = 32'h6524a2a6;
    ram_cell[   48156] = 32'he46a2cea;
    ram_cell[   48157] = 32'h024077cc;
    ram_cell[   48158] = 32'hb5857d70;
    ram_cell[   48159] = 32'h62326071;
    ram_cell[   48160] = 32'he4473bb4;
    ram_cell[   48161] = 32'hf67fa6a6;
    ram_cell[   48162] = 32'h9ec0dbcc;
    ram_cell[   48163] = 32'h7e0f3ef4;
    ram_cell[   48164] = 32'h3e745ace;
    ram_cell[   48165] = 32'hff8801c6;
    ram_cell[   48166] = 32'h21922788;
    ram_cell[   48167] = 32'haf7b2349;
    ram_cell[   48168] = 32'hedfd913f;
    ram_cell[   48169] = 32'hd307b57d;
    ram_cell[   48170] = 32'h73be42ad;
    ram_cell[   48171] = 32'h06ec6ba0;
    ram_cell[   48172] = 32'h37b339bc;
    ram_cell[   48173] = 32'hfccc9fd2;
    ram_cell[   48174] = 32'h9dd962ab;
    ram_cell[   48175] = 32'hd1847160;
    ram_cell[   48176] = 32'hde748266;
    ram_cell[   48177] = 32'hfd34d148;
    ram_cell[   48178] = 32'heed7dcc4;
    ram_cell[   48179] = 32'hd8fff752;
    ram_cell[   48180] = 32'h6a21afc8;
    ram_cell[   48181] = 32'h575c5a74;
    ram_cell[   48182] = 32'hddd86ef2;
    ram_cell[   48183] = 32'hf6eb6d7e;
    ram_cell[   48184] = 32'h60b233d9;
    ram_cell[   48185] = 32'h1be6c2b3;
    ram_cell[   48186] = 32'h9f460506;
    ram_cell[   48187] = 32'h56a582b0;
    ram_cell[   48188] = 32'h6bb99a9b;
    ram_cell[   48189] = 32'h4724d9eb;
    ram_cell[   48190] = 32'h2c8a1e25;
    ram_cell[   48191] = 32'h644c2d8b;
    ram_cell[   48192] = 32'h5cdc135b;
    ram_cell[   48193] = 32'h9c1ee8a4;
    ram_cell[   48194] = 32'h93b831b4;
    ram_cell[   48195] = 32'hbf61d4e1;
    ram_cell[   48196] = 32'h2087dc60;
    ram_cell[   48197] = 32'hf6362e7c;
    ram_cell[   48198] = 32'h529416b6;
    ram_cell[   48199] = 32'h594685e6;
    ram_cell[   48200] = 32'h967b5f16;
    ram_cell[   48201] = 32'h721fa50b;
    ram_cell[   48202] = 32'h13b6242e;
    ram_cell[   48203] = 32'h4ada5e37;
    ram_cell[   48204] = 32'h0c23e2c8;
    ram_cell[   48205] = 32'h7f25b5d7;
    ram_cell[   48206] = 32'h7a39b624;
    ram_cell[   48207] = 32'h6e7628e7;
    ram_cell[   48208] = 32'hd74d5887;
    ram_cell[   48209] = 32'h20e3b080;
    ram_cell[   48210] = 32'h2ed53274;
    ram_cell[   48211] = 32'h1390e67b;
    ram_cell[   48212] = 32'hd65d1fd1;
    ram_cell[   48213] = 32'h793768b4;
    ram_cell[   48214] = 32'hcb2f56ef;
    ram_cell[   48215] = 32'hf324564c;
    ram_cell[   48216] = 32'he685d5d6;
    ram_cell[   48217] = 32'h208efa7d;
    ram_cell[   48218] = 32'he01da0d1;
    ram_cell[   48219] = 32'hc0a3afb5;
    ram_cell[   48220] = 32'h6a69d4d5;
    ram_cell[   48221] = 32'haa785760;
    ram_cell[   48222] = 32'hc2e20bd2;
    ram_cell[   48223] = 32'hc7198052;
    ram_cell[   48224] = 32'h958be8f3;
    ram_cell[   48225] = 32'h01341c01;
    ram_cell[   48226] = 32'h68f6df80;
    ram_cell[   48227] = 32'hace95a2c;
    ram_cell[   48228] = 32'h4d5860b4;
    ram_cell[   48229] = 32'h3f332a5c;
    ram_cell[   48230] = 32'hd62c27ff;
    ram_cell[   48231] = 32'h4aa1d72a;
    ram_cell[   48232] = 32'h580d376d;
    ram_cell[   48233] = 32'h8b216ffb;
    ram_cell[   48234] = 32'h95ca2ba9;
    ram_cell[   48235] = 32'h6fca347a;
    ram_cell[   48236] = 32'hdc2516fc;
    ram_cell[   48237] = 32'h55545ced;
    ram_cell[   48238] = 32'h529c64f1;
    ram_cell[   48239] = 32'hba3ca8e9;
    ram_cell[   48240] = 32'h9e6ac4e0;
    ram_cell[   48241] = 32'he77263ce;
    ram_cell[   48242] = 32'h554e4856;
    ram_cell[   48243] = 32'h5be84c71;
    ram_cell[   48244] = 32'h33d308d3;
    ram_cell[   48245] = 32'h9af6a240;
    ram_cell[   48246] = 32'he492eea0;
    ram_cell[   48247] = 32'hf12da34f;
    ram_cell[   48248] = 32'hd5984dfe;
    ram_cell[   48249] = 32'hd480ec7a;
    ram_cell[   48250] = 32'h08ab488d;
    ram_cell[   48251] = 32'h72a1ae33;
    ram_cell[   48252] = 32'h7879eaa2;
    ram_cell[   48253] = 32'h3bd0b03c;
    ram_cell[   48254] = 32'h52475301;
    ram_cell[   48255] = 32'hd6f5793e;
    ram_cell[   48256] = 32'h683ce676;
    ram_cell[   48257] = 32'h8f691d6a;
    ram_cell[   48258] = 32'ha6312d1c;
    ram_cell[   48259] = 32'h11e3ffe9;
    ram_cell[   48260] = 32'h96058a3c;
    ram_cell[   48261] = 32'h46db1179;
    ram_cell[   48262] = 32'h6ea27b80;
    ram_cell[   48263] = 32'hf762bd9d;
    ram_cell[   48264] = 32'hdb93d59a;
    ram_cell[   48265] = 32'h3fb5c71c;
    ram_cell[   48266] = 32'h506aa2c9;
    ram_cell[   48267] = 32'hf350246b;
    ram_cell[   48268] = 32'h952994d1;
    ram_cell[   48269] = 32'h56d8cee9;
    ram_cell[   48270] = 32'h603e197f;
    ram_cell[   48271] = 32'h234f9d35;
    ram_cell[   48272] = 32'haf498ff2;
    ram_cell[   48273] = 32'h2fd1cacf;
    ram_cell[   48274] = 32'h50b17f27;
    ram_cell[   48275] = 32'h947407b1;
    ram_cell[   48276] = 32'h474cf80f;
    ram_cell[   48277] = 32'hc5dd32b0;
    ram_cell[   48278] = 32'h61cfa167;
    ram_cell[   48279] = 32'hf8d7d453;
    ram_cell[   48280] = 32'h3edbe783;
    ram_cell[   48281] = 32'hf362bd7f;
    ram_cell[   48282] = 32'h52bd2170;
    ram_cell[   48283] = 32'he892b47f;
    ram_cell[   48284] = 32'h34b1ca1d;
    ram_cell[   48285] = 32'h3a27b876;
    ram_cell[   48286] = 32'h9a911891;
    ram_cell[   48287] = 32'hb05e4928;
    ram_cell[   48288] = 32'h6772c479;
    ram_cell[   48289] = 32'h00bf7c1a;
    ram_cell[   48290] = 32'h977f12a4;
    ram_cell[   48291] = 32'h655ab8a9;
    ram_cell[   48292] = 32'h60f2d7ac;
    ram_cell[   48293] = 32'h806c95fd;
    ram_cell[   48294] = 32'h954f4fd4;
    ram_cell[   48295] = 32'hef295b3a;
    ram_cell[   48296] = 32'h80e53cb3;
    ram_cell[   48297] = 32'hed513a1f;
    ram_cell[   48298] = 32'hcb056e3f;
    ram_cell[   48299] = 32'h38ef77be;
    ram_cell[   48300] = 32'h7864d181;
    ram_cell[   48301] = 32'had15bc25;
    ram_cell[   48302] = 32'h0ece70f3;
    ram_cell[   48303] = 32'hd319a8fd;
    ram_cell[   48304] = 32'hd5562d55;
    ram_cell[   48305] = 32'he775cd24;
    ram_cell[   48306] = 32'h7efb4aad;
    ram_cell[   48307] = 32'h03327d8e;
    ram_cell[   48308] = 32'hf2be105a;
    ram_cell[   48309] = 32'hdf8040d5;
    ram_cell[   48310] = 32'h864fc6c9;
    ram_cell[   48311] = 32'h8ca05a1d;
    ram_cell[   48312] = 32'heaba5b34;
    ram_cell[   48313] = 32'h04eda4d6;
    ram_cell[   48314] = 32'h6b261694;
    ram_cell[   48315] = 32'h1991b345;
    ram_cell[   48316] = 32'hea627b0a;
    ram_cell[   48317] = 32'h2ee9e560;
    ram_cell[   48318] = 32'h782c1489;
    ram_cell[   48319] = 32'h14d29c76;
    ram_cell[   48320] = 32'hcf27b9bb;
    ram_cell[   48321] = 32'ha3d97d0d;
    ram_cell[   48322] = 32'h184ce5b6;
    ram_cell[   48323] = 32'hb0a5ab3f;
    ram_cell[   48324] = 32'h7a426cb8;
    ram_cell[   48325] = 32'ha7302cf8;
    ram_cell[   48326] = 32'hf4998dc3;
    ram_cell[   48327] = 32'hb2bffbb2;
    ram_cell[   48328] = 32'h6f88c4f9;
    ram_cell[   48329] = 32'h3d929c35;
    ram_cell[   48330] = 32'hd0ab4007;
    ram_cell[   48331] = 32'hdbc23b1e;
    ram_cell[   48332] = 32'h45ac8567;
    ram_cell[   48333] = 32'h13190d43;
    ram_cell[   48334] = 32'hda52e31a;
    ram_cell[   48335] = 32'h0b4147d7;
    ram_cell[   48336] = 32'he878f7ce;
    ram_cell[   48337] = 32'h5d51b855;
    ram_cell[   48338] = 32'he1294570;
    ram_cell[   48339] = 32'h9d3214ee;
    ram_cell[   48340] = 32'hf48d3aff;
    ram_cell[   48341] = 32'h04a8dbdb;
    ram_cell[   48342] = 32'hc254a09f;
    ram_cell[   48343] = 32'h7ef6639c;
    ram_cell[   48344] = 32'h5adae9d6;
    ram_cell[   48345] = 32'h95b39228;
    ram_cell[   48346] = 32'h7b7b3ad4;
    ram_cell[   48347] = 32'h1785b94b;
    ram_cell[   48348] = 32'had557fc5;
    ram_cell[   48349] = 32'h8701365a;
    ram_cell[   48350] = 32'h19033eed;
    ram_cell[   48351] = 32'he727372f;
    ram_cell[   48352] = 32'hb6131666;
    ram_cell[   48353] = 32'ha8f788d1;
    ram_cell[   48354] = 32'hdb9d5aad;
    ram_cell[   48355] = 32'h11350318;
    ram_cell[   48356] = 32'h5cd5b011;
    ram_cell[   48357] = 32'h5e57a110;
    ram_cell[   48358] = 32'hb73f497d;
    ram_cell[   48359] = 32'hba1c3278;
    ram_cell[   48360] = 32'h7f14f8e4;
    ram_cell[   48361] = 32'h46cf90a4;
    ram_cell[   48362] = 32'ha57e65a0;
    ram_cell[   48363] = 32'he0369545;
    ram_cell[   48364] = 32'h9c7b73f7;
    ram_cell[   48365] = 32'h876be2e9;
    ram_cell[   48366] = 32'hf2519e21;
    ram_cell[   48367] = 32'hd809bd10;
    ram_cell[   48368] = 32'h392fd6df;
    ram_cell[   48369] = 32'h39686356;
    ram_cell[   48370] = 32'h187758ad;
    ram_cell[   48371] = 32'h84c8e786;
    ram_cell[   48372] = 32'hb4374649;
    ram_cell[   48373] = 32'h03cab12f;
    ram_cell[   48374] = 32'h93285187;
    ram_cell[   48375] = 32'h23c66d88;
    ram_cell[   48376] = 32'hf9598db7;
    ram_cell[   48377] = 32'h72f4d79b;
    ram_cell[   48378] = 32'hb9f32d4f;
    ram_cell[   48379] = 32'hb3cc7bf4;
    ram_cell[   48380] = 32'h7c69d32a;
    ram_cell[   48381] = 32'hec006b8a;
    ram_cell[   48382] = 32'hbb7f03e6;
    ram_cell[   48383] = 32'he9641d43;
    ram_cell[   48384] = 32'h88258a5a;
    ram_cell[   48385] = 32'hc005fea0;
    ram_cell[   48386] = 32'h5f456992;
    ram_cell[   48387] = 32'h217b424b;
    ram_cell[   48388] = 32'h2686c443;
    ram_cell[   48389] = 32'h80c87401;
    ram_cell[   48390] = 32'h82ad77ee;
    ram_cell[   48391] = 32'h40f262c8;
    ram_cell[   48392] = 32'hae0097d2;
    ram_cell[   48393] = 32'h2e28e98c;
    ram_cell[   48394] = 32'hd1b2e75d;
    ram_cell[   48395] = 32'h4ac16634;
    ram_cell[   48396] = 32'hf7beb3f5;
    ram_cell[   48397] = 32'h056b69ce;
    ram_cell[   48398] = 32'h50dad7fb;
    ram_cell[   48399] = 32'h3235af0c;
    ram_cell[   48400] = 32'hca3a43cb;
    ram_cell[   48401] = 32'hfd2e7979;
    ram_cell[   48402] = 32'h3dcd77c0;
    ram_cell[   48403] = 32'he0eeb165;
    ram_cell[   48404] = 32'hf159f2d9;
    ram_cell[   48405] = 32'h21b92bf2;
    ram_cell[   48406] = 32'h9aa28b35;
    ram_cell[   48407] = 32'h8477c956;
    ram_cell[   48408] = 32'h15c6cbda;
    ram_cell[   48409] = 32'h1acb1da1;
    ram_cell[   48410] = 32'h86e405d1;
    ram_cell[   48411] = 32'hd5851525;
    ram_cell[   48412] = 32'hae71b9e8;
    ram_cell[   48413] = 32'h04cf8328;
    ram_cell[   48414] = 32'h80542951;
    ram_cell[   48415] = 32'h05713fc2;
    ram_cell[   48416] = 32'hbca450fd;
    ram_cell[   48417] = 32'hb604410a;
    ram_cell[   48418] = 32'h410de9ef;
    ram_cell[   48419] = 32'h116c1063;
    ram_cell[   48420] = 32'h7fc2b933;
    ram_cell[   48421] = 32'h72b2ab28;
    ram_cell[   48422] = 32'h7a8e244a;
    ram_cell[   48423] = 32'ha5b8c3b6;
    ram_cell[   48424] = 32'h06480cae;
    ram_cell[   48425] = 32'h052b3971;
    ram_cell[   48426] = 32'hb8ac967a;
    ram_cell[   48427] = 32'hd70870e1;
    ram_cell[   48428] = 32'h9d7aa48c;
    ram_cell[   48429] = 32'h2a0a63e1;
    ram_cell[   48430] = 32'h5f0fa821;
    ram_cell[   48431] = 32'h367a77b1;
    ram_cell[   48432] = 32'hd44e0124;
    ram_cell[   48433] = 32'hfc5e46da;
    ram_cell[   48434] = 32'h2bd19f1b;
    ram_cell[   48435] = 32'h1c572f07;
    ram_cell[   48436] = 32'hf545d552;
    ram_cell[   48437] = 32'h58a160f5;
    ram_cell[   48438] = 32'h593fb413;
    ram_cell[   48439] = 32'h3ae40996;
    ram_cell[   48440] = 32'hdfa7082c;
    ram_cell[   48441] = 32'h0236feb6;
    ram_cell[   48442] = 32'h138657b7;
    ram_cell[   48443] = 32'h6aca628b;
    ram_cell[   48444] = 32'hfb8bffac;
    ram_cell[   48445] = 32'he3794b34;
    ram_cell[   48446] = 32'h122f97da;
    ram_cell[   48447] = 32'ha39c7fcf;
    ram_cell[   48448] = 32'hcd5f3904;
    ram_cell[   48449] = 32'ha049dc22;
    ram_cell[   48450] = 32'hdc85dcca;
    ram_cell[   48451] = 32'he9a2e11a;
    ram_cell[   48452] = 32'h757787e4;
    ram_cell[   48453] = 32'h17769a4b;
    ram_cell[   48454] = 32'hdf68574e;
    ram_cell[   48455] = 32'h422afc19;
    ram_cell[   48456] = 32'hc5dab536;
    ram_cell[   48457] = 32'hf3d7f4da;
    ram_cell[   48458] = 32'h9c03c2b5;
    ram_cell[   48459] = 32'h38f8ef3c;
    ram_cell[   48460] = 32'he2692efb;
    ram_cell[   48461] = 32'h2c1c4c65;
    ram_cell[   48462] = 32'hef8d2ddc;
    ram_cell[   48463] = 32'hf7a6b103;
    ram_cell[   48464] = 32'ha3fa9cf4;
    ram_cell[   48465] = 32'he161706a;
    ram_cell[   48466] = 32'hbf31abb5;
    ram_cell[   48467] = 32'ha9f6954d;
    ram_cell[   48468] = 32'hb51c238b;
    ram_cell[   48469] = 32'h2b6560fd;
    ram_cell[   48470] = 32'ha1964fd6;
    ram_cell[   48471] = 32'h42c35ef6;
    ram_cell[   48472] = 32'hc0218f94;
    ram_cell[   48473] = 32'hfa56dee9;
    ram_cell[   48474] = 32'h55558ab9;
    ram_cell[   48475] = 32'h1c407a07;
    ram_cell[   48476] = 32'h103d8d65;
    ram_cell[   48477] = 32'h26d70521;
    ram_cell[   48478] = 32'hac588883;
    ram_cell[   48479] = 32'h11f5e9ce;
    ram_cell[   48480] = 32'h56194a9b;
    ram_cell[   48481] = 32'hcbaf720b;
    ram_cell[   48482] = 32'h42a559d0;
    ram_cell[   48483] = 32'h473bedc3;
    ram_cell[   48484] = 32'h0b02bd56;
    ram_cell[   48485] = 32'h6ba275a5;
    ram_cell[   48486] = 32'he79e5928;
    ram_cell[   48487] = 32'h0fd3ae78;
    ram_cell[   48488] = 32'hf14067e3;
    ram_cell[   48489] = 32'hd9156aa8;
    ram_cell[   48490] = 32'h2cfc44d6;
    ram_cell[   48491] = 32'h66c9bf04;
    ram_cell[   48492] = 32'h06383aae;
    ram_cell[   48493] = 32'hbb638b26;
    ram_cell[   48494] = 32'h63427e0f;
    ram_cell[   48495] = 32'h97c2243a;
    ram_cell[   48496] = 32'hb24664b8;
    ram_cell[   48497] = 32'hccbee035;
    ram_cell[   48498] = 32'h935ed94f;
    ram_cell[   48499] = 32'hcd69b405;
    ram_cell[   48500] = 32'h286615cf;
    ram_cell[   48501] = 32'h4b637aac;
    ram_cell[   48502] = 32'h18d37bf1;
    ram_cell[   48503] = 32'h34cf6044;
    ram_cell[   48504] = 32'h375dbece;
    ram_cell[   48505] = 32'hf907492b;
    ram_cell[   48506] = 32'hfd590c33;
    ram_cell[   48507] = 32'h00ee073a;
    ram_cell[   48508] = 32'h206400f1;
    ram_cell[   48509] = 32'h372c0c66;
    ram_cell[   48510] = 32'h9d99a264;
    ram_cell[   48511] = 32'h7f946f74;
    ram_cell[   48512] = 32'hb6778d32;
    ram_cell[   48513] = 32'h98b66eef;
    ram_cell[   48514] = 32'h4c8b4240;
    ram_cell[   48515] = 32'h5f8d6ddc;
    ram_cell[   48516] = 32'h2f3c173c;
    ram_cell[   48517] = 32'ha2d73547;
    ram_cell[   48518] = 32'h1c7d08fa;
    ram_cell[   48519] = 32'h12a269a5;
    ram_cell[   48520] = 32'hfb873d86;
    ram_cell[   48521] = 32'h0ef4c4bf;
    ram_cell[   48522] = 32'hb13b98c2;
    ram_cell[   48523] = 32'h952b3a65;
    ram_cell[   48524] = 32'h156e15ba;
    ram_cell[   48525] = 32'hde91051f;
    ram_cell[   48526] = 32'h5327bb0a;
    ram_cell[   48527] = 32'h4acdad51;
    ram_cell[   48528] = 32'h81f9ac63;
    ram_cell[   48529] = 32'hb4808b46;
    ram_cell[   48530] = 32'h65269f49;
    ram_cell[   48531] = 32'h4180dc46;
    ram_cell[   48532] = 32'h1bb60831;
    ram_cell[   48533] = 32'hb5573867;
    ram_cell[   48534] = 32'h41029b5b;
    ram_cell[   48535] = 32'h59743d72;
    ram_cell[   48536] = 32'h4ea839b2;
    ram_cell[   48537] = 32'hc6000487;
    ram_cell[   48538] = 32'h62e90220;
    ram_cell[   48539] = 32'h06a99681;
    ram_cell[   48540] = 32'h84f9bd8b;
    ram_cell[   48541] = 32'hb77dad65;
    ram_cell[   48542] = 32'h93a232a3;
    ram_cell[   48543] = 32'h0356e25c;
    ram_cell[   48544] = 32'h7f307a65;
    ram_cell[   48545] = 32'haa11235b;
    ram_cell[   48546] = 32'h4cac3e5b;
    ram_cell[   48547] = 32'h4d23c850;
    ram_cell[   48548] = 32'hd2d1e87b;
    ram_cell[   48549] = 32'h18818864;
    ram_cell[   48550] = 32'hccea5ee4;
    ram_cell[   48551] = 32'hc1c52dc0;
    ram_cell[   48552] = 32'h8a7d172c;
    ram_cell[   48553] = 32'h3b7444a4;
    ram_cell[   48554] = 32'hbfe6f36a;
    ram_cell[   48555] = 32'h8d0e4892;
    ram_cell[   48556] = 32'h00f94e1c;
    ram_cell[   48557] = 32'h64dcadf5;
    ram_cell[   48558] = 32'hec2517bb;
    ram_cell[   48559] = 32'h3b6085d9;
    ram_cell[   48560] = 32'ha6420bce;
    ram_cell[   48561] = 32'hee40cace;
    ram_cell[   48562] = 32'h6c4fec2c;
    ram_cell[   48563] = 32'hf08eec37;
    ram_cell[   48564] = 32'h8c9105a9;
    ram_cell[   48565] = 32'he811d514;
    ram_cell[   48566] = 32'h8f49b82c;
    ram_cell[   48567] = 32'haf66ecde;
    ram_cell[   48568] = 32'h49b56237;
    ram_cell[   48569] = 32'h9af829cb;
    ram_cell[   48570] = 32'h710ca31b;
    ram_cell[   48571] = 32'ha4589f5d;
    ram_cell[   48572] = 32'h2ca616cc;
    ram_cell[   48573] = 32'he42a1f5f;
    ram_cell[   48574] = 32'h361c72bb;
    ram_cell[   48575] = 32'h41fcc598;
    ram_cell[   48576] = 32'ha0eee615;
    ram_cell[   48577] = 32'h50445342;
    ram_cell[   48578] = 32'h4b49d12b;
    ram_cell[   48579] = 32'he53e0332;
    ram_cell[   48580] = 32'hcda7d290;
    ram_cell[   48581] = 32'h6362fd8a;
    ram_cell[   48582] = 32'h64bfd2db;
    ram_cell[   48583] = 32'he59ca5ba;
    ram_cell[   48584] = 32'h73d4cc2f;
    ram_cell[   48585] = 32'h6131e063;
    ram_cell[   48586] = 32'h5d463878;
    ram_cell[   48587] = 32'h478923a6;
    ram_cell[   48588] = 32'hdfad9377;
    ram_cell[   48589] = 32'ha6ddfe52;
    ram_cell[   48590] = 32'he06c2402;
    ram_cell[   48591] = 32'h7336dec8;
    ram_cell[   48592] = 32'hf9c52c57;
    ram_cell[   48593] = 32'h00d9ef50;
    ram_cell[   48594] = 32'h68403041;
    ram_cell[   48595] = 32'hac7afe41;
    ram_cell[   48596] = 32'hec71478b;
    ram_cell[   48597] = 32'hef447a5e;
    ram_cell[   48598] = 32'hf4d50bdc;
    ram_cell[   48599] = 32'h35689df5;
    ram_cell[   48600] = 32'h47609026;
    ram_cell[   48601] = 32'h2329aadb;
    ram_cell[   48602] = 32'h02b56b93;
    ram_cell[   48603] = 32'hbe0b32c2;
    ram_cell[   48604] = 32'h24cfa288;
    ram_cell[   48605] = 32'h3e4aace5;
    ram_cell[   48606] = 32'hf17a33cc;
    ram_cell[   48607] = 32'hc4d31571;
    ram_cell[   48608] = 32'h67cb1e68;
    ram_cell[   48609] = 32'h1c7865ec;
    ram_cell[   48610] = 32'h6a83f7e1;
    ram_cell[   48611] = 32'h454d66d3;
    ram_cell[   48612] = 32'h7260c683;
    ram_cell[   48613] = 32'h18841cd9;
    ram_cell[   48614] = 32'h5869077f;
    ram_cell[   48615] = 32'h950f497b;
    ram_cell[   48616] = 32'hfcd63618;
    ram_cell[   48617] = 32'hefcd0c91;
    ram_cell[   48618] = 32'h2181f1d3;
    ram_cell[   48619] = 32'ha4b6286a;
    ram_cell[   48620] = 32'h10a89566;
    ram_cell[   48621] = 32'hef8c37d2;
    ram_cell[   48622] = 32'h5ef4c39a;
    ram_cell[   48623] = 32'heec1d3ec;
    ram_cell[   48624] = 32'hb99fde0b;
    ram_cell[   48625] = 32'hc8c6c69a;
    ram_cell[   48626] = 32'h4e095eac;
    ram_cell[   48627] = 32'h07395030;
    ram_cell[   48628] = 32'h5294977d;
    ram_cell[   48629] = 32'hc9b4cc01;
    ram_cell[   48630] = 32'h9e6317a9;
    ram_cell[   48631] = 32'h64185e17;
    ram_cell[   48632] = 32'h64b5fa59;
    ram_cell[   48633] = 32'h155b9219;
    ram_cell[   48634] = 32'hfe6c61c7;
    ram_cell[   48635] = 32'h559c6519;
    ram_cell[   48636] = 32'h926557e9;
    ram_cell[   48637] = 32'hda6aa4fc;
    ram_cell[   48638] = 32'h73bd0fc8;
    ram_cell[   48639] = 32'haf0dbdc3;
    ram_cell[   48640] = 32'hb7bf79a2;
    ram_cell[   48641] = 32'h4364baef;
    ram_cell[   48642] = 32'h406a0b97;
    ram_cell[   48643] = 32'h747d1e57;
    ram_cell[   48644] = 32'h1ee5232f;
    ram_cell[   48645] = 32'hf1e36e5c;
    ram_cell[   48646] = 32'h12716453;
    ram_cell[   48647] = 32'h579c28c4;
    ram_cell[   48648] = 32'h1869feb1;
    ram_cell[   48649] = 32'hb3d63612;
    ram_cell[   48650] = 32'h49b6a9c7;
    ram_cell[   48651] = 32'h9fb1bb41;
    ram_cell[   48652] = 32'hda2a73f2;
    ram_cell[   48653] = 32'h8bb47b55;
    ram_cell[   48654] = 32'h7dd26cdd;
    ram_cell[   48655] = 32'h260615cc;
    ram_cell[   48656] = 32'had118afb;
    ram_cell[   48657] = 32'h350860e6;
    ram_cell[   48658] = 32'h0eac4ba8;
    ram_cell[   48659] = 32'h5cee552f;
    ram_cell[   48660] = 32'ha94ab6de;
    ram_cell[   48661] = 32'he63642db;
    ram_cell[   48662] = 32'hdaa436e5;
    ram_cell[   48663] = 32'he71f61a1;
    ram_cell[   48664] = 32'hed53de78;
    ram_cell[   48665] = 32'hd429d485;
    ram_cell[   48666] = 32'h6493a9e6;
    ram_cell[   48667] = 32'h6de6d31f;
    ram_cell[   48668] = 32'he01797ba;
    ram_cell[   48669] = 32'h6319e4d1;
    ram_cell[   48670] = 32'ha2f2d5b0;
    ram_cell[   48671] = 32'hb2e60a92;
    ram_cell[   48672] = 32'he801bc98;
    ram_cell[   48673] = 32'h02bea917;
    ram_cell[   48674] = 32'h3b84c139;
    ram_cell[   48675] = 32'h86a401b2;
    ram_cell[   48676] = 32'haebba0d5;
    ram_cell[   48677] = 32'h3613f5bb;
    ram_cell[   48678] = 32'h7e50e80f;
    ram_cell[   48679] = 32'h710a6861;
    ram_cell[   48680] = 32'h108031d3;
    ram_cell[   48681] = 32'h831ded18;
    ram_cell[   48682] = 32'h3c073f68;
    ram_cell[   48683] = 32'hd2a246d2;
    ram_cell[   48684] = 32'hcc92c833;
    ram_cell[   48685] = 32'h642f42d0;
    ram_cell[   48686] = 32'hb5a56f71;
    ram_cell[   48687] = 32'hfee1a5ce;
    ram_cell[   48688] = 32'h0413bc5d;
    ram_cell[   48689] = 32'h700fcae4;
    ram_cell[   48690] = 32'hca00c6f6;
    ram_cell[   48691] = 32'h65d1e8a0;
    ram_cell[   48692] = 32'hc41080d1;
    ram_cell[   48693] = 32'h9c32f6e3;
    ram_cell[   48694] = 32'had41df6b;
    ram_cell[   48695] = 32'h433df312;
    ram_cell[   48696] = 32'ha23f7c5d;
    ram_cell[   48697] = 32'h7a48dde2;
    ram_cell[   48698] = 32'h3b35db74;
    ram_cell[   48699] = 32'h22eb2cb7;
    ram_cell[   48700] = 32'h4136d3da;
    ram_cell[   48701] = 32'h946ae063;
    ram_cell[   48702] = 32'h2f6d6ad2;
    ram_cell[   48703] = 32'h2443e425;
    ram_cell[   48704] = 32'hdc67f720;
    ram_cell[   48705] = 32'hd91d8d40;
    ram_cell[   48706] = 32'he8d17117;
    ram_cell[   48707] = 32'h9097f8c1;
    ram_cell[   48708] = 32'h39d41c6f;
    ram_cell[   48709] = 32'hd817eac5;
    ram_cell[   48710] = 32'h5ff4ce42;
    ram_cell[   48711] = 32'hb82376fe;
    ram_cell[   48712] = 32'h51b7672d;
    ram_cell[   48713] = 32'he82b605d;
    ram_cell[   48714] = 32'h68f87ecb;
    ram_cell[   48715] = 32'hcfa0992a;
    ram_cell[   48716] = 32'he57764c6;
    ram_cell[   48717] = 32'h08d64a63;
    ram_cell[   48718] = 32'h629143da;
    ram_cell[   48719] = 32'h64aae6cf;
    ram_cell[   48720] = 32'h2f97ecb2;
    ram_cell[   48721] = 32'h9fa591ed;
    ram_cell[   48722] = 32'h2f092432;
    ram_cell[   48723] = 32'hb3215a6b;
    ram_cell[   48724] = 32'h8a8884c2;
    ram_cell[   48725] = 32'hfe8deae8;
    ram_cell[   48726] = 32'h44865150;
    ram_cell[   48727] = 32'h563ebd67;
    ram_cell[   48728] = 32'h68e34a80;
    ram_cell[   48729] = 32'h8b616a04;
    ram_cell[   48730] = 32'h313a72f1;
    ram_cell[   48731] = 32'hd36790b6;
    ram_cell[   48732] = 32'hc79d5bda;
    ram_cell[   48733] = 32'h6ab979f4;
    ram_cell[   48734] = 32'hb8ffde76;
    ram_cell[   48735] = 32'h57149461;
    ram_cell[   48736] = 32'h4e87d1f8;
    ram_cell[   48737] = 32'ha1aa686d;
    ram_cell[   48738] = 32'h3b57b196;
    ram_cell[   48739] = 32'h66154deb;
    ram_cell[   48740] = 32'ha1afbf21;
    ram_cell[   48741] = 32'hef801d81;
    ram_cell[   48742] = 32'h3d768fc3;
    ram_cell[   48743] = 32'h59d9434e;
    ram_cell[   48744] = 32'hf6423f6a;
    ram_cell[   48745] = 32'hbdda6c75;
    ram_cell[   48746] = 32'hcc8481a6;
    ram_cell[   48747] = 32'h378f0ba9;
    ram_cell[   48748] = 32'he0780d78;
    ram_cell[   48749] = 32'h7945afa3;
    ram_cell[   48750] = 32'hfedc0473;
    ram_cell[   48751] = 32'h7fcf973d;
    ram_cell[   48752] = 32'hde2e58de;
    ram_cell[   48753] = 32'h0e0b9af7;
    ram_cell[   48754] = 32'h2723c1ec;
    ram_cell[   48755] = 32'haf7b402c;
    ram_cell[   48756] = 32'h82ddf8cf;
    ram_cell[   48757] = 32'h74ff7e89;
    ram_cell[   48758] = 32'h3ae6b3c8;
    ram_cell[   48759] = 32'h0f12b36a;
    ram_cell[   48760] = 32'ha651aeed;
    ram_cell[   48761] = 32'h9889f848;
    ram_cell[   48762] = 32'h5e58a6a6;
    ram_cell[   48763] = 32'haf77dacc;
    ram_cell[   48764] = 32'hbf8b9c4f;
    ram_cell[   48765] = 32'h8d86a86b;
    ram_cell[   48766] = 32'h52256d2c;
    ram_cell[   48767] = 32'h1bd2b347;
    ram_cell[   48768] = 32'hd1a459fb;
    ram_cell[   48769] = 32'h0213e6d3;
    ram_cell[   48770] = 32'hc47bb98d;
    ram_cell[   48771] = 32'hcd3f487e;
    ram_cell[   48772] = 32'hf6d70e90;
    ram_cell[   48773] = 32'h796a9f11;
    ram_cell[   48774] = 32'h927825aa;
    ram_cell[   48775] = 32'he0b63f1f;
    ram_cell[   48776] = 32'h698e8ebe;
    ram_cell[   48777] = 32'h3ceeb098;
    ram_cell[   48778] = 32'hd0853654;
    ram_cell[   48779] = 32'hccbc5b85;
    ram_cell[   48780] = 32'h172c85da;
    ram_cell[   48781] = 32'hf41c3d19;
    ram_cell[   48782] = 32'h60f86c8c;
    ram_cell[   48783] = 32'he62b71aa;
    ram_cell[   48784] = 32'hbae53669;
    ram_cell[   48785] = 32'h7d21d6d4;
    ram_cell[   48786] = 32'h73ced026;
    ram_cell[   48787] = 32'h837bba06;
    ram_cell[   48788] = 32'he1637c2c;
    ram_cell[   48789] = 32'hc594c7c6;
    ram_cell[   48790] = 32'hc5986987;
    ram_cell[   48791] = 32'h43c5ff4b;
    ram_cell[   48792] = 32'h33e58008;
    ram_cell[   48793] = 32'hccbe4afb;
    ram_cell[   48794] = 32'h5bc6fc99;
    ram_cell[   48795] = 32'he9bfb5ca;
    ram_cell[   48796] = 32'h6bb19cd8;
    ram_cell[   48797] = 32'h2daf4b64;
    ram_cell[   48798] = 32'he1d2e028;
    ram_cell[   48799] = 32'h1c1ac92a;
    ram_cell[   48800] = 32'h9a645419;
    ram_cell[   48801] = 32'h5ac2eb79;
    ram_cell[   48802] = 32'h32de09b5;
    ram_cell[   48803] = 32'hbbab411f;
    ram_cell[   48804] = 32'h8020315b;
    ram_cell[   48805] = 32'h1626f50e;
    ram_cell[   48806] = 32'hf79432c5;
    ram_cell[   48807] = 32'h53ea459a;
    ram_cell[   48808] = 32'h4270c000;
    ram_cell[   48809] = 32'hd615d0d0;
    ram_cell[   48810] = 32'h20a5d52d;
    ram_cell[   48811] = 32'h7f58cde3;
    ram_cell[   48812] = 32'h21f56dfd;
    ram_cell[   48813] = 32'he9bb6c3e;
    ram_cell[   48814] = 32'he4331497;
    ram_cell[   48815] = 32'h427bbb98;
    ram_cell[   48816] = 32'ha05704ad;
    ram_cell[   48817] = 32'h13e397fc;
    ram_cell[   48818] = 32'h2457829b;
    ram_cell[   48819] = 32'hb3518250;
    ram_cell[   48820] = 32'hba206d76;
    ram_cell[   48821] = 32'h0ddfe124;
    ram_cell[   48822] = 32'h2bcb292b;
    ram_cell[   48823] = 32'h1cf12cbf;
    ram_cell[   48824] = 32'h2a0ea0fd;
    ram_cell[   48825] = 32'h3f01cd83;
    ram_cell[   48826] = 32'h538d324b;
    ram_cell[   48827] = 32'h665e9ab6;
    ram_cell[   48828] = 32'h1cd3cc0a;
    ram_cell[   48829] = 32'hd1370c94;
    ram_cell[   48830] = 32'hd2e67863;
    ram_cell[   48831] = 32'h54699195;
    ram_cell[   48832] = 32'h682125da;
    ram_cell[   48833] = 32'h46153b26;
    ram_cell[   48834] = 32'ha17ce673;
    ram_cell[   48835] = 32'h71c5bfe1;
    ram_cell[   48836] = 32'hb645eb40;
    ram_cell[   48837] = 32'h231fb354;
    ram_cell[   48838] = 32'hf22baca5;
    ram_cell[   48839] = 32'hd55454c9;
    ram_cell[   48840] = 32'hbeffe80d;
    ram_cell[   48841] = 32'h061baa0a;
    ram_cell[   48842] = 32'h414edbd8;
    ram_cell[   48843] = 32'haa938486;
    ram_cell[   48844] = 32'h193986e8;
    ram_cell[   48845] = 32'h2492e150;
    ram_cell[   48846] = 32'h7565d32e;
    ram_cell[   48847] = 32'h73a7322c;
    ram_cell[   48848] = 32'h0308e062;
    ram_cell[   48849] = 32'h1569d28e;
    ram_cell[   48850] = 32'h76a5db30;
    ram_cell[   48851] = 32'h7c5db9d0;
    ram_cell[   48852] = 32'h11d4661c;
    ram_cell[   48853] = 32'h61c4cf30;
    ram_cell[   48854] = 32'h0430e9e0;
    ram_cell[   48855] = 32'h2f0ab98d;
    ram_cell[   48856] = 32'h7e802052;
    ram_cell[   48857] = 32'h54456c71;
    ram_cell[   48858] = 32'h12e7b439;
    ram_cell[   48859] = 32'hdfdd2b0b;
    ram_cell[   48860] = 32'hfeb0b985;
    ram_cell[   48861] = 32'hf9180e86;
    ram_cell[   48862] = 32'ha7f06c4c;
    ram_cell[   48863] = 32'h4efcbe89;
    ram_cell[   48864] = 32'hae9c3803;
    ram_cell[   48865] = 32'h75243895;
    ram_cell[   48866] = 32'h7164ec72;
    ram_cell[   48867] = 32'h1dd81327;
    ram_cell[   48868] = 32'h578f4b96;
    ram_cell[   48869] = 32'hd1962e87;
    ram_cell[   48870] = 32'h21777eca;
    ram_cell[   48871] = 32'h62dd5b2c;
    ram_cell[   48872] = 32'h948c2914;
    ram_cell[   48873] = 32'h21457f8d;
    ram_cell[   48874] = 32'hdaf51f09;
    ram_cell[   48875] = 32'h2ecdb426;
    ram_cell[   48876] = 32'h1d5ae8a7;
    ram_cell[   48877] = 32'h0a414e5a;
    ram_cell[   48878] = 32'h25006be0;
    ram_cell[   48879] = 32'hc6ae5b55;
    ram_cell[   48880] = 32'h383aec49;
    ram_cell[   48881] = 32'haae9fc7f;
    ram_cell[   48882] = 32'h4ae90ae8;
    ram_cell[   48883] = 32'h23c9c219;
    ram_cell[   48884] = 32'hf3c54d11;
    ram_cell[   48885] = 32'h416f1f67;
    ram_cell[   48886] = 32'h0f68f14b;
    ram_cell[   48887] = 32'h7f920f74;
    ram_cell[   48888] = 32'h132f7e48;
    ram_cell[   48889] = 32'hb9366a65;
    ram_cell[   48890] = 32'hfcd4810b;
    ram_cell[   48891] = 32'hf186c366;
    ram_cell[   48892] = 32'ha64681ff;
    ram_cell[   48893] = 32'h4209bb55;
    ram_cell[   48894] = 32'hde964462;
    ram_cell[   48895] = 32'h0c2b846d;
    ram_cell[   48896] = 32'h46f813fd;
    ram_cell[   48897] = 32'hc0fae3da;
    ram_cell[   48898] = 32'hef505a67;
    ram_cell[   48899] = 32'h20dc0428;
    ram_cell[   48900] = 32'h4414266c;
    ram_cell[   48901] = 32'hc63e3cb9;
    ram_cell[   48902] = 32'h901e887b;
    ram_cell[   48903] = 32'h86e2ee6b;
    ram_cell[   48904] = 32'hdf78c9a1;
    ram_cell[   48905] = 32'hde2d8573;
    ram_cell[   48906] = 32'h6b1e6755;
    ram_cell[   48907] = 32'hf198d931;
    ram_cell[   48908] = 32'h0664e673;
    ram_cell[   48909] = 32'h28415551;
    ram_cell[   48910] = 32'hf7ab1dab;
    ram_cell[   48911] = 32'h2ce3ecb5;
    ram_cell[   48912] = 32'h2a41f25c;
    ram_cell[   48913] = 32'h5a57c079;
    ram_cell[   48914] = 32'h3f49f560;
    ram_cell[   48915] = 32'hf449f38f;
    ram_cell[   48916] = 32'hb854bbe4;
    ram_cell[   48917] = 32'hcce8d20a;
    ram_cell[   48918] = 32'h9caf1550;
    ram_cell[   48919] = 32'h8672e9af;
    ram_cell[   48920] = 32'h5994caa8;
    ram_cell[   48921] = 32'hc465de85;
    ram_cell[   48922] = 32'he44ca828;
    ram_cell[   48923] = 32'hab88a1b9;
    ram_cell[   48924] = 32'hb7b4c5ed;
    ram_cell[   48925] = 32'h0bc0a12c;
    ram_cell[   48926] = 32'haedc3f63;
    ram_cell[   48927] = 32'h744e5a9f;
    ram_cell[   48928] = 32'h4bf7718f;
    ram_cell[   48929] = 32'h65763617;
    ram_cell[   48930] = 32'h6c0b244b;
    ram_cell[   48931] = 32'hadd23a9c;
    ram_cell[   48932] = 32'h58700c58;
    ram_cell[   48933] = 32'h4301d752;
    ram_cell[   48934] = 32'h620b77d5;
    ram_cell[   48935] = 32'h6b853f5e;
    ram_cell[   48936] = 32'h5281f830;
    ram_cell[   48937] = 32'h1c5b5489;
    ram_cell[   48938] = 32'hf638039e;
    ram_cell[   48939] = 32'hcdb85feb;
    ram_cell[   48940] = 32'h538ae2e3;
    ram_cell[   48941] = 32'h4459f744;
    ram_cell[   48942] = 32'h471e38c6;
    ram_cell[   48943] = 32'h2ae44041;
    ram_cell[   48944] = 32'h6c6485e4;
    ram_cell[   48945] = 32'h517fa25d;
    ram_cell[   48946] = 32'hdfae8fdd;
    ram_cell[   48947] = 32'h7ab4670f;
    ram_cell[   48948] = 32'h50179072;
    ram_cell[   48949] = 32'h391ad3b2;
    ram_cell[   48950] = 32'h80439358;
    ram_cell[   48951] = 32'h36d87ecf;
    ram_cell[   48952] = 32'he2806b18;
    ram_cell[   48953] = 32'hadb58262;
    ram_cell[   48954] = 32'had3e0cf1;
    ram_cell[   48955] = 32'h07c10e11;
    ram_cell[   48956] = 32'h04e3588b;
    ram_cell[   48957] = 32'h06a515af;
    ram_cell[   48958] = 32'h18b2636f;
    ram_cell[   48959] = 32'h2ea47d43;
    ram_cell[   48960] = 32'h736dc4fe;
    ram_cell[   48961] = 32'h834fd837;
    ram_cell[   48962] = 32'hcb1dd746;
    ram_cell[   48963] = 32'h6cd5e654;
    ram_cell[   48964] = 32'h9beaed7f;
    ram_cell[   48965] = 32'h76805dee;
    ram_cell[   48966] = 32'hbfe7b9d5;
    ram_cell[   48967] = 32'h2ea232be;
    ram_cell[   48968] = 32'h37dde185;
    ram_cell[   48969] = 32'h54a5380f;
    ram_cell[   48970] = 32'he7aab967;
    ram_cell[   48971] = 32'h917aa1c5;
    ram_cell[   48972] = 32'h57ff6366;
    ram_cell[   48973] = 32'hbeabfe9d;
    ram_cell[   48974] = 32'h7789f7ca;
    ram_cell[   48975] = 32'h148d9dea;
    ram_cell[   48976] = 32'he24df9a5;
    ram_cell[   48977] = 32'hd20c564b;
    ram_cell[   48978] = 32'h49c7dc80;
    ram_cell[   48979] = 32'h16e368b5;
    ram_cell[   48980] = 32'hcfc8ed1d;
    ram_cell[   48981] = 32'hf9c3f4fd;
    ram_cell[   48982] = 32'hde8d2701;
    ram_cell[   48983] = 32'h91c32718;
    ram_cell[   48984] = 32'h851c95d4;
    ram_cell[   48985] = 32'h51afcbf5;
    ram_cell[   48986] = 32'hf2eefff4;
    ram_cell[   48987] = 32'hc49c9ee7;
    ram_cell[   48988] = 32'hed4923bb;
    ram_cell[   48989] = 32'h0d4d45d9;
    ram_cell[   48990] = 32'h283e023f;
    ram_cell[   48991] = 32'h010ea86e;
    ram_cell[   48992] = 32'h3e050440;
    ram_cell[   48993] = 32'hf6a0d912;
    ram_cell[   48994] = 32'haf1399d2;
    ram_cell[   48995] = 32'h3bb573a5;
    ram_cell[   48996] = 32'h02e508a6;
    ram_cell[   48997] = 32'hb0abd8c6;
    ram_cell[   48998] = 32'hd704f5a8;
    ram_cell[   48999] = 32'h5897e127;
    ram_cell[   49000] = 32'h85133597;
    ram_cell[   49001] = 32'h276dfb60;
    ram_cell[   49002] = 32'h208f4e03;
    ram_cell[   49003] = 32'hb496ecd4;
    ram_cell[   49004] = 32'hf69784dc;
    ram_cell[   49005] = 32'hc19a92aa;
    ram_cell[   49006] = 32'h76035bb2;
    ram_cell[   49007] = 32'h470ede37;
    ram_cell[   49008] = 32'h7e3416e0;
    ram_cell[   49009] = 32'hbe1d258a;
    ram_cell[   49010] = 32'h7eb85e31;
    ram_cell[   49011] = 32'h297a2708;
    ram_cell[   49012] = 32'h1eece695;
    ram_cell[   49013] = 32'h313e1fa8;
    ram_cell[   49014] = 32'hb4e4b805;
    ram_cell[   49015] = 32'h03d52185;
    ram_cell[   49016] = 32'h28f9135e;
    ram_cell[   49017] = 32'hc8e6f8bc;
    ram_cell[   49018] = 32'h1f8532e9;
    ram_cell[   49019] = 32'hd1a1fdfd;
    ram_cell[   49020] = 32'hb395abb9;
    ram_cell[   49021] = 32'hfb28425b;
    ram_cell[   49022] = 32'hf1b5aac0;
    ram_cell[   49023] = 32'h2e6281f1;
    ram_cell[   49024] = 32'h8cefe31b;
    ram_cell[   49025] = 32'hae52839a;
    ram_cell[   49026] = 32'h51b7ff0d;
    ram_cell[   49027] = 32'hae863854;
    ram_cell[   49028] = 32'h51e30a84;
    ram_cell[   49029] = 32'ha5d3dbae;
    ram_cell[   49030] = 32'h9fdb05f1;
    ram_cell[   49031] = 32'h1683de45;
    ram_cell[   49032] = 32'haf3f416d;
    ram_cell[   49033] = 32'h370836c0;
    ram_cell[   49034] = 32'hfb3eaa66;
    ram_cell[   49035] = 32'h1f3b75ae;
    ram_cell[   49036] = 32'h643977e5;
    ram_cell[   49037] = 32'h70f8db71;
    ram_cell[   49038] = 32'h4e580883;
    ram_cell[   49039] = 32'he6d6215c;
    ram_cell[   49040] = 32'h0b678a4e;
    ram_cell[   49041] = 32'hebbadc5f;
    ram_cell[   49042] = 32'h1445985d;
    ram_cell[   49043] = 32'h9445aaee;
    ram_cell[   49044] = 32'h98af1ea0;
    ram_cell[   49045] = 32'h4eb82aa4;
    ram_cell[   49046] = 32'h6a335fc6;
    ram_cell[   49047] = 32'hf9beca98;
    ram_cell[   49048] = 32'h52e1fa9a;
    ram_cell[   49049] = 32'h7387a508;
    ram_cell[   49050] = 32'h7eecd02e;
    ram_cell[   49051] = 32'h93adfab0;
    ram_cell[   49052] = 32'hba48bbef;
    ram_cell[   49053] = 32'h5a0f33bd;
    ram_cell[   49054] = 32'he0a8e924;
    ram_cell[   49055] = 32'h07816c90;
    ram_cell[   49056] = 32'hb3cc9584;
    ram_cell[   49057] = 32'heb978076;
    ram_cell[   49058] = 32'h6a58f039;
    ram_cell[   49059] = 32'h5d8019db;
    ram_cell[   49060] = 32'h74e9cd28;
    ram_cell[   49061] = 32'h488f9fe4;
    ram_cell[   49062] = 32'h6ee9f88f;
    ram_cell[   49063] = 32'h358a11c8;
    ram_cell[   49064] = 32'hb7b092fd;
    ram_cell[   49065] = 32'h1a3fa3af;
    ram_cell[   49066] = 32'h221ea8c8;
    ram_cell[   49067] = 32'hdd935d14;
    ram_cell[   49068] = 32'h94424511;
    ram_cell[   49069] = 32'he9ebd685;
    ram_cell[   49070] = 32'h7aae34f9;
    ram_cell[   49071] = 32'h58f93bcd;
    ram_cell[   49072] = 32'h401a11de;
    ram_cell[   49073] = 32'h47c97e82;
    ram_cell[   49074] = 32'h3eab39f9;
    ram_cell[   49075] = 32'h07e25f16;
    ram_cell[   49076] = 32'ha2c99014;
    ram_cell[   49077] = 32'h5aced5ef;
    ram_cell[   49078] = 32'h8652ffc7;
    ram_cell[   49079] = 32'h924d3434;
    ram_cell[   49080] = 32'h834764b6;
    ram_cell[   49081] = 32'h35f668b2;
    ram_cell[   49082] = 32'h0ed73feb;
    ram_cell[   49083] = 32'h4d4d3b6b;
    ram_cell[   49084] = 32'hfc3c360d;
    ram_cell[   49085] = 32'h105b04ff;
    ram_cell[   49086] = 32'hf69e7227;
    ram_cell[   49087] = 32'h1a0fb3e1;
    ram_cell[   49088] = 32'hb81d779a;
    ram_cell[   49089] = 32'h1ff56088;
    ram_cell[   49090] = 32'hcafaf8ca;
    ram_cell[   49091] = 32'h2ca8edaf;
    ram_cell[   49092] = 32'h0f463898;
    ram_cell[   49093] = 32'h19d939d7;
    ram_cell[   49094] = 32'hc1b91dfe;
    ram_cell[   49095] = 32'hf1a486c2;
    ram_cell[   49096] = 32'h3de4c850;
    ram_cell[   49097] = 32'h3180cd7a;
    ram_cell[   49098] = 32'h9a9e86f9;
    ram_cell[   49099] = 32'h73e55d32;
    ram_cell[   49100] = 32'h5a28946a;
    ram_cell[   49101] = 32'h0e87af6a;
    ram_cell[   49102] = 32'h727b96c8;
    ram_cell[   49103] = 32'h8445a308;
    ram_cell[   49104] = 32'h949aeb3c;
    ram_cell[   49105] = 32'h4c0a4ca1;
    ram_cell[   49106] = 32'h44c3c141;
    ram_cell[   49107] = 32'hc47e20a0;
    ram_cell[   49108] = 32'hef156835;
    ram_cell[   49109] = 32'h11cbeafb;
    ram_cell[   49110] = 32'h64fa61ad;
    ram_cell[   49111] = 32'ha0970007;
    ram_cell[   49112] = 32'h624e5591;
    ram_cell[   49113] = 32'he4ad5ca8;
    ram_cell[   49114] = 32'h74ff991b;
    ram_cell[   49115] = 32'he78561b2;
    ram_cell[   49116] = 32'h4979714c;
    ram_cell[   49117] = 32'h6239ed45;
    ram_cell[   49118] = 32'h51a9049a;
    ram_cell[   49119] = 32'hdc5aec9a;
    ram_cell[   49120] = 32'h36300352;
    ram_cell[   49121] = 32'hed6c2bdc;
    ram_cell[   49122] = 32'h48fb01a6;
    ram_cell[   49123] = 32'hf2463cd1;
    ram_cell[   49124] = 32'h1a3e7fb1;
    ram_cell[   49125] = 32'h33cb95cd;
    ram_cell[   49126] = 32'h7366e868;
    ram_cell[   49127] = 32'hed3f49ef;
    ram_cell[   49128] = 32'h4ecf5efc;
    ram_cell[   49129] = 32'hed671eff;
    ram_cell[   49130] = 32'hbbdaeb77;
    ram_cell[   49131] = 32'h48723519;
    ram_cell[   49132] = 32'h207ee6b2;
    ram_cell[   49133] = 32'h08cc1eec;
    ram_cell[   49134] = 32'haf5157b2;
    ram_cell[   49135] = 32'h9f1e42d7;
    ram_cell[   49136] = 32'hb2f0fed8;
    ram_cell[   49137] = 32'h42b79300;
    ram_cell[   49138] = 32'hed5bf19f;
    ram_cell[   49139] = 32'h8b09fe34;
    ram_cell[   49140] = 32'h914a8426;
    ram_cell[   49141] = 32'h7fe3d5aa;
    ram_cell[   49142] = 32'h20eddf8f;
    ram_cell[   49143] = 32'h2fdd1e5f;
    ram_cell[   49144] = 32'h82e2bd5e;
    ram_cell[   49145] = 32'hcbfdd12e;
    ram_cell[   49146] = 32'h227f5bfa;
    ram_cell[   49147] = 32'h73e8ae64;
    ram_cell[   49148] = 32'h1cb528b9;
    ram_cell[   49149] = 32'h924a81d0;
    ram_cell[   49150] = 32'h6690b5d3;
    ram_cell[   49151] = 32'h74faeac5;
end

endmodule

